VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gpio_signal_buffering
  CLASS BLOCK ;
  FOREIGN gpio_signal_buffering ;
  ORIGIN 0.000 0.000 ;
  SIZE 3588.000 BY 5188.000 ;
  PIN mgmt_io_in_unbuf[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2082.940 4983.335 2084.530 4983.535 ;
      LAYER mcon ;
        RECT 2082.940 4983.365 2084.030 4983.535 ;
      LAYER met1 ;
        RECT 2082.880 4983.315 2084.090 4983.575 ;
        RECT 2083.245 4976.235 2083.565 4976.355 ;
        RECT 2079.535 4976.095 2083.565 4976.235 ;
      LAYER via ;
        RECT 2082.940 4983.315 2084.030 4983.575 ;
        RECT 2083.275 4976.095 2083.535 4976.355 ;
      LAYER met2 ;
        RECT 2082.940 4983.285 2084.030 4983.605 ;
        RECT 2083.395 4976.385 2083.535 4983.285 ;
        RECT 2083.275 4976.065 2083.535 4976.385 ;
        RECT 2083.395 4975.645 2083.535 4976.065 ;
    END
  END mgmt_io_in_unbuf[18]
  PIN mgmt_io_out_buf[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2084.265 4986.965 2084.435 4987.445 ;
        RECT 2085.105 4986.965 2085.275 4987.445 ;
        RECT 2085.945 4986.965 2086.115 4987.445 ;
        RECT 2086.785 4986.965 2086.955 4987.445 ;
        RECT 2084.265 4986.795 2086.955 4986.965 ;
        RECT 2084.265 4986.255 2084.520 4986.795 ;
        RECT 2084.265 4986.085 2086.955 4986.255 ;
        RECT 2084.265 4985.235 2084.435 4986.085 ;
        RECT 2085.105 4985.235 2085.275 4986.085 ;
        RECT 2085.945 4985.235 2086.115 4986.085 ;
        RECT 2086.785 4985.235 2086.955 4986.085 ;
      LAYER mcon ;
        RECT 2084.350 4986.085 2084.520 4986.935 ;
      LAYER met1 ;
        RECT 2084.310 4986.025 2084.570 4986.995 ;
        RECT 2084.215 4975.955 2084.535 4976.075 ;
        RECT 2080.535 4975.815 2084.535 4975.955 ;
      LAYER via ;
        RECT 2084.310 4986.085 2084.570 4986.935 ;
        RECT 2084.245 4975.815 2084.505 4976.075 ;
      LAYER met2 ;
        RECT 2084.280 4986.085 2084.600 4986.935 ;
        RECT 2084.365 4976.105 2084.505 4986.085 ;
        RECT 2084.245 4975.785 2084.505 4976.105 ;
        RECT 2084.365 4975.645 2084.505 4975.785 ;
    END
  END mgmt_io_out_buf[18]
  PIN mgmt_io_out_buf[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3320.250 4986.555 3320.420 4987.035 ;
        RECT 3321.090 4986.555 3321.260 4987.035 ;
        RECT 3321.930 4986.555 3322.100 4987.035 ;
        RECT 3322.770 4986.555 3322.940 4987.035 ;
        RECT 3320.250 4986.385 3322.940 4986.555 ;
        RECT 3320.250 4985.845 3320.505 4986.385 ;
        RECT 3320.250 4985.675 3322.940 4985.845 ;
        RECT 3320.250 4984.825 3320.420 4985.675 ;
        RECT 3321.090 4984.825 3321.260 4985.675 ;
        RECT 3321.930 4984.825 3322.100 4985.675 ;
        RECT 3322.770 4984.825 3322.940 4985.675 ;
      LAYER mcon ;
        RECT 3320.335 4985.675 3320.505 4986.525 ;
      LAYER met1 ;
        RECT 3320.295 4985.615 3320.555 4986.585 ;
        RECT 3320.200 4975.395 3320.520 4975.515 ;
        RECT 3305.615 4975.255 3320.520 4975.395 ;
      LAYER via ;
        RECT 3320.295 4985.675 3320.555 4986.525 ;
        RECT 3320.230 4975.255 3320.490 4975.515 ;
      LAYER met2 ;
        RECT 3320.265 4985.675 3320.585 4986.525 ;
        RECT 3320.350 4975.545 3320.490 4985.675 ;
        RECT 3320.230 4975.225 3320.490 4975.545 ;
        RECT 3320.350 4973.965 3320.490 4975.225 ;
    END
  END mgmt_io_out_buf[17]
  PIN mgmt_io_out_buf[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3326.230 4986.555 3326.400 4987.035 ;
        RECT 3327.070 4986.555 3327.240 4987.035 ;
        RECT 3327.910 4986.555 3328.080 4987.035 ;
        RECT 3328.750 4986.555 3328.920 4987.035 ;
        RECT 3326.230 4986.385 3328.920 4986.555 ;
        RECT 3326.230 4985.845 3326.485 4986.385 ;
        RECT 3326.230 4985.675 3328.920 4985.845 ;
        RECT 3326.230 4984.825 3326.400 4985.675 ;
        RECT 3327.070 4984.825 3327.240 4985.675 ;
        RECT 3327.910 4984.825 3328.080 4985.675 ;
        RECT 3328.750 4984.825 3328.920 4985.675 ;
      LAYER mcon ;
        RECT 3326.315 4985.675 3326.485 4986.525 ;
      LAYER met1 ;
        RECT 3326.275 4985.615 3326.535 4986.585 ;
        RECT 3326.180 4974.835 3326.500 4974.955 ;
        RECT 3307.615 4974.695 3326.500 4974.835 ;
      LAYER via ;
        RECT 3326.275 4985.675 3326.535 4986.525 ;
        RECT 3326.210 4974.695 3326.470 4974.955 ;
      LAYER met2 ;
        RECT 3326.245 4985.675 3326.565 4986.525 ;
        RECT 3326.330 4974.985 3326.470 4985.675 ;
        RECT 3326.210 4974.665 3326.470 4974.985 ;
        RECT 3326.330 4973.965 3326.470 4974.665 ;
    END
  END mgmt_io_out_buf[16]
  PIN mgmt_io_in_unbuf[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3318.925 4982.925 3320.515 4983.125 ;
      LAYER mcon ;
        RECT 3318.925 4982.955 3320.015 4983.125 ;
      LAYER met1 ;
        RECT 3318.865 4982.905 3320.075 4983.165 ;
        RECT 3319.230 4975.675 3319.550 4975.795 ;
        RECT 3304.615 4975.535 3319.550 4975.675 ;
      LAYER via ;
        RECT 3318.925 4982.905 3320.015 4983.165 ;
        RECT 3319.260 4975.535 3319.520 4975.795 ;
      LAYER met2 ;
        RECT 3318.925 4982.875 3320.015 4983.195 ;
        RECT 3319.380 4975.825 3319.520 4982.875 ;
        RECT 3319.260 4975.505 3319.520 4975.825 ;
        RECT 3319.380 4973.965 3319.520 4975.505 ;
    END
  END mgmt_io_in_unbuf[17]
  PIN mgmt_io_in_unbuf[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3324.905 4982.925 3326.495 4983.125 ;
      LAYER mcon ;
        RECT 3324.905 4982.955 3325.995 4983.125 ;
      LAYER met1 ;
        RECT 3324.845 4982.905 3326.055 4983.165 ;
        RECT 3325.210 4975.115 3325.530 4975.235 ;
        RECT 3306.615 4974.975 3325.530 4975.115 ;
      LAYER via ;
        RECT 3324.905 4982.905 3325.995 4983.165 ;
        RECT 3325.240 4974.975 3325.500 4975.235 ;
      LAYER met2 ;
        RECT 3324.905 4982.875 3325.995 4983.195 ;
        RECT 3325.360 4975.265 3325.500 4982.875 ;
        RECT 3325.240 4974.945 3325.500 4975.265 ;
        RECT 3325.360 4973.965 3325.500 4974.945 ;
    END
  END mgmt_io_in_unbuf[16]
  PIN mgmt_io_in_unbuf[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3330.885 4982.925 3332.475 4983.125 ;
      LAYER mcon ;
        RECT 3330.885 4982.955 3331.975 4983.125 ;
      LAYER met1 ;
        RECT 3330.825 4982.905 3332.035 4983.165 ;
        RECT 3331.190 4974.555 3331.510 4974.675 ;
        RECT 3308.615 4974.415 3331.510 4974.555 ;
      LAYER via ;
        RECT 3330.885 4982.905 3331.975 4983.165 ;
        RECT 3331.220 4974.415 3331.480 4974.675 ;
      LAYER met2 ;
        RECT 3330.885 4982.875 3331.975 4983.195 ;
        RECT 3331.340 4974.705 3331.480 4982.875 ;
        RECT 3331.220 4974.385 3331.480 4974.705 ;
        RECT 3331.340 4973.965 3331.480 4974.385 ;
    END
  END mgmt_io_in_unbuf[15]
  PIN mgmt_io_out_buf[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3332.210 4986.555 3332.380 4987.035 ;
        RECT 3333.050 4986.555 3333.220 4987.035 ;
        RECT 3333.890 4986.555 3334.060 4987.035 ;
        RECT 3334.730 4986.555 3334.900 4987.035 ;
        RECT 3332.210 4986.385 3334.900 4986.555 ;
        RECT 3332.210 4985.845 3332.465 4986.385 ;
        RECT 3332.210 4985.675 3334.900 4985.845 ;
        RECT 3332.210 4984.825 3332.380 4985.675 ;
        RECT 3333.050 4984.825 3333.220 4985.675 ;
        RECT 3333.890 4984.825 3334.060 4985.675 ;
        RECT 3334.730 4984.825 3334.900 4985.675 ;
      LAYER mcon ;
        RECT 3332.295 4985.675 3332.465 4986.525 ;
      LAYER met1 ;
        RECT 3332.255 4985.615 3332.515 4986.585 ;
        RECT 3332.160 4974.275 3332.480 4974.395 ;
        RECT 3309.615 4974.135 3332.480 4974.275 ;
      LAYER via ;
        RECT 3332.255 4985.675 3332.515 4986.525 ;
        RECT 3332.190 4974.135 3332.450 4974.395 ;
      LAYER met2 ;
        RECT 3332.225 4985.675 3332.545 4986.525 ;
        RECT 3332.310 4974.425 3332.450 4985.675 ;
        RECT 3332.190 4974.105 3332.450 4974.425 ;
        RECT 3332.310 4973.965 3332.450 4974.105 ;
    END
  END mgmt_io_out_buf[15]
  PIN mgmt_io_in_unbuf[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.660 3546.780 3384.860 3548.370 ;
      LAYER mcon ;
        RECT 3384.690 3547.280 3384.860 3548.370 ;
      LAYER met1 ;
        RECT 3373.220 3548.065 3373.360 3577.605 ;
        RECT 3373.220 3547.745 3373.480 3548.065 ;
        RECT 3384.640 3547.220 3384.900 3548.430 ;
      LAYER via ;
        RECT 3373.220 3547.775 3373.480 3548.035 ;
        RECT 3384.640 3547.280 3384.900 3548.370 ;
      LAYER met2 ;
        RECT 3373.190 3547.915 3373.510 3548.035 ;
        RECT 3384.610 3547.915 3384.930 3548.370 ;
        RECT 3372.210 3547.775 3384.930 3547.915 ;
        RECT 3384.610 3547.280 3384.930 3547.775 ;
    END
  END mgmt_io_in_unbuf[14]
  PIN mgmt_io_in_unbuf[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.660 3540.800 3384.860 3542.390 ;
      LAYER mcon ;
        RECT 3384.690 3541.300 3384.860 3542.390 ;
      LAYER met1 ;
        RECT 3372.660 3542.085 3372.800 3575.605 ;
        RECT 3372.660 3541.765 3372.920 3542.085 ;
        RECT 3384.640 3541.240 3384.900 3542.450 ;
      LAYER via ;
        RECT 3372.660 3541.795 3372.920 3542.055 ;
        RECT 3384.640 3541.300 3384.900 3542.390 ;
      LAYER met2 ;
        RECT 3372.630 3541.935 3372.950 3542.055 ;
        RECT 3384.610 3541.935 3384.930 3542.390 ;
        RECT 3372.210 3541.795 3384.930 3541.935 ;
        RECT 3384.610 3541.300 3384.930 3541.795 ;
    END
  END mgmt_io_in_unbuf[13]
  PIN mgmt_io_out_buf[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3386.560 3546.875 3388.770 3547.045 ;
        RECT 3387.410 3546.790 3388.290 3546.875 ;
        RECT 3387.410 3546.205 3387.580 3546.790 ;
        RECT 3386.560 3546.035 3387.580 3546.205 ;
        RECT 3387.410 3545.365 3387.580 3546.035 ;
        RECT 3386.560 3545.195 3387.580 3545.365 ;
        RECT 3387.410 3544.525 3387.580 3545.195 ;
        RECT 3386.560 3544.355 3387.580 3544.525 ;
        RECT 3388.120 3546.205 3388.290 3546.790 ;
        RECT 3388.120 3546.035 3388.770 3546.205 ;
        RECT 3388.120 3545.365 3388.290 3546.035 ;
        RECT 3388.120 3545.195 3388.770 3545.365 ;
        RECT 3388.120 3544.525 3388.290 3545.195 ;
        RECT 3388.120 3544.355 3388.770 3544.525 ;
      LAYER met1 ;
        RECT 3372.940 3547.095 3373.080 3576.605 ;
        RECT 3372.940 3546.775 3373.200 3547.095 ;
        RECT 3387.350 3546.740 3388.320 3547.000 ;
      LAYER via ;
        RECT 3372.940 3546.805 3373.200 3547.065 ;
        RECT 3387.410 3546.740 3388.260 3547.000 ;
      LAYER met2 ;
        RECT 3372.910 3546.945 3373.230 3547.065 ;
        RECT 3387.410 3546.945 3388.260 3547.030 ;
        RECT 3372.210 3546.805 3388.260 3546.945 ;
        RECT 3387.410 3546.710 3388.260 3546.805 ;
    END
  END mgmt_io_out_buf[14]
  PIN mgmt_io_out_buf[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3386.560 3540.895 3388.770 3541.065 ;
        RECT 3387.410 3540.810 3388.290 3540.895 ;
        RECT 3387.410 3540.225 3387.580 3540.810 ;
        RECT 3386.560 3540.055 3387.580 3540.225 ;
        RECT 3387.410 3539.385 3387.580 3540.055 ;
        RECT 3386.560 3539.215 3387.580 3539.385 ;
        RECT 3387.410 3538.545 3387.580 3539.215 ;
        RECT 3386.560 3538.375 3387.580 3538.545 ;
        RECT 3388.120 3540.225 3388.290 3540.810 ;
        RECT 3388.120 3540.055 3388.770 3540.225 ;
        RECT 3388.120 3539.385 3388.290 3540.055 ;
        RECT 3388.120 3539.215 3388.770 3539.385 ;
        RECT 3388.120 3538.545 3388.290 3539.215 ;
        RECT 3388.120 3538.375 3388.770 3538.545 ;
      LAYER met1 ;
        RECT 3372.380 3541.115 3372.520 3574.605 ;
        RECT 3372.380 3540.795 3372.640 3541.115 ;
        RECT 3387.350 3540.760 3388.320 3541.020 ;
      LAYER via ;
        RECT 3372.380 3540.825 3372.640 3541.085 ;
        RECT 3387.410 3540.760 3388.260 3541.020 ;
      LAYER met2 ;
        RECT 3372.350 3540.965 3372.670 3541.085 ;
        RECT 3387.410 3540.965 3388.260 3541.050 ;
        RECT 3372.210 3540.825 3388.260 3540.965 ;
        RECT 3387.410 3540.730 3388.260 3540.825 ;
    END
  END mgmt_io_out_buf[13]
  PIN mgmt_io_in_unbuf[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.660 2230.700 3384.860 2232.290 ;
      LAYER mcon ;
        RECT 3384.690 2231.200 3384.860 2232.290 ;
      LAYER met1 ;
        RECT 3372.100 2231.985 3372.240 2281.275 ;
        RECT 3372.100 2231.665 3372.360 2231.985 ;
        RECT 3384.640 2231.140 3384.900 2232.350 ;
      LAYER via ;
        RECT 3372.100 2231.695 3372.360 2231.955 ;
        RECT 3384.640 2231.200 3384.900 2232.290 ;
      LAYER met2 ;
        RECT 3372.070 2231.835 3372.390 2231.955 ;
        RECT 3384.610 2231.835 3384.930 2232.290 ;
        RECT 3368.850 2231.695 3384.930 2231.835 ;
        RECT 3384.610 2231.200 3384.930 2231.695 ;
    END
  END mgmt_io_in_unbuf[12]
  PIN mgmt_io_in_unbuf[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.660 2224.720 3384.860 2226.310 ;
      LAYER mcon ;
        RECT 3384.690 2225.220 3384.860 2226.310 ;
      LAYER met1 ;
        RECT 3371.540 2226.005 3371.680 2279.275 ;
        RECT 3371.540 2225.685 3371.800 2226.005 ;
        RECT 3384.640 2225.160 3384.900 2226.370 ;
      LAYER via ;
        RECT 3371.540 2225.715 3371.800 2225.975 ;
        RECT 3384.640 2225.220 3384.900 2226.310 ;
      LAYER met2 ;
        RECT 3371.510 2225.855 3371.830 2225.975 ;
        RECT 3384.610 2225.855 3384.930 2226.310 ;
        RECT 3368.850 2225.715 3384.930 2225.855 ;
        RECT 3384.610 2225.220 3384.930 2225.715 ;
    END
  END mgmt_io_in_unbuf[11]
  PIN mgmt_io_in_unbuf[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.660 2218.740 3384.860 2220.330 ;
      LAYER mcon ;
        RECT 3384.690 2219.240 3384.860 2220.330 ;
      LAYER met1 ;
        RECT 3370.980 2220.025 3371.120 2277.275 ;
        RECT 3370.980 2219.705 3371.240 2220.025 ;
        RECT 3384.640 2219.180 3384.900 2220.390 ;
      LAYER via ;
        RECT 3370.980 2219.735 3371.240 2219.995 ;
        RECT 3384.640 2219.240 3384.900 2220.330 ;
      LAYER met2 ;
        RECT 3370.950 2219.875 3371.270 2219.995 ;
        RECT 3384.610 2219.875 3384.930 2220.330 ;
        RECT 3368.850 2219.735 3384.930 2219.875 ;
        RECT 3384.610 2219.240 3384.930 2219.735 ;
    END
  END mgmt_io_in_unbuf[10]
  PIN mgmt_io_in_unbuf[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.660 2212.760 3384.860 2214.350 ;
      LAYER mcon ;
        RECT 3384.690 2213.260 3384.860 2214.350 ;
      LAYER met1 ;
        RECT 3370.420 2214.045 3370.560 2275.275 ;
        RECT 3370.420 2213.725 3370.680 2214.045 ;
        RECT 3384.640 2213.200 3384.900 2214.410 ;
      LAYER via ;
        RECT 3370.420 2213.755 3370.680 2214.015 ;
        RECT 3384.640 2213.260 3384.900 2214.350 ;
      LAYER met2 ;
        RECT 3370.390 2213.895 3370.710 2214.015 ;
        RECT 3384.610 2213.895 3384.930 2214.350 ;
        RECT 3368.850 2213.755 3384.930 2213.895 ;
        RECT 3384.610 2213.260 3384.930 2213.755 ;
    END
  END mgmt_io_in_unbuf[9]
  PIN mgmt_io_in_unbuf[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.660 2206.780 3384.860 2208.370 ;
      LAYER mcon ;
        RECT 3384.690 2207.280 3384.860 2208.370 ;
      LAYER met1 ;
        RECT 3369.860 2208.065 3370.000 2273.275 ;
        RECT 3369.860 2207.745 3370.120 2208.065 ;
        RECT 3384.640 2207.220 3384.900 2208.430 ;
      LAYER via ;
        RECT 3369.860 2207.775 3370.120 2208.035 ;
        RECT 3384.640 2207.280 3384.900 2208.370 ;
      LAYER met2 ;
        RECT 3369.830 2207.915 3370.150 2208.035 ;
        RECT 3384.610 2207.915 3384.930 2208.370 ;
        RECT 3368.850 2207.775 3384.930 2207.915 ;
        RECT 3384.610 2207.280 3384.930 2207.775 ;
    END
  END mgmt_io_in_unbuf[8]
  PIN mgmt_io_in_unbuf[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3384.660 2200.800 3384.860 2202.390 ;
      LAYER mcon ;
        RECT 3384.690 2201.300 3384.860 2202.390 ;
      LAYER met1 ;
        RECT 3369.300 2202.085 3369.440 2271.275 ;
        RECT 3369.300 2201.765 3369.560 2202.085 ;
        RECT 3384.640 2201.240 3384.900 2202.450 ;
      LAYER via ;
        RECT 3369.300 2201.795 3369.560 2202.055 ;
        RECT 3384.640 2201.300 3384.900 2202.390 ;
      LAYER met2 ;
        RECT 3369.270 2201.935 3369.590 2202.055 ;
        RECT 3384.610 2201.935 3384.930 2202.390 ;
        RECT 3368.850 2201.795 3384.930 2201.935 ;
        RECT 3384.610 2201.300 3384.930 2201.795 ;
    END
  END mgmt_io_in_unbuf[7]
  PIN mgmt_io_out_buf[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3386.560 2200.895 3388.770 2201.065 ;
        RECT 3387.410 2200.810 3388.290 2200.895 ;
        RECT 3387.410 2200.225 3387.580 2200.810 ;
        RECT 3386.560 2200.055 3387.580 2200.225 ;
        RECT 3387.410 2199.385 3387.580 2200.055 ;
        RECT 3386.560 2199.215 3387.580 2199.385 ;
        RECT 3387.410 2198.545 3387.580 2199.215 ;
        RECT 3386.560 2198.375 3387.580 2198.545 ;
        RECT 3388.120 2200.225 3388.290 2200.810 ;
        RECT 3388.120 2200.055 3388.770 2200.225 ;
        RECT 3388.120 2199.385 3388.290 2200.055 ;
        RECT 3388.120 2199.215 3388.770 2199.385 ;
        RECT 3388.120 2198.545 3388.290 2199.215 ;
        RECT 3388.120 2198.375 3388.770 2198.545 ;
      LAYER met1 ;
        RECT 3369.020 2201.115 3369.160 2270.275 ;
        RECT 3369.020 2200.795 3369.280 2201.115 ;
        RECT 3387.350 2200.760 3388.320 2201.020 ;
      LAYER via ;
        RECT 3369.020 2200.825 3369.280 2201.085 ;
        RECT 3387.410 2200.760 3388.260 2201.020 ;
      LAYER met2 ;
        RECT 3368.990 2200.965 3369.310 2201.085 ;
        RECT 3387.410 2200.965 3388.260 2201.050 ;
        RECT 3368.850 2200.825 3388.260 2200.965 ;
        RECT 3387.410 2200.730 3388.260 2200.825 ;
    END
  END mgmt_io_out_buf[7]
  PIN mgmt_io_out_buf[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3386.560 2206.875 3388.770 2207.045 ;
        RECT 3387.410 2206.790 3388.290 2206.875 ;
        RECT 3387.410 2206.205 3387.580 2206.790 ;
        RECT 3386.560 2206.035 3387.580 2206.205 ;
        RECT 3387.410 2205.365 3387.580 2206.035 ;
        RECT 3386.560 2205.195 3387.580 2205.365 ;
        RECT 3387.410 2204.525 3387.580 2205.195 ;
        RECT 3386.560 2204.355 3387.580 2204.525 ;
        RECT 3388.120 2206.205 3388.290 2206.790 ;
        RECT 3388.120 2206.035 3388.770 2206.205 ;
        RECT 3388.120 2205.365 3388.290 2206.035 ;
        RECT 3388.120 2205.195 3388.770 2205.365 ;
        RECT 3388.120 2204.525 3388.290 2205.195 ;
        RECT 3388.120 2204.355 3388.770 2204.525 ;
      LAYER met1 ;
        RECT 3369.580 2207.095 3369.720 2272.275 ;
        RECT 3369.580 2206.775 3369.840 2207.095 ;
        RECT 3387.350 2206.740 3388.320 2207.000 ;
      LAYER via ;
        RECT 3369.580 2206.805 3369.840 2207.065 ;
        RECT 3387.410 2206.740 3388.260 2207.000 ;
      LAYER met2 ;
        RECT 3369.550 2206.945 3369.870 2207.065 ;
        RECT 3387.410 2206.945 3388.260 2207.030 ;
        RECT 3368.850 2206.805 3388.260 2206.945 ;
        RECT 3387.410 2206.710 3388.260 2206.805 ;
    END
  END mgmt_io_out_buf[8]
  PIN mgmt_io_out_buf[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3386.560 2212.855 3388.770 2213.025 ;
        RECT 3387.410 2212.770 3388.290 2212.855 ;
        RECT 3387.410 2212.185 3387.580 2212.770 ;
        RECT 3386.560 2212.015 3387.580 2212.185 ;
        RECT 3387.410 2211.345 3387.580 2212.015 ;
        RECT 3386.560 2211.175 3387.580 2211.345 ;
        RECT 3387.410 2210.505 3387.580 2211.175 ;
        RECT 3386.560 2210.335 3387.580 2210.505 ;
        RECT 3388.120 2212.185 3388.290 2212.770 ;
        RECT 3388.120 2212.015 3388.770 2212.185 ;
        RECT 3388.120 2211.345 3388.290 2212.015 ;
        RECT 3388.120 2211.175 3388.770 2211.345 ;
        RECT 3388.120 2210.505 3388.290 2211.175 ;
        RECT 3388.120 2210.335 3388.770 2210.505 ;
      LAYER met1 ;
        RECT 3370.140 2213.075 3370.280 2274.275 ;
        RECT 3370.140 2212.755 3370.400 2213.075 ;
        RECT 3387.350 2212.720 3388.320 2212.980 ;
      LAYER via ;
        RECT 3370.140 2212.785 3370.400 2213.045 ;
        RECT 3387.410 2212.720 3388.260 2212.980 ;
      LAYER met2 ;
        RECT 3370.110 2212.925 3370.430 2213.045 ;
        RECT 3387.410 2212.925 3388.260 2213.010 ;
        RECT 3368.850 2212.785 3388.260 2212.925 ;
        RECT 3387.410 2212.690 3388.260 2212.785 ;
    END
  END mgmt_io_out_buf[9]
  PIN mgmt_io_out_buf[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3386.560 2218.835 3388.770 2219.005 ;
        RECT 3387.410 2218.750 3388.290 2218.835 ;
        RECT 3387.410 2218.165 3387.580 2218.750 ;
        RECT 3386.560 2217.995 3387.580 2218.165 ;
        RECT 3387.410 2217.325 3387.580 2217.995 ;
        RECT 3386.560 2217.155 3387.580 2217.325 ;
        RECT 3387.410 2216.485 3387.580 2217.155 ;
        RECT 3386.560 2216.315 3387.580 2216.485 ;
        RECT 3388.120 2218.165 3388.290 2218.750 ;
        RECT 3388.120 2217.995 3388.770 2218.165 ;
        RECT 3388.120 2217.325 3388.290 2217.995 ;
        RECT 3388.120 2217.155 3388.770 2217.325 ;
        RECT 3388.120 2216.485 3388.290 2217.155 ;
        RECT 3388.120 2216.315 3388.770 2216.485 ;
      LAYER met1 ;
        RECT 3370.700 2219.055 3370.840 2276.275 ;
        RECT 3370.700 2218.735 3370.960 2219.055 ;
        RECT 3387.350 2218.700 3388.320 2218.960 ;
      LAYER via ;
        RECT 3370.700 2218.765 3370.960 2219.025 ;
        RECT 3387.410 2218.700 3388.260 2218.960 ;
      LAYER met2 ;
        RECT 3370.670 2218.905 3370.990 2219.025 ;
        RECT 3387.410 2218.905 3388.260 2218.990 ;
        RECT 3368.850 2218.765 3388.260 2218.905 ;
        RECT 3387.410 2218.670 3388.260 2218.765 ;
    END
  END mgmt_io_out_buf[10]
  PIN mgmt_io_out_buf[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3386.560 2224.815 3388.770 2224.985 ;
        RECT 3387.410 2224.730 3388.290 2224.815 ;
        RECT 3387.410 2224.145 3387.580 2224.730 ;
        RECT 3386.560 2223.975 3387.580 2224.145 ;
        RECT 3387.410 2223.305 3387.580 2223.975 ;
        RECT 3386.560 2223.135 3387.580 2223.305 ;
        RECT 3387.410 2222.465 3387.580 2223.135 ;
        RECT 3386.560 2222.295 3387.580 2222.465 ;
        RECT 3388.120 2224.145 3388.290 2224.730 ;
        RECT 3388.120 2223.975 3388.770 2224.145 ;
        RECT 3388.120 2223.305 3388.290 2223.975 ;
        RECT 3388.120 2223.135 3388.770 2223.305 ;
        RECT 3388.120 2222.465 3388.290 2223.135 ;
        RECT 3388.120 2222.295 3388.770 2222.465 ;
      LAYER met1 ;
        RECT 3371.260 2225.035 3371.400 2278.275 ;
        RECT 3371.260 2224.715 3371.520 2225.035 ;
        RECT 3387.350 2224.680 3388.320 2224.940 ;
      LAYER via ;
        RECT 3371.260 2224.745 3371.520 2225.005 ;
        RECT 3387.410 2224.680 3388.260 2224.940 ;
      LAYER met2 ;
        RECT 3371.230 2224.885 3371.550 2225.005 ;
        RECT 3387.410 2224.885 3388.260 2224.970 ;
        RECT 3368.850 2224.745 3388.260 2224.885 ;
        RECT 3387.410 2224.650 3388.260 2224.745 ;
    END
  END mgmt_io_out_buf[11]
  PIN mgmt_io_out_buf[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3386.560 2230.795 3388.770 2230.965 ;
        RECT 3387.410 2230.710 3388.290 2230.795 ;
        RECT 3387.410 2230.125 3387.580 2230.710 ;
        RECT 3386.560 2229.955 3387.580 2230.125 ;
        RECT 3387.410 2229.285 3387.580 2229.955 ;
        RECT 3386.560 2229.115 3387.580 2229.285 ;
        RECT 3387.410 2228.445 3387.580 2229.115 ;
        RECT 3386.560 2228.275 3387.580 2228.445 ;
        RECT 3388.120 2230.125 3388.290 2230.710 ;
        RECT 3388.120 2229.955 3388.770 2230.125 ;
        RECT 3388.120 2229.285 3388.290 2229.955 ;
        RECT 3388.120 2229.115 3388.770 2229.285 ;
        RECT 3388.120 2228.445 3388.290 2229.115 ;
        RECT 3388.120 2228.275 3388.770 2228.445 ;
      LAYER met1 ;
        RECT 3371.820 2231.015 3371.960 2280.275 ;
        RECT 3371.820 2230.695 3372.080 2231.015 ;
        RECT 3387.350 2230.660 3388.320 2230.920 ;
      LAYER via ;
        RECT 3371.820 2230.725 3372.080 2230.985 ;
        RECT 3387.410 2230.660 3388.260 2230.920 ;
      LAYER met2 ;
        RECT 3371.790 2230.865 3372.110 2230.985 ;
        RECT 3387.410 2230.865 3388.260 2230.950 ;
        RECT 3368.850 2230.725 3388.260 2230.865 ;
        RECT 3387.410 2230.630 3388.260 2230.725 ;
    END
  END mgmt_io_out_buf[12]
  PIN mgmt_io_out_unbuf[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3387.750 2196.660 3387.950 2197.760 ;
      LAYER mcon ;
        RECT 3387.750 2196.670 3387.920 2197.760 ;
      LAYER met1 ;
        RECT 3369.040 2196.930 3369.300 2197.250 ;
        RECT 3369.160 1075.250 3369.300 2196.930 ;
        RECT 3387.700 2196.610 3387.960 2197.820 ;
      LAYER via ;
        RECT 3369.040 2196.960 3369.300 2197.220 ;
        RECT 3387.700 2196.670 3387.960 2197.760 ;
      LAYER met2 ;
        RECT 3369.010 2197.100 3369.330 2197.220 ;
        RECT 3387.670 2197.100 3387.990 2197.760 ;
        RECT 3368.850 2196.960 3387.990 2197.100 ;
        RECT 3387.670 2196.670 3387.990 2196.960 ;
    END
  END mgmt_io_out_unbuf[7]
  PIN mgmt_io_out_unbuf[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3387.750 2202.640 3387.950 2203.740 ;
      LAYER mcon ;
        RECT 3387.750 2202.650 3387.920 2203.740 ;
      LAYER met1 ;
        RECT 3369.600 2202.910 3369.860 2203.230 ;
        RECT 3369.720 1073.250 3369.860 2202.910 ;
        RECT 3387.700 2202.590 3387.960 2203.800 ;
      LAYER via ;
        RECT 3369.600 2202.940 3369.860 2203.200 ;
        RECT 3387.700 2202.650 3387.960 2203.740 ;
      LAYER met2 ;
        RECT 3369.570 2203.080 3369.890 2203.200 ;
        RECT 3387.670 2203.080 3387.990 2203.740 ;
        RECT 3368.850 2202.940 3387.990 2203.080 ;
        RECT 3387.670 2202.650 3387.990 2202.940 ;
    END
  END mgmt_io_out_unbuf[8]
  PIN mgmt_io_out_unbuf[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3387.750 2208.620 3387.950 2209.720 ;
      LAYER mcon ;
        RECT 3387.750 2208.630 3387.920 2209.720 ;
      LAYER met1 ;
        RECT 3370.160 2208.890 3370.420 2209.210 ;
        RECT 3370.280 1071.250 3370.420 2208.890 ;
        RECT 3387.700 2208.570 3387.960 2209.780 ;
      LAYER via ;
        RECT 3370.160 2208.920 3370.420 2209.180 ;
        RECT 3387.700 2208.630 3387.960 2209.720 ;
      LAYER met2 ;
        RECT 3370.130 2209.060 3370.450 2209.180 ;
        RECT 3387.670 2209.060 3387.990 2209.720 ;
        RECT 3368.850 2208.920 3387.990 2209.060 ;
        RECT 3387.670 2208.630 3387.990 2208.920 ;
    END
  END mgmt_io_out_unbuf[9]
  PIN mgmt_io_out_unbuf[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3387.750 2214.600 3387.950 2215.700 ;
      LAYER mcon ;
        RECT 3387.750 2214.610 3387.920 2215.700 ;
      LAYER met1 ;
        RECT 3370.720 2214.870 3370.980 2215.190 ;
        RECT 3370.840 1069.250 3370.980 2214.870 ;
        RECT 3387.700 2214.550 3387.960 2215.760 ;
      LAYER via ;
        RECT 3370.720 2214.900 3370.980 2215.160 ;
        RECT 3387.700 2214.610 3387.960 2215.700 ;
      LAYER met2 ;
        RECT 3370.690 2215.040 3371.010 2215.160 ;
        RECT 3387.670 2215.040 3387.990 2215.700 ;
        RECT 3368.850 2214.900 3387.990 2215.040 ;
        RECT 3387.670 2214.610 3387.990 2214.900 ;
    END
  END mgmt_io_out_unbuf[10]
  PIN mgmt_io_out_unbuf[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3387.750 2220.580 3387.950 2221.680 ;
      LAYER mcon ;
        RECT 3387.750 2220.590 3387.920 2221.680 ;
      LAYER met1 ;
        RECT 3371.280 2220.850 3371.540 2221.170 ;
        RECT 3371.400 1067.250 3371.540 2220.850 ;
        RECT 3387.700 2220.530 3387.960 2221.740 ;
      LAYER via ;
        RECT 3371.280 2220.880 3371.540 2221.140 ;
        RECT 3387.700 2220.590 3387.960 2221.680 ;
      LAYER met2 ;
        RECT 3371.250 2221.020 3371.570 2221.140 ;
        RECT 3387.670 2221.020 3387.990 2221.680 ;
        RECT 3368.850 2220.880 3387.990 2221.020 ;
        RECT 3387.670 2220.590 3387.990 2220.880 ;
    END
  END mgmt_io_out_unbuf[11]
  PIN mgmt_io_out_unbuf[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3387.750 2226.560 3387.950 2227.660 ;
      LAYER mcon ;
        RECT 3387.750 2226.570 3387.920 2227.660 ;
      LAYER met1 ;
        RECT 3371.840 2226.830 3372.100 2227.150 ;
        RECT 3371.960 1065.250 3372.100 2226.830 ;
        RECT 3387.700 2226.510 3387.960 2227.720 ;
      LAYER via ;
        RECT 3371.840 2226.860 3372.100 2227.120 ;
        RECT 3387.700 2226.570 3387.960 2227.660 ;
      LAYER met2 ;
        RECT 3371.810 2227.000 3372.130 2227.120 ;
        RECT 3387.670 2227.000 3387.990 2227.660 ;
        RECT 3368.850 2226.860 3387.990 2227.000 ;
        RECT 3387.670 2226.570 3387.990 2226.860 ;
    END
  END mgmt_io_out_unbuf[12]
  PIN mgmt_io_out_unbuf[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3387.750 2232.540 3387.950 2233.640 ;
      LAYER mcon ;
        RECT 3387.750 2232.550 3387.920 2233.640 ;
      LAYER met1 ;
        RECT 3372.400 2232.810 3372.660 2233.130 ;
        RECT 3372.520 1063.250 3372.660 2232.810 ;
        RECT 3387.700 2232.490 3387.960 2233.700 ;
      LAYER via ;
        RECT 3372.400 2232.840 3372.660 2233.100 ;
        RECT 3387.700 2232.550 3387.960 2233.640 ;
      LAYER met2 ;
        RECT 3372.370 2232.980 3372.690 2233.100 ;
        RECT 3387.670 2232.980 3387.990 2233.640 ;
        RECT 3368.850 2232.840 3387.990 2232.980 ;
        RECT 3387.670 2232.550 3387.990 2232.840 ;
    END
  END mgmt_io_out_unbuf[13]
  PIN mgmt_io_out_unbuf[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3387.750 2238.520 3387.950 2239.620 ;
      LAYER mcon ;
        RECT 3387.750 2238.530 3387.920 2239.620 ;
      LAYER met1 ;
        RECT 3372.960 2238.790 3373.220 2239.110 ;
        RECT 3373.080 1061.250 3373.220 2238.790 ;
        RECT 3387.700 2238.470 3387.960 2239.680 ;
      LAYER via ;
        RECT 3372.960 2238.820 3373.220 2239.080 ;
        RECT 3387.700 2238.530 3387.960 2239.620 ;
      LAYER met2 ;
        RECT 3372.930 2238.960 3373.250 2239.080 ;
        RECT 3387.670 2238.960 3387.990 2239.620 ;
        RECT 3368.850 2238.820 3387.990 2238.960 ;
        RECT 3387.670 2238.530 3387.990 2238.820 ;
    END
  END mgmt_io_out_unbuf[14]
  PIN mgmt_io_out_unbuf[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3387.750 2244.500 3387.950 2245.600 ;
      LAYER mcon ;
        RECT 3387.750 2244.510 3387.920 2245.600 ;
      LAYER met1 ;
        RECT 3373.520 2244.770 3373.780 2245.090 ;
        RECT 3373.640 1059.250 3373.780 2244.770 ;
        RECT 3387.700 2244.450 3387.960 2245.660 ;
      LAYER via ;
        RECT 3373.520 2244.800 3373.780 2245.060 ;
        RECT 3387.700 2244.510 3387.960 2245.600 ;
      LAYER met2 ;
        RECT 3373.490 2244.940 3373.810 2245.060 ;
        RECT 3387.670 2244.940 3387.990 2245.600 ;
        RECT 3368.850 2244.800 3387.990 2244.940 ;
        RECT 3387.670 2244.510 3387.990 2244.800 ;
    END
  END mgmt_io_out_unbuf[15]
  PIN mgmt_io_out_unbuf[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3387.750 2250.480 3387.950 2251.580 ;
      LAYER mcon ;
        RECT 3387.750 2250.490 3387.920 2251.580 ;
      LAYER met1 ;
        RECT 3374.080 2250.750 3374.340 2251.070 ;
        RECT 3374.200 1057.250 3374.340 2250.750 ;
        RECT 3387.700 2250.430 3387.960 2251.640 ;
      LAYER via ;
        RECT 3374.080 2250.780 3374.340 2251.040 ;
        RECT 3387.700 2250.490 3387.960 2251.580 ;
      LAYER met2 ;
        RECT 3374.050 2250.920 3374.370 2251.040 ;
        RECT 3387.670 2250.920 3387.990 2251.580 ;
        RECT 3368.850 2250.780 3387.990 2250.920 ;
        RECT 3387.670 2250.490 3387.990 2250.780 ;
    END
  END mgmt_io_out_unbuf[16]
  PIN mgmt_io_out_unbuf[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3387.750 2256.460 3387.950 2257.560 ;
      LAYER mcon ;
        RECT 3387.750 2256.470 3387.920 2257.560 ;
      LAYER met1 ;
        RECT 3374.640 2256.730 3374.900 2257.050 ;
        RECT 3374.760 1055.250 3374.900 2256.730 ;
        RECT 3387.700 2256.410 3387.960 2257.620 ;
      LAYER via ;
        RECT 3374.640 2256.760 3374.900 2257.020 ;
        RECT 3387.700 2256.470 3387.960 2257.560 ;
      LAYER met2 ;
        RECT 3374.610 2256.900 3374.930 2257.020 ;
        RECT 3387.670 2256.900 3387.990 2257.560 ;
        RECT 3368.850 2256.760 3387.990 2256.900 ;
        RECT 3387.670 2256.470 3387.990 2256.760 ;
    END
  END mgmt_io_out_unbuf[17]
  PIN mgmt_io_out_unbuf[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3387.750 2262.440 3387.950 2263.540 ;
      LAYER mcon ;
        RECT 3387.750 2262.450 3387.920 2263.540 ;
      LAYER met1 ;
        RECT 3375.200 2262.710 3375.460 2263.030 ;
        RECT 3375.320 1053.250 3375.460 2262.710 ;
        RECT 3387.700 2262.390 3387.960 2263.600 ;
      LAYER via ;
        RECT 3375.200 2262.740 3375.460 2263.000 ;
        RECT 3387.700 2262.450 3387.960 2263.540 ;
      LAYER met2 ;
        RECT 3375.170 2262.880 3375.490 2263.000 ;
        RECT 3387.670 2262.880 3387.990 2263.540 ;
        RECT 3368.850 2262.740 3387.990 2262.880 ;
        RECT 3387.670 2262.450 3387.990 2262.740 ;
    END
  END mgmt_io_out_unbuf[18]
  PIN mgmt_io_in_buf[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.840 2265.795 3384.490 2265.965 ;
        RECT 3384.320 2265.125 3384.490 2265.795 ;
        RECT 3383.840 2264.955 3384.490 2265.125 ;
        RECT 3384.320 2264.285 3384.490 2264.955 ;
        RECT 3383.840 2264.115 3384.490 2264.285 ;
        RECT 3384.320 2263.530 3384.490 2264.115 ;
        RECT 3385.030 2265.795 3386.050 2265.965 ;
        RECT 3385.030 2265.125 3385.200 2265.795 ;
        RECT 3385.030 2264.955 3386.050 2265.125 ;
        RECT 3385.030 2264.285 3385.200 2264.955 ;
        RECT 3385.030 2264.115 3386.050 2264.285 ;
        RECT 3385.030 2263.530 3385.200 2264.115 ;
        RECT 3384.320 2263.445 3385.200 2263.530 ;
        RECT 3383.840 2263.275 3386.050 2263.445 ;
      LAYER mcon ;
        RECT 3384.350 2263.360 3385.200 2263.530 ;
      LAYER met1 ;
        RECT 3375.480 2263.330 3375.740 2263.650 ;
        RECT 3375.600 1052.250 3375.740 2263.330 ;
        RECT 3384.290 2263.310 3385.260 2263.570 ;
      LAYER via ;
        RECT 3375.480 2263.360 3375.740 2263.620 ;
        RECT 3384.350 2263.310 3385.200 2263.570 ;
      LAYER met2 ;
        RECT 3375.450 2263.500 3375.770 2263.620 ;
        RECT 3384.350 2263.500 3385.200 2263.600 ;
        RECT 3368.850 2263.360 3385.200 2263.500 ;
        RECT 3384.350 2263.280 3385.200 2263.360 ;
    END
  END mgmt_io_in_buf[18]
  PIN mgmt_io_in_buf[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.840 2259.815 3384.490 2259.985 ;
        RECT 3384.320 2259.145 3384.490 2259.815 ;
        RECT 3383.840 2258.975 3384.490 2259.145 ;
        RECT 3384.320 2258.305 3384.490 2258.975 ;
        RECT 3383.840 2258.135 3384.490 2258.305 ;
        RECT 3384.320 2257.550 3384.490 2258.135 ;
        RECT 3385.030 2259.815 3386.050 2259.985 ;
        RECT 3385.030 2259.145 3385.200 2259.815 ;
        RECT 3385.030 2258.975 3386.050 2259.145 ;
        RECT 3385.030 2258.305 3385.200 2258.975 ;
        RECT 3385.030 2258.135 3386.050 2258.305 ;
        RECT 3385.030 2257.550 3385.200 2258.135 ;
        RECT 3384.320 2257.465 3385.200 2257.550 ;
        RECT 3383.840 2257.295 3386.050 2257.465 ;
      LAYER mcon ;
        RECT 3384.350 2257.380 3385.200 2257.550 ;
      LAYER met1 ;
        RECT 3374.920 2257.350 3375.180 2257.670 ;
        RECT 3375.040 1054.250 3375.180 2257.350 ;
        RECT 3384.290 2257.330 3385.260 2257.590 ;
      LAYER via ;
        RECT 3374.920 2257.380 3375.180 2257.640 ;
        RECT 3384.350 2257.330 3385.200 2257.590 ;
      LAYER met2 ;
        RECT 3374.890 2257.520 3375.210 2257.640 ;
        RECT 3384.350 2257.520 3385.200 2257.620 ;
        RECT 3368.850 2257.380 3385.200 2257.520 ;
        RECT 3384.350 2257.300 3385.200 2257.380 ;
    END
  END mgmt_io_in_buf[17]
  PIN mgmt_io_in_buf[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.840 2253.835 3384.490 2254.005 ;
        RECT 3384.320 2253.165 3384.490 2253.835 ;
        RECT 3383.840 2252.995 3384.490 2253.165 ;
        RECT 3384.320 2252.325 3384.490 2252.995 ;
        RECT 3383.840 2252.155 3384.490 2252.325 ;
        RECT 3384.320 2251.570 3384.490 2252.155 ;
        RECT 3385.030 2253.835 3386.050 2254.005 ;
        RECT 3385.030 2253.165 3385.200 2253.835 ;
        RECT 3385.030 2252.995 3386.050 2253.165 ;
        RECT 3385.030 2252.325 3385.200 2252.995 ;
        RECT 3385.030 2252.155 3386.050 2252.325 ;
        RECT 3385.030 2251.570 3385.200 2252.155 ;
        RECT 3384.320 2251.485 3385.200 2251.570 ;
        RECT 3383.840 2251.315 3386.050 2251.485 ;
      LAYER mcon ;
        RECT 3384.350 2251.400 3385.200 2251.570 ;
      LAYER met1 ;
        RECT 3374.360 2251.370 3374.620 2251.690 ;
        RECT 3374.480 1056.250 3374.620 2251.370 ;
        RECT 3384.290 2251.350 3385.260 2251.610 ;
      LAYER via ;
        RECT 3374.360 2251.400 3374.620 2251.660 ;
        RECT 3384.350 2251.350 3385.200 2251.610 ;
      LAYER met2 ;
        RECT 3374.330 2251.540 3374.650 2251.660 ;
        RECT 3384.350 2251.540 3385.200 2251.640 ;
        RECT 3368.850 2251.400 3385.200 2251.540 ;
        RECT 3384.350 2251.320 3385.200 2251.400 ;
    END
  END mgmt_io_in_buf[16]
  PIN mgmt_io_in_buf[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.840 2247.855 3384.490 2248.025 ;
        RECT 3384.320 2247.185 3384.490 2247.855 ;
        RECT 3383.840 2247.015 3384.490 2247.185 ;
        RECT 3384.320 2246.345 3384.490 2247.015 ;
        RECT 3383.840 2246.175 3384.490 2246.345 ;
        RECT 3384.320 2245.590 3384.490 2246.175 ;
        RECT 3385.030 2247.855 3386.050 2248.025 ;
        RECT 3385.030 2247.185 3385.200 2247.855 ;
        RECT 3385.030 2247.015 3386.050 2247.185 ;
        RECT 3385.030 2246.345 3385.200 2247.015 ;
        RECT 3385.030 2246.175 3386.050 2246.345 ;
        RECT 3385.030 2245.590 3385.200 2246.175 ;
        RECT 3384.320 2245.505 3385.200 2245.590 ;
        RECT 3383.840 2245.335 3386.050 2245.505 ;
      LAYER mcon ;
        RECT 3384.350 2245.420 3385.200 2245.590 ;
      LAYER met1 ;
        RECT 3373.800 2245.390 3374.060 2245.710 ;
        RECT 3373.920 1058.250 3374.060 2245.390 ;
        RECT 3384.290 2245.370 3385.260 2245.630 ;
      LAYER via ;
        RECT 3373.800 2245.420 3374.060 2245.680 ;
        RECT 3384.350 2245.370 3385.200 2245.630 ;
      LAYER met2 ;
        RECT 3373.770 2245.560 3374.090 2245.680 ;
        RECT 3384.350 2245.560 3385.200 2245.660 ;
        RECT 3368.850 2245.420 3385.200 2245.560 ;
        RECT 3384.350 2245.340 3385.200 2245.420 ;
    END
  END mgmt_io_in_buf[15]
  PIN mgmt_io_in_buf[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.840 2241.875 3384.490 2242.045 ;
        RECT 3384.320 2241.205 3384.490 2241.875 ;
        RECT 3383.840 2241.035 3384.490 2241.205 ;
        RECT 3384.320 2240.365 3384.490 2241.035 ;
        RECT 3383.840 2240.195 3384.490 2240.365 ;
        RECT 3384.320 2239.610 3384.490 2240.195 ;
        RECT 3385.030 2241.875 3386.050 2242.045 ;
        RECT 3385.030 2241.205 3385.200 2241.875 ;
        RECT 3385.030 2241.035 3386.050 2241.205 ;
        RECT 3385.030 2240.365 3385.200 2241.035 ;
        RECT 3385.030 2240.195 3386.050 2240.365 ;
        RECT 3385.030 2239.610 3385.200 2240.195 ;
        RECT 3384.320 2239.525 3385.200 2239.610 ;
        RECT 3383.840 2239.355 3386.050 2239.525 ;
      LAYER mcon ;
        RECT 3384.350 2239.440 3385.200 2239.610 ;
      LAYER met1 ;
        RECT 3373.240 2239.410 3373.500 2239.730 ;
        RECT 3373.360 1060.250 3373.500 2239.410 ;
        RECT 3384.290 2239.390 3385.260 2239.650 ;
      LAYER via ;
        RECT 3373.240 2239.440 3373.500 2239.700 ;
        RECT 3384.350 2239.390 3385.200 2239.650 ;
      LAYER met2 ;
        RECT 3373.210 2239.580 3373.530 2239.700 ;
        RECT 3384.350 2239.580 3385.200 2239.680 ;
        RECT 3368.850 2239.440 3385.200 2239.580 ;
        RECT 3384.350 2239.360 3385.200 2239.440 ;
    END
  END mgmt_io_in_buf[14]
  PIN mgmt_io_in_buf[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.840 2235.895 3384.490 2236.065 ;
        RECT 3384.320 2235.225 3384.490 2235.895 ;
        RECT 3383.840 2235.055 3384.490 2235.225 ;
        RECT 3384.320 2234.385 3384.490 2235.055 ;
        RECT 3383.840 2234.215 3384.490 2234.385 ;
        RECT 3384.320 2233.630 3384.490 2234.215 ;
        RECT 3385.030 2235.895 3386.050 2236.065 ;
        RECT 3385.030 2235.225 3385.200 2235.895 ;
        RECT 3385.030 2235.055 3386.050 2235.225 ;
        RECT 3385.030 2234.385 3385.200 2235.055 ;
        RECT 3385.030 2234.215 3386.050 2234.385 ;
        RECT 3385.030 2233.630 3385.200 2234.215 ;
        RECT 3384.320 2233.545 3385.200 2233.630 ;
        RECT 3383.840 2233.375 3386.050 2233.545 ;
      LAYER mcon ;
        RECT 3384.350 2233.460 3385.200 2233.630 ;
      LAYER met1 ;
        RECT 3372.680 2233.430 3372.940 2233.750 ;
        RECT 3372.800 1062.250 3372.940 2233.430 ;
        RECT 3384.290 2233.410 3385.260 2233.670 ;
      LAYER via ;
        RECT 3372.680 2233.460 3372.940 2233.720 ;
        RECT 3384.350 2233.410 3385.200 2233.670 ;
      LAYER met2 ;
        RECT 3372.650 2233.600 3372.970 2233.720 ;
        RECT 3384.350 2233.600 3385.200 2233.700 ;
        RECT 3368.850 2233.460 3385.200 2233.600 ;
        RECT 3384.350 2233.380 3385.200 2233.460 ;
    END
  END mgmt_io_in_buf[13]
  PIN mgmt_io_in_buf[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.840 2229.915 3384.490 2230.085 ;
        RECT 3384.320 2229.245 3384.490 2229.915 ;
        RECT 3383.840 2229.075 3384.490 2229.245 ;
        RECT 3384.320 2228.405 3384.490 2229.075 ;
        RECT 3383.840 2228.235 3384.490 2228.405 ;
        RECT 3384.320 2227.650 3384.490 2228.235 ;
        RECT 3385.030 2229.915 3386.050 2230.085 ;
        RECT 3385.030 2229.245 3385.200 2229.915 ;
        RECT 3385.030 2229.075 3386.050 2229.245 ;
        RECT 3385.030 2228.405 3385.200 2229.075 ;
        RECT 3385.030 2228.235 3386.050 2228.405 ;
        RECT 3385.030 2227.650 3385.200 2228.235 ;
        RECT 3384.320 2227.565 3385.200 2227.650 ;
        RECT 3383.840 2227.395 3386.050 2227.565 ;
      LAYER mcon ;
        RECT 3384.350 2227.480 3385.200 2227.650 ;
      LAYER met1 ;
        RECT 3372.120 2227.450 3372.380 2227.770 ;
        RECT 3372.240 1064.250 3372.380 2227.450 ;
        RECT 3384.290 2227.430 3385.260 2227.690 ;
      LAYER via ;
        RECT 3372.120 2227.480 3372.380 2227.740 ;
        RECT 3384.350 2227.430 3385.200 2227.690 ;
      LAYER met2 ;
        RECT 3372.090 2227.620 3372.410 2227.740 ;
        RECT 3384.350 2227.620 3385.200 2227.720 ;
        RECT 3368.850 2227.480 3385.200 2227.620 ;
        RECT 3384.350 2227.400 3385.200 2227.480 ;
    END
  END mgmt_io_in_buf[12]
  PIN mgmt_io_in_buf[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.840 2223.935 3384.490 2224.105 ;
        RECT 3384.320 2223.265 3384.490 2223.935 ;
        RECT 3383.840 2223.095 3384.490 2223.265 ;
        RECT 3384.320 2222.425 3384.490 2223.095 ;
        RECT 3383.840 2222.255 3384.490 2222.425 ;
        RECT 3384.320 2221.670 3384.490 2222.255 ;
        RECT 3385.030 2223.935 3386.050 2224.105 ;
        RECT 3385.030 2223.265 3385.200 2223.935 ;
        RECT 3385.030 2223.095 3386.050 2223.265 ;
        RECT 3385.030 2222.425 3385.200 2223.095 ;
        RECT 3385.030 2222.255 3386.050 2222.425 ;
        RECT 3385.030 2221.670 3385.200 2222.255 ;
        RECT 3384.320 2221.585 3385.200 2221.670 ;
        RECT 3383.840 2221.415 3386.050 2221.585 ;
      LAYER mcon ;
        RECT 3384.350 2221.500 3385.200 2221.670 ;
      LAYER met1 ;
        RECT 3371.560 2221.470 3371.820 2221.790 ;
        RECT 3371.680 1066.250 3371.820 2221.470 ;
        RECT 3384.290 2221.450 3385.260 2221.710 ;
      LAYER via ;
        RECT 3371.560 2221.500 3371.820 2221.760 ;
        RECT 3384.350 2221.450 3385.200 2221.710 ;
      LAYER met2 ;
        RECT 3371.530 2221.640 3371.850 2221.760 ;
        RECT 3384.350 2221.640 3385.200 2221.740 ;
        RECT 3368.850 2221.500 3385.200 2221.640 ;
        RECT 3384.350 2221.420 3385.200 2221.500 ;
    END
  END mgmt_io_in_buf[11]
  PIN mgmt_io_in_buf[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.840 2217.955 3384.490 2218.125 ;
        RECT 3384.320 2217.285 3384.490 2217.955 ;
        RECT 3383.840 2217.115 3384.490 2217.285 ;
        RECT 3384.320 2216.445 3384.490 2217.115 ;
        RECT 3383.840 2216.275 3384.490 2216.445 ;
        RECT 3384.320 2215.690 3384.490 2216.275 ;
        RECT 3385.030 2217.955 3386.050 2218.125 ;
        RECT 3385.030 2217.285 3385.200 2217.955 ;
        RECT 3385.030 2217.115 3386.050 2217.285 ;
        RECT 3385.030 2216.445 3385.200 2217.115 ;
        RECT 3385.030 2216.275 3386.050 2216.445 ;
        RECT 3385.030 2215.690 3385.200 2216.275 ;
        RECT 3384.320 2215.605 3385.200 2215.690 ;
        RECT 3383.840 2215.435 3386.050 2215.605 ;
      LAYER mcon ;
        RECT 3384.350 2215.520 3385.200 2215.690 ;
      LAYER met1 ;
        RECT 3371.000 2215.490 3371.260 2215.810 ;
        RECT 3371.120 1068.250 3371.260 2215.490 ;
        RECT 3384.290 2215.470 3385.260 2215.730 ;
      LAYER via ;
        RECT 3371.000 2215.520 3371.260 2215.780 ;
        RECT 3384.350 2215.470 3385.200 2215.730 ;
      LAYER met2 ;
        RECT 3370.970 2215.660 3371.290 2215.780 ;
        RECT 3384.350 2215.660 3385.200 2215.760 ;
        RECT 3368.850 2215.520 3385.200 2215.660 ;
        RECT 3384.350 2215.440 3385.200 2215.520 ;
    END
  END mgmt_io_in_buf[10]
  PIN mgmt_io_in_buf[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.840 2211.975 3384.490 2212.145 ;
        RECT 3384.320 2211.305 3384.490 2211.975 ;
        RECT 3383.840 2211.135 3384.490 2211.305 ;
        RECT 3384.320 2210.465 3384.490 2211.135 ;
        RECT 3383.840 2210.295 3384.490 2210.465 ;
        RECT 3384.320 2209.710 3384.490 2210.295 ;
        RECT 3385.030 2211.975 3386.050 2212.145 ;
        RECT 3385.030 2211.305 3385.200 2211.975 ;
        RECT 3385.030 2211.135 3386.050 2211.305 ;
        RECT 3385.030 2210.465 3385.200 2211.135 ;
        RECT 3385.030 2210.295 3386.050 2210.465 ;
        RECT 3385.030 2209.710 3385.200 2210.295 ;
        RECT 3384.320 2209.625 3385.200 2209.710 ;
        RECT 3383.840 2209.455 3386.050 2209.625 ;
      LAYER mcon ;
        RECT 3384.350 2209.540 3385.200 2209.710 ;
      LAYER met1 ;
        RECT 3370.440 2209.510 3370.700 2209.830 ;
        RECT 3370.560 1070.250 3370.700 2209.510 ;
        RECT 3384.290 2209.490 3385.260 2209.750 ;
      LAYER via ;
        RECT 3370.440 2209.540 3370.700 2209.800 ;
        RECT 3384.350 2209.490 3385.200 2209.750 ;
      LAYER met2 ;
        RECT 3370.410 2209.680 3370.730 2209.800 ;
        RECT 3384.350 2209.680 3385.200 2209.780 ;
        RECT 3368.850 2209.540 3385.200 2209.680 ;
        RECT 3384.350 2209.460 3385.200 2209.540 ;
    END
  END mgmt_io_in_buf[9]
  PIN mgmt_io_in_buf[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.840 2205.995 3384.490 2206.165 ;
        RECT 3384.320 2205.325 3384.490 2205.995 ;
        RECT 3383.840 2205.155 3384.490 2205.325 ;
        RECT 3384.320 2204.485 3384.490 2205.155 ;
        RECT 3383.840 2204.315 3384.490 2204.485 ;
        RECT 3384.320 2203.730 3384.490 2204.315 ;
        RECT 3385.030 2205.995 3386.050 2206.165 ;
        RECT 3385.030 2205.325 3385.200 2205.995 ;
        RECT 3385.030 2205.155 3386.050 2205.325 ;
        RECT 3385.030 2204.485 3385.200 2205.155 ;
        RECT 3385.030 2204.315 3386.050 2204.485 ;
        RECT 3385.030 2203.730 3385.200 2204.315 ;
        RECT 3384.320 2203.645 3385.200 2203.730 ;
        RECT 3383.840 2203.475 3386.050 2203.645 ;
      LAYER mcon ;
        RECT 3384.350 2203.560 3385.200 2203.730 ;
      LAYER met1 ;
        RECT 3369.880 2203.530 3370.140 2203.850 ;
        RECT 3370.000 1072.250 3370.140 2203.530 ;
        RECT 3384.290 2203.510 3385.260 2203.770 ;
      LAYER via ;
        RECT 3369.880 2203.560 3370.140 2203.820 ;
        RECT 3384.350 2203.510 3385.200 2203.770 ;
      LAYER met2 ;
        RECT 3369.850 2203.700 3370.170 2203.820 ;
        RECT 3384.350 2203.700 3385.200 2203.800 ;
        RECT 3368.850 2203.560 3385.200 2203.700 ;
        RECT 3384.350 2203.480 3385.200 2203.560 ;
    END
  END mgmt_io_in_buf[8]
  PIN mgmt_io_in_buf[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3383.840 2200.015 3384.490 2200.185 ;
        RECT 3384.320 2199.345 3384.490 2200.015 ;
        RECT 3383.840 2199.175 3384.490 2199.345 ;
        RECT 3384.320 2198.505 3384.490 2199.175 ;
        RECT 3383.840 2198.335 3384.490 2198.505 ;
        RECT 3384.320 2197.750 3384.490 2198.335 ;
        RECT 3385.030 2200.015 3386.050 2200.185 ;
        RECT 3385.030 2199.345 3385.200 2200.015 ;
        RECT 3385.030 2199.175 3386.050 2199.345 ;
        RECT 3385.030 2198.505 3385.200 2199.175 ;
        RECT 3385.030 2198.335 3386.050 2198.505 ;
        RECT 3385.030 2197.750 3385.200 2198.335 ;
        RECT 3384.320 2197.665 3385.200 2197.750 ;
        RECT 3383.840 2197.495 3386.050 2197.665 ;
      LAYER mcon ;
        RECT 3384.350 2197.580 3385.200 2197.750 ;
      LAYER met1 ;
        RECT 3369.320 2197.550 3369.580 2197.870 ;
        RECT 3369.440 1074.250 3369.580 2197.550 ;
        RECT 3384.290 2197.530 3385.260 2197.790 ;
      LAYER via ;
        RECT 3369.320 2197.580 3369.580 2197.840 ;
        RECT 3384.350 2197.530 3385.200 2197.790 ;
      LAYER met2 ;
        RECT 3369.290 2197.720 3369.610 2197.840 ;
        RECT 3384.350 2197.720 3385.200 2197.820 ;
        RECT 3368.850 2197.580 3385.200 2197.720 ;
        RECT 3384.350 2197.500 3385.200 2197.580 ;
    END
  END mgmt_io_in_buf[7]
  PIN mgmt_io_in_unbuf[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 851.350 4981.710 852.940 4981.910 ;
      LAYER mcon ;
        RECT 851.850 4981.740 852.940 4981.910 ;
      LAYER met1 ;
        RECT 851.790 4981.690 853.000 4981.950 ;
        RECT 852.315 4977.145 852.635 4977.265 ;
        RECT 852.315 4977.005 860.545 4977.145 ;
      LAYER via ;
        RECT 851.850 4981.690 852.940 4981.950 ;
        RECT 852.345 4977.005 852.605 4977.265 ;
      LAYER met2 ;
        RECT 851.850 4981.660 852.940 4981.980 ;
        RECT 852.345 4977.295 852.485 4981.660 ;
        RECT 852.345 4976.975 852.605 4977.295 ;
        RECT 852.345 4975.520 852.485 4976.975 ;
    END
  END mgmt_io_in_unbuf[19]
  PIN mgmt_io_in_unbuf[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 845.370 4981.710 846.960 4981.910 ;
      LAYER mcon ;
        RECT 845.870 4981.740 846.960 4981.910 ;
      LAYER met1 ;
        RECT 845.810 4981.690 847.020 4981.950 ;
        RECT 846.215 4976.585 846.535 4976.705 ;
        RECT 846.215 4976.445 858.555 4976.585 ;
      LAYER via ;
        RECT 845.870 4981.690 846.960 4981.950 ;
        RECT 846.245 4976.445 846.505 4976.705 ;
      LAYER met2 ;
        RECT 845.870 4981.660 846.960 4981.980 ;
        RECT 846.365 4976.735 846.505 4981.660 ;
        RECT 846.245 4976.415 846.505 4976.735 ;
        RECT 846.365 4975.520 846.505 4976.415 ;
    END
  END mgmt_io_in_unbuf[20]
  PIN mgmt_io_in_unbuf[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 839.390 4981.710 840.980 4981.910 ;
      LAYER mcon ;
        RECT 839.890 4981.740 840.980 4981.910 ;
      LAYER met1 ;
        RECT 839.830 4981.690 841.040 4981.950 ;
        RECT 840.355 4976.025 840.675 4976.145 ;
        RECT 840.355 4975.885 856.550 4976.025 ;
      LAYER via ;
        RECT 839.890 4981.690 840.980 4981.950 ;
        RECT 840.385 4975.885 840.645 4976.145 ;
      LAYER met2 ;
        RECT 839.890 4981.660 840.980 4981.980 ;
        RECT 840.385 4976.175 840.525 4981.660 ;
        RECT 840.385 4975.855 840.645 4976.175 ;
        RECT 840.385 4975.520 840.525 4975.855 ;
    END
  END mgmt_io_in_unbuf[21]
  PIN mgmt_io_out_buf[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 836.965 4985.340 837.135 4985.820 ;
        RECT 837.805 4985.340 837.975 4985.820 ;
        RECT 838.645 4985.340 838.815 4985.820 ;
        RECT 839.485 4985.340 839.655 4985.820 ;
        RECT 836.965 4985.170 839.655 4985.340 ;
        RECT 839.400 4984.630 839.655 4985.170 ;
        RECT 836.965 4984.460 839.655 4984.630 ;
        RECT 836.965 4983.610 837.135 4984.460 ;
        RECT 837.805 4983.610 837.975 4984.460 ;
        RECT 838.645 4983.610 838.815 4984.460 ;
        RECT 839.485 4983.610 839.655 4984.460 ;
      LAYER mcon ;
        RECT 839.400 4984.460 839.570 4985.310 ;
      LAYER met1 ;
        RECT 839.350 4984.400 839.610 4985.370 ;
        RECT 839.385 4975.745 839.705 4975.865 ;
        RECT 839.385 4975.605 855.550 4975.745 ;
      LAYER via ;
        RECT 839.350 4984.460 839.610 4985.310 ;
        RECT 839.415 4975.605 839.675 4975.865 ;
      LAYER met2 ;
        RECT 839.320 4984.460 839.640 4985.310 ;
        RECT 839.415 4975.895 839.555 4984.460 ;
        RECT 839.415 4975.575 839.675 4975.895 ;
        RECT 839.415 4975.520 839.555 4975.575 ;
    END
  END mgmt_io_out_buf[21]
  PIN mgmt_io_out_buf[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 842.945 4985.340 843.115 4985.820 ;
        RECT 843.785 4985.340 843.955 4985.820 ;
        RECT 844.625 4985.340 844.795 4985.820 ;
        RECT 845.465 4985.340 845.635 4985.820 ;
        RECT 842.945 4985.170 845.635 4985.340 ;
        RECT 845.380 4984.630 845.635 4985.170 ;
        RECT 842.945 4984.460 845.635 4984.630 ;
        RECT 842.945 4983.610 843.115 4984.460 ;
        RECT 843.785 4983.610 843.955 4984.460 ;
        RECT 844.625 4983.610 844.795 4984.460 ;
        RECT 845.465 4983.610 845.635 4984.460 ;
      LAYER mcon ;
        RECT 845.380 4984.460 845.550 4985.310 ;
      LAYER met1 ;
        RECT 845.330 4984.400 845.590 4985.370 ;
        RECT 845.365 4976.305 845.685 4976.425 ;
        RECT 845.365 4976.165 857.555 4976.305 ;
      LAYER via ;
        RECT 845.330 4984.460 845.590 4985.310 ;
        RECT 845.395 4976.165 845.655 4976.425 ;
      LAYER met2 ;
        RECT 845.300 4984.460 845.620 4985.310 ;
        RECT 845.395 4976.455 845.535 4984.460 ;
        RECT 845.395 4976.135 845.655 4976.455 ;
        RECT 845.395 4975.520 845.535 4976.135 ;
    END
  END mgmt_io_out_buf[20]
  PIN mgmt_io_out_buf[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 848.925 4985.340 849.095 4985.820 ;
        RECT 849.765 4985.340 849.935 4985.820 ;
        RECT 850.605 4985.340 850.775 4985.820 ;
        RECT 851.445 4985.340 851.615 4985.820 ;
        RECT 848.925 4985.170 851.615 4985.340 ;
        RECT 851.360 4984.630 851.615 4985.170 ;
        RECT 848.925 4984.460 851.615 4984.630 ;
        RECT 848.925 4983.610 849.095 4984.460 ;
        RECT 849.765 4983.610 849.935 4984.460 ;
        RECT 850.605 4983.610 850.775 4984.460 ;
        RECT 851.445 4983.610 851.615 4984.460 ;
      LAYER mcon ;
        RECT 851.360 4984.460 851.530 4985.310 ;
      LAYER met1 ;
        RECT 851.310 4984.400 851.570 4985.370 ;
        RECT 851.345 4976.865 851.665 4976.985 ;
        RECT 851.345 4976.725 859.545 4976.865 ;
      LAYER via ;
        RECT 851.310 4984.460 851.570 4985.310 ;
        RECT 851.375 4976.725 851.635 4976.985 ;
      LAYER met2 ;
        RECT 851.280 4984.460 851.600 4985.310 ;
        RECT 851.375 4977.015 851.515 4984.460 ;
        RECT 851.375 4976.695 851.635 4977.015 ;
        RECT 851.375 4975.520 851.515 4976.695 ;
    END
  END mgmt_io_out_buf[19]
  PIN mgmt_io_out_buf[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 198.900 4437.655 201.110 4437.825 ;
        RECT 199.380 4437.570 200.260 4437.655 ;
        RECT 199.380 4436.985 199.550 4437.570 ;
        RECT 198.900 4436.815 199.550 4436.985 ;
        RECT 199.380 4436.145 199.550 4436.815 ;
        RECT 198.900 4435.975 199.550 4436.145 ;
        RECT 199.380 4435.305 199.550 4435.975 ;
        RECT 198.900 4435.135 199.550 4435.305 ;
        RECT 200.090 4436.985 200.260 4437.570 ;
        RECT 200.090 4436.815 201.110 4436.985 ;
        RECT 200.090 4436.145 200.260 4436.815 ;
        RECT 200.090 4435.975 201.110 4436.145 ;
        RECT 200.090 4435.305 200.260 4435.975 ;
        RECT 200.090 4435.135 201.110 4435.305 ;
      LAYER mcon ;
        RECT 199.410 4437.570 200.260 4437.740 ;
      LAYER met1 ;
        RECT 214.415 4437.875 214.555 4461.585 ;
        RECT 199.350 4437.520 200.320 4437.780 ;
        RECT 214.295 4437.555 214.555 4437.875 ;
      LAYER via ;
        RECT 199.410 4437.520 200.260 4437.780 ;
        RECT 214.295 4437.585 214.555 4437.845 ;
      LAYER met2 ;
        RECT 199.410 4437.725 200.260 4437.810 ;
        RECT 214.265 4437.725 214.585 4437.845 ;
        RECT 199.410 4437.585 215.175 4437.725 ;
        RECT 199.410 4437.490 200.260 4437.585 ;
    END
  END mgmt_io_out_buf[22]
  PIN mgmt_io_out_buf[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 198.900 4431.675 201.110 4431.845 ;
        RECT 199.380 4431.590 200.260 4431.675 ;
        RECT 199.380 4431.005 199.550 4431.590 ;
        RECT 198.900 4430.835 199.550 4431.005 ;
        RECT 199.380 4430.165 199.550 4430.835 ;
        RECT 198.900 4429.995 199.550 4430.165 ;
        RECT 199.380 4429.325 199.550 4429.995 ;
        RECT 198.900 4429.155 199.550 4429.325 ;
        RECT 200.090 4431.005 200.260 4431.590 ;
        RECT 200.090 4430.835 201.110 4431.005 ;
        RECT 200.090 4430.165 200.260 4430.835 ;
        RECT 200.090 4429.995 201.110 4430.165 ;
        RECT 200.090 4429.325 200.260 4429.995 ;
        RECT 200.090 4429.155 201.110 4429.325 ;
      LAYER mcon ;
        RECT 199.410 4431.590 200.260 4431.760 ;
      LAYER met1 ;
        RECT 214.975 4431.895 215.115 4459.585 ;
        RECT 199.350 4431.540 200.320 4431.800 ;
        RECT 214.855 4431.575 215.115 4431.895 ;
      LAYER via ;
        RECT 199.410 4431.540 200.260 4431.800 ;
        RECT 214.855 4431.605 215.115 4431.865 ;
      LAYER met2 ;
        RECT 199.410 4431.745 200.260 4431.830 ;
        RECT 214.825 4431.745 215.145 4431.865 ;
        RECT 199.410 4431.605 215.175 4431.745 ;
        RECT 199.410 4431.510 200.260 4431.605 ;
    END
  END mgmt_io_out_buf[23]
  PIN mgmt_io_in_unbuf[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.810 4431.580 203.010 4433.170 ;
      LAYER mcon ;
        RECT 202.810 4432.080 202.980 4433.170 ;
      LAYER met1 ;
        RECT 202.770 4432.020 203.030 4433.230 ;
        RECT 214.695 4432.865 214.835 4460.585 ;
        RECT 214.575 4432.545 214.835 4432.865 ;
      LAYER via ;
        RECT 202.770 4432.080 203.030 4433.170 ;
        RECT 214.575 4432.575 214.835 4432.835 ;
      LAYER met2 ;
        RECT 202.740 4432.715 203.060 4433.170 ;
        RECT 214.545 4432.715 214.865 4432.835 ;
        RECT 202.740 4432.575 215.175 4432.715 ;
        RECT 202.740 4432.080 203.060 4432.575 ;
    END
  END mgmt_io_in_unbuf[23]
  PIN mgmt_io_in_unbuf[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.810 4437.560 203.010 4439.150 ;
      LAYER mcon ;
        RECT 202.810 4438.060 202.980 4439.150 ;
      LAYER met1 ;
        RECT 202.770 4438.000 203.030 4439.210 ;
        RECT 214.135 4438.725 214.275 4462.585 ;
        RECT 214.015 4438.405 214.275 4438.725 ;
      LAYER via ;
        RECT 202.770 4438.060 203.030 4439.150 ;
        RECT 214.015 4438.435 214.275 4438.695 ;
      LAYER met2 ;
        RECT 202.740 4438.695 203.060 4439.150 ;
        RECT 202.740 4438.555 215.175 4438.695 ;
        RECT 202.740 4438.060 203.060 4438.555 ;
        RECT 213.985 4438.435 214.305 4438.555 ;
    END
  END mgmt_io_in_unbuf[22]
  PIN mgmt_io_out_buf[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 199.025 3022.465 201.235 3022.635 ;
        RECT 199.505 3022.380 200.385 3022.465 ;
        RECT 199.505 3021.795 199.675 3022.380 ;
        RECT 199.025 3021.625 199.675 3021.795 ;
        RECT 199.505 3020.955 199.675 3021.625 ;
        RECT 199.025 3020.785 199.675 3020.955 ;
        RECT 199.505 3020.115 199.675 3020.785 ;
        RECT 199.025 3019.945 199.675 3020.115 ;
        RECT 200.215 3021.795 200.385 3022.380 ;
        RECT 200.215 3021.625 201.235 3021.795 ;
        RECT 200.215 3020.955 200.385 3021.625 ;
        RECT 200.215 3020.785 201.235 3020.955 ;
        RECT 200.215 3020.115 200.385 3020.785 ;
        RECT 200.215 3019.945 201.235 3020.115 ;
      LAYER mcon ;
        RECT 199.535 3022.380 200.385 3022.550 ;
      LAYER met1 ;
        RECT 215.395 3022.685 215.535 3066.780 ;
        RECT 199.475 3022.330 200.445 3022.590 ;
        RECT 215.275 3022.365 215.535 3022.685 ;
      LAYER via ;
        RECT 199.535 3022.330 200.385 3022.590 ;
        RECT 215.275 3022.395 215.535 3022.655 ;
      LAYER met2 ;
        RECT 199.535 3022.535 200.385 3022.620 ;
        RECT 215.245 3022.535 215.565 3022.655 ;
        RECT 199.535 3022.395 218.400 3022.535 ;
        RECT 199.535 3022.300 200.385 3022.395 ;
    END
  END mgmt_io_out_buf[24]
  PIN mgmt_io_out_buf[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 199.025 3016.485 201.235 3016.655 ;
        RECT 199.505 3016.400 200.385 3016.485 ;
        RECT 199.505 3015.815 199.675 3016.400 ;
        RECT 199.025 3015.645 199.675 3015.815 ;
        RECT 199.505 3014.975 199.675 3015.645 ;
        RECT 199.025 3014.805 199.675 3014.975 ;
        RECT 199.505 3014.135 199.675 3014.805 ;
        RECT 199.025 3013.965 199.675 3014.135 ;
        RECT 200.215 3015.815 200.385 3016.400 ;
        RECT 200.215 3015.645 201.235 3015.815 ;
        RECT 200.215 3014.975 200.385 3015.645 ;
        RECT 200.215 3014.805 201.235 3014.975 ;
        RECT 200.215 3014.135 200.385 3014.805 ;
        RECT 200.215 3013.965 201.235 3014.135 ;
      LAYER mcon ;
        RECT 199.535 3016.400 200.385 3016.570 ;
      LAYER met1 ;
        RECT 215.955 3016.705 216.095 3064.780 ;
        RECT 199.475 3016.350 200.445 3016.610 ;
        RECT 215.835 3016.385 216.095 3016.705 ;
      LAYER via ;
        RECT 199.535 3016.350 200.385 3016.610 ;
        RECT 215.835 3016.415 216.095 3016.675 ;
      LAYER met2 ;
        RECT 199.535 3016.555 200.385 3016.640 ;
        RECT 215.805 3016.555 216.125 3016.675 ;
        RECT 199.535 3016.415 218.400 3016.555 ;
        RECT 199.535 3016.320 200.385 3016.415 ;
    END
  END mgmt_io_out_buf[25]
  PIN mgmt_io_out_buf[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 199.025 3010.505 201.235 3010.675 ;
        RECT 199.505 3010.420 200.385 3010.505 ;
        RECT 199.505 3009.835 199.675 3010.420 ;
        RECT 199.025 3009.665 199.675 3009.835 ;
        RECT 199.505 3008.995 199.675 3009.665 ;
        RECT 199.025 3008.825 199.675 3008.995 ;
        RECT 199.505 3008.155 199.675 3008.825 ;
        RECT 199.025 3007.985 199.675 3008.155 ;
        RECT 200.215 3009.835 200.385 3010.420 ;
        RECT 200.215 3009.665 201.235 3009.835 ;
        RECT 200.215 3008.995 200.385 3009.665 ;
        RECT 200.215 3008.825 201.235 3008.995 ;
        RECT 200.215 3008.155 200.385 3008.825 ;
        RECT 200.215 3007.985 201.235 3008.155 ;
      LAYER mcon ;
        RECT 199.535 3010.420 200.385 3010.590 ;
      LAYER met1 ;
        RECT 216.515 3010.725 216.655 3062.780 ;
        RECT 199.475 3010.370 200.445 3010.630 ;
        RECT 216.395 3010.405 216.655 3010.725 ;
      LAYER via ;
        RECT 199.535 3010.370 200.385 3010.630 ;
        RECT 216.395 3010.435 216.655 3010.695 ;
      LAYER met2 ;
        RECT 199.535 3010.575 200.385 3010.660 ;
        RECT 216.365 3010.575 216.685 3010.695 ;
        RECT 199.535 3010.435 218.400 3010.575 ;
        RECT 199.535 3010.340 200.385 3010.435 ;
    END
  END mgmt_io_out_buf[26]
  PIN mgmt_io_out_buf[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 199.025 3004.525 201.235 3004.695 ;
        RECT 199.505 3004.440 200.385 3004.525 ;
        RECT 199.505 3003.855 199.675 3004.440 ;
        RECT 199.025 3003.685 199.675 3003.855 ;
        RECT 199.505 3003.015 199.675 3003.685 ;
        RECT 199.025 3002.845 199.675 3003.015 ;
        RECT 199.505 3002.175 199.675 3002.845 ;
        RECT 199.025 3002.005 199.675 3002.175 ;
        RECT 200.215 3003.855 200.385 3004.440 ;
        RECT 200.215 3003.685 201.235 3003.855 ;
        RECT 200.215 3003.015 200.385 3003.685 ;
        RECT 200.215 3002.845 201.235 3003.015 ;
        RECT 200.215 3002.175 200.385 3002.845 ;
        RECT 200.215 3002.005 201.235 3002.175 ;
      LAYER mcon ;
        RECT 199.535 3004.440 200.385 3004.610 ;
      LAYER met1 ;
        RECT 217.075 3004.745 217.215 3060.780 ;
        RECT 199.475 3004.390 200.445 3004.650 ;
        RECT 216.955 3004.425 217.215 3004.745 ;
      LAYER via ;
        RECT 199.535 3004.390 200.385 3004.650 ;
        RECT 216.955 3004.455 217.215 3004.715 ;
      LAYER met2 ;
        RECT 199.535 3004.595 200.385 3004.680 ;
        RECT 216.925 3004.595 217.245 3004.715 ;
        RECT 199.535 3004.455 218.400 3004.595 ;
        RECT 199.535 3004.360 200.385 3004.455 ;
    END
  END mgmt_io_out_buf[27]
  PIN mgmt_io_out_buf[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 199.025 2998.545 201.235 2998.715 ;
        RECT 199.505 2998.460 200.385 2998.545 ;
        RECT 199.505 2997.875 199.675 2998.460 ;
        RECT 199.025 2997.705 199.675 2997.875 ;
        RECT 199.505 2997.035 199.675 2997.705 ;
        RECT 199.025 2996.865 199.675 2997.035 ;
        RECT 199.505 2996.195 199.675 2996.865 ;
        RECT 199.025 2996.025 199.675 2996.195 ;
        RECT 200.215 2997.875 200.385 2998.460 ;
        RECT 200.215 2997.705 201.235 2997.875 ;
        RECT 200.215 2997.035 200.385 2997.705 ;
        RECT 200.215 2996.865 201.235 2997.035 ;
        RECT 200.215 2996.195 200.385 2996.865 ;
        RECT 200.215 2996.025 201.235 2996.195 ;
      LAYER mcon ;
        RECT 199.535 2998.460 200.385 2998.630 ;
      LAYER met1 ;
        RECT 217.635 2998.765 217.775 3058.780 ;
        RECT 199.475 2998.410 200.445 2998.670 ;
        RECT 217.515 2998.445 217.775 2998.765 ;
      LAYER via ;
        RECT 199.535 2998.410 200.385 2998.670 ;
        RECT 217.515 2998.475 217.775 2998.735 ;
      LAYER met2 ;
        RECT 199.535 2998.615 200.385 2998.700 ;
        RECT 217.485 2998.615 217.805 2998.735 ;
        RECT 199.535 2998.475 218.400 2998.615 ;
        RECT 199.535 2998.380 200.385 2998.475 ;
    END
  END mgmt_io_out_buf[28]
  PIN mgmt_io_out_buf[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 199.025 2992.565 201.235 2992.735 ;
        RECT 199.505 2992.480 200.385 2992.565 ;
        RECT 199.505 2991.895 199.675 2992.480 ;
        RECT 199.025 2991.725 199.675 2991.895 ;
        RECT 199.505 2991.055 199.675 2991.725 ;
        RECT 199.025 2990.885 199.675 2991.055 ;
        RECT 199.505 2990.215 199.675 2990.885 ;
        RECT 199.025 2990.045 199.675 2990.215 ;
        RECT 200.215 2991.895 200.385 2992.480 ;
        RECT 200.215 2991.725 201.235 2991.895 ;
        RECT 200.215 2991.055 200.385 2991.725 ;
        RECT 200.215 2990.885 201.235 2991.055 ;
        RECT 200.215 2990.215 200.385 2990.885 ;
        RECT 200.215 2990.045 201.235 2990.215 ;
      LAYER mcon ;
        RECT 199.535 2992.480 200.385 2992.650 ;
      LAYER met1 ;
        RECT 218.195 2992.785 218.335 3056.780 ;
        RECT 199.475 2992.430 200.445 2992.690 ;
        RECT 218.075 2992.465 218.335 2992.785 ;
      LAYER via ;
        RECT 199.535 2992.430 200.385 2992.690 ;
        RECT 218.075 2992.495 218.335 2992.755 ;
      LAYER met2 ;
        RECT 199.535 2992.635 200.385 2992.720 ;
        RECT 218.045 2992.635 218.365 2992.755 ;
        RECT 199.535 2992.495 218.400 2992.635 ;
        RECT 199.535 2992.400 200.385 2992.495 ;
    END
  END mgmt_io_out_buf[29]
  PIN mgmt_io_in_unbuf[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.935 2992.470 203.135 2994.060 ;
      LAYER mcon ;
        RECT 202.935 2992.970 203.105 2994.060 ;
      LAYER met1 ;
        RECT 202.895 2992.910 203.155 2994.120 ;
        RECT 217.915 2993.755 218.055 3057.780 ;
        RECT 217.795 2993.435 218.055 2993.755 ;
      LAYER via ;
        RECT 202.895 2992.970 203.155 2994.060 ;
        RECT 217.795 2993.465 218.055 2993.725 ;
      LAYER met2 ;
        RECT 202.865 2993.605 203.185 2994.060 ;
        RECT 217.765 2993.605 218.085 2993.725 ;
        RECT 202.865 2993.465 218.400 2993.605 ;
        RECT 202.865 2992.970 203.185 2993.465 ;
    END
  END mgmt_io_in_unbuf[29]
  PIN mgmt_io_in_unbuf[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.935 2998.450 203.135 3000.040 ;
      LAYER mcon ;
        RECT 202.935 2998.950 203.105 3000.040 ;
      LAYER met1 ;
        RECT 202.895 2998.890 203.155 3000.100 ;
        RECT 217.355 2999.735 217.495 3059.780 ;
        RECT 217.235 2999.415 217.495 2999.735 ;
      LAYER via ;
        RECT 202.895 2998.950 203.155 3000.040 ;
        RECT 217.235 2999.445 217.495 2999.705 ;
      LAYER met2 ;
        RECT 202.865 2999.585 203.185 3000.040 ;
        RECT 217.205 2999.585 217.525 2999.705 ;
        RECT 202.865 2999.445 218.400 2999.585 ;
        RECT 202.865 2998.950 203.185 2999.445 ;
    END
  END mgmt_io_in_unbuf[28]
  PIN mgmt_io_in_unbuf[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.935 3004.430 203.135 3006.020 ;
      LAYER mcon ;
        RECT 202.935 3004.930 203.105 3006.020 ;
      LAYER met1 ;
        RECT 202.895 3004.870 203.155 3006.080 ;
        RECT 216.795 3005.715 216.935 3061.780 ;
        RECT 216.675 3005.395 216.935 3005.715 ;
      LAYER via ;
        RECT 202.895 3004.930 203.155 3006.020 ;
        RECT 216.675 3005.425 216.935 3005.685 ;
      LAYER met2 ;
        RECT 202.865 3005.565 203.185 3006.020 ;
        RECT 216.645 3005.565 216.965 3005.685 ;
        RECT 202.865 3005.425 218.400 3005.565 ;
        RECT 202.865 3004.930 203.185 3005.425 ;
    END
  END mgmt_io_in_unbuf[27]
  PIN mgmt_io_in_unbuf[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.935 3010.410 203.135 3012.000 ;
      LAYER mcon ;
        RECT 202.935 3010.910 203.105 3012.000 ;
      LAYER met1 ;
        RECT 202.895 3010.850 203.155 3012.060 ;
        RECT 216.235 3011.695 216.375 3063.780 ;
        RECT 216.115 3011.375 216.375 3011.695 ;
      LAYER via ;
        RECT 202.895 3010.910 203.155 3012.000 ;
        RECT 216.115 3011.405 216.375 3011.665 ;
      LAYER met2 ;
        RECT 202.865 3011.545 203.185 3012.000 ;
        RECT 216.085 3011.545 216.405 3011.665 ;
        RECT 202.865 3011.405 218.400 3011.545 ;
        RECT 202.865 3010.910 203.185 3011.405 ;
    END
  END mgmt_io_in_unbuf[26]
  PIN mgmt_io_in_unbuf[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.935 3016.390 203.135 3017.980 ;
      LAYER mcon ;
        RECT 202.935 3016.890 203.105 3017.980 ;
      LAYER met1 ;
        RECT 202.895 3016.830 203.155 3018.040 ;
        RECT 215.675 3017.675 215.815 3065.780 ;
        RECT 215.555 3017.355 215.815 3017.675 ;
      LAYER via ;
        RECT 202.895 3016.890 203.155 3017.980 ;
        RECT 215.555 3017.385 215.815 3017.645 ;
      LAYER met2 ;
        RECT 202.865 3017.525 203.185 3017.980 ;
        RECT 215.525 3017.525 215.845 3017.645 ;
        RECT 202.865 3017.385 218.400 3017.525 ;
        RECT 202.865 3016.890 203.185 3017.385 ;
    END
  END mgmt_io_in_unbuf[25]
  PIN mgmt_io_in_unbuf[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 202.935 3022.370 203.135 3023.960 ;
      LAYER mcon ;
        RECT 202.935 3022.870 203.105 3023.960 ;
      LAYER met1 ;
        RECT 202.895 3022.810 203.155 3024.020 ;
        RECT 215.115 3023.655 215.255 3067.780 ;
        RECT 214.995 3023.335 215.255 3023.655 ;
      LAYER via ;
        RECT 202.895 3022.870 203.155 3023.960 ;
        RECT 214.995 3023.365 215.255 3023.625 ;
      LAYER met2 ;
        RECT 202.865 3023.505 203.185 3023.960 ;
        RECT 214.965 3023.505 215.285 3023.625 ;
        RECT 202.865 3023.365 218.400 3023.505 ;
        RECT 202.865 3022.870 203.185 3023.365 ;
    END
  END mgmt_io_in_unbuf[24]
  PIN mgmt_io_out_buf[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 199.135 1695.680 201.345 1695.850 ;
        RECT 199.615 1695.595 200.495 1695.680 ;
        RECT 199.615 1695.010 199.785 1695.595 ;
        RECT 199.135 1694.840 199.785 1695.010 ;
        RECT 199.615 1694.170 199.785 1694.840 ;
        RECT 199.135 1694.000 199.785 1694.170 ;
        RECT 199.615 1693.330 199.785 1694.000 ;
        RECT 199.135 1693.160 199.785 1693.330 ;
        RECT 200.325 1695.010 200.495 1695.595 ;
        RECT 200.325 1694.840 201.345 1695.010 ;
        RECT 200.325 1694.170 200.495 1694.840 ;
        RECT 200.325 1694.000 201.345 1694.170 ;
        RECT 200.325 1693.330 200.495 1694.000 ;
        RECT 200.325 1693.160 201.345 1693.330 ;
      LAYER mcon ;
        RECT 199.645 1695.595 200.495 1695.765 ;
      LAYER met1 ;
        RECT 218.615 1695.900 218.755 1772.650 ;
        RECT 199.585 1695.545 200.555 1695.805 ;
        RECT 218.495 1695.580 218.755 1695.900 ;
      LAYER via ;
        RECT 199.645 1695.545 200.495 1695.805 ;
        RECT 218.495 1695.610 218.755 1695.870 ;
      LAYER met2 ;
        RECT 199.645 1695.750 200.495 1695.835 ;
        RECT 218.465 1695.750 218.785 1695.870 ;
        RECT 199.645 1695.610 220.540 1695.750 ;
        RECT 199.645 1695.515 200.495 1695.610 ;
    END
  END mgmt_io_out_buf[30]
  PIN mgmt_io_out_buf[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 199.135 1689.700 201.345 1689.870 ;
        RECT 199.615 1689.615 200.495 1689.700 ;
        RECT 199.615 1689.030 199.785 1689.615 ;
        RECT 199.135 1688.860 199.785 1689.030 ;
        RECT 199.615 1688.190 199.785 1688.860 ;
        RECT 199.135 1688.020 199.785 1688.190 ;
        RECT 199.615 1687.350 199.785 1688.020 ;
        RECT 199.135 1687.180 199.785 1687.350 ;
        RECT 200.325 1689.030 200.495 1689.615 ;
        RECT 200.325 1688.860 201.345 1689.030 ;
        RECT 200.325 1688.190 200.495 1688.860 ;
        RECT 200.325 1688.020 201.345 1688.190 ;
        RECT 200.325 1687.350 200.495 1688.020 ;
        RECT 200.325 1687.180 201.345 1687.350 ;
      LAYER mcon ;
        RECT 199.645 1689.615 200.495 1689.785 ;
      LAYER met1 ;
        RECT 219.175 1689.920 219.315 1770.650 ;
        RECT 199.585 1689.565 200.555 1689.825 ;
        RECT 219.055 1689.600 219.315 1689.920 ;
      LAYER via ;
        RECT 199.645 1689.565 200.495 1689.825 ;
        RECT 219.055 1689.630 219.315 1689.890 ;
      LAYER met2 ;
        RECT 199.645 1689.770 200.495 1689.855 ;
        RECT 219.025 1689.770 219.345 1689.890 ;
        RECT 199.645 1689.630 220.540 1689.770 ;
        RECT 199.645 1689.535 200.495 1689.630 ;
    END
  END mgmt_io_out_buf[31]
  PIN mgmt_io_out_buf[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 199.135 1683.720 201.345 1683.890 ;
        RECT 199.615 1683.635 200.495 1683.720 ;
        RECT 199.615 1683.050 199.785 1683.635 ;
        RECT 199.135 1682.880 199.785 1683.050 ;
        RECT 199.615 1682.210 199.785 1682.880 ;
        RECT 199.135 1682.040 199.785 1682.210 ;
        RECT 199.615 1681.370 199.785 1682.040 ;
        RECT 199.135 1681.200 199.785 1681.370 ;
        RECT 200.325 1683.050 200.495 1683.635 ;
        RECT 200.325 1682.880 201.345 1683.050 ;
        RECT 200.325 1682.210 200.495 1682.880 ;
        RECT 200.325 1682.040 201.345 1682.210 ;
        RECT 200.325 1681.370 200.495 1682.040 ;
        RECT 200.325 1681.200 201.345 1681.370 ;
      LAYER mcon ;
        RECT 199.645 1683.635 200.495 1683.805 ;
      LAYER met1 ;
        RECT 219.735 1683.940 219.875 1768.650 ;
        RECT 199.585 1683.585 200.555 1683.845 ;
        RECT 219.615 1683.620 219.875 1683.940 ;
      LAYER via ;
        RECT 199.645 1683.585 200.495 1683.845 ;
        RECT 219.615 1683.650 219.875 1683.910 ;
      LAYER met2 ;
        RECT 199.645 1683.790 200.495 1683.875 ;
        RECT 219.585 1683.790 219.905 1683.910 ;
        RECT 199.645 1683.650 220.540 1683.790 ;
        RECT 199.645 1683.555 200.495 1683.650 ;
    END
  END mgmt_io_out_buf[32]
  PIN mgmt_io_out_buf[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 199.135 1677.740 201.345 1677.910 ;
        RECT 199.615 1677.655 200.495 1677.740 ;
        RECT 199.615 1677.070 199.785 1677.655 ;
        RECT 199.135 1676.900 199.785 1677.070 ;
        RECT 199.615 1676.230 199.785 1676.900 ;
        RECT 199.135 1676.060 199.785 1676.230 ;
        RECT 199.615 1675.390 199.785 1676.060 ;
        RECT 199.135 1675.220 199.785 1675.390 ;
        RECT 200.325 1677.070 200.495 1677.655 ;
        RECT 200.325 1676.900 201.345 1677.070 ;
        RECT 200.325 1676.230 200.495 1676.900 ;
        RECT 200.325 1676.060 201.345 1676.230 ;
        RECT 200.325 1675.390 200.495 1676.060 ;
        RECT 200.325 1675.220 201.345 1675.390 ;
      LAYER mcon ;
        RECT 199.645 1677.655 200.495 1677.825 ;
      LAYER met1 ;
        RECT 220.295 1677.960 220.435 1766.650 ;
        RECT 199.585 1677.605 200.555 1677.865 ;
        RECT 220.175 1677.640 220.435 1677.960 ;
      LAYER via ;
        RECT 199.645 1677.605 200.495 1677.865 ;
        RECT 220.175 1677.670 220.435 1677.930 ;
      LAYER met2 ;
        RECT 199.645 1677.810 200.495 1677.895 ;
        RECT 220.145 1677.810 220.465 1677.930 ;
        RECT 199.645 1677.670 220.540 1677.810 ;
        RECT 199.645 1677.575 200.495 1677.670 ;
    END
  END mgmt_io_out_buf[33]
  PIN mgmt_io_in_unbuf[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 203.045 1677.645 203.245 1679.235 ;
      LAYER mcon ;
        RECT 203.045 1678.145 203.215 1679.235 ;
      LAYER met1 ;
        RECT 203.005 1678.085 203.265 1679.295 ;
        RECT 220.015 1678.930 220.155 1767.650 ;
        RECT 219.895 1678.610 220.155 1678.930 ;
      LAYER via ;
        RECT 203.005 1678.145 203.265 1679.235 ;
        RECT 219.895 1678.640 220.155 1678.900 ;
      LAYER met2 ;
        RECT 202.975 1678.780 203.295 1679.235 ;
        RECT 219.865 1678.780 220.185 1678.900 ;
        RECT 202.975 1678.640 220.540 1678.780 ;
        RECT 202.975 1678.145 203.295 1678.640 ;
    END
  END mgmt_io_in_unbuf[33]
  PIN mgmt_io_in_unbuf[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 203.045 1683.625 203.245 1685.215 ;
      LAYER mcon ;
        RECT 203.045 1684.125 203.215 1685.215 ;
      LAYER met1 ;
        RECT 203.005 1684.065 203.265 1685.275 ;
        RECT 219.455 1684.790 219.595 1769.650 ;
        RECT 219.335 1684.470 219.595 1684.790 ;
      LAYER via ;
        RECT 203.005 1684.125 203.265 1685.215 ;
        RECT 219.335 1684.500 219.595 1684.760 ;
      LAYER met2 ;
        RECT 202.975 1684.760 203.295 1685.215 ;
        RECT 202.975 1684.620 220.540 1684.760 ;
        RECT 202.975 1684.125 203.295 1684.620 ;
        RECT 219.305 1684.500 219.625 1684.620 ;
    END
  END mgmt_io_in_unbuf[32]
  PIN mgmt_io_in_unbuf[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 203.045 1689.605 203.245 1691.195 ;
      LAYER mcon ;
        RECT 203.045 1690.105 203.215 1691.195 ;
      LAYER met1 ;
        RECT 203.005 1690.045 203.265 1691.255 ;
        RECT 218.895 1690.890 219.035 1771.650 ;
        RECT 218.775 1690.570 219.035 1690.890 ;
      LAYER via ;
        RECT 203.005 1690.105 203.265 1691.195 ;
        RECT 218.775 1690.600 219.035 1690.860 ;
      LAYER met2 ;
        RECT 202.975 1690.740 203.295 1691.195 ;
        RECT 218.745 1690.740 219.065 1690.860 ;
        RECT 202.975 1690.600 220.540 1690.740 ;
        RECT 202.975 1690.105 203.295 1690.600 ;
    END
  END mgmt_io_in_unbuf[31]
  PIN mgmt_io_in_unbuf[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 203.045 1695.585 203.245 1697.175 ;
      LAYER mcon ;
        RECT 203.045 1696.085 203.215 1697.175 ;
      LAYER met1 ;
        RECT 203.005 1696.025 203.265 1697.235 ;
        RECT 218.335 1696.870 218.475 1773.650 ;
        RECT 218.215 1696.550 218.475 1696.870 ;
      LAYER via ;
        RECT 203.005 1696.085 203.265 1697.175 ;
        RECT 218.215 1696.580 218.475 1696.840 ;
      LAYER met2 ;
        RECT 202.975 1696.720 203.295 1697.175 ;
        RECT 218.185 1696.720 218.505 1696.840 ;
        RECT 202.975 1696.580 220.540 1696.720 ;
        RECT 202.975 1696.085 203.295 1696.580 ;
    END
  END mgmt_io_in_unbuf[30]
  PIN mgmt_io_out_buf[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 760.135 1116.390 760.305 1116.870 ;
        RECT 760.975 1116.390 761.145 1116.870 ;
        RECT 761.815 1116.390 761.985 1116.870 ;
        RECT 762.655 1116.390 762.825 1116.870 ;
        RECT 760.135 1116.220 762.825 1116.390 ;
        RECT 760.135 1115.680 760.390 1116.220 ;
        RECT 760.135 1115.510 762.825 1115.680 ;
        RECT 760.135 1114.660 760.305 1115.510 ;
        RECT 760.975 1114.660 761.145 1115.510 ;
        RECT 761.815 1114.660 761.985 1115.510 ;
        RECT 762.655 1114.660 762.825 1115.510 ;
      LAYER mcon ;
        RECT 760.220 1115.510 760.390 1116.360 ;
      LAYER met1 ;
        RECT 760.190 1120.980 760.510 1121.100 ;
        RECT 655.615 1120.840 760.510 1120.980 ;
        RECT 760.170 1115.450 760.430 1116.420 ;
      LAYER via ;
        RECT 760.220 1120.840 760.480 1121.100 ;
        RECT 760.170 1115.510 760.430 1116.360 ;
      LAYER met2 ;
        RECT 760.220 1121.130 760.360 1129.625 ;
        RECT 760.220 1120.810 760.480 1121.130 ;
        RECT 760.220 1116.360 760.360 1120.810 ;
        RECT 760.140 1115.510 760.460 1116.360 ;
    END
  END mgmt_io_out_buf[34]
  PIN mgmt_io_out_buf[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 766.115 1116.390 766.285 1116.870 ;
        RECT 766.955 1116.390 767.125 1116.870 ;
        RECT 767.795 1116.390 767.965 1116.870 ;
        RECT 768.635 1116.390 768.805 1116.870 ;
        RECT 766.115 1116.220 768.805 1116.390 ;
        RECT 766.115 1115.680 766.370 1116.220 ;
        RECT 766.115 1115.510 768.805 1115.680 ;
        RECT 766.115 1114.660 766.285 1115.510 ;
        RECT 766.955 1114.660 767.125 1115.510 ;
        RECT 767.795 1114.660 767.965 1115.510 ;
        RECT 768.635 1114.660 768.805 1115.510 ;
      LAYER mcon ;
        RECT 766.200 1115.510 766.370 1116.360 ;
      LAYER met1 ;
        RECT 766.170 1120.420 766.490 1120.540 ;
        RECT 657.615 1120.280 766.490 1120.420 ;
        RECT 766.150 1115.450 766.410 1116.420 ;
      LAYER via ;
        RECT 766.200 1120.280 766.460 1120.540 ;
        RECT 766.150 1115.510 766.410 1116.360 ;
      LAYER met2 ;
        RECT 766.200 1120.570 766.340 1129.625 ;
        RECT 766.200 1120.250 766.460 1120.570 ;
        RECT 766.200 1116.360 766.340 1120.250 ;
        RECT 766.120 1115.510 766.440 1116.360 ;
    END
  END mgmt_io_out_buf[35]
  PIN mgmt_io_out_buf[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 772.095 1116.390 772.265 1116.870 ;
        RECT 772.935 1116.390 773.105 1116.870 ;
        RECT 773.775 1116.390 773.945 1116.870 ;
        RECT 774.615 1116.390 774.785 1116.870 ;
        RECT 772.095 1116.220 774.785 1116.390 ;
        RECT 772.095 1115.680 772.350 1116.220 ;
        RECT 772.095 1115.510 774.785 1115.680 ;
        RECT 772.095 1114.660 772.265 1115.510 ;
        RECT 772.935 1114.660 773.105 1115.510 ;
        RECT 773.775 1114.660 773.945 1115.510 ;
        RECT 774.615 1114.660 774.785 1115.510 ;
      LAYER mcon ;
        RECT 772.180 1115.510 772.350 1116.360 ;
      LAYER met1 ;
        RECT 772.150 1119.860 772.470 1119.980 ;
        RECT 659.615 1119.720 772.470 1119.860 ;
        RECT 772.130 1115.450 772.390 1116.420 ;
      LAYER via ;
        RECT 772.180 1119.720 772.440 1119.980 ;
        RECT 772.130 1115.510 772.390 1116.360 ;
      LAYER met2 ;
        RECT 772.180 1120.010 772.320 1129.625 ;
        RECT 772.180 1119.690 772.440 1120.010 ;
        RECT 772.180 1116.360 772.320 1119.690 ;
        RECT 772.100 1115.510 772.420 1116.360 ;
    END
  END mgmt_io_out_buf[36]
  PIN mgmt_io_out_buf[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 778.075 1116.390 778.245 1116.870 ;
        RECT 778.915 1116.390 779.085 1116.870 ;
        RECT 779.755 1116.390 779.925 1116.870 ;
        RECT 780.595 1116.390 780.765 1116.870 ;
        RECT 778.075 1116.220 780.765 1116.390 ;
        RECT 778.075 1115.680 778.330 1116.220 ;
        RECT 778.075 1115.510 780.765 1115.680 ;
        RECT 778.075 1114.660 778.245 1115.510 ;
        RECT 778.915 1114.660 779.085 1115.510 ;
        RECT 779.755 1114.660 779.925 1115.510 ;
        RECT 780.595 1114.660 780.765 1115.510 ;
      LAYER mcon ;
        RECT 778.160 1115.510 778.330 1116.360 ;
      LAYER met1 ;
        RECT 778.130 1119.300 778.450 1119.420 ;
        RECT 661.615 1119.160 778.450 1119.300 ;
        RECT 778.110 1115.450 778.370 1116.420 ;
      LAYER via ;
        RECT 778.160 1119.160 778.420 1119.420 ;
        RECT 778.110 1115.510 778.370 1116.360 ;
      LAYER met2 ;
        RECT 778.160 1119.450 778.300 1129.625 ;
        RECT 778.160 1119.130 778.420 1119.450 ;
        RECT 778.160 1116.360 778.300 1119.130 ;
        RECT 778.080 1115.510 778.400 1116.360 ;
    END
  END mgmt_io_out_buf[37]
  PIN mgmt_io_in_unbuf[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 783.220 1112.760 784.320 1112.960 ;
      LAYER mcon ;
        RECT 783.230 1112.790 784.320 1112.960 ;
      LAYER met1 ;
        RECT 783.490 1119.020 783.810 1119.140 ;
        RECT 662.615 1118.880 783.810 1119.020 ;
        RECT 783.170 1112.750 784.380 1113.010 ;
      LAYER via ;
        RECT 783.520 1118.880 783.780 1119.140 ;
        RECT 783.230 1112.750 784.320 1113.010 ;
      LAYER met2 ;
        RECT 783.520 1119.170 783.660 1129.625 ;
        RECT 783.520 1118.850 783.780 1119.170 ;
        RECT 783.520 1113.040 783.660 1118.850 ;
        RECT 783.230 1112.720 784.320 1113.040 ;
    END
  END mgmt_io_in_unbuf[37]
  PIN mgmt_io_in_unbuf[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 777.240 1112.760 778.340 1112.960 ;
      LAYER mcon ;
        RECT 777.250 1112.790 778.340 1112.960 ;
      LAYER met1 ;
        RECT 777.510 1119.580 777.830 1119.700 ;
        RECT 660.615 1119.440 777.830 1119.580 ;
        RECT 777.190 1112.750 778.400 1113.010 ;
      LAYER via ;
        RECT 777.540 1119.440 777.800 1119.700 ;
        RECT 777.250 1112.750 778.340 1113.010 ;
      LAYER met2 ;
        RECT 777.540 1119.730 777.680 1129.625 ;
        RECT 777.540 1119.410 777.800 1119.730 ;
        RECT 777.540 1113.040 777.680 1119.410 ;
        RECT 777.250 1112.720 778.340 1113.040 ;
    END
  END mgmt_io_in_unbuf[36]
  PIN mgmt_io_in_unbuf[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 771.260 1112.760 772.360 1112.960 ;
      LAYER mcon ;
        RECT 771.270 1112.790 772.360 1112.960 ;
      LAYER met1 ;
        RECT 771.530 1120.140 771.850 1120.260 ;
        RECT 658.615 1120.000 771.850 1120.140 ;
        RECT 771.210 1112.750 772.420 1113.010 ;
      LAYER via ;
        RECT 771.560 1120.000 771.820 1120.260 ;
        RECT 771.270 1112.750 772.360 1113.010 ;
      LAYER met2 ;
        RECT 771.560 1120.290 771.700 1129.625 ;
        RECT 771.560 1119.970 771.820 1120.290 ;
        RECT 771.560 1113.040 771.700 1119.970 ;
        RECT 771.270 1112.720 772.360 1113.040 ;
    END
  END mgmt_io_in_unbuf[35]
  PIN mgmt_io_in_unbuf[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 765.280 1112.760 766.380 1112.960 ;
      LAYER mcon ;
        RECT 765.290 1112.790 766.380 1112.960 ;
      LAYER met1 ;
        RECT 765.550 1120.700 765.870 1120.820 ;
        RECT 656.615 1120.560 765.870 1120.700 ;
        RECT 765.230 1112.750 766.440 1113.010 ;
      LAYER via ;
        RECT 765.580 1120.560 765.840 1120.820 ;
        RECT 765.290 1112.750 766.380 1113.010 ;
      LAYER met2 ;
        RECT 765.580 1120.850 765.720 1129.625 ;
        RECT 765.580 1120.530 765.840 1120.850 ;
        RECT 765.580 1113.040 765.720 1120.530 ;
        RECT 765.290 1112.720 766.380 1113.040 ;
    END
  END mgmt_io_in_unbuf[34]
  PIN mgmt_io_oeb_buf[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 784.055 1116.390 784.225 1116.870 ;
        RECT 784.895 1116.390 785.065 1116.870 ;
        RECT 785.735 1116.390 785.905 1116.870 ;
        RECT 786.575 1116.390 786.745 1116.870 ;
        RECT 784.055 1116.220 786.745 1116.390 ;
        RECT 784.055 1115.680 784.310 1116.220 ;
        RECT 784.055 1115.510 786.745 1115.680 ;
        RECT 784.055 1114.660 784.225 1115.510 ;
        RECT 784.895 1114.660 785.065 1115.510 ;
        RECT 785.735 1114.660 785.905 1115.510 ;
        RECT 786.575 1114.660 786.745 1115.510 ;
      LAYER mcon ;
        RECT 784.140 1115.510 784.310 1116.360 ;
      LAYER met1 ;
        RECT 784.110 1118.740 784.430 1118.860 ;
        RECT 663.615 1118.600 784.430 1118.740 ;
        RECT 784.090 1115.450 784.350 1116.420 ;
      LAYER via ;
        RECT 784.140 1118.600 784.400 1118.860 ;
        RECT 784.090 1115.510 784.350 1116.360 ;
      LAYER met2 ;
        RECT 784.140 1118.890 784.280 1129.625 ;
        RECT 784.140 1118.570 784.400 1118.890 ;
        RECT 784.140 1116.360 784.280 1118.570 ;
        RECT 784.060 1115.510 784.380 1116.360 ;
    END
  END mgmt_io_oeb_buf[35]
  PIN mgmt_io_oeb_buf[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 790.035 1113.300 790.205 1114.150 ;
        RECT 790.875 1113.300 791.045 1114.150 ;
        RECT 791.715 1113.300 791.885 1114.150 ;
        RECT 792.555 1113.300 792.725 1114.150 ;
        RECT 790.035 1113.130 792.725 1113.300 ;
        RECT 790.035 1112.590 790.290 1113.130 ;
        RECT 790.035 1112.420 792.725 1112.590 ;
        RECT 790.035 1111.940 790.205 1112.420 ;
        RECT 790.875 1111.940 791.045 1112.420 ;
        RECT 791.715 1111.940 791.885 1112.420 ;
        RECT 792.555 1111.940 792.725 1112.420 ;
      LAYER mcon ;
        RECT 790.120 1112.450 790.290 1113.300 ;
      LAYER met1 ;
        RECT 789.470 1118.460 789.790 1118.580 ;
        RECT 664.615 1118.320 789.790 1118.460 ;
        RECT 790.080 1112.390 790.340 1113.360 ;
      LAYER via ;
        RECT 789.500 1118.320 789.760 1118.580 ;
        RECT 790.080 1112.450 790.340 1113.300 ;
      LAYER met2 ;
        RECT 789.500 1118.610 789.640 1129.625 ;
        RECT 789.500 1118.290 789.760 1118.610 ;
        RECT 789.500 1114.240 789.640 1118.290 ;
        RECT 789.500 1114.100 790.275 1114.240 ;
        RECT 790.135 1113.300 790.275 1114.100 ;
        RECT 790.050 1112.450 790.370 1113.300 ;
    END
  END mgmt_io_oeb_buf[36]
  PIN mgmt_io_oeb_buf[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 790.035 1116.390 790.205 1116.870 ;
        RECT 790.875 1116.390 791.045 1116.870 ;
        RECT 791.715 1116.390 791.885 1116.870 ;
        RECT 792.555 1116.390 792.725 1116.870 ;
        RECT 790.035 1116.220 792.725 1116.390 ;
        RECT 790.035 1115.680 790.290 1116.220 ;
        RECT 790.035 1115.510 792.725 1115.680 ;
        RECT 790.035 1114.660 790.205 1115.510 ;
        RECT 790.875 1114.660 791.045 1115.510 ;
        RECT 791.715 1114.660 791.885 1115.510 ;
        RECT 792.555 1114.660 792.725 1115.510 ;
      LAYER mcon ;
        RECT 790.120 1115.510 790.290 1116.360 ;
      LAYER met1 ;
        RECT 790.090 1118.180 790.410 1118.300 ;
        RECT 665.615 1118.040 790.410 1118.180 ;
        RECT 790.070 1115.450 790.330 1116.420 ;
      LAYER via ;
        RECT 790.120 1118.040 790.380 1118.300 ;
        RECT 790.070 1115.510 790.330 1116.360 ;
      LAYER met2 ;
        RECT 790.120 1118.330 790.260 1129.625 ;
        RECT 790.120 1118.010 790.380 1118.330 ;
        RECT 790.120 1116.360 790.260 1118.010 ;
        RECT 790.040 1115.510 790.360 1116.360 ;
    END
  END mgmt_io_oeb_buf[37]
  PIN mgmt_io_oeb_unbuf[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2093.340 1115.850 2094.930 1116.050 ;
      LAYER mcon ;
        RECT 2093.840 1115.850 2094.930 1116.020 ;
      LAYER met1 ;
        RECT 2094.305 1118.320 3357.540 1118.460 ;
        RECT 2094.305 1118.200 2094.625 1118.320 ;
        RECT 2093.780 1115.810 2094.990 1116.070 ;
        RECT 3357.400 1115.250 3357.540 1118.320 ;
      LAYER via ;
        RECT 2094.335 1118.200 2094.595 1118.460 ;
        RECT 2093.840 1115.810 2094.930 1116.070 ;
      LAYER met2 ;
        RECT 2094.335 1118.490 2094.475 1129.765 ;
        RECT 2094.335 1118.170 2094.595 1118.490 ;
        RECT 2094.335 1116.100 2094.475 1118.170 ;
        RECT 2093.840 1115.780 2094.930 1116.100 ;
    END
  END mgmt_io_oeb_unbuf[37]
  PIN mgmt_io_oeb_unbuf[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2093.340 1112.760 2094.440 1112.960 ;
      LAYER mcon ;
        RECT 2093.340 1112.790 2094.430 1112.960 ;
      LAYER met1 ;
        RECT 2093.335 1118.600 3357.820 1118.740 ;
        RECT 2093.335 1118.480 2093.655 1118.600 ;
        RECT 3357.680 1114.250 3357.820 1118.600 ;
        RECT 2093.280 1112.750 2094.490 1113.010 ;
      LAYER via ;
        RECT 2093.365 1118.480 2093.625 1118.740 ;
        RECT 2093.340 1112.750 2094.430 1113.010 ;
      LAYER met2 ;
        RECT 2093.365 1118.770 2093.505 1129.765 ;
        RECT 2093.365 1118.450 2093.625 1118.770 ;
        RECT 2093.365 1114.170 2093.505 1118.450 ;
        RECT 2093.365 1114.030 2094.140 1114.170 ;
        RECT 2094.000 1113.040 2094.140 1114.030 ;
        RECT 2093.340 1112.720 2094.430 1113.040 ;
    END
  END mgmt_io_oeb_unbuf[36]
  PIN mgmt_io_oeb_unbuf[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2087.360 1115.850 2088.950 1116.050 ;
      LAYER mcon ;
        RECT 2087.860 1115.850 2088.950 1116.020 ;
      LAYER met1 ;
        RECT 2088.205 1118.880 3358.100 1119.020 ;
        RECT 2088.205 1118.760 2088.525 1118.880 ;
        RECT 2087.800 1115.810 2089.010 1116.070 ;
        RECT 3357.960 1113.250 3358.100 1118.880 ;
      LAYER via ;
        RECT 2088.235 1118.760 2088.495 1119.020 ;
        RECT 2087.860 1115.810 2088.950 1116.070 ;
      LAYER met2 ;
        RECT 2088.355 1119.050 2088.495 1129.765 ;
        RECT 2088.235 1118.730 2088.495 1119.050 ;
        RECT 2088.355 1116.100 2088.495 1118.730 ;
        RECT 2087.860 1115.780 2088.950 1116.100 ;
    END
  END mgmt_io_oeb_unbuf[35]
  PIN mgmt_io_in_buf[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2084.935 1113.300 2085.105 1114.150 ;
        RECT 2085.775 1113.300 2085.945 1114.150 ;
        RECT 2086.615 1113.300 2086.785 1114.150 ;
        RECT 2087.455 1113.300 2087.625 1114.150 ;
        RECT 2084.935 1113.130 2087.625 1113.300 ;
        RECT 2087.370 1112.590 2087.625 1113.130 ;
        RECT 2084.935 1112.420 2087.625 1112.590 ;
        RECT 2084.935 1111.940 2085.105 1112.420 ;
        RECT 2085.775 1111.940 2085.945 1112.420 ;
        RECT 2086.615 1111.940 2086.785 1112.420 ;
        RECT 2087.455 1111.940 2087.625 1112.420 ;
      LAYER mcon ;
        RECT 2087.370 1112.450 2087.540 1113.300 ;
      LAYER met1 ;
        RECT 2087.355 1119.160 3358.380 1119.300 ;
        RECT 2087.355 1119.040 2087.675 1119.160 ;
        RECT 2087.320 1112.390 2087.580 1113.360 ;
        RECT 3358.240 1112.250 3358.380 1119.160 ;
      LAYER via ;
        RECT 2087.385 1119.040 2087.645 1119.300 ;
        RECT 2087.320 1112.450 2087.580 1113.300 ;
      LAYER met2 ;
        RECT 2087.385 1119.330 2087.525 1129.765 ;
        RECT 2087.385 1119.010 2087.645 1119.330 ;
        RECT 2087.385 1113.300 2087.525 1119.010 ;
        RECT 2087.290 1112.450 2087.610 1113.300 ;
    END
  END mgmt_io_in_buf[37]
  PIN mgmt_io_in_buf[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2078.955 1113.300 2079.125 1114.150 ;
        RECT 2079.795 1113.300 2079.965 1114.150 ;
        RECT 2080.635 1113.300 2080.805 1114.150 ;
        RECT 2081.475 1113.300 2081.645 1114.150 ;
        RECT 2078.955 1113.130 2081.645 1113.300 ;
        RECT 2081.390 1112.590 2081.645 1113.130 ;
        RECT 2078.955 1112.420 2081.645 1112.590 ;
        RECT 2078.955 1111.940 2079.125 1112.420 ;
        RECT 2079.795 1111.940 2079.965 1112.420 ;
        RECT 2080.635 1111.940 2080.805 1112.420 ;
        RECT 2081.475 1111.940 2081.645 1112.420 ;
      LAYER mcon ;
        RECT 2081.390 1112.450 2081.560 1113.300 ;
      LAYER met1 ;
        RECT 2081.375 1119.720 3358.940 1119.860 ;
        RECT 2081.375 1119.600 2081.695 1119.720 ;
        RECT 2081.340 1112.390 2081.600 1113.360 ;
        RECT 3358.800 1110.250 3358.940 1119.720 ;
      LAYER via ;
        RECT 2081.405 1119.600 2081.665 1119.860 ;
        RECT 2081.340 1112.450 2081.600 1113.300 ;
      LAYER met2 ;
        RECT 2081.405 1119.890 2081.545 1129.765 ;
        RECT 2081.405 1119.570 2081.665 1119.890 ;
        RECT 2081.405 1113.300 2081.545 1119.570 ;
        RECT 2081.310 1112.450 2081.630 1113.300 ;
    END
  END mgmt_io_in_buf[36]
  PIN mgmt_io_in_buf[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2072.975 1113.300 2073.145 1114.150 ;
        RECT 2073.815 1113.300 2073.985 1114.150 ;
        RECT 2074.655 1113.300 2074.825 1114.150 ;
        RECT 2075.495 1113.300 2075.665 1114.150 ;
        RECT 2072.975 1113.130 2075.665 1113.300 ;
        RECT 2075.410 1112.590 2075.665 1113.130 ;
        RECT 2072.975 1112.420 2075.665 1112.590 ;
        RECT 2072.975 1111.940 2073.145 1112.420 ;
        RECT 2073.815 1111.940 2073.985 1112.420 ;
        RECT 2074.655 1111.940 2074.825 1112.420 ;
        RECT 2075.495 1111.940 2075.665 1112.420 ;
      LAYER mcon ;
        RECT 2075.410 1112.450 2075.580 1113.300 ;
      LAYER met1 ;
        RECT 2075.395 1120.280 3359.500 1120.420 ;
        RECT 2075.395 1120.160 2075.715 1120.280 ;
        RECT 2075.360 1112.390 2075.620 1113.360 ;
        RECT 3359.360 1108.250 3359.500 1120.280 ;
      LAYER via ;
        RECT 2075.425 1120.160 2075.685 1120.420 ;
        RECT 2075.360 1112.450 2075.620 1113.300 ;
      LAYER met2 ;
        RECT 2075.425 1120.450 2075.565 1129.765 ;
        RECT 2075.425 1120.130 2075.685 1120.450 ;
        RECT 2075.425 1113.300 2075.565 1120.130 ;
        RECT 2075.330 1112.450 2075.650 1113.300 ;
    END
  END mgmt_io_in_buf[35]
  PIN mgmt_io_in_buf[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2066.995 1113.300 2067.165 1114.150 ;
        RECT 2067.835 1113.300 2068.005 1114.150 ;
        RECT 2068.675 1113.300 2068.845 1114.150 ;
        RECT 2069.515 1113.300 2069.685 1114.150 ;
        RECT 2066.995 1113.130 2069.685 1113.300 ;
        RECT 2069.430 1112.590 2069.685 1113.130 ;
        RECT 2066.995 1112.420 2069.685 1112.590 ;
        RECT 2066.995 1111.940 2067.165 1112.420 ;
        RECT 2067.835 1111.940 2068.005 1112.420 ;
        RECT 2068.675 1111.940 2068.845 1112.420 ;
        RECT 2069.515 1111.940 2069.685 1112.420 ;
      LAYER mcon ;
        RECT 2069.430 1112.450 2069.600 1113.300 ;
      LAYER met1 ;
        RECT 2069.415 1120.840 3360.060 1120.980 ;
        RECT 2069.415 1120.720 2069.735 1120.840 ;
        RECT 2069.380 1112.390 2069.640 1113.360 ;
        RECT 3359.920 1106.250 3360.060 1120.840 ;
      LAYER via ;
        RECT 2069.445 1120.720 2069.705 1120.980 ;
        RECT 2069.380 1112.450 2069.640 1113.300 ;
      LAYER met2 ;
        RECT 2069.445 1121.010 2069.585 1129.765 ;
        RECT 2069.445 1120.690 2069.705 1121.010 ;
        RECT 2069.445 1113.300 2069.585 1120.690 ;
        RECT 2069.350 1112.450 2069.670 1113.300 ;
    END
  END mgmt_io_in_buf[34]
  PIN mgmt_io_out_unbuf[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2063.440 1115.850 2065.030 1116.050 ;
      LAYER mcon ;
        RECT 2063.940 1115.850 2065.030 1116.020 ;
      LAYER met1 ;
        RECT 2064.405 1121.120 3360.340 1121.260 ;
        RECT 2064.405 1121.000 2064.725 1121.120 ;
        RECT 2063.880 1115.810 2065.090 1116.070 ;
        RECT 3360.200 1105.250 3360.340 1121.120 ;
      LAYER via ;
        RECT 2064.435 1121.000 2064.695 1121.260 ;
        RECT 2063.940 1115.810 2065.030 1116.070 ;
      LAYER met2 ;
        RECT 2064.435 1121.290 2064.575 1129.765 ;
        RECT 2064.435 1120.970 2064.695 1121.290 ;
        RECT 2064.435 1116.100 2064.575 1120.970 ;
        RECT 2063.940 1115.780 2065.030 1116.100 ;
    END
  END mgmt_io_out_unbuf[34]
  PIN mgmt_io_out_unbuf[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2069.420 1115.850 2071.010 1116.050 ;
      LAYER mcon ;
        RECT 2069.920 1115.850 2071.010 1116.020 ;
      LAYER met1 ;
        RECT 2070.385 1120.560 3359.780 1120.700 ;
        RECT 2070.385 1120.440 2070.705 1120.560 ;
        RECT 2069.860 1115.810 2071.070 1116.070 ;
        RECT 3359.640 1107.250 3359.780 1120.560 ;
      LAYER via ;
        RECT 2070.415 1120.440 2070.675 1120.700 ;
        RECT 2069.920 1115.810 2071.010 1116.070 ;
      LAYER met2 ;
        RECT 2070.415 1120.730 2070.555 1129.765 ;
        RECT 2070.415 1120.410 2070.675 1120.730 ;
        RECT 2070.415 1116.100 2070.555 1120.410 ;
        RECT 2069.920 1115.780 2071.010 1116.100 ;
    END
  END mgmt_io_out_unbuf[35]
  PIN mgmt_io_out_unbuf[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2075.400 1115.850 2076.990 1116.050 ;
      LAYER mcon ;
        RECT 2075.900 1115.850 2076.990 1116.020 ;
      LAYER met1 ;
        RECT 2076.245 1120.000 3359.220 1120.140 ;
        RECT 2076.245 1119.880 2076.565 1120.000 ;
        RECT 2075.840 1115.810 2077.050 1116.070 ;
        RECT 3359.080 1109.250 3359.220 1120.000 ;
      LAYER via ;
        RECT 2076.275 1119.880 2076.535 1120.140 ;
        RECT 2075.900 1115.810 2076.990 1116.070 ;
      LAYER met2 ;
        RECT 2076.395 1120.170 2076.535 1129.765 ;
        RECT 2076.275 1119.850 2076.535 1120.170 ;
        RECT 2076.395 1116.100 2076.535 1119.850 ;
        RECT 2075.900 1115.780 2076.990 1116.100 ;
    END
  END mgmt_io_out_unbuf[36]
  PIN mgmt_io_out_unbuf[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2081.380 1115.850 2082.970 1116.050 ;
      LAYER mcon ;
        RECT 2081.880 1115.850 2082.970 1116.020 ;
      LAYER met1 ;
        RECT 2082.345 1119.440 3358.660 1119.580 ;
        RECT 2082.345 1119.320 2082.665 1119.440 ;
        RECT 2081.820 1115.810 2083.030 1116.070 ;
        RECT 3358.520 1111.250 3358.660 1119.440 ;
      LAYER via ;
        RECT 2082.375 1119.320 2082.635 1119.580 ;
        RECT 2081.880 1115.810 2082.970 1116.070 ;
      LAYER met2 ;
        RECT 2082.375 1119.610 2082.515 1129.765 ;
        RECT 2082.375 1119.290 2082.635 1119.610 ;
        RECT 2082.375 1116.100 2082.515 1119.290 ;
        RECT 2081.880 1115.780 2082.970 1116.100 ;
    END
  END mgmt_io_out_unbuf[37]
  PIN mgmt_io_out_unbuf[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1973.740 1115.850 1975.330 1116.050 ;
      LAYER mcon ;
        RECT 1974.240 1115.850 1975.330 1116.020 ;
      LAYER met1 ;
        RECT 1974.705 1129.520 3368.740 1129.660 ;
        RECT 1974.705 1129.400 1975.025 1129.520 ;
        RECT 1974.180 1115.810 1975.390 1116.070 ;
        RECT 3368.600 1075.250 3368.740 1129.520 ;
      LAYER via ;
        RECT 1974.735 1129.400 1974.995 1129.660 ;
        RECT 1974.240 1115.810 1975.330 1116.070 ;
      LAYER met2 ;
        RECT 1974.735 1129.690 1974.875 1129.765 ;
        RECT 1974.735 1129.370 1974.995 1129.690 ;
        RECT 1974.735 1116.100 1974.875 1129.370 ;
        RECT 1974.240 1115.780 1975.330 1116.100 ;
    END
  END mgmt_io_out_unbuf[33]
  PIN mgmt_io_out_unbuf[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1979.720 1115.850 1981.310 1116.050 ;
      LAYER mcon ;
        RECT 1980.220 1115.850 1981.310 1116.020 ;
      LAYER met1 ;
        RECT 1980.685 1128.960 3368.180 1129.100 ;
        RECT 1980.685 1128.840 1981.005 1128.960 ;
        RECT 1980.160 1115.810 1981.370 1116.070 ;
        RECT 3368.040 1077.250 3368.180 1128.960 ;
      LAYER via ;
        RECT 1980.715 1128.840 1980.975 1129.100 ;
        RECT 1980.220 1115.810 1981.310 1116.070 ;
      LAYER met2 ;
        RECT 1980.715 1129.130 1980.855 1129.765 ;
        RECT 1980.715 1128.810 1980.975 1129.130 ;
        RECT 1980.715 1116.100 1980.855 1128.810 ;
        RECT 1980.220 1115.780 1981.310 1116.100 ;
    END
  END mgmt_io_out_unbuf[32]
  PIN mgmt_io_out_unbuf[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1985.700 1115.850 1987.290 1116.050 ;
      LAYER mcon ;
        RECT 1986.200 1115.850 1987.290 1116.020 ;
      LAYER met1 ;
        RECT 1986.665 1128.400 3367.620 1128.540 ;
        RECT 1986.665 1128.280 1986.985 1128.400 ;
        RECT 1986.140 1115.810 1987.350 1116.070 ;
        RECT 3367.480 1079.250 3367.620 1128.400 ;
      LAYER via ;
        RECT 1986.695 1128.280 1986.955 1128.540 ;
        RECT 1986.200 1115.810 1987.290 1116.070 ;
      LAYER met2 ;
        RECT 1986.695 1128.570 1986.835 1129.765 ;
        RECT 1986.695 1128.250 1986.955 1128.570 ;
        RECT 1986.695 1116.100 1986.835 1128.250 ;
        RECT 1986.200 1115.780 1987.290 1116.100 ;
    END
  END mgmt_io_out_unbuf[31]
  PIN mgmt_io_out_unbuf[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1991.680 1115.850 1993.270 1116.050 ;
      LAYER mcon ;
        RECT 1992.180 1115.850 1993.270 1116.020 ;
      LAYER met1 ;
        RECT 1992.645 1127.840 3367.060 1127.980 ;
        RECT 1992.645 1127.720 1992.965 1127.840 ;
        RECT 1992.120 1115.810 1993.330 1116.070 ;
        RECT 3366.920 1081.250 3367.060 1127.840 ;
      LAYER via ;
        RECT 1992.675 1127.720 1992.935 1127.980 ;
        RECT 1992.180 1115.810 1993.270 1116.070 ;
      LAYER met2 ;
        RECT 1992.675 1128.010 1992.815 1129.765 ;
        RECT 1992.675 1127.690 1992.935 1128.010 ;
        RECT 1992.675 1116.100 1992.815 1127.690 ;
        RECT 1992.180 1115.780 1993.270 1116.100 ;
    END
  END mgmt_io_out_unbuf[30]
  PIN mgmt_io_out_unbuf[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1997.660 1115.850 1999.250 1116.050 ;
      LAYER mcon ;
        RECT 1998.160 1115.850 1999.250 1116.020 ;
      LAYER met1 ;
        RECT 1998.625 1127.280 3366.500 1127.420 ;
        RECT 1998.625 1127.160 1998.945 1127.280 ;
        RECT 1998.100 1115.810 1999.310 1116.070 ;
        RECT 3366.360 1083.250 3366.500 1127.280 ;
      LAYER via ;
        RECT 1998.655 1127.160 1998.915 1127.420 ;
        RECT 1998.160 1115.810 1999.250 1116.070 ;
      LAYER met2 ;
        RECT 1998.655 1127.450 1998.795 1129.765 ;
        RECT 1998.655 1127.130 1998.915 1127.450 ;
        RECT 1998.655 1116.100 1998.795 1127.130 ;
        RECT 1998.160 1115.780 1999.250 1116.100 ;
    END
  END mgmt_io_out_unbuf[29]
  PIN mgmt_io_out_unbuf[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2003.640 1115.850 2005.230 1116.050 ;
      LAYER mcon ;
        RECT 2004.140 1115.850 2005.230 1116.020 ;
      LAYER met1 ;
        RECT 2004.485 1126.720 3365.940 1126.860 ;
        RECT 2004.485 1126.600 2004.805 1126.720 ;
        RECT 2004.080 1115.810 2005.290 1116.070 ;
        RECT 3365.800 1085.250 3365.940 1126.720 ;
      LAYER via ;
        RECT 2004.515 1126.600 2004.775 1126.860 ;
        RECT 2004.140 1115.810 2005.230 1116.070 ;
      LAYER met2 ;
        RECT 2004.635 1126.890 2004.775 1129.765 ;
        RECT 2004.515 1126.570 2004.775 1126.890 ;
        RECT 2004.635 1116.100 2004.775 1126.570 ;
        RECT 2004.140 1115.780 2005.230 1116.100 ;
    END
  END mgmt_io_out_unbuf[28]
  PIN mgmt_io_out_unbuf[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2009.620 1115.850 2011.210 1116.050 ;
      LAYER mcon ;
        RECT 2010.120 1115.850 2011.210 1116.020 ;
      LAYER met1 ;
        RECT 2010.585 1126.160 3365.380 1126.300 ;
        RECT 2010.585 1126.040 2010.905 1126.160 ;
        RECT 2010.060 1115.810 2011.270 1116.070 ;
        RECT 3365.240 1087.250 3365.380 1126.160 ;
      LAYER via ;
        RECT 2010.615 1126.040 2010.875 1126.300 ;
        RECT 2010.120 1115.810 2011.210 1116.070 ;
      LAYER met2 ;
        RECT 2010.615 1126.330 2010.755 1129.765 ;
        RECT 2010.615 1126.010 2010.875 1126.330 ;
        RECT 2010.615 1116.100 2010.755 1126.010 ;
        RECT 2010.120 1115.780 2011.210 1116.100 ;
    END
  END mgmt_io_out_unbuf[27]
  PIN mgmt_io_out_unbuf[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2015.600 1115.850 2017.190 1116.050 ;
      LAYER mcon ;
        RECT 2016.100 1115.850 2017.190 1116.020 ;
      LAYER met1 ;
        RECT 2016.445 1125.600 3364.820 1125.740 ;
        RECT 2016.445 1125.480 2016.765 1125.600 ;
        RECT 2016.040 1115.810 2017.250 1116.070 ;
        RECT 3364.680 1089.250 3364.820 1125.600 ;
      LAYER via ;
        RECT 2016.475 1125.480 2016.735 1125.740 ;
        RECT 2016.100 1115.810 2017.190 1116.070 ;
      LAYER met2 ;
        RECT 2016.595 1125.770 2016.735 1129.765 ;
        RECT 2016.475 1125.450 2016.735 1125.770 ;
        RECT 2016.595 1116.100 2016.735 1125.450 ;
        RECT 2016.100 1115.780 2017.190 1116.100 ;
    END
  END mgmt_io_out_unbuf[26]
  PIN mgmt_io_out_unbuf[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2021.580 1115.850 2023.170 1116.050 ;
      LAYER mcon ;
        RECT 2022.080 1115.850 2023.170 1116.020 ;
      LAYER met1 ;
        RECT 2022.545 1125.040 3364.260 1125.180 ;
        RECT 2022.545 1124.920 2022.865 1125.040 ;
        RECT 2022.020 1115.810 2023.230 1116.070 ;
        RECT 3364.120 1091.250 3364.260 1125.040 ;
      LAYER via ;
        RECT 2022.575 1124.920 2022.835 1125.180 ;
        RECT 2022.080 1115.810 2023.170 1116.070 ;
      LAYER met2 ;
        RECT 2022.575 1125.210 2022.715 1129.765 ;
        RECT 2022.575 1124.890 2022.835 1125.210 ;
        RECT 2022.575 1116.100 2022.715 1124.890 ;
        RECT 2022.080 1115.780 2023.170 1116.100 ;
    END
  END mgmt_io_out_unbuf[25]
  PIN mgmt_io_out_unbuf[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2027.560 1115.850 2029.150 1116.050 ;
      LAYER mcon ;
        RECT 2028.060 1115.850 2029.150 1116.020 ;
      LAYER met1 ;
        RECT 2028.525 1124.480 3363.700 1124.620 ;
        RECT 2028.525 1124.360 2028.845 1124.480 ;
        RECT 2028.000 1115.810 2029.210 1116.070 ;
        RECT 3363.560 1093.250 3363.700 1124.480 ;
      LAYER via ;
        RECT 2028.555 1124.360 2028.815 1124.620 ;
        RECT 2028.060 1115.810 2029.150 1116.070 ;
      LAYER met2 ;
        RECT 2028.555 1124.650 2028.695 1129.765 ;
        RECT 2028.555 1124.330 2028.815 1124.650 ;
        RECT 2028.555 1116.100 2028.695 1124.330 ;
        RECT 2028.060 1115.780 2029.150 1116.100 ;
    END
  END mgmt_io_out_unbuf[24]
  PIN mgmt_io_out_unbuf[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2033.540 1115.850 2035.130 1116.050 ;
      LAYER mcon ;
        RECT 2034.040 1115.850 2035.130 1116.020 ;
      LAYER met1 ;
        RECT 2034.505 1123.920 3363.140 1124.060 ;
        RECT 2034.505 1123.800 2034.825 1123.920 ;
        RECT 2033.980 1115.810 2035.190 1116.070 ;
        RECT 3363.000 1095.250 3363.140 1123.920 ;
      LAYER via ;
        RECT 2034.535 1123.800 2034.795 1124.060 ;
        RECT 2034.040 1115.810 2035.130 1116.070 ;
      LAYER met2 ;
        RECT 2034.535 1124.090 2034.675 1129.765 ;
        RECT 2034.535 1123.770 2034.795 1124.090 ;
        RECT 2034.535 1116.100 2034.675 1123.770 ;
        RECT 2034.040 1115.780 2035.130 1116.100 ;
    END
  END mgmt_io_out_unbuf[23]
  PIN mgmt_io_out_unbuf[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2039.520 1115.850 2041.110 1116.050 ;
      LAYER mcon ;
        RECT 2040.020 1115.850 2041.110 1116.020 ;
      LAYER met1 ;
        RECT 2040.485 1123.360 3362.580 1123.500 ;
        RECT 2040.485 1123.240 2040.805 1123.360 ;
        RECT 2039.960 1115.810 2041.170 1116.070 ;
        RECT 3362.440 1097.250 3362.580 1123.360 ;
      LAYER via ;
        RECT 2040.515 1123.240 2040.775 1123.500 ;
        RECT 2040.020 1115.810 2041.110 1116.070 ;
      LAYER met2 ;
        RECT 2040.515 1123.530 2040.655 1129.765 ;
        RECT 2040.515 1123.210 2040.775 1123.530 ;
        RECT 2040.515 1116.100 2040.655 1123.210 ;
        RECT 2040.020 1115.780 2041.110 1116.100 ;
    END
  END mgmt_io_out_unbuf[22]
  PIN mgmt_io_out_unbuf[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2045.500 1115.850 2047.090 1116.050 ;
      LAYER mcon ;
        RECT 2046.000 1115.850 2047.090 1116.020 ;
      LAYER met1 ;
        RECT 2046.465 1122.800 3362.020 1122.940 ;
        RECT 2046.465 1122.680 2046.785 1122.800 ;
        RECT 2045.940 1115.810 2047.150 1116.070 ;
        RECT 3361.880 1099.250 3362.020 1122.800 ;
      LAYER via ;
        RECT 2046.495 1122.680 2046.755 1122.940 ;
        RECT 2046.000 1115.810 2047.090 1116.070 ;
      LAYER met2 ;
        RECT 2046.495 1122.970 2046.635 1129.765 ;
        RECT 2046.495 1122.650 2046.755 1122.970 ;
        RECT 2046.495 1116.100 2046.635 1122.650 ;
        RECT 2046.000 1115.780 2047.090 1116.100 ;
    END
  END mgmt_io_out_unbuf[21]
  PIN mgmt_io_out_unbuf[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2051.480 1115.850 2053.070 1116.050 ;
      LAYER mcon ;
        RECT 2051.980 1115.850 2053.070 1116.020 ;
      LAYER met1 ;
        RECT 2052.445 1122.240 3361.460 1122.380 ;
        RECT 2052.445 1122.120 2052.765 1122.240 ;
        RECT 2051.920 1115.810 2053.130 1116.070 ;
        RECT 3361.320 1101.250 3361.460 1122.240 ;
      LAYER via ;
        RECT 2052.475 1122.120 2052.735 1122.380 ;
        RECT 2051.980 1115.810 2053.070 1116.070 ;
      LAYER met2 ;
        RECT 2052.475 1122.410 2052.615 1129.765 ;
        RECT 2052.475 1122.090 2052.735 1122.410 ;
        RECT 2052.475 1116.100 2052.615 1122.090 ;
        RECT 2051.980 1115.780 2053.070 1116.100 ;
    END
  END mgmt_io_out_unbuf[20]
  PIN mgmt_io_out_unbuf[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2057.460 1115.850 2059.050 1116.050 ;
      LAYER mcon ;
        RECT 2057.960 1115.850 2059.050 1116.020 ;
      LAYER met1 ;
        RECT 2058.425 1121.680 3360.900 1121.820 ;
        RECT 2058.425 1121.560 2058.745 1121.680 ;
        RECT 2057.900 1115.810 2059.110 1116.070 ;
        RECT 3360.760 1103.250 3360.900 1121.680 ;
      LAYER via ;
        RECT 2058.455 1121.560 2058.715 1121.820 ;
        RECT 2057.960 1115.810 2059.050 1116.070 ;
      LAYER met2 ;
        RECT 2058.455 1121.850 2058.595 1129.765 ;
        RECT 2058.455 1121.530 2058.715 1121.850 ;
        RECT 2058.455 1116.100 2058.595 1121.530 ;
        RECT 2057.960 1115.780 2059.050 1116.100 ;
    END
  END mgmt_io_out_unbuf[19]
  PIN mgmt_io_in_buf[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2061.015 1113.300 2061.185 1114.150 ;
        RECT 2061.855 1113.300 2062.025 1114.150 ;
        RECT 2062.695 1113.300 2062.865 1114.150 ;
        RECT 2063.535 1113.300 2063.705 1114.150 ;
        RECT 2061.015 1113.130 2063.705 1113.300 ;
        RECT 2063.450 1112.590 2063.705 1113.130 ;
        RECT 2061.015 1112.420 2063.705 1112.590 ;
        RECT 2061.015 1111.940 2061.185 1112.420 ;
        RECT 2061.855 1111.940 2062.025 1112.420 ;
        RECT 2062.695 1111.940 2062.865 1112.420 ;
        RECT 2063.535 1111.940 2063.705 1112.420 ;
      LAYER mcon ;
        RECT 2063.450 1112.450 2063.620 1113.300 ;
      LAYER met1 ;
        RECT 2063.435 1121.400 3360.620 1121.540 ;
        RECT 2063.435 1121.280 2063.755 1121.400 ;
        RECT 2063.400 1112.390 2063.660 1113.360 ;
        RECT 3360.480 1104.250 3360.620 1121.400 ;
      LAYER via ;
        RECT 2063.465 1121.280 2063.725 1121.540 ;
        RECT 2063.400 1112.450 2063.660 1113.300 ;
      LAYER met2 ;
        RECT 2063.465 1121.570 2063.605 1129.765 ;
        RECT 2063.465 1121.250 2063.725 1121.570 ;
        RECT 2063.465 1113.300 2063.605 1121.250 ;
        RECT 2063.370 1112.450 2063.690 1113.300 ;
    END
  END mgmt_io_in_buf[19]
  PIN mgmt_io_in_buf[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2055.035 1113.300 2055.205 1114.150 ;
        RECT 2055.875 1113.300 2056.045 1114.150 ;
        RECT 2056.715 1113.300 2056.885 1114.150 ;
        RECT 2057.555 1113.300 2057.725 1114.150 ;
        RECT 2055.035 1113.130 2057.725 1113.300 ;
        RECT 2057.470 1112.590 2057.725 1113.130 ;
        RECT 2055.035 1112.420 2057.725 1112.590 ;
        RECT 2055.035 1111.940 2055.205 1112.420 ;
        RECT 2055.875 1111.940 2056.045 1112.420 ;
        RECT 2056.715 1111.940 2056.885 1112.420 ;
        RECT 2057.555 1111.940 2057.725 1112.420 ;
      LAYER mcon ;
        RECT 2057.470 1112.450 2057.640 1113.300 ;
      LAYER met1 ;
        RECT 2057.455 1121.960 3361.180 1122.100 ;
        RECT 2057.455 1121.840 2057.775 1121.960 ;
        RECT 2057.420 1112.390 2057.680 1113.360 ;
        RECT 3361.040 1102.250 3361.180 1121.960 ;
      LAYER via ;
        RECT 2057.485 1121.840 2057.745 1122.100 ;
        RECT 2057.420 1112.450 2057.680 1113.300 ;
      LAYER met2 ;
        RECT 2057.485 1122.130 2057.625 1129.765 ;
        RECT 2057.485 1121.810 2057.745 1122.130 ;
        RECT 2057.485 1113.300 2057.625 1121.810 ;
        RECT 2057.390 1112.450 2057.710 1113.300 ;
    END
  END mgmt_io_in_buf[20]
  PIN mgmt_io_in_buf[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2049.055 1113.300 2049.225 1114.150 ;
        RECT 2049.895 1113.300 2050.065 1114.150 ;
        RECT 2050.735 1113.300 2050.905 1114.150 ;
        RECT 2051.575 1113.300 2051.745 1114.150 ;
        RECT 2049.055 1113.130 2051.745 1113.300 ;
        RECT 2051.490 1112.590 2051.745 1113.130 ;
        RECT 2049.055 1112.420 2051.745 1112.590 ;
        RECT 2049.055 1111.940 2049.225 1112.420 ;
        RECT 2049.895 1111.940 2050.065 1112.420 ;
        RECT 2050.735 1111.940 2050.905 1112.420 ;
        RECT 2051.575 1111.940 2051.745 1112.420 ;
      LAYER mcon ;
        RECT 2051.490 1112.450 2051.660 1113.300 ;
      LAYER met1 ;
        RECT 2051.475 1122.520 3361.740 1122.660 ;
        RECT 2051.475 1122.400 2051.795 1122.520 ;
        RECT 2051.440 1112.390 2051.700 1113.360 ;
        RECT 3361.600 1100.250 3361.740 1122.520 ;
      LAYER via ;
        RECT 2051.505 1122.400 2051.765 1122.660 ;
        RECT 2051.440 1112.450 2051.700 1113.300 ;
      LAYER met2 ;
        RECT 2051.505 1122.690 2051.645 1129.765 ;
        RECT 2051.505 1122.370 2051.765 1122.690 ;
        RECT 2051.505 1113.300 2051.645 1122.370 ;
        RECT 2051.410 1112.450 2051.730 1113.300 ;
    END
  END mgmt_io_in_buf[21]
  PIN mgmt_io_in_buf[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2043.075 1113.300 2043.245 1114.150 ;
        RECT 2043.915 1113.300 2044.085 1114.150 ;
        RECT 2044.755 1113.300 2044.925 1114.150 ;
        RECT 2045.595 1113.300 2045.765 1114.150 ;
        RECT 2043.075 1113.130 2045.765 1113.300 ;
        RECT 2045.510 1112.590 2045.765 1113.130 ;
        RECT 2043.075 1112.420 2045.765 1112.590 ;
        RECT 2043.075 1111.940 2043.245 1112.420 ;
        RECT 2043.915 1111.940 2044.085 1112.420 ;
        RECT 2044.755 1111.940 2044.925 1112.420 ;
        RECT 2045.595 1111.940 2045.765 1112.420 ;
      LAYER mcon ;
        RECT 2045.510 1112.450 2045.680 1113.300 ;
      LAYER met1 ;
        RECT 2045.495 1123.080 3362.300 1123.220 ;
        RECT 2045.495 1122.960 2045.815 1123.080 ;
        RECT 2045.460 1112.390 2045.720 1113.360 ;
        RECT 3362.160 1098.250 3362.300 1123.080 ;
      LAYER via ;
        RECT 2045.525 1122.960 2045.785 1123.220 ;
        RECT 2045.460 1112.450 2045.720 1113.300 ;
      LAYER met2 ;
        RECT 2045.525 1123.250 2045.665 1129.765 ;
        RECT 2045.525 1122.930 2045.785 1123.250 ;
        RECT 2045.525 1113.300 2045.665 1122.930 ;
        RECT 2045.430 1112.450 2045.750 1113.300 ;
    END
  END mgmt_io_in_buf[22]
  PIN mgmt_io_in_buf[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2037.095 1113.300 2037.265 1114.150 ;
        RECT 2037.935 1113.300 2038.105 1114.150 ;
        RECT 2038.775 1113.300 2038.945 1114.150 ;
        RECT 2039.615 1113.300 2039.785 1114.150 ;
        RECT 2037.095 1113.130 2039.785 1113.300 ;
        RECT 2039.530 1112.590 2039.785 1113.130 ;
        RECT 2037.095 1112.420 2039.785 1112.590 ;
        RECT 2037.095 1111.940 2037.265 1112.420 ;
        RECT 2037.935 1111.940 2038.105 1112.420 ;
        RECT 2038.775 1111.940 2038.945 1112.420 ;
        RECT 2039.615 1111.940 2039.785 1112.420 ;
      LAYER mcon ;
        RECT 2039.530 1112.450 2039.700 1113.300 ;
      LAYER met1 ;
        RECT 2039.515 1123.640 3362.860 1123.780 ;
        RECT 2039.515 1123.520 2039.835 1123.640 ;
        RECT 2039.480 1112.390 2039.740 1113.360 ;
        RECT 3362.720 1096.250 3362.860 1123.640 ;
      LAYER via ;
        RECT 2039.545 1123.520 2039.805 1123.780 ;
        RECT 2039.480 1112.450 2039.740 1113.300 ;
      LAYER met2 ;
        RECT 2039.545 1123.810 2039.685 1129.765 ;
        RECT 2039.545 1123.490 2039.805 1123.810 ;
        RECT 2039.545 1113.300 2039.685 1123.490 ;
        RECT 2039.450 1112.450 2039.770 1113.300 ;
    END
  END mgmt_io_in_buf[23]
  PIN mgmt_io_in_buf[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2031.115 1113.300 2031.285 1114.150 ;
        RECT 2031.955 1113.300 2032.125 1114.150 ;
        RECT 2032.795 1113.300 2032.965 1114.150 ;
        RECT 2033.635 1113.300 2033.805 1114.150 ;
        RECT 2031.115 1113.130 2033.805 1113.300 ;
        RECT 2033.550 1112.590 2033.805 1113.130 ;
        RECT 2031.115 1112.420 2033.805 1112.590 ;
        RECT 2031.115 1111.940 2031.285 1112.420 ;
        RECT 2031.955 1111.940 2032.125 1112.420 ;
        RECT 2032.795 1111.940 2032.965 1112.420 ;
        RECT 2033.635 1111.940 2033.805 1112.420 ;
      LAYER mcon ;
        RECT 2033.550 1112.450 2033.720 1113.300 ;
      LAYER met1 ;
        RECT 2033.535 1124.200 3363.420 1124.340 ;
        RECT 2033.535 1124.080 2033.855 1124.200 ;
        RECT 2033.500 1112.390 2033.760 1113.360 ;
        RECT 3363.280 1094.250 3363.420 1124.200 ;
      LAYER via ;
        RECT 2033.565 1124.080 2033.825 1124.340 ;
        RECT 2033.500 1112.450 2033.760 1113.300 ;
      LAYER met2 ;
        RECT 2033.565 1124.370 2033.705 1129.765 ;
        RECT 2033.565 1124.050 2033.825 1124.370 ;
        RECT 2033.565 1113.300 2033.705 1124.050 ;
        RECT 2033.470 1112.450 2033.790 1113.300 ;
    END
  END mgmt_io_in_buf[24]
  PIN mgmt_io_in_buf[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2025.135 1113.300 2025.305 1114.150 ;
        RECT 2025.975 1113.300 2026.145 1114.150 ;
        RECT 2026.815 1113.300 2026.985 1114.150 ;
        RECT 2027.655 1113.300 2027.825 1114.150 ;
        RECT 2025.135 1113.130 2027.825 1113.300 ;
        RECT 2027.570 1112.590 2027.825 1113.130 ;
        RECT 2025.135 1112.420 2027.825 1112.590 ;
        RECT 2025.135 1111.940 2025.305 1112.420 ;
        RECT 2025.975 1111.940 2026.145 1112.420 ;
        RECT 2026.815 1111.940 2026.985 1112.420 ;
        RECT 2027.655 1111.940 2027.825 1112.420 ;
      LAYER mcon ;
        RECT 2027.570 1112.450 2027.740 1113.300 ;
      LAYER met1 ;
        RECT 2027.555 1124.760 3363.980 1124.900 ;
        RECT 2027.555 1124.640 2027.875 1124.760 ;
        RECT 2027.520 1112.390 2027.780 1113.360 ;
        RECT 3363.840 1092.250 3363.980 1124.760 ;
      LAYER via ;
        RECT 2027.585 1124.640 2027.845 1124.900 ;
        RECT 2027.520 1112.450 2027.780 1113.300 ;
      LAYER met2 ;
        RECT 2027.585 1124.930 2027.725 1129.765 ;
        RECT 2027.585 1124.610 2027.845 1124.930 ;
        RECT 2027.585 1113.300 2027.725 1124.610 ;
        RECT 2027.490 1112.450 2027.810 1113.300 ;
    END
  END mgmt_io_in_buf[25]
  PIN mgmt_io_in_buf[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2019.155 1113.300 2019.325 1114.150 ;
        RECT 2019.995 1113.300 2020.165 1114.150 ;
        RECT 2020.835 1113.300 2021.005 1114.150 ;
        RECT 2021.675 1113.300 2021.845 1114.150 ;
        RECT 2019.155 1113.130 2021.845 1113.300 ;
        RECT 2021.590 1112.590 2021.845 1113.130 ;
        RECT 2019.155 1112.420 2021.845 1112.590 ;
        RECT 2019.155 1111.940 2019.325 1112.420 ;
        RECT 2019.995 1111.940 2020.165 1112.420 ;
        RECT 2020.835 1111.940 2021.005 1112.420 ;
        RECT 2021.675 1111.940 2021.845 1112.420 ;
      LAYER mcon ;
        RECT 2021.590 1112.450 2021.760 1113.300 ;
      LAYER met1 ;
        RECT 2021.575 1125.320 3364.540 1125.460 ;
        RECT 2021.575 1125.200 2021.895 1125.320 ;
        RECT 2021.540 1112.390 2021.800 1113.360 ;
        RECT 3364.400 1090.250 3364.540 1125.320 ;
      LAYER via ;
        RECT 2021.605 1125.200 2021.865 1125.460 ;
        RECT 2021.540 1112.450 2021.800 1113.300 ;
      LAYER met2 ;
        RECT 2021.605 1125.490 2021.745 1129.765 ;
        RECT 2021.605 1125.170 2021.865 1125.490 ;
        RECT 2021.605 1113.300 2021.745 1125.170 ;
        RECT 2021.510 1112.450 2021.830 1113.300 ;
    END
  END mgmt_io_in_buf[26]
  PIN mgmt_io_in_buf[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2013.175 1113.300 2013.345 1114.150 ;
        RECT 2014.015 1113.300 2014.185 1114.150 ;
        RECT 2014.855 1113.300 2015.025 1114.150 ;
        RECT 2015.695 1113.300 2015.865 1114.150 ;
        RECT 2013.175 1113.130 2015.865 1113.300 ;
        RECT 2015.610 1112.590 2015.865 1113.130 ;
        RECT 2013.175 1112.420 2015.865 1112.590 ;
        RECT 2013.175 1111.940 2013.345 1112.420 ;
        RECT 2014.015 1111.940 2014.185 1112.420 ;
        RECT 2014.855 1111.940 2015.025 1112.420 ;
        RECT 2015.695 1111.940 2015.865 1112.420 ;
      LAYER mcon ;
        RECT 2015.610 1112.450 2015.780 1113.300 ;
      LAYER met1 ;
        RECT 2015.595 1125.880 3365.100 1126.020 ;
        RECT 2015.595 1125.760 2015.915 1125.880 ;
        RECT 2015.560 1112.390 2015.820 1113.360 ;
        RECT 3364.960 1088.250 3365.100 1125.880 ;
      LAYER via ;
        RECT 2015.625 1125.760 2015.885 1126.020 ;
        RECT 2015.560 1112.450 2015.820 1113.300 ;
      LAYER met2 ;
        RECT 2015.625 1126.050 2015.765 1129.765 ;
        RECT 2015.625 1125.730 2015.885 1126.050 ;
        RECT 2015.625 1113.300 2015.765 1125.730 ;
        RECT 2015.530 1112.450 2015.850 1113.300 ;
    END
  END mgmt_io_in_buf[27]
  PIN mgmt_io_in_buf[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2007.195 1113.300 2007.365 1114.150 ;
        RECT 2008.035 1113.300 2008.205 1114.150 ;
        RECT 2008.875 1113.300 2009.045 1114.150 ;
        RECT 2009.715 1113.300 2009.885 1114.150 ;
        RECT 2007.195 1113.130 2009.885 1113.300 ;
        RECT 2009.630 1112.590 2009.885 1113.130 ;
        RECT 2007.195 1112.420 2009.885 1112.590 ;
        RECT 2007.195 1111.940 2007.365 1112.420 ;
        RECT 2008.035 1111.940 2008.205 1112.420 ;
        RECT 2008.875 1111.940 2009.045 1112.420 ;
        RECT 2009.715 1111.940 2009.885 1112.420 ;
      LAYER mcon ;
        RECT 2009.630 1112.450 2009.800 1113.300 ;
      LAYER met1 ;
        RECT 2009.615 1126.440 3365.660 1126.580 ;
        RECT 2009.615 1126.320 2009.935 1126.440 ;
        RECT 2009.580 1112.390 2009.840 1113.360 ;
        RECT 3365.520 1086.250 3365.660 1126.440 ;
      LAYER via ;
        RECT 2009.645 1126.320 2009.905 1126.580 ;
        RECT 2009.580 1112.450 2009.840 1113.300 ;
      LAYER met2 ;
        RECT 2009.645 1126.610 2009.785 1129.765 ;
        RECT 2009.645 1126.290 2009.905 1126.610 ;
        RECT 2009.645 1113.300 2009.785 1126.290 ;
        RECT 2009.550 1112.450 2009.870 1113.300 ;
    END
  END mgmt_io_in_buf[28]
  PIN mgmt_io_in_buf[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2001.215 1113.300 2001.385 1114.150 ;
        RECT 2002.055 1113.300 2002.225 1114.150 ;
        RECT 2002.895 1113.300 2003.065 1114.150 ;
        RECT 2003.735 1113.300 2003.905 1114.150 ;
        RECT 2001.215 1113.130 2003.905 1113.300 ;
        RECT 2003.650 1112.590 2003.905 1113.130 ;
        RECT 2001.215 1112.420 2003.905 1112.590 ;
        RECT 2001.215 1111.940 2001.385 1112.420 ;
        RECT 2002.055 1111.940 2002.225 1112.420 ;
        RECT 2002.895 1111.940 2003.065 1112.420 ;
        RECT 2003.735 1111.940 2003.905 1112.420 ;
      LAYER mcon ;
        RECT 2003.650 1112.450 2003.820 1113.300 ;
      LAYER met1 ;
        RECT 2003.635 1127.000 3366.220 1127.140 ;
        RECT 2003.635 1126.880 2003.955 1127.000 ;
        RECT 2003.600 1112.390 2003.860 1113.360 ;
        RECT 3366.080 1084.250 3366.220 1127.000 ;
      LAYER via ;
        RECT 2003.665 1126.880 2003.925 1127.140 ;
        RECT 2003.600 1112.450 2003.860 1113.300 ;
      LAYER met2 ;
        RECT 2003.665 1127.170 2003.805 1129.765 ;
        RECT 2003.665 1126.850 2003.925 1127.170 ;
        RECT 2003.665 1113.300 2003.805 1126.850 ;
        RECT 2003.570 1112.450 2003.890 1113.300 ;
    END
  END mgmt_io_in_buf[29]
  PIN mgmt_io_in_buf[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1995.235 1113.300 1995.405 1114.150 ;
        RECT 1996.075 1113.300 1996.245 1114.150 ;
        RECT 1996.915 1113.300 1997.085 1114.150 ;
        RECT 1997.755 1113.300 1997.925 1114.150 ;
        RECT 1995.235 1113.130 1997.925 1113.300 ;
        RECT 1997.670 1112.590 1997.925 1113.130 ;
        RECT 1995.235 1112.420 1997.925 1112.590 ;
        RECT 1995.235 1111.940 1995.405 1112.420 ;
        RECT 1996.075 1111.940 1996.245 1112.420 ;
        RECT 1996.915 1111.940 1997.085 1112.420 ;
        RECT 1997.755 1111.940 1997.925 1112.420 ;
      LAYER mcon ;
        RECT 1997.670 1112.450 1997.840 1113.300 ;
      LAYER met1 ;
        RECT 1997.655 1127.560 3366.780 1127.700 ;
        RECT 1997.655 1127.440 1997.975 1127.560 ;
        RECT 1997.620 1112.390 1997.880 1113.360 ;
        RECT 3366.640 1082.250 3366.780 1127.560 ;
      LAYER via ;
        RECT 1997.685 1127.440 1997.945 1127.700 ;
        RECT 1997.620 1112.450 1997.880 1113.300 ;
      LAYER met2 ;
        RECT 1997.685 1127.730 1997.825 1129.765 ;
        RECT 1997.685 1127.410 1997.945 1127.730 ;
        RECT 1997.685 1113.300 1997.825 1127.410 ;
        RECT 1997.590 1112.450 1997.910 1113.300 ;
    END
  END mgmt_io_in_buf[30]
  PIN mgmt_io_in_buf[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1989.255 1113.300 1989.425 1114.150 ;
        RECT 1990.095 1113.300 1990.265 1114.150 ;
        RECT 1990.935 1113.300 1991.105 1114.150 ;
        RECT 1991.775 1113.300 1991.945 1114.150 ;
        RECT 1989.255 1113.130 1991.945 1113.300 ;
        RECT 1991.690 1112.590 1991.945 1113.130 ;
        RECT 1989.255 1112.420 1991.945 1112.590 ;
        RECT 1989.255 1111.940 1989.425 1112.420 ;
        RECT 1990.095 1111.940 1990.265 1112.420 ;
        RECT 1990.935 1111.940 1991.105 1112.420 ;
        RECT 1991.775 1111.940 1991.945 1112.420 ;
      LAYER mcon ;
        RECT 1991.690 1112.450 1991.860 1113.300 ;
      LAYER met1 ;
        RECT 1991.675 1128.120 3367.340 1128.260 ;
        RECT 1991.675 1128.000 1991.995 1128.120 ;
        RECT 1991.640 1112.390 1991.900 1113.360 ;
        RECT 3367.200 1080.250 3367.340 1128.120 ;
      LAYER via ;
        RECT 1991.705 1128.000 1991.965 1128.260 ;
        RECT 1991.640 1112.450 1991.900 1113.300 ;
      LAYER met2 ;
        RECT 1991.705 1128.290 1991.845 1129.765 ;
        RECT 1991.705 1127.970 1991.965 1128.290 ;
        RECT 1991.705 1113.300 1991.845 1127.970 ;
        RECT 1991.610 1112.450 1991.930 1113.300 ;
    END
  END mgmt_io_in_buf[31]
  PIN mgmt_io_in_buf[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1983.275 1113.300 1983.445 1114.150 ;
        RECT 1984.115 1113.300 1984.285 1114.150 ;
        RECT 1984.955 1113.300 1985.125 1114.150 ;
        RECT 1985.795 1113.300 1985.965 1114.150 ;
        RECT 1983.275 1113.130 1985.965 1113.300 ;
        RECT 1985.710 1112.590 1985.965 1113.130 ;
        RECT 1983.275 1112.420 1985.965 1112.590 ;
        RECT 1983.275 1111.940 1983.445 1112.420 ;
        RECT 1984.115 1111.940 1984.285 1112.420 ;
        RECT 1984.955 1111.940 1985.125 1112.420 ;
        RECT 1985.795 1111.940 1985.965 1112.420 ;
      LAYER mcon ;
        RECT 1985.710 1112.450 1985.880 1113.300 ;
      LAYER met1 ;
        RECT 1985.695 1128.680 3367.900 1128.820 ;
        RECT 1985.695 1128.560 1986.015 1128.680 ;
        RECT 1985.660 1112.390 1985.920 1113.360 ;
        RECT 3367.760 1078.250 3367.900 1128.680 ;
      LAYER via ;
        RECT 1985.725 1128.560 1985.985 1128.820 ;
        RECT 1985.660 1112.450 1985.920 1113.300 ;
      LAYER met2 ;
        RECT 1985.725 1128.850 1985.865 1129.765 ;
        RECT 1985.725 1128.530 1985.985 1128.850 ;
        RECT 1985.725 1113.300 1985.865 1128.530 ;
        RECT 1985.630 1112.450 1985.950 1113.300 ;
    END
  END mgmt_io_in_buf[32]
  PIN mgmt_io_in_buf[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1977.295 1113.300 1977.465 1114.150 ;
        RECT 1978.135 1113.300 1978.305 1114.150 ;
        RECT 1978.975 1113.300 1979.145 1114.150 ;
        RECT 1979.815 1113.300 1979.985 1114.150 ;
        RECT 1977.295 1113.130 1979.985 1113.300 ;
        RECT 1979.730 1112.590 1979.985 1113.130 ;
        RECT 1977.295 1112.420 1979.985 1112.590 ;
        RECT 1977.295 1111.940 1977.465 1112.420 ;
        RECT 1978.135 1111.940 1978.305 1112.420 ;
        RECT 1978.975 1111.940 1979.145 1112.420 ;
        RECT 1979.815 1111.940 1979.985 1112.420 ;
      LAYER mcon ;
        RECT 1979.730 1112.450 1979.900 1113.300 ;
      LAYER met1 ;
        RECT 1979.715 1129.240 3368.460 1129.380 ;
        RECT 1979.715 1129.120 1980.035 1129.240 ;
        RECT 1979.680 1112.390 1979.940 1113.360 ;
        RECT 3368.320 1076.250 3368.460 1129.240 ;
      LAYER via ;
        RECT 1979.745 1129.120 1980.005 1129.380 ;
        RECT 1979.680 1112.450 1979.940 1113.300 ;
      LAYER met2 ;
        RECT 1979.745 1129.410 1979.885 1129.765 ;
        RECT 1979.745 1129.090 1980.005 1129.410 ;
        RECT 1979.745 1113.300 1979.885 1129.090 ;
        RECT 1979.650 1112.450 1979.970 1113.300 ;
    END
  END mgmt_io_in_buf[33]
  PIN vssd
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 3312.980 4987.205 3313.150 4987.375 ;
        RECT 3313.440 4987.205 3313.610 4987.375 ;
        RECT 3313.900 4987.205 3314.070 4987.375 ;
        RECT 3314.360 4987.205 3314.530 4987.375 ;
        RECT 3314.820 4987.205 3314.990 4987.375 ;
        RECT 3315.280 4987.205 3315.450 4987.375 ;
        RECT 3315.740 4987.205 3315.910 4987.375 ;
        RECT 3316.200 4987.205 3316.370 4987.375 ;
        RECT 3316.660 4987.205 3316.830 4987.375 ;
        RECT 3317.120 4987.205 3317.290 4987.375 ;
        RECT 3317.580 4987.205 3317.750 4987.375 ;
        RECT 3318.040 4987.205 3318.210 4987.375 ;
        RECT 3318.500 4987.205 3318.670 4987.375 ;
        RECT 3318.960 4987.205 3319.130 4987.375 ;
        RECT 3319.420 4987.205 3319.590 4987.375 ;
        RECT 3319.880 4987.205 3320.050 4987.375 ;
        RECT 3320.340 4987.205 3320.510 4987.375 ;
        RECT 3320.800 4987.205 3320.970 4987.375 ;
        RECT 3321.260 4987.205 3321.430 4987.375 ;
        RECT 3321.720 4987.205 3321.890 4987.375 ;
        RECT 3322.180 4987.205 3322.350 4987.375 ;
        RECT 3322.640 4987.205 3322.810 4987.375 ;
        RECT 3323.100 4987.205 3323.270 4987.375 ;
        RECT 3323.560 4987.205 3323.730 4987.375 ;
        RECT 3324.020 4987.205 3324.190 4987.375 ;
        RECT 3324.480 4987.205 3324.650 4987.375 ;
        RECT 3324.940 4987.205 3325.110 4987.375 ;
        RECT 3325.400 4987.205 3325.570 4987.375 ;
        RECT 3325.860 4987.205 3326.030 4987.375 ;
        RECT 3326.320 4987.205 3326.490 4987.375 ;
        RECT 3326.780 4987.205 3326.950 4987.375 ;
        RECT 3327.240 4987.205 3327.410 4987.375 ;
        RECT 3327.700 4987.205 3327.870 4987.375 ;
        RECT 3328.160 4987.205 3328.330 4987.375 ;
        RECT 3328.620 4987.205 3328.790 4987.375 ;
        RECT 3329.080 4987.205 3329.250 4987.375 ;
        RECT 3329.540 4987.205 3329.710 4987.375 ;
        RECT 3330.000 4987.205 3330.170 4987.375 ;
        RECT 3330.460 4987.205 3330.630 4987.375 ;
        RECT 3330.920 4987.205 3331.090 4987.375 ;
        RECT 3331.380 4987.205 3331.550 4987.375 ;
        RECT 3331.840 4987.205 3332.010 4987.375 ;
        RECT 3332.300 4987.205 3332.470 4987.375 ;
        RECT 3332.760 4987.205 3332.930 4987.375 ;
        RECT 3333.220 4987.205 3333.390 4987.375 ;
        RECT 3333.680 4987.205 3333.850 4987.375 ;
        RECT 3334.140 4987.205 3334.310 4987.375 ;
        RECT 3334.600 4987.205 3334.770 4987.375 ;
        RECT 3335.060 4987.205 3335.230 4987.375 ;
        RECT 3335.520 4987.205 3335.690 4987.375 ;
        RECT 3335.980 4987.205 3336.150 4987.375 ;
        RECT 3336.440 4987.205 3336.610 4987.375 ;
        RECT 3336.900 4987.205 3337.070 4987.375 ;
        RECT 3312.980 4981.765 3313.150 4981.935 ;
        RECT 3313.440 4981.765 3313.610 4981.935 ;
        RECT 3313.900 4981.765 3314.070 4981.935 ;
        RECT 3314.360 4981.765 3314.530 4981.935 ;
        RECT 3314.820 4981.765 3314.990 4981.935 ;
        RECT 3315.280 4981.765 3315.450 4981.935 ;
        RECT 3315.740 4981.765 3315.910 4981.935 ;
        RECT 3316.200 4981.765 3316.370 4981.935 ;
        RECT 3316.660 4981.765 3316.830 4981.935 ;
        RECT 3317.120 4981.765 3317.290 4981.935 ;
        RECT 3317.580 4981.765 3317.750 4981.935 ;
        RECT 3318.040 4981.765 3318.210 4981.935 ;
        RECT 3318.500 4981.765 3318.670 4981.935 ;
        RECT 3318.960 4981.765 3319.130 4981.935 ;
        RECT 3319.420 4981.765 3319.590 4981.935 ;
        RECT 3319.880 4981.765 3320.050 4981.935 ;
        RECT 3320.340 4981.765 3320.510 4981.935 ;
        RECT 3320.800 4981.765 3320.970 4981.935 ;
        RECT 3321.260 4981.765 3321.430 4981.935 ;
        RECT 3321.720 4981.765 3321.890 4981.935 ;
        RECT 3322.180 4981.765 3322.350 4981.935 ;
        RECT 3322.640 4981.765 3322.810 4981.935 ;
        RECT 3323.100 4981.765 3323.270 4981.935 ;
        RECT 3323.560 4981.765 3323.730 4981.935 ;
        RECT 3324.020 4981.765 3324.190 4981.935 ;
        RECT 3324.480 4981.765 3324.650 4981.935 ;
        RECT 3324.940 4981.765 3325.110 4981.935 ;
        RECT 3325.400 4981.765 3325.570 4981.935 ;
        RECT 3325.860 4981.765 3326.030 4981.935 ;
        RECT 3326.320 4981.765 3326.490 4981.935 ;
        RECT 3326.780 4981.765 3326.950 4981.935 ;
        RECT 3327.240 4981.765 3327.410 4981.935 ;
        RECT 3327.700 4981.765 3327.870 4981.935 ;
        RECT 3328.160 4981.765 3328.330 4981.935 ;
        RECT 3328.620 4981.765 3328.790 4981.935 ;
        RECT 3329.080 4981.765 3329.250 4981.935 ;
        RECT 3329.540 4981.765 3329.710 4981.935 ;
        RECT 3330.000 4981.765 3330.170 4981.935 ;
        RECT 3330.460 4981.765 3330.630 4981.935 ;
        RECT 3330.920 4981.765 3331.090 4981.935 ;
        RECT 3331.380 4981.765 3331.550 4981.935 ;
        RECT 3331.840 4981.765 3332.010 4981.935 ;
        RECT 3332.300 4981.765 3332.470 4981.935 ;
        RECT 3332.760 4981.765 3332.930 4981.935 ;
        RECT 3333.220 4981.765 3333.390 4981.935 ;
        RECT 3333.680 4981.765 3333.850 4981.935 ;
        RECT 3334.140 4981.765 3334.310 4981.935 ;
        RECT 3334.600 4981.765 3334.770 4981.935 ;
        RECT 3335.060 4981.765 3335.230 4981.935 ;
        RECT 3335.520 4981.765 3335.690 4981.935 ;
        RECT 3335.980 4981.765 3336.150 4981.935 ;
        RECT 3336.440 4981.765 3336.610 4981.935 ;
        RECT 3336.900 4981.765 3337.070 4981.935 ;
      LAYER met1 ;
        RECT 3312.835 4987.050 3337.215 4987.530 ;
        RECT 3312.835 4981.610 3337.215 4982.090 ;
      LAYER via ;
        RECT 3321.185 4987.125 3322.970 4987.425 ;
        RECT 3321.185 4981.715 3322.970 4982.015 ;
      LAYER met2 ;
        RECT 3321.145 4987.080 3323.010 4987.510 ;
        RECT 3321.145 4981.655 3323.010 4982.085 ;
      LAYER via2 ;
        RECT 3321.185 4987.125 3322.970 4987.425 ;
        RECT 3321.185 4981.715 3322.970 4982.015 ;
      LAYER met3 ;
        RECT 3321.140 4981.640 3323.005 4989.165 ;
    END
    PORT
      LAYER li1 ;
        RECT 2082.975 4987.615 2083.145 4987.785 ;
        RECT 2083.435 4987.615 2083.605 4987.785 ;
        RECT 2083.895 4987.615 2084.065 4987.785 ;
        RECT 2084.355 4987.615 2084.525 4987.785 ;
        RECT 2084.815 4987.615 2084.985 4987.785 ;
        RECT 2085.275 4987.615 2085.445 4987.785 ;
        RECT 2085.735 4987.615 2085.905 4987.785 ;
        RECT 2086.195 4987.615 2086.365 4987.785 ;
        RECT 2086.655 4987.615 2086.825 4987.785 ;
        RECT 2087.115 4987.615 2087.285 4987.785 ;
        RECT 2087.575 4987.615 2087.745 4987.785 ;
        RECT 2088.035 4987.615 2088.205 4987.785 ;
        RECT 2088.495 4987.615 2088.665 4987.785 ;
        RECT 2088.955 4987.615 2089.125 4987.785 ;
        RECT 2082.975 4982.175 2083.145 4982.345 ;
        RECT 2083.435 4982.175 2083.605 4982.345 ;
        RECT 2083.895 4982.175 2084.065 4982.345 ;
        RECT 2084.355 4982.175 2084.525 4982.345 ;
        RECT 2084.815 4982.175 2084.985 4982.345 ;
        RECT 2085.275 4982.175 2085.445 4982.345 ;
        RECT 2085.735 4982.175 2085.905 4982.345 ;
        RECT 2086.195 4982.175 2086.365 4982.345 ;
        RECT 2086.655 4982.175 2086.825 4982.345 ;
        RECT 2087.115 4982.175 2087.285 4982.345 ;
        RECT 2087.575 4982.175 2087.745 4982.345 ;
        RECT 2088.035 4982.175 2088.205 4982.345 ;
        RECT 2088.495 4982.175 2088.665 4982.345 ;
        RECT 2088.955 4982.175 2089.125 4982.345 ;
      LAYER met1 ;
        RECT 2082.830 4987.460 2089.270 4987.940 ;
        RECT 2082.830 4982.020 2089.270 4982.500 ;
      LAYER via ;
        RECT 2085.135 4987.535 2086.920 4987.835 ;
        RECT 2085.135 4982.125 2086.920 4982.425 ;
      LAYER met2 ;
        RECT 2085.095 4987.490 2086.960 4987.920 ;
        RECT 2085.095 4982.065 2086.960 4982.495 ;
      LAYER via2 ;
        RECT 2085.135 4987.535 2086.920 4987.835 ;
        RECT 2085.135 4982.125 2086.920 4982.425 ;
      LAYER met3 ;
        RECT 2085.090 4982.050 2086.955 4989.575 ;
    END
    PORT
      LAYER li1 ;
        RECT 834.795 4985.990 834.965 4986.160 ;
        RECT 835.255 4985.990 835.425 4986.160 ;
        RECT 835.715 4985.990 835.885 4986.160 ;
        RECT 836.175 4985.990 836.345 4986.160 ;
        RECT 836.635 4985.990 836.805 4986.160 ;
        RECT 837.095 4985.990 837.265 4986.160 ;
        RECT 837.555 4985.990 837.725 4986.160 ;
        RECT 838.015 4985.990 838.185 4986.160 ;
        RECT 838.475 4985.990 838.645 4986.160 ;
        RECT 838.935 4985.990 839.105 4986.160 ;
        RECT 839.395 4985.990 839.565 4986.160 ;
        RECT 839.855 4985.990 840.025 4986.160 ;
        RECT 840.315 4985.990 840.485 4986.160 ;
        RECT 840.775 4985.990 840.945 4986.160 ;
        RECT 841.235 4985.990 841.405 4986.160 ;
        RECT 841.695 4985.990 841.865 4986.160 ;
        RECT 842.155 4985.990 842.325 4986.160 ;
        RECT 842.615 4985.990 842.785 4986.160 ;
        RECT 843.075 4985.990 843.245 4986.160 ;
        RECT 843.535 4985.990 843.705 4986.160 ;
        RECT 843.995 4985.990 844.165 4986.160 ;
        RECT 844.455 4985.990 844.625 4986.160 ;
        RECT 844.915 4985.990 845.085 4986.160 ;
        RECT 845.375 4985.990 845.545 4986.160 ;
        RECT 845.835 4985.990 846.005 4986.160 ;
        RECT 846.295 4985.990 846.465 4986.160 ;
        RECT 846.755 4985.990 846.925 4986.160 ;
        RECT 847.215 4985.990 847.385 4986.160 ;
        RECT 847.675 4985.990 847.845 4986.160 ;
        RECT 848.135 4985.990 848.305 4986.160 ;
        RECT 848.595 4985.990 848.765 4986.160 ;
        RECT 849.055 4985.990 849.225 4986.160 ;
        RECT 849.515 4985.990 849.685 4986.160 ;
        RECT 849.975 4985.990 850.145 4986.160 ;
        RECT 850.435 4985.990 850.605 4986.160 ;
        RECT 850.895 4985.990 851.065 4986.160 ;
        RECT 851.355 4985.990 851.525 4986.160 ;
        RECT 851.815 4985.990 851.985 4986.160 ;
        RECT 852.275 4985.990 852.445 4986.160 ;
        RECT 852.735 4985.990 852.905 4986.160 ;
        RECT 834.795 4980.550 834.965 4980.720 ;
        RECT 835.255 4980.550 835.425 4980.720 ;
        RECT 835.715 4980.550 835.885 4980.720 ;
        RECT 836.175 4980.550 836.345 4980.720 ;
        RECT 836.635 4980.550 836.805 4980.720 ;
        RECT 837.095 4980.550 837.265 4980.720 ;
        RECT 837.555 4980.550 837.725 4980.720 ;
        RECT 838.015 4980.550 838.185 4980.720 ;
        RECT 838.475 4980.550 838.645 4980.720 ;
        RECT 838.935 4980.550 839.105 4980.720 ;
        RECT 839.395 4980.550 839.565 4980.720 ;
        RECT 839.855 4980.550 840.025 4980.720 ;
        RECT 840.315 4980.550 840.485 4980.720 ;
        RECT 840.775 4980.550 840.945 4980.720 ;
        RECT 841.235 4980.550 841.405 4980.720 ;
        RECT 841.695 4980.550 841.865 4980.720 ;
        RECT 842.155 4980.550 842.325 4980.720 ;
        RECT 842.615 4980.550 842.785 4980.720 ;
        RECT 843.075 4980.550 843.245 4980.720 ;
        RECT 843.535 4980.550 843.705 4980.720 ;
        RECT 843.995 4980.550 844.165 4980.720 ;
        RECT 844.455 4980.550 844.625 4980.720 ;
        RECT 844.915 4980.550 845.085 4980.720 ;
        RECT 845.375 4980.550 845.545 4980.720 ;
        RECT 845.835 4980.550 846.005 4980.720 ;
        RECT 846.295 4980.550 846.465 4980.720 ;
        RECT 846.755 4980.550 846.925 4980.720 ;
        RECT 847.215 4980.550 847.385 4980.720 ;
        RECT 847.675 4980.550 847.845 4980.720 ;
        RECT 848.135 4980.550 848.305 4980.720 ;
        RECT 848.595 4980.550 848.765 4980.720 ;
        RECT 849.055 4980.550 849.225 4980.720 ;
        RECT 849.515 4980.550 849.685 4980.720 ;
        RECT 849.975 4980.550 850.145 4980.720 ;
        RECT 850.435 4980.550 850.605 4980.720 ;
        RECT 850.895 4980.550 851.065 4980.720 ;
        RECT 851.355 4980.550 851.525 4980.720 ;
        RECT 851.815 4980.550 851.985 4980.720 ;
        RECT 852.275 4980.550 852.445 4980.720 ;
        RECT 852.735 4980.550 852.905 4980.720 ;
      LAYER met1 ;
        RECT 834.650 4985.835 853.050 4986.315 ;
        RECT 834.650 4980.395 853.050 4980.875 ;
      LAYER via ;
        RECT 842.950 4985.890 844.735 4986.190 ;
        RECT 842.950 4980.480 844.735 4980.780 ;
      LAYER met2 ;
        RECT 842.910 4985.845 844.775 4986.275 ;
        RECT 842.910 4980.420 844.775 4980.850 ;
      LAYER via2 ;
        RECT 842.950 4985.890 844.735 4986.190 ;
        RECT 842.950 4980.480 844.735 4980.780 ;
      LAYER met3 ;
        RECT 842.905 4980.405 844.770 4987.930 ;
    END
    PORT
      LAYER li1 ;
        RECT 669.145 1117.040 669.315 1117.210 ;
        RECT 669.605 1117.040 669.775 1117.210 ;
        RECT 670.065 1117.040 670.235 1117.210 ;
        RECT 670.525 1117.040 670.695 1117.210 ;
        RECT 670.985 1117.040 671.155 1117.210 ;
        RECT 671.445 1117.040 671.615 1117.210 ;
        RECT 671.905 1117.040 672.075 1117.210 ;
        RECT 672.365 1117.040 672.535 1117.210 ;
        RECT 672.825 1117.040 672.995 1117.210 ;
        RECT 673.285 1117.040 673.455 1117.210 ;
        RECT 673.745 1117.040 673.915 1117.210 ;
        RECT 674.205 1117.040 674.375 1117.210 ;
        RECT 674.665 1117.040 674.835 1117.210 ;
        RECT 675.125 1117.040 675.295 1117.210 ;
        RECT 675.585 1117.040 675.755 1117.210 ;
        RECT 676.045 1117.040 676.215 1117.210 ;
        RECT 676.505 1117.040 676.675 1117.210 ;
        RECT 676.965 1117.040 677.135 1117.210 ;
        RECT 677.425 1117.040 677.595 1117.210 ;
        RECT 677.885 1117.040 678.055 1117.210 ;
        RECT 678.345 1117.040 678.515 1117.210 ;
        RECT 678.805 1117.040 678.975 1117.210 ;
        RECT 679.265 1117.040 679.435 1117.210 ;
        RECT 679.725 1117.040 679.895 1117.210 ;
        RECT 680.185 1117.040 680.355 1117.210 ;
        RECT 680.645 1117.040 680.815 1117.210 ;
        RECT 681.105 1117.040 681.275 1117.210 ;
        RECT 681.565 1117.040 681.735 1117.210 ;
        RECT 682.025 1117.040 682.195 1117.210 ;
        RECT 682.485 1117.040 682.655 1117.210 ;
        RECT 682.945 1117.040 683.115 1117.210 ;
        RECT 683.405 1117.040 683.575 1117.210 ;
        RECT 683.865 1117.040 684.035 1117.210 ;
        RECT 684.325 1117.040 684.495 1117.210 ;
        RECT 684.785 1117.040 684.955 1117.210 ;
        RECT 685.245 1117.040 685.415 1117.210 ;
        RECT 685.705 1117.040 685.875 1117.210 ;
        RECT 686.165 1117.040 686.335 1117.210 ;
        RECT 686.625 1117.040 686.795 1117.210 ;
        RECT 687.085 1117.040 687.255 1117.210 ;
        RECT 687.545 1117.040 687.715 1117.210 ;
        RECT 688.005 1117.040 688.175 1117.210 ;
        RECT 688.465 1117.040 688.635 1117.210 ;
        RECT 688.925 1117.040 689.095 1117.210 ;
        RECT 689.385 1117.040 689.555 1117.210 ;
        RECT 689.845 1117.040 690.015 1117.210 ;
        RECT 690.305 1117.040 690.475 1117.210 ;
        RECT 690.765 1117.040 690.935 1117.210 ;
        RECT 691.225 1117.040 691.395 1117.210 ;
        RECT 691.685 1117.040 691.855 1117.210 ;
        RECT 692.145 1117.040 692.315 1117.210 ;
        RECT 692.605 1117.040 692.775 1117.210 ;
        RECT 693.065 1117.040 693.235 1117.210 ;
        RECT 693.525 1117.040 693.695 1117.210 ;
        RECT 693.985 1117.040 694.155 1117.210 ;
        RECT 694.445 1117.040 694.615 1117.210 ;
        RECT 694.905 1117.040 695.075 1117.210 ;
        RECT 695.365 1117.040 695.535 1117.210 ;
        RECT 695.825 1117.040 695.995 1117.210 ;
        RECT 696.285 1117.040 696.455 1117.210 ;
        RECT 696.745 1117.040 696.915 1117.210 ;
        RECT 697.205 1117.040 697.375 1117.210 ;
        RECT 697.665 1117.040 697.835 1117.210 ;
        RECT 698.125 1117.040 698.295 1117.210 ;
        RECT 698.585 1117.040 698.755 1117.210 ;
        RECT 699.045 1117.040 699.215 1117.210 ;
        RECT 699.505 1117.040 699.675 1117.210 ;
        RECT 699.965 1117.040 700.135 1117.210 ;
        RECT 700.425 1117.040 700.595 1117.210 ;
        RECT 700.885 1117.040 701.055 1117.210 ;
        RECT 701.345 1117.040 701.515 1117.210 ;
        RECT 701.805 1117.040 701.975 1117.210 ;
        RECT 702.265 1117.040 702.435 1117.210 ;
        RECT 702.725 1117.040 702.895 1117.210 ;
        RECT 703.185 1117.040 703.355 1117.210 ;
        RECT 703.645 1117.040 703.815 1117.210 ;
        RECT 704.105 1117.040 704.275 1117.210 ;
        RECT 704.565 1117.040 704.735 1117.210 ;
        RECT 705.025 1117.040 705.195 1117.210 ;
        RECT 705.485 1117.040 705.655 1117.210 ;
        RECT 705.945 1117.040 706.115 1117.210 ;
        RECT 706.405 1117.040 706.575 1117.210 ;
        RECT 706.865 1117.040 707.035 1117.210 ;
        RECT 707.325 1117.040 707.495 1117.210 ;
        RECT 707.785 1117.040 707.955 1117.210 ;
        RECT 708.245 1117.040 708.415 1117.210 ;
        RECT 708.705 1117.040 708.875 1117.210 ;
        RECT 709.165 1117.040 709.335 1117.210 ;
        RECT 709.625 1117.040 709.795 1117.210 ;
        RECT 710.085 1117.040 710.255 1117.210 ;
        RECT 710.545 1117.040 710.715 1117.210 ;
        RECT 711.005 1117.040 711.175 1117.210 ;
        RECT 711.465 1117.040 711.635 1117.210 ;
        RECT 711.925 1117.040 712.095 1117.210 ;
        RECT 712.385 1117.040 712.555 1117.210 ;
        RECT 712.845 1117.040 713.015 1117.210 ;
        RECT 713.305 1117.040 713.475 1117.210 ;
        RECT 713.765 1117.040 713.935 1117.210 ;
        RECT 714.225 1117.040 714.395 1117.210 ;
        RECT 714.685 1117.040 714.855 1117.210 ;
        RECT 715.145 1117.040 715.315 1117.210 ;
        RECT 715.605 1117.040 715.775 1117.210 ;
        RECT 716.065 1117.040 716.235 1117.210 ;
        RECT 716.525 1117.040 716.695 1117.210 ;
        RECT 716.985 1117.040 717.155 1117.210 ;
        RECT 717.445 1117.040 717.615 1117.210 ;
        RECT 717.905 1117.040 718.075 1117.210 ;
        RECT 718.365 1117.040 718.535 1117.210 ;
        RECT 718.825 1117.040 718.995 1117.210 ;
        RECT 719.285 1117.040 719.455 1117.210 ;
        RECT 719.745 1117.040 719.915 1117.210 ;
        RECT 720.205 1117.040 720.375 1117.210 ;
        RECT 720.665 1117.040 720.835 1117.210 ;
        RECT 721.125 1117.040 721.295 1117.210 ;
        RECT 721.585 1117.040 721.755 1117.210 ;
        RECT 722.045 1117.040 722.215 1117.210 ;
        RECT 722.505 1117.040 722.675 1117.210 ;
        RECT 722.965 1117.040 723.135 1117.210 ;
        RECT 723.425 1117.040 723.595 1117.210 ;
        RECT 723.885 1117.040 724.055 1117.210 ;
        RECT 724.345 1117.040 724.515 1117.210 ;
        RECT 724.805 1117.040 724.975 1117.210 ;
        RECT 725.265 1117.040 725.435 1117.210 ;
        RECT 725.725 1117.040 725.895 1117.210 ;
        RECT 726.185 1117.040 726.355 1117.210 ;
        RECT 726.645 1117.040 726.815 1117.210 ;
        RECT 727.105 1117.040 727.275 1117.210 ;
        RECT 727.565 1117.040 727.735 1117.210 ;
        RECT 728.025 1117.040 728.195 1117.210 ;
        RECT 728.485 1117.040 728.655 1117.210 ;
        RECT 728.945 1117.040 729.115 1117.210 ;
        RECT 729.405 1117.040 729.575 1117.210 ;
        RECT 729.865 1117.040 730.035 1117.210 ;
        RECT 730.325 1117.040 730.495 1117.210 ;
        RECT 730.785 1117.040 730.955 1117.210 ;
        RECT 731.245 1117.040 731.415 1117.210 ;
        RECT 731.705 1117.040 731.875 1117.210 ;
        RECT 732.165 1117.040 732.335 1117.210 ;
        RECT 732.625 1117.040 732.795 1117.210 ;
        RECT 733.085 1117.040 733.255 1117.210 ;
        RECT 733.545 1117.040 733.715 1117.210 ;
        RECT 734.005 1117.040 734.175 1117.210 ;
        RECT 734.465 1117.040 734.635 1117.210 ;
        RECT 734.925 1117.040 735.095 1117.210 ;
        RECT 735.385 1117.040 735.555 1117.210 ;
        RECT 735.845 1117.040 736.015 1117.210 ;
        RECT 736.305 1117.040 736.475 1117.210 ;
        RECT 736.765 1117.040 736.935 1117.210 ;
        RECT 737.225 1117.040 737.395 1117.210 ;
        RECT 737.685 1117.040 737.855 1117.210 ;
        RECT 738.145 1117.040 738.315 1117.210 ;
        RECT 738.605 1117.040 738.775 1117.210 ;
        RECT 739.065 1117.040 739.235 1117.210 ;
        RECT 739.525 1117.040 739.695 1117.210 ;
        RECT 739.985 1117.040 740.155 1117.210 ;
        RECT 740.445 1117.040 740.615 1117.210 ;
        RECT 740.905 1117.040 741.075 1117.210 ;
        RECT 741.365 1117.040 741.535 1117.210 ;
        RECT 741.825 1117.040 741.995 1117.210 ;
        RECT 742.285 1117.040 742.455 1117.210 ;
        RECT 742.745 1117.040 742.915 1117.210 ;
        RECT 743.205 1117.040 743.375 1117.210 ;
        RECT 743.665 1117.040 743.835 1117.210 ;
        RECT 744.125 1117.040 744.295 1117.210 ;
        RECT 744.585 1117.040 744.755 1117.210 ;
        RECT 745.045 1117.040 745.215 1117.210 ;
        RECT 745.505 1117.040 745.675 1117.210 ;
        RECT 745.965 1117.040 746.135 1117.210 ;
        RECT 746.425 1117.040 746.595 1117.210 ;
        RECT 746.885 1117.040 747.055 1117.210 ;
        RECT 747.345 1117.040 747.515 1117.210 ;
        RECT 747.805 1117.040 747.975 1117.210 ;
        RECT 748.265 1117.040 748.435 1117.210 ;
        RECT 748.725 1117.040 748.895 1117.210 ;
        RECT 749.185 1117.040 749.355 1117.210 ;
        RECT 749.645 1117.040 749.815 1117.210 ;
        RECT 750.105 1117.040 750.275 1117.210 ;
        RECT 750.565 1117.040 750.735 1117.210 ;
        RECT 751.025 1117.040 751.195 1117.210 ;
        RECT 751.485 1117.040 751.655 1117.210 ;
        RECT 751.945 1117.040 752.115 1117.210 ;
        RECT 752.405 1117.040 752.575 1117.210 ;
        RECT 752.865 1117.040 753.035 1117.210 ;
        RECT 753.325 1117.040 753.495 1117.210 ;
        RECT 753.785 1117.040 753.955 1117.210 ;
        RECT 754.245 1117.040 754.415 1117.210 ;
        RECT 754.705 1117.040 754.875 1117.210 ;
        RECT 755.165 1117.040 755.335 1117.210 ;
        RECT 755.625 1117.040 755.795 1117.210 ;
        RECT 756.085 1117.040 756.255 1117.210 ;
        RECT 756.545 1117.040 756.715 1117.210 ;
        RECT 757.005 1117.040 757.175 1117.210 ;
        RECT 757.465 1117.040 757.635 1117.210 ;
        RECT 757.925 1117.040 758.095 1117.210 ;
        RECT 758.385 1117.040 758.555 1117.210 ;
        RECT 758.845 1117.040 759.015 1117.210 ;
        RECT 759.305 1117.040 759.475 1117.210 ;
        RECT 759.765 1117.040 759.935 1117.210 ;
        RECT 760.225 1117.040 760.395 1117.210 ;
        RECT 760.685 1117.040 760.855 1117.210 ;
        RECT 761.145 1117.040 761.315 1117.210 ;
        RECT 761.605 1117.040 761.775 1117.210 ;
        RECT 762.065 1117.040 762.235 1117.210 ;
        RECT 762.525 1117.040 762.695 1117.210 ;
        RECT 762.985 1117.040 763.155 1117.210 ;
        RECT 763.445 1117.040 763.615 1117.210 ;
        RECT 763.905 1117.040 764.075 1117.210 ;
        RECT 764.365 1117.040 764.535 1117.210 ;
        RECT 764.825 1117.040 764.995 1117.210 ;
        RECT 765.285 1117.040 765.455 1117.210 ;
        RECT 765.745 1117.040 765.915 1117.210 ;
        RECT 766.205 1117.040 766.375 1117.210 ;
        RECT 766.665 1117.040 766.835 1117.210 ;
        RECT 767.125 1117.040 767.295 1117.210 ;
        RECT 767.585 1117.040 767.755 1117.210 ;
        RECT 768.045 1117.040 768.215 1117.210 ;
        RECT 768.505 1117.040 768.675 1117.210 ;
        RECT 768.965 1117.040 769.135 1117.210 ;
        RECT 769.425 1117.040 769.595 1117.210 ;
        RECT 769.885 1117.040 770.055 1117.210 ;
        RECT 770.345 1117.040 770.515 1117.210 ;
        RECT 770.805 1117.040 770.975 1117.210 ;
        RECT 771.265 1117.040 771.435 1117.210 ;
        RECT 771.725 1117.040 771.895 1117.210 ;
        RECT 772.185 1117.040 772.355 1117.210 ;
        RECT 772.645 1117.040 772.815 1117.210 ;
        RECT 773.105 1117.040 773.275 1117.210 ;
        RECT 773.565 1117.040 773.735 1117.210 ;
        RECT 774.025 1117.040 774.195 1117.210 ;
        RECT 774.485 1117.040 774.655 1117.210 ;
        RECT 774.945 1117.040 775.115 1117.210 ;
        RECT 775.405 1117.040 775.575 1117.210 ;
        RECT 775.865 1117.040 776.035 1117.210 ;
        RECT 776.325 1117.040 776.495 1117.210 ;
        RECT 776.785 1117.040 776.955 1117.210 ;
        RECT 777.245 1117.040 777.415 1117.210 ;
        RECT 777.705 1117.040 777.875 1117.210 ;
        RECT 778.165 1117.040 778.335 1117.210 ;
        RECT 778.625 1117.040 778.795 1117.210 ;
        RECT 779.085 1117.040 779.255 1117.210 ;
        RECT 779.545 1117.040 779.715 1117.210 ;
        RECT 780.005 1117.040 780.175 1117.210 ;
        RECT 780.465 1117.040 780.635 1117.210 ;
        RECT 780.925 1117.040 781.095 1117.210 ;
        RECT 781.385 1117.040 781.555 1117.210 ;
        RECT 781.845 1117.040 782.015 1117.210 ;
        RECT 782.305 1117.040 782.475 1117.210 ;
        RECT 782.765 1117.040 782.935 1117.210 ;
        RECT 783.225 1117.040 783.395 1117.210 ;
        RECT 783.685 1117.040 783.855 1117.210 ;
        RECT 784.145 1117.040 784.315 1117.210 ;
        RECT 784.605 1117.040 784.775 1117.210 ;
        RECT 785.065 1117.040 785.235 1117.210 ;
        RECT 785.525 1117.040 785.695 1117.210 ;
        RECT 785.985 1117.040 786.155 1117.210 ;
        RECT 786.445 1117.040 786.615 1117.210 ;
        RECT 786.905 1117.040 787.075 1117.210 ;
        RECT 787.365 1117.040 787.535 1117.210 ;
        RECT 787.825 1117.040 787.995 1117.210 ;
        RECT 788.285 1117.040 788.455 1117.210 ;
        RECT 788.745 1117.040 788.915 1117.210 ;
        RECT 789.205 1117.040 789.375 1117.210 ;
        RECT 789.665 1117.040 789.835 1117.210 ;
        RECT 790.125 1117.040 790.295 1117.210 ;
        RECT 790.585 1117.040 790.755 1117.210 ;
        RECT 791.045 1117.040 791.215 1117.210 ;
        RECT 791.505 1117.040 791.675 1117.210 ;
        RECT 791.965 1117.040 792.135 1117.210 ;
        RECT 792.425 1117.040 792.595 1117.210 ;
        RECT 792.885 1117.040 793.055 1117.210 ;
        RECT 793.345 1117.040 793.515 1117.210 ;
        RECT 793.805 1117.040 793.975 1117.210 ;
        RECT 794.265 1117.040 794.435 1117.210 ;
        RECT 794.725 1117.040 794.895 1117.210 ;
        RECT 675.125 1111.600 675.295 1111.770 ;
        RECT 675.585 1111.600 675.755 1111.770 ;
        RECT 676.045 1111.600 676.215 1111.770 ;
        RECT 676.505 1111.600 676.675 1111.770 ;
        RECT 676.965 1111.600 677.135 1111.770 ;
        RECT 677.425 1111.600 677.595 1111.770 ;
        RECT 677.885 1111.600 678.055 1111.770 ;
        RECT 678.345 1111.600 678.515 1111.770 ;
        RECT 678.805 1111.600 678.975 1111.770 ;
        RECT 679.265 1111.600 679.435 1111.770 ;
        RECT 679.725 1111.600 679.895 1111.770 ;
        RECT 680.185 1111.600 680.355 1111.770 ;
        RECT 680.645 1111.600 680.815 1111.770 ;
        RECT 681.105 1111.600 681.275 1111.770 ;
        RECT 681.565 1111.600 681.735 1111.770 ;
        RECT 682.025 1111.600 682.195 1111.770 ;
        RECT 682.485 1111.600 682.655 1111.770 ;
        RECT 682.945 1111.600 683.115 1111.770 ;
        RECT 683.405 1111.600 683.575 1111.770 ;
        RECT 683.865 1111.600 684.035 1111.770 ;
        RECT 684.325 1111.600 684.495 1111.770 ;
        RECT 684.785 1111.600 684.955 1111.770 ;
        RECT 685.245 1111.600 685.415 1111.770 ;
        RECT 685.705 1111.600 685.875 1111.770 ;
        RECT 686.165 1111.600 686.335 1111.770 ;
        RECT 686.625 1111.600 686.795 1111.770 ;
        RECT 687.085 1111.600 687.255 1111.770 ;
        RECT 687.545 1111.600 687.715 1111.770 ;
        RECT 688.005 1111.600 688.175 1111.770 ;
        RECT 688.465 1111.600 688.635 1111.770 ;
        RECT 688.925 1111.600 689.095 1111.770 ;
        RECT 689.385 1111.600 689.555 1111.770 ;
        RECT 689.845 1111.600 690.015 1111.770 ;
        RECT 690.305 1111.600 690.475 1111.770 ;
        RECT 690.765 1111.600 690.935 1111.770 ;
        RECT 691.225 1111.600 691.395 1111.770 ;
        RECT 691.685 1111.600 691.855 1111.770 ;
        RECT 692.145 1111.600 692.315 1111.770 ;
        RECT 692.605 1111.600 692.775 1111.770 ;
        RECT 693.065 1111.600 693.235 1111.770 ;
        RECT 693.525 1111.600 693.695 1111.770 ;
        RECT 693.985 1111.600 694.155 1111.770 ;
        RECT 694.445 1111.600 694.615 1111.770 ;
        RECT 694.905 1111.600 695.075 1111.770 ;
        RECT 695.365 1111.600 695.535 1111.770 ;
        RECT 695.825 1111.600 695.995 1111.770 ;
        RECT 696.285 1111.600 696.455 1111.770 ;
        RECT 696.745 1111.600 696.915 1111.770 ;
        RECT 697.205 1111.600 697.375 1111.770 ;
        RECT 697.665 1111.600 697.835 1111.770 ;
        RECT 698.125 1111.600 698.295 1111.770 ;
        RECT 698.585 1111.600 698.755 1111.770 ;
        RECT 699.045 1111.600 699.215 1111.770 ;
        RECT 699.505 1111.600 699.675 1111.770 ;
        RECT 699.965 1111.600 700.135 1111.770 ;
        RECT 700.425 1111.600 700.595 1111.770 ;
        RECT 700.885 1111.600 701.055 1111.770 ;
        RECT 701.345 1111.600 701.515 1111.770 ;
        RECT 701.805 1111.600 701.975 1111.770 ;
        RECT 702.265 1111.600 702.435 1111.770 ;
        RECT 702.725 1111.600 702.895 1111.770 ;
        RECT 703.185 1111.600 703.355 1111.770 ;
        RECT 703.645 1111.600 703.815 1111.770 ;
        RECT 704.105 1111.600 704.275 1111.770 ;
        RECT 704.565 1111.600 704.735 1111.770 ;
        RECT 705.025 1111.600 705.195 1111.770 ;
        RECT 705.485 1111.600 705.655 1111.770 ;
        RECT 705.945 1111.600 706.115 1111.770 ;
        RECT 706.405 1111.600 706.575 1111.770 ;
        RECT 706.865 1111.600 707.035 1111.770 ;
        RECT 707.325 1111.600 707.495 1111.770 ;
        RECT 707.785 1111.600 707.955 1111.770 ;
        RECT 708.245 1111.600 708.415 1111.770 ;
        RECT 708.705 1111.600 708.875 1111.770 ;
        RECT 709.165 1111.600 709.335 1111.770 ;
        RECT 709.625 1111.600 709.795 1111.770 ;
        RECT 710.085 1111.600 710.255 1111.770 ;
        RECT 710.545 1111.600 710.715 1111.770 ;
        RECT 711.005 1111.600 711.175 1111.770 ;
        RECT 711.465 1111.600 711.635 1111.770 ;
        RECT 711.925 1111.600 712.095 1111.770 ;
        RECT 712.385 1111.600 712.555 1111.770 ;
        RECT 712.845 1111.600 713.015 1111.770 ;
        RECT 713.305 1111.600 713.475 1111.770 ;
        RECT 713.765 1111.600 713.935 1111.770 ;
        RECT 714.225 1111.600 714.395 1111.770 ;
        RECT 714.685 1111.600 714.855 1111.770 ;
        RECT 715.145 1111.600 715.315 1111.770 ;
        RECT 715.605 1111.600 715.775 1111.770 ;
        RECT 716.065 1111.600 716.235 1111.770 ;
        RECT 716.525 1111.600 716.695 1111.770 ;
        RECT 716.985 1111.600 717.155 1111.770 ;
        RECT 717.445 1111.600 717.615 1111.770 ;
        RECT 717.905 1111.600 718.075 1111.770 ;
        RECT 718.365 1111.600 718.535 1111.770 ;
        RECT 718.825 1111.600 718.995 1111.770 ;
        RECT 719.285 1111.600 719.455 1111.770 ;
        RECT 719.745 1111.600 719.915 1111.770 ;
        RECT 720.205 1111.600 720.375 1111.770 ;
        RECT 720.665 1111.600 720.835 1111.770 ;
        RECT 721.125 1111.600 721.295 1111.770 ;
        RECT 721.585 1111.600 721.755 1111.770 ;
        RECT 722.045 1111.600 722.215 1111.770 ;
        RECT 722.505 1111.600 722.675 1111.770 ;
        RECT 722.965 1111.600 723.135 1111.770 ;
        RECT 723.425 1111.600 723.595 1111.770 ;
        RECT 723.885 1111.600 724.055 1111.770 ;
        RECT 724.345 1111.600 724.515 1111.770 ;
        RECT 724.805 1111.600 724.975 1111.770 ;
        RECT 725.265 1111.600 725.435 1111.770 ;
        RECT 725.725 1111.600 725.895 1111.770 ;
        RECT 726.185 1111.600 726.355 1111.770 ;
        RECT 726.645 1111.600 726.815 1111.770 ;
        RECT 727.105 1111.600 727.275 1111.770 ;
        RECT 727.565 1111.600 727.735 1111.770 ;
        RECT 728.025 1111.600 728.195 1111.770 ;
        RECT 728.485 1111.600 728.655 1111.770 ;
        RECT 728.945 1111.600 729.115 1111.770 ;
        RECT 729.405 1111.600 729.575 1111.770 ;
        RECT 729.865 1111.600 730.035 1111.770 ;
        RECT 730.325 1111.600 730.495 1111.770 ;
        RECT 730.785 1111.600 730.955 1111.770 ;
        RECT 731.245 1111.600 731.415 1111.770 ;
        RECT 731.705 1111.600 731.875 1111.770 ;
        RECT 732.165 1111.600 732.335 1111.770 ;
        RECT 732.625 1111.600 732.795 1111.770 ;
        RECT 733.085 1111.600 733.255 1111.770 ;
        RECT 733.545 1111.600 733.715 1111.770 ;
        RECT 734.005 1111.600 734.175 1111.770 ;
        RECT 734.465 1111.600 734.635 1111.770 ;
        RECT 734.925 1111.600 735.095 1111.770 ;
        RECT 735.385 1111.600 735.555 1111.770 ;
        RECT 735.845 1111.600 736.015 1111.770 ;
        RECT 736.305 1111.600 736.475 1111.770 ;
        RECT 736.765 1111.600 736.935 1111.770 ;
        RECT 737.225 1111.600 737.395 1111.770 ;
        RECT 737.685 1111.600 737.855 1111.770 ;
        RECT 738.145 1111.600 738.315 1111.770 ;
        RECT 738.605 1111.600 738.775 1111.770 ;
        RECT 739.065 1111.600 739.235 1111.770 ;
        RECT 739.525 1111.600 739.695 1111.770 ;
        RECT 739.985 1111.600 740.155 1111.770 ;
        RECT 740.445 1111.600 740.615 1111.770 ;
        RECT 740.905 1111.600 741.075 1111.770 ;
        RECT 741.365 1111.600 741.535 1111.770 ;
        RECT 741.825 1111.600 741.995 1111.770 ;
        RECT 742.285 1111.600 742.455 1111.770 ;
        RECT 742.745 1111.600 742.915 1111.770 ;
        RECT 743.205 1111.600 743.375 1111.770 ;
        RECT 743.665 1111.600 743.835 1111.770 ;
        RECT 744.125 1111.600 744.295 1111.770 ;
        RECT 744.585 1111.600 744.755 1111.770 ;
        RECT 745.045 1111.600 745.215 1111.770 ;
        RECT 745.505 1111.600 745.675 1111.770 ;
        RECT 745.965 1111.600 746.135 1111.770 ;
        RECT 746.425 1111.600 746.595 1111.770 ;
        RECT 746.885 1111.600 747.055 1111.770 ;
        RECT 747.345 1111.600 747.515 1111.770 ;
        RECT 747.805 1111.600 747.975 1111.770 ;
        RECT 748.265 1111.600 748.435 1111.770 ;
        RECT 748.725 1111.600 748.895 1111.770 ;
        RECT 749.185 1111.600 749.355 1111.770 ;
        RECT 749.645 1111.600 749.815 1111.770 ;
        RECT 750.105 1111.600 750.275 1111.770 ;
        RECT 750.565 1111.600 750.735 1111.770 ;
        RECT 751.025 1111.600 751.195 1111.770 ;
        RECT 751.485 1111.600 751.655 1111.770 ;
        RECT 751.945 1111.600 752.115 1111.770 ;
        RECT 752.405 1111.600 752.575 1111.770 ;
        RECT 752.865 1111.600 753.035 1111.770 ;
        RECT 753.325 1111.600 753.495 1111.770 ;
        RECT 753.785 1111.600 753.955 1111.770 ;
        RECT 754.245 1111.600 754.415 1111.770 ;
        RECT 754.705 1111.600 754.875 1111.770 ;
        RECT 755.165 1111.600 755.335 1111.770 ;
        RECT 755.625 1111.600 755.795 1111.770 ;
        RECT 756.085 1111.600 756.255 1111.770 ;
        RECT 756.545 1111.600 756.715 1111.770 ;
        RECT 757.005 1111.600 757.175 1111.770 ;
        RECT 757.465 1111.600 757.635 1111.770 ;
        RECT 757.925 1111.600 758.095 1111.770 ;
        RECT 758.385 1111.600 758.555 1111.770 ;
        RECT 758.845 1111.600 759.015 1111.770 ;
        RECT 759.305 1111.600 759.475 1111.770 ;
        RECT 759.765 1111.600 759.935 1111.770 ;
        RECT 760.225 1111.600 760.395 1111.770 ;
        RECT 760.685 1111.600 760.855 1111.770 ;
        RECT 761.145 1111.600 761.315 1111.770 ;
        RECT 761.605 1111.600 761.775 1111.770 ;
        RECT 762.065 1111.600 762.235 1111.770 ;
        RECT 762.525 1111.600 762.695 1111.770 ;
        RECT 762.985 1111.600 763.155 1111.770 ;
        RECT 763.445 1111.600 763.615 1111.770 ;
        RECT 763.905 1111.600 764.075 1111.770 ;
        RECT 764.365 1111.600 764.535 1111.770 ;
        RECT 764.825 1111.600 764.995 1111.770 ;
        RECT 765.285 1111.600 765.455 1111.770 ;
        RECT 765.745 1111.600 765.915 1111.770 ;
        RECT 766.205 1111.600 766.375 1111.770 ;
        RECT 766.665 1111.600 766.835 1111.770 ;
        RECT 767.125 1111.600 767.295 1111.770 ;
        RECT 767.585 1111.600 767.755 1111.770 ;
        RECT 768.045 1111.600 768.215 1111.770 ;
        RECT 768.505 1111.600 768.675 1111.770 ;
        RECT 768.965 1111.600 769.135 1111.770 ;
        RECT 769.425 1111.600 769.595 1111.770 ;
        RECT 769.885 1111.600 770.055 1111.770 ;
        RECT 770.345 1111.600 770.515 1111.770 ;
        RECT 770.805 1111.600 770.975 1111.770 ;
        RECT 771.265 1111.600 771.435 1111.770 ;
        RECT 771.725 1111.600 771.895 1111.770 ;
        RECT 772.185 1111.600 772.355 1111.770 ;
        RECT 772.645 1111.600 772.815 1111.770 ;
        RECT 773.105 1111.600 773.275 1111.770 ;
        RECT 773.565 1111.600 773.735 1111.770 ;
        RECT 774.025 1111.600 774.195 1111.770 ;
        RECT 774.485 1111.600 774.655 1111.770 ;
        RECT 774.945 1111.600 775.115 1111.770 ;
        RECT 775.405 1111.600 775.575 1111.770 ;
        RECT 775.865 1111.600 776.035 1111.770 ;
        RECT 776.325 1111.600 776.495 1111.770 ;
        RECT 776.785 1111.600 776.955 1111.770 ;
        RECT 777.245 1111.600 777.415 1111.770 ;
        RECT 777.705 1111.600 777.875 1111.770 ;
        RECT 778.165 1111.600 778.335 1111.770 ;
        RECT 778.625 1111.600 778.795 1111.770 ;
        RECT 779.085 1111.600 779.255 1111.770 ;
        RECT 779.545 1111.600 779.715 1111.770 ;
        RECT 780.005 1111.600 780.175 1111.770 ;
        RECT 780.465 1111.600 780.635 1111.770 ;
        RECT 780.925 1111.600 781.095 1111.770 ;
        RECT 781.385 1111.600 781.555 1111.770 ;
        RECT 781.845 1111.600 782.015 1111.770 ;
        RECT 782.305 1111.600 782.475 1111.770 ;
        RECT 782.765 1111.600 782.935 1111.770 ;
        RECT 783.225 1111.600 783.395 1111.770 ;
        RECT 783.685 1111.600 783.855 1111.770 ;
        RECT 784.145 1111.600 784.315 1111.770 ;
        RECT 784.605 1111.600 784.775 1111.770 ;
        RECT 785.065 1111.600 785.235 1111.770 ;
        RECT 785.525 1111.600 785.695 1111.770 ;
        RECT 785.985 1111.600 786.155 1111.770 ;
        RECT 786.445 1111.600 786.615 1111.770 ;
        RECT 786.905 1111.600 787.075 1111.770 ;
        RECT 787.365 1111.600 787.535 1111.770 ;
        RECT 787.825 1111.600 787.995 1111.770 ;
        RECT 788.285 1111.600 788.455 1111.770 ;
        RECT 788.745 1111.600 788.915 1111.770 ;
        RECT 789.205 1111.600 789.375 1111.770 ;
        RECT 789.665 1111.600 789.835 1111.770 ;
        RECT 790.125 1111.600 790.295 1111.770 ;
        RECT 790.585 1111.600 790.755 1111.770 ;
        RECT 791.045 1111.600 791.215 1111.770 ;
        RECT 791.505 1111.600 791.675 1111.770 ;
        RECT 791.965 1111.600 792.135 1111.770 ;
        RECT 792.425 1111.600 792.595 1111.770 ;
        RECT 792.885 1111.600 793.055 1111.770 ;
        RECT 793.345 1111.600 793.515 1111.770 ;
        RECT 793.805 1111.600 793.975 1111.770 ;
        RECT 794.265 1111.600 794.435 1111.770 ;
        RECT 794.725 1111.600 794.895 1111.770 ;
      LAYER met1 ;
        RECT 669.000 1116.885 795.040 1117.365 ;
        RECT 674.980 1111.445 795.040 1111.925 ;
      LAYER via ;
        RECT 736.975 1116.985 738.760 1117.285 ;
        RECT 736.975 1111.575 738.760 1111.875 ;
      LAYER met2 ;
        RECT 736.935 1116.915 738.800 1117.345 ;
        RECT 736.935 1111.490 738.800 1111.920 ;
      LAYER via2 ;
        RECT 736.975 1116.985 738.760 1117.285 ;
        RECT 736.975 1111.575 738.760 1111.875 ;
      LAYER met3 ;
        RECT 736.940 1109.835 738.805 1117.360 ;
    END
    PORT
      LAYER li1 ;
        RECT 1969.145 1117.040 1969.315 1117.210 ;
        RECT 1969.605 1117.040 1969.775 1117.210 ;
        RECT 1970.065 1117.040 1970.235 1117.210 ;
        RECT 1970.525 1117.040 1970.695 1117.210 ;
        RECT 1970.985 1117.040 1971.155 1117.210 ;
        RECT 1971.445 1117.040 1971.615 1117.210 ;
        RECT 1971.905 1117.040 1972.075 1117.210 ;
        RECT 1972.365 1117.040 1972.535 1117.210 ;
        RECT 1972.825 1117.040 1972.995 1117.210 ;
        RECT 1973.285 1117.040 1973.455 1117.210 ;
        RECT 1973.745 1117.040 1973.915 1117.210 ;
        RECT 1974.205 1117.040 1974.375 1117.210 ;
        RECT 1974.665 1117.040 1974.835 1117.210 ;
        RECT 1975.125 1117.040 1975.295 1117.210 ;
        RECT 1975.585 1117.040 1975.755 1117.210 ;
        RECT 1976.045 1117.040 1976.215 1117.210 ;
        RECT 1976.505 1117.040 1976.675 1117.210 ;
        RECT 1976.965 1117.040 1977.135 1117.210 ;
        RECT 1977.425 1117.040 1977.595 1117.210 ;
        RECT 1977.885 1117.040 1978.055 1117.210 ;
        RECT 1978.345 1117.040 1978.515 1117.210 ;
        RECT 1978.805 1117.040 1978.975 1117.210 ;
        RECT 1979.265 1117.040 1979.435 1117.210 ;
        RECT 1979.725 1117.040 1979.895 1117.210 ;
        RECT 1980.185 1117.040 1980.355 1117.210 ;
        RECT 1980.645 1117.040 1980.815 1117.210 ;
        RECT 1981.105 1117.040 1981.275 1117.210 ;
        RECT 1981.565 1117.040 1981.735 1117.210 ;
        RECT 1982.025 1117.040 1982.195 1117.210 ;
        RECT 1982.485 1117.040 1982.655 1117.210 ;
        RECT 1982.945 1117.040 1983.115 1117.210 ;
        RECT 1983.405 1117.040 1983.575 1117.210 ;
        RECT 1983.865 1117.040 1984.035 1117.210 ;
        RECT 1984.325 1117.040 1984.495 1117.210 ;
        RECT 1984.785 1117.040 1984.955 1117.210 ;
        RECT 1985.245 1117.040 1985.415 1117.210 ;
        RECT 1985.705 1117.040 1985.875 1117.210 ;
        RECT 1986.165 1117.040 1986.335 1117.210 ;
        RECT 1986.625 1117.040 1986.795 1117.210 ;
        RECT 1987.085 1117.040 1987.255 1117.210 ;
        RECT 1987.545 1117.040 1987.715 1117.210 ;
        RECT 1988.005 1117.040 1988.175 1117.210 ;
        RECT 1988.465 1117.040 1988.635 1117.210 ;
        RECT 1988.925 1117.040 1989.095 1117.210 ;
        RECT 1989.385 1117.040 1989.555 1117.210 ;
        RECT 1989.845 1117.040 1990.015 1117.210 ;
        RECT 1990.305 1117.040 1990.475 1117.210 ;
        RECT 1990.765 1117.040 1990.935 1117.210 ;
        RECT 1991.225 1117.040 1991.395 1117.210 ;
        RECT 1991.685 1117.040 1991.855 1117.210 ;
        RECT 1992.145 1117.040 1992.315 1117.210 ;
        RECT 1992.605 1117.040 1992.775 1117.210 ;
        RECT 1993.065 1117.040 1993.235 1117.210 ;
        RECT 1993.525 1117.040 1993.695 1117.210 ;
        RECT 1993.985 1117.040 1994.155 1117.210 ;
        RECT 1994.445 1117.040 1994.615 1117.210 ;
        RECT 1994.905 1117.040 1995.075 1117.210 ;
        RECT 1995.365 1117.040 1995.535 1117.210 ;
        RECT 1995.825 1117.040 1995.995 1117.210 ;
        RECT 1996.285 1117.040 1996.455 1117.210 ;
        RECT 1996.745 1117.040 1996.915 1117.210 ;
        RECT 1997.205 1117.040 1997.375 1117.210 ;
        RECT 1997.665 1117.040 1997.835 1117.210 ;
        RECT 1998.125 1117.040 1998.295 1117.210 ;
        RECT 1998.585 1117.040 1998.755 1117.210 ;
        RECT 1999.045 1117.040 1999.215 1117.210 ;
        RECT 1999.505 1117.040 1999.675 1117.210 ;
        RECT 1999.965 1117.040 2000.135 1117.210 ;
        RECT 2000.425 1117.040 2000.595 1117.210 ;
        RECT 2000.885 1117.040 2001.055 1117.210 ;
        RECT 2001.345 1117.040 2001.515 1117.210 ;
        RECT 2001.805 1117.040 2001.975 1117.210 ;
        RECT 2002.265 1117.040 2002.435 1117.210 ;
        RECT 2002.725 1117.040 2002.895 1117.210 ;
        RECT 2003.185 1117.040 2003.355 1117.210 ;
        RECT 2003.645 1117.040 2003.815 1117.210 ;
        RECT 2004.105 1117.040 2004.275 1117.210 ;
        RECT 2004.565 1117.040 2004.735 1117.210 ;
        RECT 2005.025 1117.040 2005.195 1117.210 ;
        RECT 2005.485 1117.040 2005.655 1117.210 ;
        RECT 2005.945 1117.040 2006.115 1117.210 ;
        RECT 2006.405 1117.040 2006.575 1117.210 ;
        RECT 2006.865 1117.040 2007.035 1117.210 ;
        RECT 2007.325 1117.040 2007.495 1117.210 ;
        RECT 2007.785 1117.040 2007.955 1117.210 ;
        RECT 2008.245 1117.040 2008.415 1117.210 ;
        RECT 2008.705 1117.040 2008.875 1117.210 ;
        RECT 2009.165 1117.040 2009.335 1117.210 ;
        RECT 2009.625 1117.040 2009.795 1117.210 ;
        RECT 2010.085 1117.040 2010.255 1117.210 ;
        RECT 2010.545 1117.040 2010.715 1117.210 ;
        RECT 2011.005 1117.040 2011.175 1117.210 ;
        RECT 2011.465 1117.040 2011.635 1117.210 ;
        RECT 2011.925 1117.040 2012.095 1117.210 ;
        RECT 2012.385 1117.040 2012.555 1117.210 ;
        RECT 2012.845 1117.040 2013.015 1117.210 ;
        RECT 2013.305 1117.040 2013.475 1117.210 ;
        RECT 2013.765 1117.040 2013.935 1117.210 ;
        RECT 2014.225 1117.040 2014.395 1117.210 ;
        RECT 2014.685 1117.040 2014.855 1117.210 ;
        RECT 2015.145 1117.040 2015.315 1117.210 ;
        RECT 2015.605 1117.040 2015.775 1117.210 ;
        RECT 2016.065 1117.040 2016.235 1117.210 ;
        RECT 2016.525 1117.040 2016.695 1117.210 ;
        RECT 2016.985 1117.040 2017.155 1117.210 ;
        RECT 2017.445 1117.040 2017.615 1117.210 ;
        RECT 2017.905 1117.040 2018.075 1117.210 ;
        RECT 2018.365 1117.040 2018.535 1117.210 ;
        RECT 2018.825 1117.040 2018.995 1117.210 ;
        RECT 2019.285 1117.040 2019.455 1117.210 ;
        RECT 2019.745 1117.040 2019.915 1117.210 ;
        RECT 2020.205 1117.040 2020.375 1117.210 ;
        RECT 2020.665 1117.040 2020.835 1117.210 ;
        RECT 2021.125 1117.040 2021.295 1117.210 ;
        RECT 2021.585 1117.040 2021.755 1117.210 ;
        RECT 2022.045 1117.040 2022.215 1117.210 ;
        RECT 2022.505 1117.040 2022.675 1117.210 ;
        RECT 2022.965 1117.040 2023.135 1117.210 ;
        RECT 2023.425 1117.040 2023.595 1117.210 ;
        RECT 2023.885 1117.040 2024.055 1117.210 ;
        RECT 2024.345 1117.040 2024.515 1117.210 ;
        RECT 2024.805 1117.040 2024.975 1117.210 ;
        RECT 2025.265 1117.040 2025.435 1117.210 ;
        RECT 2025.725 1117.040 2025.895 1117.210 ;
        RECT 2026.185 1117.040 2026.355 1117.210 ;
        RECT 2026.645 1117.040 2026.815 1117.210 ;
        RECT 2027.105 1117.040 2027.275 1117.210 ;
        RECT 2027.565 1117.040 2027.735 1117.210 ;
        RECT 2028.025 1117.040 2028.195 1117.210 ;
        RECT 2028.485 1117.040 2028.655 1117.210 ;
        RECT 2028.945 1117.040 2029.115 1117.210 ;
        RECT 2029.405 1117.040 2029.575 1117.210 ;
        RECT 2029.865 1117.040 2030.035 1117.210 ;
        RECT 2030.325 1117.040 2030.495 1117.210 ;
        RECT 2030.785 1117.040 2030.955 1117.210 ;
        RECT 2031.245 1117.040 2031.415 1117.210 ;
        RECT 2031.705 1117.040 2031.875 1117.210 ;
        RECT 2032.165 1117.040 2032.335 1117.210 ;
        RECT 2032.625 1117.040 2032.795 1117.210 ;
        RECT 2033.085 1117.040 2033.255 1117.210 ;
        RECT 2033.545 1117.040 2033.715 1117.210 ;
        RECT 2034.005 1117.040 2034.175 1117.210 ;
        RECT 2034.465 1117.040 2034.635 1117.210 ;
        RECT 2034.925 1117.040 2035.095 1117.210 ;
        RECT 2035.385 1117.040 2035.555 1117.210 ;
        RECT 2035.845 1117.040 2036.015 1117.210 ;
        RECT 2036.305 1117.040 2036.475 1117.210 ;
        RECT 2036.765 1117.040 2036.935 1117.210 ;
        RECT 2037.225 1117.040 2037.395 1117.210 ;
        RECT 2037.685 1117.040 2037.855 1117.210 ;
        RECT 2038.145 1117.040 2038.315 1117.210 ;
        RECT 2038.605 1117.040 2038.775 1117.210 ;
        RECT 2039.065 1117.040 2039.235 1117.210 ;
        RECT 2039.525 1117.040 2039.695 1117.210 ;
        RECT 2039.985 1117.040 2040.155 1117.210 ;
        RECT 2040.445 1117.040 2040.615 1117.210 ;
        RECT 2040.905 1117.040 2041.075 1117.210 ;
        RECT 2041.365 1117.040 2041.535 1117.210 ;
        RECT 2041.825 1117.040 2041.995 1117.210 ;
        RECT 2042.285 1117.040 2042.455 1117.210 ;
        RECT 2042.745 1117.040 2042.915 1117.210 ;
        RECT 2043.205 1117.040 2043.375 1117.210 ;
        RECT 2043.665 1117.040 2043.835 1117.210 ;
        RECT 2044.125 1117.040 2044.295 1117.210 ;
        RECT 2044.585 1117.040 2044.755 1117.210 ;
        RECT 2045.045 1117.040 2045.215 1117.210 ;
        RECT 2045.505 1117.040 2045.675 1117.210 ;
        RECT 2045.965 1117.040 2046.135 1117.210 ;
        RECT 2046.425 1117.040 2046.595 1117.210 ;
        RECT 2046.885 1117.040 2047.055 1117.210 ;
        RECT 2047.345 1117.040 2047.515 1117.210 ;
        RECT 2047.805 1117.040 2047.975 1117.210 ;
        RECT 2048.265 1117.040 2048.435 1117.210 ;
        RECT 2048.725 1117.040 2048.895 1117.210 ;
        RECT 2049.185 1117.040 2049.355 1117.210 ;
        RECT 2049.645 1117.040 2049.815 1117.210 ;
        RECT 2050.105 1117.040 2050.275 1117.210 ;
        RECT 2050.565 1117.040 2050.735 1117.210 ;
        RECT 2051.025 1117.040 2051.195 1117.210 ;
        RECT 2051.485 1117.040 2051.655 1117.210 ;
        RECT 2051.945 1117.040 2052.115 1117.210 ;
        RECT 2052.405 1117.040 2052.575 1117.210 ;
        RECT 2052.865 1117.040 2053.035 1117.210 ;
        RECT 2053.325 1117.040 2053.495 1117.210 ;
        RECT 2053.785 1117.040 2053.955 1117.210 ;
        RECT 2054.245 1117.040 2054.415 1117.210 ;
        RECT 2054.705 1117.040 2054.875 1117.210 ;
        RECT 2055.165 1117.040 2055.335 1117.210 ;
        RECT 2055.625 1117.040 2055.795 1117.210 ;
        RECT 2056.085 1117.040 2056.255 1117.210 ;
        RECT 2056.545 1117.040 2056.715 1117.210 ;
        RECT 2057.005 1117.040 2057.175 1117.210 ;
        RECT 2057.465 1117.040 2057.635 1117.210 ;
        RECT 2057.925 1117.040 2058.095 1117.210 ;
        RECT 2058.385 1117.040 2058.555 1117.210 ;
        RECT 2058.845 1117.040 2059.015 1117.210 ;
        RECT 2059.305 1117.040 2059.475 1117.210 ;
        RECT 2059.765 1117.040 2059.935 1117.210 ;
        RECT 2060.225 1117.040 2060.395 1117.210 ;
        RECT 2060.685 1117.040 2060.855 1117.210 ;
        RECT 2061.145 1117.040 2061.315 1117.210 ;
        RECT 2061.605 1117.040 2061.775 1117.210 ;
        RECT 2062.065 1117.040 2062.235 1117.210 ;
        RECT 2062.525 1117.040 2062.695 1117.210 ;
        RECT 2062.985 1117.040 2063.155 1117.210 ;
        RECT 2063.445 1117.040 2063.615 1117.210 ;
        RECT 2063.905 1117.040 2064.075 1117.210 ;
        RECT 2064.365 1117.040 2064.535 1117.210 ;
        RECT 2064.825 1117.040 2064.995 1117.210 ;
        RECT 2065.285 1117.040 2065.455 1117.210 ;
        RECT 2065.745 1117.040 2065.915 1117.210 ;
        RECT 2066.205 1117.040 2066.375 1117.210 ;
        RECT 2066.665 1117.040 2066.835 1117.210 ;
        RECT 2067.125 1117.040 2067.295 1117.210 ;
        RECT 2067.585 1117.040 2067.755 1117.210 ;
        RECT 2068.045 1117.040 2068.215 1117.210 ;
        RECT 2068.505 1117.040 2068.675 1117.210 ;
        RECT 2068.965 1117.040 2069.135 1117.210 ;
        RECT 2069.425 1117.040 2069.595 1117.210 ;
        RECT 2069.885 1117.040 2070.055 1117.210 ;
        RECT 2070.345 1117.040 2070.515 1117.210 ;
        RECT 2070.805 1117.040 2070.975 1117.210 ;
        RECT 2071.265 1117.040 2071.435 1117.210 ;
        RECT 2071.725 1117.040 2071.895 1117.210 ;
        RECT 2072.185 1117.040 2072.355 1117.210 ;
        RECT 2072.645 1117.040 2072.815 1117.210 ;
        RECT 2073.105 1117.040 2073.275 1117.210 ;
        RECT 2073.565 1117.040 2073.735 1117.210 ;
        RECT 2074.025 1117.040 2074.195 1117.210 ;
        RECT 2074.485 1117.040 2074.655 1117.210 ;
        RECT 2074.945 1117.040 2075.115 1117.210 ;
        RECT 2075.405 1117.040 2075.575 1117.210 ;
        RECT 2075.865 1117.040 2076.035 1117.210 ;
        RECT 2076.325 1117.040 2076.495 1117.210 ;
        RECT 2076.785 1117.040 2076.955 1117.210 ;
        RECT 2077.245 1117.040 2077.415 1117.210 ;
        RECT 2077.705 1117.040 2077.875 1117.210 ;
        RECT 2078.165 1117.040 2078.335 1117.210 ;
        RECT 2078.625 1117.040 2078.795 1117.210 ;
        RECT 2079.085 1117.040 2079.255 1117.210 ;
        RECT 2079.545 1117.040 2079.715 1117.210 ;
        RECT 2080.005 1117.040 2080.175 1117.210 ;
        RECT 2080.465 1117.040 2080.635 1117.210 ;
        RECT 2080.925 1117.040 2081.095 1117.210 ;
        RECT 2081.385 1117.040 2081.555 1117.210 ;
        RECT 2081.845 1117.040 2082.015 1117.210 ;
        RECT 2082.305 1117.040 2082.475 1117.210 ;
        RECT 2082.765 1117.040 2082.935 1117.210 ;
        RECT 2083.225 1117.040 2083.395 1117.210 ;
        RECT 2083.685 1117.040 2083.855 1117.210 ;
        RECT 2084.145 1117.040 2084.315 1117.210 ;
        RECT 2084.605 1117.040 2084.775 1117.210 ;
        RECT 2085.065 1117.040 2085.235 1117.210 ;
        RECT 2085.525 1117.040 2085.695 1117.210 ;
        RECT 2085.985 1117.040 2086.155 1117.210 ;
        RECT 2086.445 1117.040 2086.615 1117.210 ;
        RECT 2086.905 1117.040 2087.075 1117.210 ;
        RECT 2087.365 1117.040 2087.535 1117.210 ;
        RECT 2087.825 1117.040 2087.995 1117.210 ;
        RECT 2088.285 1117.040 2088.455 1117.210 ;
        RECT 2088.745 1117.040 2088.915 1117.210 ;
        RECT 2089.205 1117.040 2089.375 1117.210 ;
        RECT 2089.665 1117.040 2089.835 1117.210 ;
        RECT 2090.125 1117.040 2090.295 1117.210 ;
        RECT 2090.585 1117.040 2090.755 1117.210 ;
        RECT 2091.045 1117.040 2091.215 1117.210 ;
        RECT 2091.505 1117.040 2091.675 1117.210 ;
        RECT 2091.965 1117.040 2092.135 1117.210 ;
        RECT 2092.425 1117.040 2092.595 1117.210 ;
        RECT 2092.885 1117.040 2093.055 1117.210 ;
        RECT 2093.345 1117.040 2093.515 1117.210 ;
        RECT 2093.805 1117.040 2093.975 1117.210 ;
        RECT 2094.265 1117.040 2094.435 1117.210 ;
        RECT 2094.725 1117.040 2094.895 1117.210 ;
        RECT 1975.125 1111.600 1975.295 1111.770 ;
        RECT 1975.585 1111.600 1975.755 1111.770 ;
        RECT 1976.045 1111.600 1976.215 1111.770 ;
        RECT 1976.505 1111.600 1976.675 1111.770 ;
        RECT 1976.965 1111.600 1977.135 1111.770 ;
        RECT 1977.425 1111.600 1977.595 1111.770 ;
        RECT 1977.885 1111.600 1978.055 1111.770 ;
        RECT 1978.345 1111.600 1978.515 1111.770 ;
        RECT 1978.805 1111.600 1978.975 1111.770 ;
        RECT 1979.265 1111.600 1979.435 1111.770 ;
        RECT 1979.725 1111.600 1979.895 1111.770 ;
        RECT 1980.185 1111.600 1980.355 1111.770 ;
        RECT 1980.645 1111.600 1980.815 1111.770 ;
        RECT 1981.105 1111.600 1981.275 1111.770 ;
        RECT 1981.565 1111.600 1981.735 1111.770 ;
        RECT 1982.025 1111.600 1982.195 1111.770 ;
        RECT 1982.485 1111.600 1982.655 1111.770 ;
        RECT 1982.945 1111.600 1983.115 1111.770 ;
        RECT 1983.405 1111.600 1983.575 1111.770 ;
        RECT 1983.865 1111.600 1984.035 1111.770 ;
        RECT 1984.325 1111.600 1984.495 1111.770 ;
        RECT 1984.785 1111.600 1984.955 1111.770 ;
        RECT 1985.245 1111.600 1985.415 1111.770 ;
        RECT 1985.705 1111.600 1985.875 1111.770 ;
        RECT 1986.165 1111.600 1986.335 1111.770 ;
        RECT 1986.625 1111.600 1986.795 1111.770 ;
        RECT 1987.085 1111.600 1987.255 1111.770 ;
        RECT 1987.545 1111.600 1987.715 1111.770 ;
        RECT 1988.005 1111.600 1988.175 1111.770 ;
        RECT 1988.465 1111.600 1988.635 1111.770 ;
        RECT 1988.925 1111.600 1989.095 1111.770 ;
        RECT 1989.385 1111.600 1989.555 1111.770 ;
        RECT 1989.845 1111.600 1990.015 1111.770 ;
        RECT 1990.305 1111.600 1990.475 1111.770 ;
        RECT 1990.765 1111.600 1990.935 1111.770 ;
        RECT 1991.225 1111.600 1991.395 1111.770 ;
        RECT 1991.685 1111.600 1991.855 1111.770 ;
        RECT 1992.145 1111.600 1992.315 1111.770 ;
        RECT 1992.605 1111.600 1992.775 1111.770 ;
        RECT 1993.065 1111.600 1993.235 1111.770 ;
        RECT 1993.525 1111.600 1993.695 1111.770 ;
        RECT 1993.985 1111.600 1994.155 1111.770 ;
        RECT 1994.445 1111.600 1994.615 1111.770 ;
        RECT 1994.905 1111.600 1995.075 1111.770 ;
        RECT 1995.365 1111.600 1995.535 1111.770 ;
        RECT 1995.825 1111.600 1995.995 1111.770 ;
        RECT 1996.285 1111.600 1996.455 1111.770 ;
        RECT 1996.745 1111.600 1996.915 1111.770 ;
        RECT 1997.205 1111.600 1997.375 1111.770 ;
        RECT 1997.665 1111.600 1997.835 1111.770 ;
        RECT 1998.125 1111.600 1998.295 1111.770 ;
        RECT 1998.585 1111.600 1998.755 1111.770 ;
        RECT 1999.045 1111.600 1999.215 1111.770 ;
        RECT 1999.505 1111.600 1999.675 1111.770 ;
        RECT 1999.965 1111.600 2000.135 1111.770 ;
        RECT 2000.425 1111.600 2000.595 1111.770 ;
        RECT 2000.885 1111.600 2001.055 1111.770 ;
        RECT 2001.345 1111.600 2001.515 1111.770 ;
        RECT 2001.805 1111.600 2001.975 1111.770 ;
        RECT 2002.265 1111.600 2002.435 1111.770 ;
        RECT 2002.725 1111.600 2002.895 1111.770 ;
        RECT 2003.185 1111.600 2003.355 1111.770 ;
        RECT 2003.645 1111.600 2003.815 1111.770 ;
        RECT 2004.105 1111.600 2004.275 1111.770 ;
        RECT 2004.565 1111.600 2004.735 1111.770 ;
        RECT 2005.025 1111.600 2005.195 1111.770 ;
        RECT 2005.485 1111.600 2005.655 1111.770 ;
        RECT 2005.945 1111.600 2006.115 1111.770 ;
        RECT 2006.405 1111.600 2006.575 1111.770 ;
        RECT 2006.865 1111.600 2007.035 1111.770 ;
        RECT 2007.325 1111.600 2007.495 1111.770 ;
        RECT 2007.785 1111.600 2007.955 1111.770 ;
        RECT 2008.245 1111.600 2008.415 1111.770 ;
        RECT 2008.705 1111.600 2008.875 1111.770 ;
        RECT 2009.165 1111.600 2009.335 1111.770 ;
        RECT 2009.625 1111.600 2009.795 1111.770 ;
        RECT 2010.085 1111.600 2010.255 1111.770 ;
        RECT 2010.545 1111.600 2010.715 1111.770 ;
        RECT 2011.005 1111.600 2011.175 1111.770 ;
        RECT 2011.465 1111.600 2011.635 1111.770 ;
        RECT 2011.925 1111.600 2012.095 1111.770 ;
        RECT 2012.385 1111.600 2012.555 1111.770 ;
        RECT 2012.845 1111.600 2013.015 1111.770 ;
        RECT 2013.305 1111.600 2013.475 1111.770 ;
        RECT 2013.765 1111.600 2013.935 1111.770 ;
        RECT 2014.225 1111.600 2014.395 1111.770 ;
        RECT 2014.685 1111.600 2014.855 1111.770 ;
        RECT 2015.145 1111.600 2015.315 1111.770 ;
        RECT 2015.605 1111.600 2015.775 1111.770 ;
        RECT 2016.065 1111.600 2016.235 1111.770 ;
        RECT 2016.525 1111.600 2016.695 1111.770 ;
        RECT 2016.985 1111.600 2017.155 1111.770 ;
        RECT 2017.445 1111.600 2017.615 1111.770 ;
        RECT 2017.905 1111.600 2018.075 1111.770 ;
        RECT 2018.365 1111.600 2018.535 1111.770 ;
        RECT 2018.825 1111.600 2018.995 1111.770 ;
        RECT 2019.285 1111.600 2019.455 1111.770 ;
        RECT 2019.745 1111.600 2019.915 1111.770 ;
        RECT 2020.205 1111.600 2020.375 1111.770 ;
        RECT 2020.665 1111.600 2020.835 1111.770 ;
        RECT 2021.125 1111.600 2021.295 1111.770 ;
        RECT 2021.585 1111.600 2021.755 1111.770 ;
        RECT 2022.045 1111.600 2022.215 1111.770 ;
        RECT 2022.505 1111.600 2022.675 1111.770 ;
        RECT 2022.965 1111.600 2023.135 1111.770 ;
        RECT 2023.425 1111.600 2023.595 1111.770 ;
        RECT 2023.885 1111.600 2024.055 1111.770 ;
        RECT 2024.345 1111.600 2024.515 1111.770 ;
        RECT 2024.805 1111.600 2024.975 1111.770 ;
        RECT 2025.265 1111.600 2025.435 1111.770 ;
        RECT 2025.725 1111.600 2025.895 1111.770 ;
        RECT 2026.185 1111.600 2026.355 1111.770 ;
        RECT 2026.645 1111.600 2026.815 1111.770 ;
        RECT 2027.105 1111.600 2027.275 1111.770 ;
        RECT 2027.565 1111.600 2027.735 1111.770 ;
        RECT 2028.025 1111.600 2028.195 1111.770 ;
        RECT 2028.485 1111.600 2028.655 1111.770 ;
        RECT 2028.945 1111.600 2029.115 1111.770 ;
        RECT 2029.405 1111.600 2029.575 1111.770 ;
        RECT 2029.865 1111.600 2030.035 1111.770 ;
        RECT 2030.325 1111.600 2030.495 1111.770 ;
        RECT 2030.785 1111.600 2030.955 1111.770 ;
        RECT 2031.245 1111.600 2031.415 1111.770 ;
        RECT 2031.705 1111.600 2031.875 1111.770 ;
        RECT 2032.165 1111.600 2032.335 1111.770 ;
        RECT 2032.625 1111.600 2032.795 1111.770 ;
        RECT 2033.085 1111.600 2033.255 1111.770 ;
        RECT 2033.545 1111.600 2033.715 1111.770 ;
        RECT 2034.005 1111.600 2034.175 1111.770 ;
        RECT 2034.465 1111.600 2034.635 1111.770 ;
        RECT 2034.925 1111.600 2035.095 1111.770 ;
        RECT 2035.385 1111.600 2035.555 1111.770 ;
        RECT 2035.845 1111.600 2036.015 1111.770 ;
        RECT 2036.305 1111.600 2036.475 1111.770 ;
        RECT 2036.765 1111.600 2036.935 1111.770 ;
        RECT 2037.225 1111.600 2037.395 1111.770 ;
        RECT 2037.685 1111.600 2037.855 1111.770 ;
        RECT 2038.145 1111.600 2038.315 1111.770 ;
        RECT 2038.605 1111.600 2038.775 1111.770 ;
        RECT 2039.065 1111.600 2039.235 1111.770 ;
        RECT 2039.525 1111.600 2039.695 1111.770 ;
        RECT 2039.985 1111.600 2040.155 1111.770 ;
        RECT 2040.445 1111.600 2040.615 1111.770 ;
        RECT 2040.905 1111.600 2041.075 1111.770 ;
        RECT 2041.365 1111.600 2041.535 1111.770 ;
        RECT 2041.825 1111.600 2041.995 1111.770 ;
        RECT 2042.285 1111.600 2042.455 1111.770 ;
        RECT 2042.745 1111.600 2042.915 1111.770 ;
        RECT 2043.205 1111.600 2043.375 1111.770 ;
        RECT 2043.665 1111.600 2043.835 1111.770 ;
        RECT 2044.125 1111.600 2044.295 1111.770 ;
        RECT 2044.585 1111.600 2044.755 1111.770 ;
        RECT 2045.045 1111.600 2045.215 1111.770 ;
        RECT 2045.505 1111.600 2045.675 1111.770 ;
        RECT 2045.965 1111.600 2046.135 1111.770 ;
        RECT 2046.425 1111.600 2046.595 1111.770 ;
        RECT 2046.885 1111.600 2047.055 1111.770 ;
        RECT 2047.345 1111.600 2047.515 1111.770 ;
        RECT 2047.805 1111.600 2047.975 1111.770 ;
        RECT 2048.265 1111.600 2048.435 1111.770 ;
        RECT 2048.725 1111.600 2048.895 1111.770 ;
        RECT 2049.185 1111.600 2049.355 1111.770 ;
        RECT 2049.645 1111.600 2049.815 1111.770 ;
        RECT 2050.105 1111.600 2050.275 1111.770 ;
        RECT 2050.565 1111.600 2050.735 1111.770 ;
        RECT 2051.025 1111.600 2051.195 1111.770 ;
        RECT 2051.485 1111.600 2051.655 1111.770 ;
        RECT 2051.945 1111.600 2052.115 1111.770 ;
        RECT 2052.405 1111.600 2052.575 1111.770 ;
        RECT 2052.865 1111.600 2053.035 1111.770 ;
        RECT 2053.325 1111.600 2053.495 1111.770 ;
        RECT 2053.785 1111.600 2053.955 1111.770 ;
        RECT 2054.245 1111.600 2054.415 1111.770 ;
        RECT 2054.705 1111.600 2054.875 1111.770 ;
        RECT 2055.165 1111.600 2055.335 1111.770 ;
        RECT 2055.625 1111.600 2055.795 1111.770 ;
        RECT 2056.085 1111.600 2056.255 1111.770 ;
        RECT 2056.545 1111.600 2056.715 1111.770 ;
        RECT 2057.005 1111.600 2057.175 1111.770 ;
        RECT 2057.465 1111.600 2057.635 1111.770 ;
        RECT 2057.925 1111.600 2058.095 1111.770 ;
        RECT 2058.385 1111.600 2058.555 1111.770 ;
        RECT 2058.845 1111.600 2059.015 1111.770 ;
        RECT 2059.305 1111.600 2059.475 1111.770 ;
        RECT 2059.765 1111.600 2059.935 1111.770 ;
        RECT 2060.225 1111.600 2060.395 1111.770 ;
        RECT 2060.685 1111.600 2060.855 1111.770 ;
        RECT 2061.145 1111.600 2061.315 1111.770 ;
        RECT 2061.605 1111.600 2061.775 1111.770 ;
        RECT 2062.065 1111.600 2062.235 1111.770 ;
        RECT 2062.525 1111.600 2062.695 1111.770 ;
        RECT 2062.985 1111.600 2063.155 1111.770 ;
        RECT 2063.445 1111.600 2063.615 1111.770 ;
        RECT 2063.905 1111.600 2064.075 1111.770 ;
        RECT 2064.365 1111.600 2064.535 1111.770 ;
        RECT 2064.825 1111.600 2064.995 1111.770 ;
        RECT 2065.285 1111.600 2065.455 1111.770 ;
        RECT 2065.745 1111.600 2065.915 1111.770 ;
        RECT 2066.205 1111.600 2066.375 1111.770 ;
        RECT 2066.665 1111.600 2066.835 1111.770 ;
        RECT 2067.125 1111.600 2067.295 1111.770 ;
        RECT 2067.585 1111.600 2067.755 1111.770 ;
        RECT 2068.045 1111.600 2068.215 1111.770 ;
        RECT 2068.505 1111.600 2068.675 1111.770 ;
        RECT 2068.965 1111.600 2069.135 1111.770 ;
        RECT 2069.425 1111.600 2069.595 1111.770 ;
        RECT 2069.885 1111.600 2070.055 1111.770 ;
        RECT 2070.345 1111.600 2070.515 1111.770 ;
        RECT 2070.805 1111.600 2070.975 1111.770 ;
        RECT 2071.265 1111.600 2071.435 1111.770 ;
        RECT 2071.725 1111.600 2071.895 1111.770 ;
        RECT 2072.185 1111.600 2072.355 1111.770 ;
        RECT 2072.645 1111.600 2072.815 1111.770 ;
        RECT 2073.105 1111.600 2073.275 1111.770 ;
        RECT 2073.565 1111.600 2073.735 1111.770 ;
        RECT 2074.025 1111.600 2074.195 1111.770 ;
        RECT 2074.485 1111.600 2074.655 1111.770 ;
        RECT 2074.945 1111.600 2075.115 1111.770 ;
        RECT 2075.405 1111.600 2075.575 1111.770 ;
        RECT 2075.865 1111.600 2076.035 1111.770 ;
        RECT 2076.325 1111.600 2076.495 1111.770 ;
        RECT 2076.785 1111.600 2076.955 1111.770 ;
        RECT 2077.245 1111.600 2077.415 1111.770 ;
        RECT 2077.705 1111.600 2077.875 1111.770 ;
        RECT 2078.165 1111.600 2078.335 1111.770 ;
        RECT 2078.625 1111.600 2078.795 1111.770 ;
        RECT 2079.085 1111.600 2079.255 1111.770 ;
        RECT 2079.545 1111.600 2079.715 1111.770 ;
        RECT 2080.005 1111.600 2080.175 1111.770 ;
        RECT 2080.465 1111.600 2080.635 1111.770 ;
        RECT 2080.925 1111.600 2081.095 1111.770 ;
        RECT 2081.385 1111.600 2081.555 1111.770 ;
        RECT 2081.845 1111.600 2082.015 1111.770 ;
        RECT 2082.305 1111.600 2082.475 1111.770 ;
        RECT 2082.765 1111.600 2082.935 1111.770 ;
        RECT 2083.225 1111.600 2083.395 1111.770 ;
        RECT 2083.685 1111.600 2083.855 1111.770 ;
        RECT 2084.145 1111.600 2084.315 1111.770 ;
        RECT 2084.605 1111.600 2084.775 1111.770 ;
        RECT 2085.065 1111.600 2085.235 1111.770 ;
        RECT 2085.525 1111.600 2085.695 1111.770 ;
        RECT 2085.985 1111.600 2086.155 1111.770 ;
        RECT 2086.445 1111.600 2086.615 1111.770 ;
        RECT 2086.905 1111.600 2087.075 1111.770 ;
        RECT 2087.365 1111.600 2087.535 1111.770 ;
        RECT 2087.825 1111.600 2087.995 1111.770 ;
        RECT 2088.285 1111.600 2088.455 1111.770 ;
        RECT 2088.745 1111.600 2088.915 1111.770 ;
        RECT 2089.205 1111.600 2089.375 1111.770 ;
        RECT 2089.665 1111.600 2089.835 1111.770 ;
        RECT 2090.125 1111.600 2090.295 1111.770 ;
        RECT 2090.585 1111.600 2090.755 1111.770 ;
        RECT 2091.045 1111.600 2091.215 1111.770 ;
        RECT 2091.505 1111.600 2091.675 1111.770 ;
        RECT 2091.965 1111.600 2092.135 1111.770 ;
        RECT 2092.425 1111.600 2092.595 1111.770 ;
        RECT 2092.885 1111.600 2093.055 1111.770 ;
        RECT 2093.345 1111.600 2093.515 1111.770 ;
        RECT 2093.805 1111.600 2093.975 1111.770 ;
        RECT 2094.265 1111.600 2094.435 1111.770 ;
        RECT 2094.725 1111.600 2094.895 1111.770 ;
      LAYER met1 ;
        RECT 1969.000 1116.885 2095.040 1117.365 ;
        RECT 1974.980 1111.445 2095.040 1111.925 ;
      LAYER via ;
        RECT 2031.130 1116.950 2032.915 1117.250 ;
        RECT 2031.130 1111.540 2032.915 1111.840 ;
      LAYER met2 ;
        RECT 2031.090 1116.880 2032.955 1117.310 ;
        RECT 2031.090 1111.455 2032.955 1111.885 ;
      LAYER via2 ;
        RECT 2031.130 1116.950 2032.915 1117.250 ;
        RECT 2031.130 1111.540 2032.915 1111.840 ;
      LAYER met3 ;
        RECT 2031.095 1109.800 2032.960 1117.325 ;
    END
    PORT
      LAYER li1 ;
        RECT 198.795 1762.750 198.965 1762.920 ;
        RECT 204.235 1762.750 204.405 1762.920 ;
        RECT 198.795 1762.290 198.965 1762.460 ;
        RECT 204.235 1762.290 204.405 1762.460 ;
        RECT 198.795 1761.830 198.965 1762.000 ;
        RECT 204.235 1761.830 204.405 1762.000 ;
        RECT 198.795 1761.370 198.965 1761.540 ;
        RECT 204.235 1761.370 204.405 1761.540 ;
        RECT 198.795 1760.910 198.965 1761.080 ;
        RECT 204.235 1760.910 204.405 1761.080 ;
        RECT 198.795 1760.450 198.965 1760.620 ;
        RECT 204.235 1760.450 204.405 1760.620 ;
        RECT 198.795 1759.990 198.965 1760.160 ;
        RECT 204.235 1759.990 204.405 1760.160 ;
        RECT 198.795 1759.530 198.965 1759.700 ;
        RECT 204.235 1759.530 204.405 1759.700 ;
        RECT 198.795 1759.070 198.965 1759.240 ;
        RECT 204.235 1759.070 204.405 1759.240 ;
        RECT 198.795 1758.610 198.965 1758.780 ;
        RECT 204.235 1758.610 204.405 1758.780 ;
        RECT 198.795 1758.150 198.965 1758.320 ;
        RECT 204.235 1758.150 204.405 1758.320 ;
        RECT 198.795 1757.690 198.965 1757.860 ;
        RECT 204.235 1757.690 204.405 1757.860 ;
        RECT 198.795 1757.230 198.965 1757.400 ;
        RECT 204.235 1757.230 204.405 1757.400 ;
        RECT 198.795 1756.770 198.965 1756.940 ;
        RECT 204.235 1756.770 204.405 1756.940 ;
        RECT 198.795 1756.310 198.965 1756.480 ;
        RECT 204.235 1756.310 204.405 1756.480 ;
        RECT 198.795 1755.850 198.965 1756.020 ;
        RECT 204.235 1755.850 204.405 1756.020 ;
        RECT 198.795 1755.390 198.965 1755.560 ;
        RECT 204.235 1755.390 204.405 1755.560 ;
        RECT 198.795 1754.930 198.965 1755.100 ;
        RECT 204.235 1754.930 204.405 1755.100 ;
        RECT 198.795 1754.470 198.965 1754.640 ;
        RECT 204.235 1754.470 204.405 1754.640 ;
        RECT 198.795 1754.010 198.965 1754.180 ;
        RECT 204.235 1754.010 204.405 1754.180 ;
        RECT 198.795 1753.550 198.965 1753.720 ;
        RECT 204.235 1753.550 204.405 1753.720 ;
        RECT 198.795 1753.090 198.965 1753.260 ;
        RECT 204.235 1753.090 204.405 1753.260 ;
        RECT 198.795 1752.630 198.965 1752.800 ;
        RECT 204.235 1752.630 204.405 1752.800 ;
        RECT 198.795 1752.170 198.965 1752.340 ;
        RECT 204.235 1752.170 204.405 1752.340 ;
        RECT 198.795 1751.710 198.965 1751.880 ;
        RECT 204.235 1751.710 204.405 1751.880 ;
        RECT 198.795 1751.250 198.965 1751.420 ;
        RECT 204.235 1751.250 204.405 1751.420 ;
        RECT 198.795 1750.790 198.965 1750.960 ;
        RECT 204.235 1750.790 204.405 1750.960 ;
        RECT 198.795 1750.330 198.965 1750.500 ;
        RECT 204.235 1750.330 204.405 1750.500 ;
        RECT 198.795 1749.870 198.965 1750.040 ;
        RECT 204.235 1749.870 204.405 1750.040 ;
        RECT 198.795 1749.410 198.965 1749.580 ;
        RECT 204.235 1749.410 204.405 1749.580 ;
        RECT 198.795 1748.950 198.965 1749.120 ;
        RECT 204.235 1748.950 204.405 1749.120 ;
        RECT 198.795 1748.490 198.965 1748.660 ;
        RECT 204.235 1748.490 204.405 1748.660 ;
        RECT 198.795 1748.030 198.965 1748.200 ;
        RECT 204.235 1748.030 204.405 1748.200 ;
        RECT 198.795 1747.570 198.965 1747.740 ;
        RECT 204.235 1747.570 204.405 1747.740 ;
        RECT 198.795 1747.110 198.965 1747.280 ;
        RECT 204.235 1747.110 204.405 1747.280 ;
        RECT 198.795 1746.650 198.965 1746.820 ;
        RECT 204.235 1746.650 204.405 1746.820 ;
        RECT 198.795 1746.190 198.965 1746.360 ;
        RECT 204.235 1746.190 204.405 1746.360 ;
        RECT 198.795 1745.730 198.965 1745.900 ;
        RECT 204.235 1745.730 204.405 1745.900 ;
        RECT 198.795 1745.270 198.965 1745.440 ;
        RECT 204.235 1745.270 204.405 1745.440 ;
        RECT 198.795 1744.810 198.965 1744.980 ;
        RECT 204.235 1744.810 204.405 1744.980 ;
        RECT 198.795 1744.350 198.965 1744.520 ;
        RECT 204.235 1744.350 204.405 1744.520 ;
        RECT 198.795 1743.890 198.965 1744.060 ;
        RECT 204.235 1743.890 204.405 1744.060 ;
        RECT 198.795 1743.430 198.965 1743.600 ;
        RECT 204.235 1743.430 204.405 1743.600 ;
        RECT 198.795 1742.970 198.965 1743.140 ;
        RECT 204.235 1742.970 204.405 1743.140 ;
        RECT 198.795 1742.510 198.965 1742.680 ;
        RECT 204.235 1742.510 204.405 1742.680 ;
        RECT 198.795 1742.050 198.965 1742.220 ;
        RECT 204.235 1742.050 204.405 1742.220 ;
        RECT 198.795 1741.590 198.965 1741.760 ;
        RECT 204.235 1741.590 204.405 1741.760 ;
        RECT 198.795 1741.130 198.965 1741.300 ;
        RECT 204.235 1741.130 204.405 1741.300 ;
        RECT 198.795 1740.670 198.965 1740.840 ;
        RECT 204.235 1740.670 204.405 1740.840 ;
        RECT 198.795 1740.210 198.965 1740.380 ;
        RECT 204.235 1740.210 204.405 1740.380 ;
        RECT 198.795 1739.750 198.965 1739.920 ;
        RECT 204.235 1739.750 204.405 1739.920 ;
        RECT 198.795 1739.290 198.965 1739.460 ;
        RECT 204.235 1739.290 204.405 1739.460 ;
        RECT 198.795 1738.830 198.965 1739.000 ;
        RECT 204.235 1738.830 204.405 1739.000 ;
        RECT 198.795 1738.370 198.965 1738.540 ;
        RECT 204.235 1738.370 204.405 1738.540 ;
        RECT 198.795 1737.910 198.965 1738.080 ;
        RECT 204.235 1737.910 204.405 1738.080 ;
        RECT 198.795 1737.450 198.965 1737.620 ;
        RECT 204.235 1737.450 204.405 1737.620 ;
        RECT 198.795 1736.990 198.965 1737.160 ;
        RECT 204.235 1736.990 204.405 1737.160 ;
        RECT 198.795 1736.530 198.965 1736.700 ;
        RECT 204.235 1736.530 204.405 1736.700 ;
        RECT 198.795 1736.070 198.965 1736.240 ;
        RECT 204.235 1736.070 204.405 1736.240 ;
        RECT 198.795 1735.610 198.965 1735.780 ;
        RECT 204.235 1735.610 204.405 1735.780 ;
        RECT 198.795 1735.150 198.965 1735.320 ;
        RECT 204.235 1735.150 204.405 1735.320 ;
        RECT 198.795 1734.690 198.965 1734.860 ;
        RECT 204.235 1734.690 204.405 1734.860 ;
        RECT 198.795 1734.230 198.965 1734.400 ;
        RECT 204.235 1734.230 204.405 1734.400 ;
        RECT 198.795 1733.770 198.965 1733.940 ;
        RECT 204.235 1733.770 204.405 1733.940 ;
        RECT 198.795 1733.310 198.965 1733.480 ;
        RECT 204.235 1733.310 204.405 1733.480 ;
        RECT 198.795 1732.850 198.965 1733.020 ;
        RECT 204.235 1732.850 204.405 1733.020 ;
        RECT 198.795 1732.390 198.965 1732.560 ;
        RECT 204.235 1732.390 204.405 1732.560 ;
        RECT 198.795 1731.930 198.965 1732.100 ;
        RECT 204.235 1731.930 204.405 1732.100 ;
        RECT 198.795 1731.470 198.965 1731.640 ;
        RECT 204.235 1731.470 204.405 1731.640 ;
        RECT 198.795 1731.010 198.965 1731.180 ;
        RECT 204.235 1731.010 204.405 1731.180 ;
        RECT 198.795 1730.550 198.965 1730.720 ;
        RECT 204.235 1730.550 204.405 1730.720 ;
        RECT 198.795 1730.090 198.965 1730.260 ;
        RECT 204.235 1730.090 204.405 1730.260 ;
        RECT 198.795 1729.630 198.965 1729.800 ;
        RECT 204.235 1729.630 204.405 1729.800 ;
        RECT 198.795 1729.170 198.965 1729.340 ;
        RECT 204.235 1729.170 204.405 1729.340 ;
        RECT 198.795 1728.710 198.965 1728.880 ;
        RECT 204.235 1728.710 204.405 1728.880 ;
        RECT 198.795 1728.250 198.965 1728.420 ;
        RECT 204.235 1728.250 204.405 1728.420 ;
        RECT 198.795 1727.790 198.965 1727.960 ;
        RECT 204.235 1727.790 204.405 1727.960 ;
        RECT 198.795 1727.330 198.965 1727.500 ;
        RECT 204.235 1727.330 204.405 1727.500 ;
        RECT 198.795 1726.870 198.965 1727.040 ;
        RECT 204.235 1726.870 204.405 1727.040 ;
        RECT 198.795 1726.410 198.965 1726.580 ;
        RECT 204.235 1726.410 204.405 1726.580 ;
        RECT 198.795 1725.950 198.965 1726.120 ;
        RECT 204.235 1725.950 204.405 1726.120 ;
        RECT 198.795 1725.490 198.965 1725.660 ;
        RECT 204.235 1725.490 204.405 1725.660 ;
        RECT 198.795 1725.030 198.965 1725.200 ;
        RECT 204.235 1725.030 204.405 1725.200 ;
        RECT 198.795 1724.570 198.965 1724.740 ;
        RECT 204.235 1724.570 204.405 1724.740 ;
        RECT 198.795 1724.110 198.965 1724.280 ;
        RECT 204.235 1724.110 204.405 1724.280 ;
        RECT 198.795 1723.650 198.965 1723.820 ;
        RECT 204.235 1723.650 204.405 1723.820 ;
        RECT 198.795 1723.190 198.965 1723.360 ;
        RECT 204.235 1723.190 204.405 1723.360 ;
        RECT 198.795 1722.730 198.965 1722.900 ;
        RECT 204.235 1722.730 204.405 1722.900 ;
        RECT 198.795 1722.270 198.965 1722.440 ;
        RECT 204.235 1722.270 204.405 1722.440 ;
        RECT 198.795 1721.810 198.965 1721.980 ;
        RECT 204.235 1721.810 204.405 1721.980 ;
        RECT 198.795 1721.350 198.965 1721.520 ;
        RECT 204.235 1721.350 204.405 1721.520 ;
        RECT 198.795 1720.890 198.965 1721.060 ;
        RECT 204.235 1720.890 204.405 1721.060 ;
        RECT 198.795 1720.430 198.965 1720.600 ;
        RECT 204.235 1720.430 204.405 1720.600 ;
        RECT 198.795 1719.970 198.965 1720.140 ;
        RECT 204.235 1719.970 204.405 1720.140 ;
        RECT 198.795 1719.510 198.965 1719.680 ;
        RECT 204.235 1719.510 204.405 1719.680 ;
        RECT 198.795 1719.050 198.965 1719.220 ;
        RECT 204.235 1719.050 204.405 1719.220 ;
        RECT 198.795 1718.590 198.965 1718.760 ;
        RECT 204.235 1718.590 204.405 1718.760 ;
        RECT 198.795 1718.130 198.965 1718.300 ;
        RECT 204.235 1718.130 204.405 1718.300 ;
        RECT 198.795 1717.670 198.965 1717.840 ;
        RECT 204.235 1717.670 204.405 1717.840 ;
        RECT 198.795 1717.210 198.965 1717.380 ;
        RECT 204.235 1717.210 204.405 1717.380 ;
        RECT 198.795 1716.750 198.965 1716.920 ;
        RECT 204.235 1716.750 204.405 1716.920 ;
        RECT 198.795 1716.290 198.965 1716.460 ;
        RECT 204.235 1716.290 204.405 1716.460 ;
        RECT 198.795 1715.830 198.965 1716.000 ;
        RECT 204.235 1715.830 204.405 1716.000 ;
        RECT 198.795 1715.370 198.965 1715.540 ;
        RECT 204.235 1715.370 204.405 1715.540 ;
        RECT 198.795 1714.910 198.965 1715.080 ;
        RECT 204.235 1714.910 204.405 1715.080 ;
        RECT 198.795 1714.450 198.965 1714.620 ;
        RECT 204.235 1714.450 204.405 1714.620 ;
        RECT 198.795 1713.990 198.965 1714.160 ;
        RECT 204.235 1713.990 204.405 1714.160 ;
        RECT 198.795 1713.530 198.965 1713.700 ;
        RECT 204.235 1713.530 204.405 1713.700 ;
        RECT 198.795 1713.070 198.965 1713.240 ;
        RECT 204.235 1713.070 204.405 1713.240 ;
        RECT 198.795 1712.610 198.965 1712.780 ;
        RECT 204.235 1712.610 204.405 1712.780 ;
        RECT 198.795 1712.150 198.965 1712.320 ;
        RECT 204.235 1712.150 204.405 1712.320 ;
        RECT 198.795 1711.690 198.965 1711.860 ;
        RECT 204.235 1711.690 204.405 1711.860 ;
        RECT 198.795 1711.230 198.965 1711.400 ;
        RECT 204.235 1711.230 204.405 1711.400 ;
        RECT 198.795 1710.770 198.965 1710.940 ;
        RECT 204.235 1710.770 204.405 1710.940 ;
        RECT 198.795 1710.310 198.965 1710.480 ;
        RECT 204.235 1710.310 204.405 1710.480 ;
        RECT 198.795 1709.850 198.965 1710.020 ;
        RECT 204.235 1709.850 204.405 1710.020 ;
        RECT 198.795 1709.390 198.965 1709.560 ;
        RECT 204.235 1709.390 204.405 1709.560 ;
        RECT 198.795 1708.930 198.965 1709.100 ;
        RECT 204.235 1708.930 204.405 1709.100 ;
        RECT 198.795 1708.470 198.965 1708.640 ;
        RECT 204.235 1708.470 204.405 1708.640 ;
        RECT 198.795 1708.010 198.965 1708.180 ;
        RECT 204.235 1708.010 204.405 1708.180 ;
        RECT 198.795 1707.550 198.965 1707.720 ;
        RECT 204.235 1707.550 204.405 1707.720 ;
        RECT 198.795 1707.090 198.965 1707.260 ;
        RECT 204.235 1707.090 204.405 1707.260 ;
        RECT 198.795 1706.630 198.965 1706.800 ;
        RECT 204.235 1706.630 204.405 1706.800 ;
        RECT 198.795 1706.170 198.965 1706.340 ;
        RECT 204.235 1706.170 204.405 1706.340 ;
        RECT 198.795 1705.710 198.965 1705.880 ;
        RECT 204.235 1705.710 204.405 1705.880 ;
        RECT 198.795 1705.250 198.965 1705.420 ;
        RECT 204.235 1705.250 204.405 1705.420 ;
        RECT 198.795 1704.790 198.965 1704.960 ;
        RECT 204.235 1704.790 204.405 1704.960 ;
        RECT 198.795 1704.330 198.965 1704.500 ;
        RECT 204.235 1704.330 204.405 1704.500 ;
        RECT 198.795 1703.870 198.965 1704.040 ;
        RECT 204.235 1703.870 204.405 1704.040 ;
        RECT 198.795 1703.410 198.965 1703.580 ;
        RECT 204.235 1703.410 204.405 1703.580 ;
        RECT 198.795 1702.950 198.965 1703.120 ;
        RECT 204.235 1702.950 204.405 1703.120 ;
        RECT 198.795 1702.490 198.965 1702.660 ;
        RECT 204.235 1702.490 204.405 1702.660 ;
        RECT 198.795 1702.030 198.965 1702.200 ;
        RECT 204.235 1702.030 204.405 1702.200 ;
        RECT 198.795 1701.570 198.965 1701.740 ;
        RECT 204.235 1701.570 204.405 1701.740 ;
        RECT 198.795 1701.110 198.965 1701.280 ;
        RECT 204.235 1701.110 204.405 1701.280 ;
        RECT 198.795 1700.650 198.965 1700.820 ;
        RECT 204.235 1700.650 204.405 1700.820 ;
        RECT 198.795 1700.190 198.965 1700.360 ;
        RECT 204.235 1700.190 204.405 1700.360 ;
        RECT 198.795 1699.730 198.965 1699.900 ;
        RECT 204.235 1699.730 204.405 1699.900 ;
        RECT 198.795 1699.270 198.965 1699.440 ;
        RECT 204.235 1699.270 204.405 1699.440 ;
        RECT 198.795 1698.810 198.965 1698.980 ;
        RECT 204.235 1698.810 204.405 1698.980 ;
        RECT 198.795 1698.350 198.965 1698.520 ;
        RECT 204.235 1698.350 204.405 1698.520 ;
        RECT 198.795 1697.890 198.965 1698.060 ;
        RECT 204.235 1697.890 204.405 1698.060 ;
        RECT 198.795 1697.430 198.965 1697.600 ;
        RECT 204.235 1697.430 204.405 1697.600 ;
        RECT 198.795 1696.970 198.965 1697.140 ;
        RECT 204.235 1696.970 204.405 1697.140 ;
        RECT 198.795 1696.510 198.965 1696.680 ;
        RECT 204.235 1696.510 204.405 1696.680 ;
        RECT 198.795 1696.050 198.965 1696.220 ;
        RECT 204.235 1696.050 204.405 1696.220 ;
        RECT 198.795 1695.590 198.965 1695.760 ;
        RECT 204.235 1695.590 204.405 1695.760 ;
        RECT 198.795 1695.130 198.965 1695.300 ;
        RECT 204.235 1695.130 204.405 1695.300 ;
        RECT 198.795 1694.670 198.965 1694.840 ;
        RECT 204.235 1694.670 204.405 1694.840 ;
        RECT 198.795 1694.210 198.965 1694.380 ;
        RECT 204.235 1694.210 204.405 1694.380 ;
        RECT 198.795 1693.750 198.965 1693.920 ;
        RECT 204.235 1693.750 204.405 1693.920 ;
        RECT 198.795 1693.290 198.965 1693.460 ;
        RECT 204.235 1693.290 204.405 1693.460 ;
        RECT 198.795 1692.830 198.965 1693.000 ;
        RECT 204.235 1692.830 204.405 1693.000 ;
        RECT 198.795 1692.370 198.965 1692.540 ;
        RECT 204.235 1692.370 204.405 1692.540 ;
        RECT 198.795 1691.910 198.965 1692.080 ;
        RECT 204.235 1691.910 204.405 1692.080 ;
        RECT 198.795 1691.450 198.965 1691.620 ;
        RECT 204.235 1691.450 204.405 1691.620 ;
        RECT 198.795 1690.990 198.965 1691.160 ;
        RECT 204.235 1690.990 204.405 1691.160 ;
        RECT 198.795 1690.530 198.965 1690.700 ;
        RECT 204.235 1690.530 204.405 1690.700 ;
        RECT 198.795 1690.070 198.965 1690.240 ;
        RECT 204.235 1690.070 204.405 1690.240 ;
        RECT 198.795 1689.610 198.965 1689.780 ;
        RECT 204.235 1689.610 204.405 1689.780 ;
        RECT 198.795 1689.150 198.965 1689.320 ;
        RECT 204.235 1689.150 204.405 1689.320 ;
        RECT 198.795 1688.690 198.965 1688.860 ;
        RECT 204.235 1688.690 204.405 1688.860 ;
        RECT 198.795 1688.230 198.965 1688.400 ;
        RECT 204.235 1688.230 204.405 1688.400 ;
        RECT 198.795 1687.770 198.965 1687.940 ;
        RECT 204.235 1687.770 204.405 1687.940 ;
        RECT 198.795 1687.310 198.965 1687.480 ;
        RECT 204.235 1687.310 204.405 1687.480 ;
        RECT 198.795 1686.850 198.965 1687.020 ;
        RECT 204.235 1686.850 204.405 1687.020 ;
        RECT 198.795 1686.390 198.965 1686.560 ;
        RECT 204.235 1686.390 204.405 1686.560 ;
        RECT 198.795 1685.930 198.965 1686.100 ;
        RECT 204.235 1685.930 204.405 1686.100 ;
        RECT 198.795 1685.470 198.965 1685.640 ;
        RECT 204.235 1685.470 204.405 1685.640 ;
        RECT 198.795 1685.010 198.965 1685.180 ;
        RECT 204.235 1685.010 204.405 1685.180 ;
        RECT 198.795 1684.550 198.965 1684.720 ;
        RECT 204.235 1684.550 204.405 1684.720 ;
        RECT 198.795 1684.090 198.965 1684.260 ;
        RECT 204.235 1684.090 204.405 1684.260 ;
        RECT 198.795 1683.630 198.965 1683.800 ;
        RECT 204.235 1683.630 204.405 1683.800 ;
        RECT 198.795 1683.170 198.965 1683.340 ;
        RECT 204.235 1683.170 204.405 1683.340 ;
        RECT 198.795 1682.710 198.965 1682.880 ;
        RECT 204.235 1682.710 204.405 1682.880 ;
        RECT 198.795 1682.250 198.965 1682.420 ;
        RECT 204.235 1682.250 204.405 1682.420 ;
        RECT 198.795 1681.790 198.965 1681.960 ;
        RECT 204.235 1681.790 204.405 1681.960 ;
        RECT 198.795 1681.330 198.965 1681.500 ;
        RECT 204.235 1681.330 204.405 1681.500 ;
        RECT 198.795 1680.870 198.965 1681.040 ;
        RECT 204.235 1680.870 204.405 1681.040 ;
        RECT 198.795 1680.410 198.965 1680.580 ;
        RECT 204.235 1680.410 204.405 1680.580 ;
        RECT 198.795 1679.950 198.965 1680.120 ;
        RECT 204.235 1679.950 204.405 1680.120 ;
        RECT 198.795 1679.490 198.965 1679.660 ;
        RECT 204.235 1679.490 204.405 1679.660 ;
        RECT 198.795 1679.030 198.965 1679.200 ;
        RECT 204.235 1679.030 204.405 1679.200 ;
        RECT 198.795 1678.570 198.965 1678.740 ;
        RECT 204.235 1678.570 204.405 1678.740 ;
        RECT 198.795 1678.110 198.965 1678.280 ;
        RECT 204.235 1678.110 204.405 1678.280 ;
        RECT 198.795 1677.650 198.965 1677.820 ;
        RECT 204.235 1677.650 204.405 1677.820 ;
        RECT 198.795 1677.190 198.965 1677.360 ;
        RECT 204.235 1677.190 204.405 1677.360 ;
        RECT 198.795 1676.730 198.965 1676.900 ;
        RECT 204.235 1676.730 204.405 1676.900 ;
        RECT 198.795 1676.270 198.965 1676.440 ;
        RECT 204.235 1676.270 204.405 1676.440 ;
        RECT 198.795 1675.810 198.965 1675.980 ;
        RECT 204.235 1675.810 204.405 1675.980 ;
        RECT 198.795 1675.350 198.965 1675.520 ;
        RECT 204.235 1675.350 204.405 1675.520 ;
        RECT 198.795 1674.890 198.965 1675.060 ;
        RECT 204.235 1674.890 204.405 1675.060 ;
        RECT 198.795 1674.430 198.965 1674.600 ;
        RECT 204.235 1674.430 204.405 1674.600 ;
        RECT 198.795 1673.970 198.965 1674.140 ;
        RECT 204.235 1673.970 204.405 1674.140 ;
        RECT 198.795 1673.510 198.965 1673.680 ;
        RECT 204.235 1673.510 204.405 1673.680 ;
        RECT 198.795 1673.050 198.965 1673.220 ;
        RECT 204.235 1673.050 204.405 1673.220 ;
      LAYER met1 ;
        RECT 198.640 1672.905 199.120 1763.065 ;
        RECT 204.080 1672.905 204.560 1763.065 ;
      LAYER via ;
        RECT 198.750 1710.875 199.050 1712.660 ;
        RECT 204.160 1710.875 204.460 1712.660 ;
      LAYER met2 ;
        RECT 198.665 1710.835 199.095 1712.700 ;
        RECT 204.090 1710.835 204.520 1712.700 ;
      LAYER via2 ;
        RECT 198.750 1710.875 199.050 1712.660 ;
        RECT 204.160 1710.875 204.460 1712.660 ;
      LAYER met3 ;
        RECT 197.010 1710.830 204.535 1712.695 ;
    END
    PORT
      LAYER li1 ;
        RECT 198.685 3053.655 198.855 3053.825 ;
        RECT 204.125 3053.655 204.295 3053.825 ;
        RECT 198.685 3053.195 198.855 3053.365 ;
        RECT 204.125 3053.195 204.295 3053.365 ;
        RECT 198.685 3052.735 198.855 3052.905 ;
        RECT 204.125 3052.735 204.295 3052.905 ;
        RECT 198.685 3052.275 198.855 3052.445 ;
        RECT 204.125 3052.275 204.295 3052.445 ;
        RECT 198.685 3051.815 198.855 3051.985 ;
        RECT 204.125 3051.815 204.295 3051.985 ;
        RECT 198.685 3051.355 198.855 3051.525 ;
        RECT 204.125 3051.355 204.295 3051.525 ;
        RECT 198.685 3050.895 198.855 3051.065 ;
        RECT 204.125 3050.895 204.295 3051.065 ;
        RECT 198.685 3050.435 198.855 3050.605 ;
        RECT 204.125 3050.435 204.295 3050.605 ;
        RECT 198.685 3049.975 198.855 3050.145 ;
        RECT 204.125 3049.975 204.295 3050.145 ;
        RECT 198.685 3049.515 198.855 3049.685 ;
        RECT 204.125 3049.515 204.295 3049.685 ;
        RECT 198.685 3049.055 198.855 3049.225 ;
        RECT 204.125 3049.055 204.295 3049.225 ;
        RECT 198.685 3048.595 198.855 3048.765 ;
        RECT 204.125 3048.595 204.295 3048.765 ;
        RECT 198.685 3048.135 198.855 3048.305 ;
        RECT 204.125 3048.135 204.295 3048.305 ;
        RECT 198.685 3047.675 198.855 3047.845 ;
        RECT 204.125 3047.675 204.295 3047.845 ;
        RECT 198.685 3047.215 198.855 3047.385 ;
        RECT 204.125 3047.215 204.295 3047.385 ;
        RECT 198.685 3046.755 198.855 3046.925 ;
        RECT 204.125 3046.755 204.295 3046.925 ;
        RECT 198.685 3046.295 198.855 3046.465 ;
        RECT 204.125 3046.295 204.295 3046.465 ;
        RECT 198.685 3045.835 198.855 3046.005 ;
        RECT 204.125 3045.835 204.295 3046.005 ;
        RECT 198.685 3045.375 198.855 3045.545 ;
        RECT 204.125 3045.375 204.295 3045.545 ;
        RECT 198.685 3044.915 198.855 3045.085 ;
        RECT 204.125 3044.915 204.295 3045.085 ;
        RECT 198.685 3044.455 198.855 3044.625 ;
        RECT 204.125 3044.455 204.295 3044.625 ;
        RECT 198.685 3043.995 198.855 3044.165 ;
        RECT 204.125 3043.995 204.295 3044.165 ;
        RECT 198.685 3043.535 198.855 3043.705 ;
        RECT 204.125 3043.535 204.295 3043.705 ;
        RECT 198.685 3043.075 198.855 3043.245 ;
        RECT 204.125 3043.075 204.295 3043.245 ;
        RECT 198.685 3042.615 198.855 3042.785 ;
        RECT 204.125 3042.615 204.295 3042.785 ;
        RECT 198.685 3042.155 198.855 3042.325 ;
        RECT 204.125 3042.155 204.295 3042.325 ;
        RECT 198.685 3041.695 198.855 3041.865 ;
        RECT 204.125 3041.695 204.295 3041.865 ;
        RECT 198.685 3041.235 198.855 3041.405 ;
        RECT 204.125 3041.235 204.295 3041.405 ;
        RECT 198.685 3040.775 198.855 3040.945 ;
        RECT 204.125 3040.775 204.295 3040.945 ;
        RECT 198.685 3040.315 198.855 3040.485 ;
        RECT 204.125 3040.315 204.295 3040.485 ;
        RECT 198.685 3039.855 198.855 3040.025 ;
        RECT 204.125 3039.855 204.295 3040.025 ;
        RECT 198.685 3039.395 198.855 3039.565 ;
        RECT 204.125 3039.395 204.295 3039.565 ;
        RECT 198.685 3038.935 198.855 3039.105 ;
        RECT 204.125 3038.935 204.295 3039.105 ;
        RECT 198.685 3038.475 198.855 3038.645 ;
        RECT 204.125 3038.475 204.295 3038.645 ;
        RECT 198.685 3038.015 198.855 3038.185 ;
        RECT 204.125 3038.015 204.295 3038.185 ;
        RECT 198.685 3037.555 198.855 3037.725 ;
        RECT 204.125 3037.555 204.295 3037.725 ;
        RECT 198.685 3037.095 198.855 3037.265 ;
        RECT 204.125 3037.095 204.295 3037.265 ;
        RECT 198.685 3036.635 198.855 3036.805 ;
        RECT 204.125 3036.635 204.295 3036.805 ;
        RECT 198.685 3036.175 198.855 3036.345 ;
        RECT 204.125 3036.175 204.295 3036.345 ;
        RECT 198.685 3035.715 198.855 3035.885 ;
        RECT 204.125 3035.715 204.295 3035.885 ;
        RECT 198.685 3035.255 198.855 3035.425 ;
        RECT 204.125 3035.255 204.295 3035.425 ;
        RECT 198.685 3034.795 198.855 3034.965 ;
        RECT 204.125 3034.795 204.295 3034.965 ;
        RECT 198.685 3034.335 198.855 3034.505 ;
        RECT 204.125 3034.335 204.295 3034.505 ;
        RECT 198.685 3033.875 198.855 3034.045 ;
        RECT 204.125 3033.875 204.295 3034.045 ;
        RECT 198.685 3033.415 198.855 3033.585 ;
        RECT 204.125 3033.415 204.295 3033.585 ;
        RECT 198.685 3032.955 198.855 3033.125 ;
        RECT 204.125 3032.955 204.295 3033.125 ;
        RECT 198.685 3032.495 198.855 3032.665 ;
        RECT 204.125 3032.495 204.295 3032.665 ;
        RECT 198.685 3032.035 198.855 3032.205 ;
        RECT 204.125 3032.035 204.295 3032.205 ;
        RECT 198.685 3031.575 198.855 3031.745 ;
        RECT 204.125 3031.575 204.295 3031.745 ;
        RECT 198.685 3031.115 198.855 3031.285 ;
        RECT 204.125 3031.115 204.295 3031.285 ;
        RECT 198.685 3030.655 198.855 3030.825 ;
        RECT 204.125 3030.655 204.295 3030.825 ;
        RECT 198.685 3030.195 198.855 3030.365 ;
        RECT 204.125 3030.195 204.295 3030.365 ;
        RECT 198.685 3029.735 198.855 3029.905 ;
        RECT 204.125 3029.735 204.295 3029.905 ;
        RECT 198.685 3029.275 198.855 3029.445 ;
        RECT 204.125 3029.275 204.295 3029.445 ;
        RECT 198.685 3028.815 198.855 3028.985 ;
        RECT 204.125 3028.815 204.295 3028.985 ;
        RECT 198.685 3028.355 198.855 3028.525 ;
        RECT 204.125 3028.355 204.295 3028.525 ;
        RECT 198.685 3027.895 198.855 3028.065 ;
        RECT 204.125 3027.895 204.295 3028.065 ;
        RECT 198.685 3027.435 198.855 3027.605 ;
        RECT 204.125 3027.435 204.295 3027.605 ;
        RECT 198.685 3026.975 198.855 3027.145 ;
        RECT 204.125 3026.975 204.295 3027.145 ;
        RECT 198.685 3026.515 198.855 3026.685 ;
        RECT 204.125 3026.515 204.295 3026.685 ;
        RECT 198.685 3026.055 198.855 3026.225 ;
        RECT 204.125 3026.055 204.295 3026.225 ;
        RECT 198.685 3025.595 198.855 3025.765 ;
        RECT 204.125 3025.595 204.295 3025.765 ;
        RECT 198.685 3025.135 198.855 3025.305 ;
        RECT 204.125 3025.135 204.295 3025.305 ;
        RECT 198.685 3024.675 198.855 3024.845 ;
        RECT 204.125 3024.675 204.295 3024.845 ;
        RECT 198.685 3024.215 198.855 3024.385 ;
        RECT 204.125 3024.215 204.295 3024.385 ;
        RECT 198.685 3023.755 198.855 3023.925 ;
        RECT 204.125 3023.755 204.295 3023.925 ;
        RECT 198.685 3023.295 198.855 3023.465 ;
        RECT 204.125 3023.295 204.295 3023.465 ;
        RECT 198.685 3022.835 198.855 3023.005 ;
        RECT 204.125 3022.835 204.295 3023.005 ;
        RECT 198.685 3022.375 198.855 3022.545 ;
        RECT 204.125 3022.375 204.295 3022.545 ;
        RECT 198.685 3021.915 198.855 3022.085 ;
        RECT 204.125 3021.915 204.295 3022.085 ;
        RECT 198.685 3021.455 198.855 3021.625 ;
        RECT 204.125 3021.455 204.295 3021.625 ;
        RECT 198.685 3020.995 198.855 3021.165 ;
        RECT 204.125 3020.995 204.295 3021.165 ;
        RECT 198.685 3020.535 198.855 3020.705 ;
        RECT 204.125 3020.535 204.295 3020.705 ;
        RECT 198.685 3020.075 198.855 3020.245 ;
        RECT 204.125 3020.075 204.295 3020.245 ;
        RECT 198.685 3019.615 198.855 3019.785 ;
        RECT 204.125 3019.615 204.295 3019.785 ;
        RECT 198.685 3019.155 198.855 3019.325 ;
        RECT 204.125 3019.155 204.295 3019.325 ;
        RECT 198.685 3018.695 198.855 3018.865 ;
        RECT 204.125 3018.695 204.295 3018.865 ;
        RECT 198.685 3018.235 198.855 3018.405 ;
        RECT 204.125 3018.235 204.295 3018.405 ;
        RECT 198.685 3017.775 198.855 3017.945 ;
        RECT 204.125 3017.775 204.295 3017.945 ;
        RECT 198.685 3017.315 198.855 3017.485 ;
        RECT 204.125 3017.315 204.295 3017.485 ;
        RECT 198.685 3016.855 198.855 3017.025 ;
        RECT 204.125 3016.855 204.295 3017.025 ;
        RECT 198.685 3016.395 198.855 3016.565 ;
        RECT 204.125 3016.395 204.295 3016.565 ;
        RECT 198.685 3015.935 198.855 3016.105 ;
        RECT 204.125 3015.935 204.295 3016.105 ;
        RECT 198.685 3015.475 198.855 3015.645 ;
        RECT 204.125 3015.475 204.295 3015.645 ;
        RECT 198.685 3015.015 198.855 3015.185 ;
        RECT 204.125 3015.015 204.295 3015.185 ;
        RECT 198.685 3014.555 198.855 3014.725 ;
        RECT 204.125 3014.555 204.295 3014.725 ;
        RECT 198.685 3014.095 198.855 3014.265 ;
        RECT 204.125 3014.095 204.295 3014.265 ;
        RECT 198.685 3013.635 198.855 3013.805 ;
        RECT 204.125 3013.635 204.295 3013.805 ;
        RECT 198.685 3013.175 198.855 3013.345 ;
        RECT 204.125 3013.175 204.295 3013.345 ;
        RECT 198.685 3012.715 198.855 3012.885 ;
        RECT 204.125 3012.715 204.295 3012.885 ;
        RECT 198.685 3012.255 198.855 3012.425 ;
        RECT 204.125 3012.255 204.295 3012.425 ;
        RECT 198.685 3011.795 198.855 3011.965 ;
        RECT 204.125 3011.795 204.295 3011.965 ;
        RECT 198.685 3011.335 198.855 3011.505 ;
        RECT 204.125 3011.335 204.295 3011.505 ;
        RECT 198.685 3010.875 198.855 3011.045 ;
        RECT 204.125 3010.875 204.295 3011.045 ;
        RECT 198.685 3010.415 198.855 3010.585 ;
        RECT 204.125 3010.415 204.295 3010.585 ;
        RECT 198.685 3009.955 198.855 3010.125 ;
        RECT 204.125 3009.955 204.295 3010.125 ;
        RECT 198.685 3009.495 198.855 3009.665 ;
        RECT 204.125 3009.495 204.295 3009.665 ;
        RECT 198.685 3009.035 198.855 3009.205 ;
        RECT 204.125 3009.035 204.295 3009.205 ;
        RECT 198.685 3008.575 198.855 3008.745 ;
        RECT 204.125 3008.575 204.295 3008.745 ;
        RECT 198.685 3008.115 198.855 3008.285 ;
        RECT 204.125 3008.115 204.295 3008.285 ;
        RECT 198.685 3007.655 198.855 3007.825 ;
        RECT 204.125 3007.655 204.295 3007.825 ;
        RECT 198.685 3007.195 198.855 3007.365 ;
        RECT 204.125 3007.195 204.295 3007.365 ;
        RECT 198.685 3006.735 198.855 3006.905 ;
        RECT 204.125 3006.735 204.295 3006.905 ;
        RECT 198.685 3006.275 198.855 3006.445 ;
        RECT 204.125 3006.275 204.295 3006.445 ;
        RECT 198.685 3005.815 198.855 3005.985 ;
        RECT 204.125 3005.815 204.295 3005.985 ;
        RECT 198.685 3005.355 198.855 3005.525 ;
        RECT 204.125 3005.355 204.295 3005.525 ;
        RECT 198.685 3004.895 198.855 3005.065 ;
        RECT 204.125 3004.895 204.295 3005.065 ;
        RECT 198.685 3004.435 198.855 3004.605 ;
        RECT 204.125 3004.435 204.295 3004.605 ;
        RECT 198.685 3003.975 198.855 3004.145 ;
        RECT 204.125 3003.975 204.295 3004.145 ;
        RECT 198.685 3003.515 198.855 3003.685 ;
        RECT 204.125 3003.515 204.295 3003.685 ;
        RECT 198.685 3003.055 198.855 3003.225 ;
        RECT 204.125 3003.055 204.295 3003.225 ;
        RECT 198.685 3002.595 198.855 3002.765 ;
        RECT 204.125 3002.595 204.295 3002.765 ;
        RECT 198.685 3002.135 198.855 3002.305 ;
        RECT 204.125 3002.135 204.295 3002.305 ;
        RECT 198.685 3001.675 198.855 3001.845 ;
        RECT 204.125 3001.675 204.295 3001.845 ;
        RECT 198.685 3001.215 198.855 3001.385 ;
        RECT 204.125 3001.215 204.295 3001.385 ;
        RECT 198.685 3000.755 198.855 3000.925 ;
        RECT 204.125 3000.755 204.295 3000.925 ;
        RECT 198.685 3000.295 198.855 3000.465 ;
        RECT 204.125 3000.295 204.295 3000.465 ;
        RECT 198.685 2999.835 198.855 3000.005 ;
        RECT 204.125 2999.835 204.295 3000.005 ;
        RECT 198.685 2999.375 198.855 2999.545 ;
        RECT 204.125 2999.375 204.295 2999.545 ;
        RECT 198.685 2998.915 198.855 2999.085 ;
        RECT 204.125 2998.915 204.295 2999.085 ;
        RECT 198.685 2998.455 198.855 2998.625 ;
        RECT 204.125 2998.455 204.295 2998.625 ;
        RECT 198.685 2997.995 198.855 2998.165 ;
        RECT 204.125 2997.995 204.295 2998.165 ;
        RECT 198.685 2997.535 198.855 2997.705 ;
        RECT 204.125 2997.535 204.295 2997.705 ;
        RECT 198.685 2997.075 198.855 2997.245 ;
        RECT 204.125 2997.075 204.295 2997.245 ;
        RECT 198.685 2996.615 198.855 2996.785 ;
        RECT 204.125 2996.615 204.295 2996.785 ;
        RECT 198.685 2996.155 198.855 2996.325 ;
        RECT 204.125 2996.155 204.295 2996.325 ;
        RECT 198.685 2995.695 198.855 2995.865 ;
        RECT 204.125 2995.695 204.295 2995.865 ;
        RECT 198.685 2995.235 198.855 2995.405 ;
        RECT 204.125 2995.235 204.295 2995.405 ;
        RECT 198.685 2994.775 198.855 2994.945 ;
        RECT 204.125 2994.775 204.295 2994.945 ;
        RECT 198.685 2994.315 198.855 2994.485 ;
        RECT 204.125 2994.315 204.295 2994.485 ;
        RECT 198.685 2993.855 198.855 2994.025 ;
        RECT 204.125 2993.855 204.295 2994.025 ;
        RECT 198.685 2993.395 198.855 2993.565 ;
        RECT 204.125 2993.395 204.295 2993.565 ;
        RECT 198.685 2992.935 198.855 2993.105 ;
        RECT 204.125 2992.935 204.295 2993.105 ;
        RECT 198.685 2992.475 198.855 2992.645 ;
        RECT 204.125 2992.475 204.295 2992.645 ;
        RECT 198.685 2992.015 198.855 2992.185 ;
        RECT 204.125 2992.015 204.295 2992.185 ;
        RECT 198.685 2991.555 198.855 2991.725 ;
        RECT 204.125 2991.555 204.295 2991.725 ;
        RECT 198.685 2991.095 198.855 2991.265 ;
        RECT 204.125 2991.095 204.295 2991.265 ;
        RECT 198.685 2990.635 198.855 2990.805 ;
        RECT 204.125 2990.635 204.295 2990.805 ;
        RECT 198.685 2990.175 198.855 2990.345 ;
        RECT 204.125 2990.175 204.295 2990.345 ;
        RECT 198.685 2989.715 198.855 2989.885 ;
        RECT 204.125 2989.715 204.295 2989.885 ;
        RECT 198.685 2989.255 198.855 2989.425 ;
        RECT 204.125 2989.255 204.295 2989.425 ;
        RECT 198.685 2988.795 198.855 2988.965 ;
        RECT 204.125 2988.795 204.295 2988.965 ;
        RECT 198.685 2988.335 198.855 2988.505 ;
        RECT 204.125 2988.335 204.295 2988.505 ;
        RECT 198.685 2987.875 198.855 2988.045 ;
        RECT 204.125 2987.875 204.295 2988.045 ;
      LAYER met1 ;
        RECT 198.530 2987.730 199.010 3053.970 ;
        RECT 203.970 2987.730 204.450 3053.970 ;
      LAYER via ;
        RECT 198.655 3020.070 198.955 3021.855 ;
        RECT 204.065 3020.070 204.365 3021.855 ;
      LAYER met2 ;
        RECT 198.570 3020.030 199.000 3021.895 ;
        RECT 203.995 3020.030 204.425 3021.895 ;
      LAYER via2 ;
        RECT 198.655 3020.070 198.955 3021.855 ;
        RECT 204.065 3020.070 204.365 3021.855 ;
      LAYER met3 ;
        RECT 196.915 3020.025 204.440 3021.890 ;
    END
    PORT
      LAYER li1 ;
        RECT 198.560 4456.885 198.730 4457.055 ;
        RECT 204.000 4456.885 204.170 4457.055 ;
        RECT 198.560 4456.425 198.730 4456.595 ;
        RECT 204.000 4456.425 204.170 4456.595 ;
        RECT 198.560 4455.965 198.730 4456.135 ;
        RECT 204.000 4455.965 204.170 4456.135 ;
        RECT 198.560 4455.505 198.730 4455.675 ;
        RECT 204.000 4455.505 204.170 4455.675 ;
        RECT 198.560 4455.045 198.730 4455.215 ;
        RECT 204.000 4455.045 204.170 4455.215 ;
        RECT 198.560 4454.585 198.730 4454.755 ;
        RECT 204.000 4454.585 204.170 4454.755 ;
        RECT 198.560 4454.125 198.730 4454.295 ;
        RECT 204.000 4454.125 204.170 4454.295 ;
        RECT 198.560 4453.665 198.730 4453.835 ;
        RECT 204.000 4453.665 204.170 4453.835 ;
        RECT 198.560 4453.205 198.730 4453.375 ;
        RECT 204.000 4453.205 204.170 4453.375 ;
        RECT 198.560 4452.745 198.730 4452.915 ;
        RECT 204.000 4452.745 204.170 4452.915 ;
        RECT 198.560 4452.285 198.730 4452.455 ;
        RECT 204.000 4452.285 204.170 4452.455 ;
        RECT 198.560 4451.825 198.730 4451.995 ;
        RECT 204.000 4451.825 204.170 4451.995 ;
        RECT 198.560 4451.365 198.730 4451.535 ;
        RECT 204.000 4451.365 204.170 4451.535 ;
        RECT 198.560 4450.905 198.730 4451.075 ;
        RECT 204.000 4450.905 204.170 4451.075 ;
        RECT 198.560 4450.445 198.730 4450.615 ;
        RECT 204.000 4450.445 204.170 4450.615 ;
        RECT 198.560 4449.985 198.730 4450.155 ;
        RECT 204.000 4449.985 204.170 4450.155 ;
        RECT 198.560 4449.525 198.730 4449.695 ;
        RECT 204.000 4449.525 204.170 4449.695 ;
        RECT 198.560 4449.065 198.730 4449.235 ;
        RECT 204.000 4449.065 204.170 4449.235 ;
        RECT 198.560 4448.605 198.730 4448.775 ;
        RECT 204.000 4448.605 204.170 4448.775 ;
        RECT 198.560 4448.145 198.730 4448.315 ;
        RECT 204.000 4448.145 204.170 4448.315 ;
        RECT 198.560 4447.685 198.730 4447.855 ;
        RECT 204.000 4447.685 204.170 4447.855 ;
        RECT 198.560 4447.225 198.730 4447.395 ;
        RECT 204.000 4447.225 204.170 4447.395 ;
        RECT 198.560 4446.765 198.730 4446.935 ;
        RECT 204.000 4446.765 204.170 4446.935 ;
        RECT 198.560 4446.305 198.730 4446.475 ;
        RECT 204.000 4446.305 204.170 4446.475 ;
        RECT 198.560 4445.845 198.730 4446.015 ;
        RECT 204.000 4445.845 204.170 4446.015 ;
        RECT 198.560 4445.385 198.730 4445.555 ;
        RECT 204.000 4445.385 204.170 4445.555 ;
        RECT 198.560 4444.925 198.730 4445.095 ;
        RECT 204.000 4444.925 204.170 4445.095 ;
        RECT 198.560 4444.465 198.730 4444.635 ;
        RECT 204.000 4444.465 204.170 4444.635 ;
        RECT 198.560 4444.005 198.730 4444.175 ;
        RECT 204.000 4444.005 204.170 4444.175 ;
        RECT 198.560 4443.545 198.730 4443.715 ;
        RECT 204.000 4443.545 204.170 4443.715 ;
        RECT 198.560 4443.085 198.730 4443.255 ;
        RECT 204.000 4443.085 204.170 4443.255 ;
        RECT 198.560 4442.625 198.730 4442.795 ;
        RECT 204.000 4442.625 204.170 4442.795 ;
        RECT 198.560 4442.165 198.730 4442.335 ;
        RECT 204.000 4442.165 204.170 4442.335 ;
        RECT 198.560 4441.705 198.730 4441.875 ;
        RECT 204.000 4441.705 204.170 4441.875 ;
        RECT 198.560 4441.245 198.730 4441.415 ;
        RECT 204.000 4441.245 204.170 4441.415 ;
        RECT 198.560 4440.785 198.730 4440.955 ;
        RECT 204.000 4440.785 204.170 4440.955 ;
        RECT 198.560 4440.325 198.730 4440.495 ;
        RECT 204.000 4440.325 204.170 4440.495 ;
        RECT 198.560 4439.865 198.730 4440.035 ;
        RECT 204.000 4439.865 204.170 4440.035 ;
        RECT 198.560 4439.405 198.730 4439.575 ;
        RECT 204.000 4439.405 204.170 4439.575 ;
        RECT 198.560 4438.945 198.730 4439.115 ;
        RECT 204.000 4438.945 204.170 4439.115 ;
        RECT 198.560 4438.485 198.730 4438.655 ;
        RECT 204.000 4438.485 204.170 4438.655 ;
        RECT 198.560 4438.025 198.730 4438.195 ;
        RECT 204.000 4438.025 204.170 4438.195 ;
        RECT 198.560 4437.565 198.730 4437.735 ;
        RECT 204.000 4437.565 204.170 4437.735 ;
        RECT 198.560 4437.105 198.730 4437.275 ;
        RECT 204.000 4437.105 204.170 4437.275 ;
        RECT 198.560 4436.645 198.730 4436.815 ;
        RECT 204.000 4436.645 204.170 4436.815 ;
        RECT 198.560 4436.185 198.730 4436.355 ;
        RECT 204.000 4436.185 204.170 4436.355 ;
        RECT 198.560 4435.725 198.730 4435.895 ;
        RECT 204.000 4435.725 204.170 4435.895 ;
        RECT 198.560 4435.265 198.730 4435.435 ;
        RECT 204.000 4435.265 204.170 4435.435 ;
        RECT 198.560 4434.805 198.730 4434.975 ;
        RECT 204.000 4434.805 204.170 4434.975 ;
        RECT 198.560 4434.345 198.730 4434.515 ;
        RECT 204.000 4434.345 204.170 4434.515 ;
        RECT 198.560 4433.885 198.730 4434.055 ;
        RECT 204.000 4433.885 204.170 4434.055 ;
        RECT 198.560 4433.425 198.730 4433.595 ;
        RECT 204.000 4433.425 204.170 4433.595 ;
        RECT 198.560 4432.965 198.730 4433.135 ;
        RECT 204.000 4432.965 204.170 4433.135 ;
        RECT 198.560 4432.505 198.730 4432.675 ;
        RECT 204.000 4432.505 204.170 4432.675 ;
        RECT 198.560 4432.045 198.730 4432.215 ;
        RECT 204.000 4432.045 204.170 4432.215 ;
        RECT 198.560 4431.585 198.730 4431.755 ;
        RECT 204.000 4431.585 204.170 4431.755 ;
        RECT 198.560 4431.125 198.730 4431.295 ;
        RECT 204.000 4431.125 204.170 4431.295 ;
        RECT 198.560 4430.665 198.730 4430.835 ;
        RECT 204.000 4430.665 204.170 4430.835 ;
        RECT 198.560 4430.205 198.730 4430.375 ;
        RECT 204.000 4430.205 204.170 4430.375 ;
        RECT 198.560 4429.745 198.730 4429.915 ;
        RECT 204.000 4429.745 204.170 4429.915 ;
        RECT 198.560 4429.285 198.730 4429.455 ;
        RECT 204.000 4429.285 204.170 4429.455 ;
        RECT 198.560 4428.825 198.730 4428.995 ;
        RECT 204.000 4428.825 204.170 4428.995 ;
        RECT 198.560 4428.365 198.730 4428.535 ;
        RECT 204.000 4428.365 204.170 4428.535 ;
        RECT 198.560 4427.905 198.730 4428.075 ;
        RECT 204.000 4427.905 204.170 4428.075 ;
        RECT 198.560 4427.445 198.730 4427.615 ;
        RECT 204.000 4427.445 204.170 4427.615 ;
        RECT 198.560 4426.985 198.730 4427.155 ;
        RECT 204.000 4426.985 204.170 4427.155 ;
      LAYER met1 ;
        RECT 198.405 4426.840 198.885 4457.200 ;
        RECT 203.845 4426.840 204.325 4457.200 ;
      LAYER via ;
        RECT 198.500 4440.940 198.800 4442.725 ;
        RECT 203.910 4440.940 204.210 4442.725 ;
      LAYER met2 ;
        RECT 198.415 4440.900 198.845 4442.765 ;
        RECT 203.840 4440.900 204.270 4442.765 ;
      LAYER via2 ;
        RECT 198.500 4440.940 198.800 4442.725 ;
        RECT 203.910 4440.940 204.210 4442.725 ;
      LAYER met3 ;
        RECT 196.760 4440.895 204.285 4442.760 ;
    END
    PORT
      LAYER li1 ;
        RECT 3383.500 3572.085 3383.670 3572.255 ;
        RECT 3388.940 3572.085 3389.110 3572.255 ;
        RECT 3383.500 3571.625 3383.670 3571.795 ;
        RECT 3388.940 3571.625 3389.110 3571.795 ;
        RECT 3383.500 3571.165 3383.670 3571.335 ;
        RECT 3388.940 3571.165 3389.110 3571.335 ;
        RECT 3383.500 3570.705 3383.670 3570.875 ;
        RECT 3388.940 3570.705 3389.110 3570.875 ;
        RECT 3383.500 3570.245 3383.670 3570.415 ;
        RECT 3388.940 3570.245 3389.110 3570.415 ;
        RECT 3383.500 3569.785 3383.670 3569.955 ;
        RECT 3388.940 3569.785 3389.110 3569.955 ;
        RECT 3383.500 3569.325 3383.670 3569.495 ;
        RECT 3388.940 3569.325 3389.110 3569.495 ;
        RECT 3383.500 3568.865 3383.670 3569.035 ;
        RECT 3388.940 3568.865 3389.110 3569.035 ;
        RECT 3383.500 3568.405 3383.670 3568.575 ;
        RECT 3388.940 3568.405 3389.110 3568.575 ;
        RECT 3383.500 3567.945 3383.670 3568.115 ;
        RECT 3388.940 3567.945 3389.110 3568.115 ;
        RECT 3383.500 3567.485 3383.670 3567.655 ;
        RECT 3388.940 3567.485 3389.110 3567.655 ;
        RECT 3383.500 3567.025 3383.670 3567.195 ;
        RECT 3388.940 3567.025 3389.110 3567.195 ;
        RECT 3383.500 3566.565 3383.670 3566.735 ;
        RECT 3388.940 3566.565 3389.110 3566.735 ;
        RECT 3383.500 3566.105 3383.670 3566.275 ;
        RECT 3388.940 3566.105 3389.110 3566.275 ;
        RECT 3383.500 3565.645 3383.670 3565.815 ;
        RECT 3388.940 3565.645 3389.110 3565.815 ;
        RECT 3383.500 3565.185 3383.670 3565.355 ;
        RECT 3388.940 3565.185 3389.110 3565.355 ;
        RECT 3383.500 3564.725 3383.670 3564.895 ;
        RECT 3388.940 3564.725 3389.110 3564.895 ;
        RECT 3383.500 3564.265 3383.670 3564.435 ;
        RECT 3388.940 3564.265 3389.110 3564.435 ;
        RECT 3383.500 3563.805 3383.670 3563.975 ;
        RECT 3388.940 3563.805 3389.110 3563.975 ;
        RECT 3383.500 3563.345 3383.670 3563.515 ;
        RECT 3388.940 3563.345 3389.110 3563.515 ;
        RECT 3383.500 3562.885 3383.670 3563.055 ;
        RECT 3388.940 3562.885 3389.110 3563.055 ;
        RECT 3383.500 3562.425 3383.670 3562.595 ;
        RECT 3388.940 3562.425 3389.110 3562.595 ;
        RECT 3383.500 3561.965 3383.670 3562.135 ;
        RECT 3388.940 3561.965 3389.110 3562.135 ;
        RECT 3383.500 3561.505 3383.670 3561.675 ;
        RECT 3388.940 3561.505 3389.110 3561.675 ;
        RECT 3383.500 3561.045 3383.670 3561.215 ;
        RECT 3388.940 3561.045 3389.110 3561.215 ;
        RECT 3383.500 3560.585 3383.670 3560.755 ;
        RECT 3388.940 3560.585 3389.110 3560.755 ;
        RECT 3383.500 3560.125 3383.670 3560.295 ;
        RECT 3388.940 3560.125 3389.110 3560.295 ;
        RECT 3383.500 3559.665 3383.670 3559.835 ;
        RECT 3388.940 3559.665 3389.110 3559.835 ;
        RECT 3383.500 3559.205 3383.670 3559.375 ;
        RECT 3388.940 3559.205 3389.110 3559.375 ;
        RECT 3383.500 3558.745 3383.670 3558.915 ;
        RECT 3388.940 3558.745 3389.110 3558.915 ;
        RECT 3383.500 3558.285 3383.670 3558.455 ;
        RECT 3388.940 3558.285 3389.110 3558.455 ;
        RECT 3383.500 3557.825 3383.670 3557.995 ;
        RECT 3388.940 3557.825 3389.110 3557.995 ;
        RECT 3383.500 3557.365 3383.670 3557.535 ;
        RECT 3388.940 3557.365 3389.110 3557.535 ;
        RECT 3383.500 3556.905 3383.670 3557.075 ;
        RECT 3388.940 3556.905 3389.110 3557.075 ;
        RECT 3383.500 3556.445 3383.670 3556.615 ;
        RECT 3388.940 3556.445 3389.110 3556.615 ;
        RECT 3383.500 3555.985 3383.670 3556.155 ;
        RECT 3388.940 3555.985 3389.110 3556.155 ;
        RECT 3383.500 3555.525 3383.670 3555.695 ;
        RECT 3388.940 3555.525 3389.110 3555.695 ;
        RECT 3383.500 3555.065 3383.670 3555.235 ;
        RECT 3388.940 3555.065 3389.110 3555.235 ;
        RECT 3383.500 3554.605 3383.670 3554.775 ;
        RECT 3388.940 3554.605 3389.110 3554.775 ;
        RECT 3383.500 3554.145 3383.670 3554.315 ;
        RECT 3388.940 3554.145 3389.110 3554.315 ;
        RECT 3383.500 3553.685 3383.670 3553.855 ;
        RECT 3388.940 3553.685 3389.110 3553.855 ;
        RECT 3383.500 3553.225 3383.670 3553.395 ;
        RECT 3388.940 3553.225 3389.110 3553.395 ;
        RECT 3383.500 3552.765 3383.670 3552.935 ;
        RECT 3388.940 3552.765 3389.110 3552.935 ;
        RECT 3383.500 3552.305 3383.670 3552.475 ;
        RECT 3388.940 3552.305 3389.110 3552.475 ;
        RECT 3383.500 3551.845 3383.670 3552.015 ;
        RECT 3388.940 3551.845 3389.110 3552.015 ;
        RECT 3383.500 3551.385 3383.670 3551.555 ;
        RECT 3388.940 3551.385 3389.110 3551.555 ;
        RECT 3383.500 3550.925 3383.670 3551.095 ;
        RECT 3388.940 3550.925 3389.110 3551.095 ;
        RECT 3383.500 3550.465 3383.670 3550.635 ;
        RECT 3388.940 3550.465 3389.110 3550.635 ;
        RECT 3383.500 3550.005 3383.670 3550.175 ;
        RECT 3388.940 3550.005 3389.110 3550.175 ;
        RECT 3383.500 3549.545 3383.670 3549.715 ;
        RECT 3388.940 3549.545 3389.110 3549.715 ;
        RECT 3383.500 3549.085 3383.670 3549.255 ;
        RECT 3388.940 3549.085 3389.110 3549.255 ;
        RECT 3383.500 3548.625 3383.670 3548.795 ;
        RECT 3388.940 3548.625 3389.110 3548.795 ;
        RECT 3383.500 3548.165 3383.670 3548.335 ;
        RECT 3388.940 3548.165 3389.110 3548.335 ;
        RECT 3383.500 3547.705 3383.670 3547.875 ;
        RECT 3388.940 3547.705 3389.110 3547.875 ;
        RECT 3383.500 3547.245 3383.670 3547.415 ;
        RECT 3388.940 3547.245 3389.110 3547.415 ;
        RECT 3383.500 3546.785 3383.670 3546.955 ;
        RECT 3388.940 3546.785 3389.110 3546.955 ;
        RECT 3383.500 3546.325 3383.670 3546.495 ;
        RECT 3388.940 3546.325 3389.110 3546.495 ;
        RECT 3383.500 3545.865 3383.670 3546.035 ;
        RECT 3388.940 3545.865 3389.110 3546.035 ;
        RECT 3383.500 3545.405 3383.670 3545.575 ;
        RECT 3388.940 3545.405 3389.110 3545.575 ;
        RECT 3383.500 3544.945 3383.670 3545.115 ;
        RECT 3388.940 3544.945 3389.110 3545.115 ;
        RECT 3383.500 3544.485 3383.670 3544.655 ;
        RECT 3388.940 3544.485 3389.110 3544.655 ;
        RECT 3383.500 3544.025 3383.670 3544.195 ;
        RECT 3388.940 3544.025 3389.110 3544.195 ;
        RECT 3383.500 3543.565 3383.670 3543.735 ;
        RECT 3388.940 3543.565 3389.110 3543.735 ;
        RECT 3383.500 3543.105 3383.670 3543.275 ;
        RECT 3388.940 3543.105 3389.110 3543.275 ;
        RECT 3383.500 3542.645 3383.670 3542.815 ;
        RECT 3388.940 3542.645 3389.110 3542.815 ;
        RECT 3383.500 3542.185 3383.670 3542.355 ;
        RECT 3388.940 3542.185 3389.110 3542.355 ;
        RECT 3383.500 3541.725 3383.670 3541.895 ;
        RECT 3388.940 3541.725 3389.110 3541.895 ;
        RECT 3383.500 3541.265 3383.670 3541.435 ;
        RECT 3388.940 3541.265 3389.110 3541.435 ;
        RECT 3383.500 3540.805 3383.670 3540.975 ;
        RECT 3388.940 3540.805 3389.110 3540.975 ;
        RECT 3383.500 3540.345 3383.670 3540.515 ;
        RECT 3388.940 3540.345 3389.110 3540.515 ;
        RECT 3383.500 3539.885 3383.670 3540.055 ;
        RECT 3388.940 3539.885 3389.110 3540.055 ;
        RECT 3383.500 3539.425 3383.670 3539.595 ;
        RECT 3388.940 3539.425 3389.110 3539.595 ;
        RECT 3383.500 3538.965 3383.670 3539.135 ;
        RECT 3388.940 3538.965 3389.110 3539.135 ;
        RECT 3383.500 3538.505 3383.670 3538.675 ;
        RECT 3388.940 3538.505 3389.110 3538.675 ;
        RECT 3383.500 3538.045 3383.670 3538.215 ;
        RECT 3388.940 3538.045 3389.110 3538.215 ;
        RECT 3383.500 3537.585 3383.670 3537.755 ;
        RECT 3388.940 3537.585 3389.110 3537.755 ;
        RECT 3383.500 3537.125 3383.670 3537.295 ;
        RECT 3388.940 3537.125 3389.110 3537.295 ;
        RECT 3383.500 3536.665 3383.670 3536.835 ;
        RECT 3388.940 3536.665 3389.110 3536.835 ;
        RECT 3383.500 3536.205 3383.670 3536.375 ;
        RECT 3388.940 3536.205 3389.110 3536.375 ;
      LAYER met1 ;
        RECT 3383.345 3536.060 3383.825 3572.400 ;
        RECT 3388.785 3536.060 3389.265 3572.400 ;
      LAYER via ;
        RECT 3383.465 3556.480 3383.765 3558.265 ;
        RECT 3388.875 3556.480 3389.175 3558.265 ;
      LAYER met2 ;
        RECT 3383.405 3556.440 3383.835 3558.305 ;
        RECT 3388.830 3556.440 3389.260 3558.305 ;
      LAYER via2 ;
        RECT 3383.465 3556.480 3383.765 3558.265 ;
        RECT 3388.875 3556.480 3389.175 3558.265 ;
      LAYER met3 ;
        RECT 3383.390 3556.445 3390.915 3558.310 ;
    END
    PORT
      LAYER li1 ;
        RECT 3383.500 2267.965 3383.670 2268.135 ;
        RECT 3388.940 2267.965 3389.110 2268.135 ;
        RECT 3383.500 2267.505 3383.670 2267.675 ;
        RECT 3388.940 2267.505 3389.110 2267.675 ;
        RECT 3383.500 2267.045 3383.670 2267.215 ;
        RECT 3388.940 2267.045 3389.110 2267.215 ;
        RECT 3383.500 2266.585 3383.670 2266.755 ;
        RECT 3388.940 2266.585 3389.110 2266.755 ;
        RECT 3383.500 2266.125 3383.670 2266.295 ;
        RECT 3388.940 2266.125 3389.110 2266.295 ;
        RECT 3383.500 2265.665 3383.670 2265.835 ;
        RECT 3388.940 2265.665 3389.110 2265.835 ;
        RECT 3383.500 2265.205 3383.670 2265.375 ;
        RECT 3388.940 2265.205 3389.110 2265.375 ;
        RECT 3383.500 2264.745 3383.670 2264.915 ;
        RECT 3388.940 2264.745 3389.110 2264.915 ;
        RECT 3383.500 2264.285 3383.670 2264.455 ;
        RECT 3388.940 2264.285 3389.110 2264.455 ;
        RECT 3383.500 2263.825 3383.670 2263.995 ;
        RECT 3388.940 2263.825 3389.110 2263.995 ;
        RECT 3383.500 2263.365 3383.670 2263.535 ;
        RECT 3388.940 2263.365 3389.110 2263.535 ;
        RECT 3383.500 2262.905 3383.670 2263.075 ;
        RECT 3388.940 2262.905 3389.110 2263.075 ;
        RECT 3383.500 2262.445 3383.670 2262.615 ;
        RECT 3388.940 2262.445 3389.110 2262.615 ;
        RECT 3383.500 2261.985 3383.670 2262.155 ;
        RECT 3388.940 2261.985 3389.110 2262.155 ;
        RECT 3383.500 2261.525 3383.670 2261.695 ;
        RECT 3388.940 2261.525 3389.110 2261.695 ;
        RECT 3383.500 2261.065 3383.670 2261.235 ;
        RECT 3388.940 2261.065 3389.110 2261.235 ;
        RECT 3383.500 2260.605 3383.670 2260.775 ;
        RECT 3388.940 2260.605 3389.110 2260.775 ;
        RECT 3383.500 2260.145 3383.670 2260.315 ;
        RECT 3388.940 2260.145 3389.110 2260.315 ;
        RECT 3383.500 2259.685 3383.670 2259.855 ;
        RECT 3388.940 2259.685 3389.110 2259.855 ;
        RECT 3383.500 2259.225 3383.670 2259.395 ;
        RECT 3388.940 2259.225 3389.110 2259.395 ;
        RECT 3383.500 2258.765 3383.670 2258.935 ;
        RECT 3388.940 2258.765 3389.110 2258.935 ;
        RECT 3383.500 2258.305 3383.670 2258.475 ;
        RECT 3388.940 2258.305 3389.110 2258.475 ;
        RECT 3383.500 2257.845 3383.670 2258.015 ;
        RECT 3388.940 2257.845 3389.110 2258.015 ;
        RECT 3383.500 2257.385 3383.670 2257.555 ;
        RECT 3388.940 2257.385 3389.110 2257.555 ;
        RECT 3383.500 2256.925 3383.670 2257.095 ;
        RECT 3388.940 2256.925 3389.110 2257.095 ;
        RECT 3383.500 2256.465 3383.670 2256.635 ;
        RECT 3388.940 2256.465 3389.110 2256.635 ;
        RECT 3383.500 2256.005 3383.670 2256.175 ;
        RECT 3388.940 2256.005 3389.110 2256.175 ;
        RECT 3383.500 2255.545 3383.670 2255.715 ;
        RECT 3388.940 2255.545 3389.110 2255.715 ;
        RECT 3383.500 2255.085 3383.670 2255.255 ;
        RECT 3388.940 2255.085 3389.110 2255.255 ;
        RECT 3383.500 2254.625 3383.670 2254.795 ;
        RECT 3388.940 2254.625 3389.110 2254.795 ;
        RECT 3383.500 2254.165 3383.670 2254.335 ;
        RECT 3388.940 2254.165 3389.110 2254.335 ;
        RECT 3383.500 2253.705 3383.670 2253.875 ;
        RECT 3388.940 2253.705 3389.110 2253.875 ;
        RECT 3383.500 2253.245 3383.670 2253.415 ;
        RECT 3388.940 2253.245 3389.110 2253.415 ;
        RECT 3383.500 2252.785 3383.670 2252.955 ;
        RECT 3388.940 2252.785 3389.110 2252.955 ;
        RECT 3383.500 2252.325 3383.670 2252.495 ;
        RECT 3388.940 2252.325 3389.110 2252.495 ;
        RECT 3383.500 2251.865 3383.670 2252.035 ;
        RECT 3388.940 2251.865 3389.110 2252.035 ;
        RECT 3383.500 2251.405 3383.670 2251.575 ;
        RECT 3388.940 2251.405 3389.110 2251.575 ;
        RECT 3383.500 2250.945 3383.670 2251.115 ;
        RECT 3388.940 2250.945 3389.110 2251.115 ;
        RECT 3383.500 2250.485 3383.670 2250.655 ;
        RECT 3388.940 2250.485 3389.110 2250.655 ;
        RECT 3383.500 2250.025 3383.670 2250.195 ;
        RECT 3388.940 2250.025 3389.110 2250.195 ;
        RECT 3383.500 2249.565 3383.670 2249.735 ;
        RECT 3388.940 2249.565 3389.110 2249.735 ;
        RECT 3383.500 2249.105 3383.670 2249.275 ;
        RECT 3388.940 2249.105 3389.110 2249.275 ;
        RECT 3383.500 2248.645 3383.670 2248.815 ;
        RECT 3388.940 2248.645 3389.110 2248.815 ;
        RECT 3383.500 2248.185 3383.670 2248.355 ;
        RECT 3388.940 2248.185 3389.110 2248.355 ;
        RECT 3383.500 2247.725 3383.670 2247.895 ;
        RECT 3388.940 2247.725 3389.110 2247.895 ;
        RECT 3383.500 2247.265 3383.670 2247.435 ;
        RECT 3388.940 2247.265 3389.110 2247.435 ;
        RECT 3383.500 2246.805 3383.670 2246.975 ;
        RECT 3388.940 2246.805 3389.110 2246.975 ;
        RECT 3383.500 2246.345 3383.670 2246.515 ;
        RECT 3388.940 2246.345 3389.110 2246.515 ;
        RECT 3383.500 2245.885 3383.670 2246.055 ;
        RECT 3388.940 2245.885 3389.110 2246.055 ;
        RECT 3383.500 2245.425 3383.670 2245.595 ;
        RECT 3388.940 2245.425 3389.110 2245.595 ;
        RECT 3383.500 2244.965 3383.670 2245.135 ;
        RECT 3388.940 2244.965 3389.110 2245.135 ;
        RECT 3383.500 2244.505 3383.670 2244.675 ;
        RECT 3388.940 2244.505 3389.110 2244.675 ;
        RECT 3383.500 2244.045 3383.670 2244.215 ;
        RECT 3388.940 2244.045 3389.110 2244.215 ;
        RECT 3383.500 2243.585 3383.670 2243.755 ;
        RECT 3388.940 2243.585 3389.110 2243.755 ;
        RECT 3383.500 2243.125 3383.670 2243.295 ;
        RECT 3388.940 2243.125 3389.110 2243.295 ;
        RECT 3383.500 2242.665 3383.670 2242.835 ;
        RECT 3388.940 2242.665 3389.110 2242.835 ;
        RECT 3383.500 2242.205 3383.670 2242.375 ;
        RECT 3388.940 2242.205 3389.110 2242.375 ;
        RECT 3383.500 2241.745 3383.670 2241.915 ;
        RECT 3388.940 2241.745 3389.110 2241.915 ;
        RECT 3383.500 2241.285 3383.670 2241.455 ;
        RECT 3388.940 2241.285 3389.110 2241.455 ;
        RECT 3383.500 2240.825 3383.670 2240.995 ;
        RECT 3388.940 2240.825 3389.110 2240.995 ;
        RECT 3383.500 2240.365 3383.670 2240.535 ;
        RECT 3388.940 2240.365 3389.110 2240.535 ;
        RECT 3383.500 2239.905 3383.670 2240.075 ;
        RECT 3388.940 2239.905 3389.110 2240.075 ;
        RECT 3383.500 2239.445 3383.670 2239.615 ;
        RECT 3388.940 2239.445 3389.110 2239.615 ;
        RECT 3383.500 2238.985 3383.670 2239.155 ;
        RECT 3388.940 2238.985 3389.110 2239.155 ;
        RECT 3383.500 2238.525 3383.670 2238.695 ;
        RECT 3388.940 2238.525 3389.110 2238.695 ;
        RECT 3383.500 2238.065 3383.670 2238.235 ;
        RECT 3388.940 2238.065 3389.110 2238.235 ;
        RECT 3383.500 2237.605 3383.670 2237.775 ;
        RECT 3388.940 2237.605 3389.110 2237.775 ;
        RECT 3383.500 2237.145 3383.670 2237.315 ;
        RECT 3388.940 2237.145 3389.110 2237.315 ;
        RECT 3383.500 2236.685 3383.670 2236.855 ;
        RECT 3388.940 2236.685 3389.110 2236.855 ;
        RECT 3383.500 2236.225 3383.670 2236.395 ;
        RECT 3388.940 2236.225 3389.110 2236.395 ;
        RECT 3383.500 2235.765 3383.670 2235.935 ;
        RECT 3388.940 2235.765 3389.110 2235.935 ;
        RECT 3383.500 2235.305 3383.670 2235.475 ;
        RECT 3388.940 2235.305 3389.110 2235.475 ;
        RECT 3383.500 2234.845 3383.670 2235.015 ;
        RECT 3388.940 2234.845 3389.110 2235.015 ;
        RECT 3383.500 2234.385 3383.670 2234.555 ;
        RECT 3388.940 2234.385 3389.110 2234.555 ;
        RECT 3383.500 2233.925 3383.670 2234.095 ;
        RECT 3388.940 2233.925 3389.110 2234.095 ;
        RECT 3383.500 2233.465 3383.670 2233.635 ;
        RECT 3388.940 2233.465 3389.110 2233.635 ;
        RECT 3383.500 2233.005 3383.670 2233.175 ;
        RECT 3388.940 2233.005 3389.110 2233.175 ;
        RECT 3383.500 2232.545 3383.670 2232.715 ;
        RECT 3388.940 2232.545 3389.110 2232.715 ;
        RECT 3383.500 2232.085 3383.670 2232.255 ;
        RECT 3388.940 2232.085 3389.110 2232.255 ;
        RECT 3383.500 2231.625 3383.670 2231.795 ;
        RECT 3388.940 2231.625 3389.110 2231.795 ;
        RECT 3383.500 2231.165 3383.670 2231.335 ;
        RECT 3388.940 2231.165 3389.110 2231.335 ;
        RECT 3383.500 2230.705 3383.670 2230.875 ;
        RECT 3388.940 2230.705 3389.110 2230.875 ;
        RECT 3383.500 2230.245 3383.670 2230.415 ;
        RECT 3388.940 2230.245 3389.110 2230.415 ;
        RECT 3383.500 2229.785 3383.670 2229.955 ;
        RECT 3388.940 2229.785 3389.110 2229.955 ;
        RECT 3383.500 2229.325 3383.670 2229.495 ;
        RECT 3388.940 2229.325 3389.110 2229.495 ;
        RECT 3383.500 2228.865 3383.670 2229.035 ;
        RECT 3388.940 2228.865 3389.110 2229.035 ;
        RECT 3383.500 2228.405 3383.670 2228.575 ;
        RECT 3388.940 2228.405 3389.110 2228.575 ;
        RECT 3383.500 2227.945 3383.670 2228.115 ;
        RECT 3388.940 2227.945 3389.110 2228.115 ;
        RECT 3383.500 2227.485 3383.670 2227.655 ;
        RECT 3388.940 2227.485 3389.110 2227.655 ;
        RECT 3383.500 2227.025 3383.670 2227.195 ;
        RECT 3388.940 2227.025 3389.110 2227.195 ;
        RECT 3383.500 2226.565 3383.670 2226.735 ;
        RECT 3388.940 2226.565 3389.110 2226.735 ;
        RECT 3383.500 2226.105 3383.670 2226.275 ;
        RECT 3388.940 2226.105 3389.110 2226.275 ;
        RECT 3383.500 2225.645 3383.670 2225.815 ;
        RECT 3388.940 2225.645 3389.110 2225.815 ;
        RECT 3383.500 2225.185 3383.670 2225.355 ;
        RECT 3388.940 2225.185 3389.110 2225.355 ;
        RECT 3383.500 2224.725 3383.670 2224.895 ;
        RECT 3388.940 2224.725 3389.110 2224.895 ;
        RECT 3383.500 2224.265 3383.670 2224.435 ;
        RECT 3388.940 2224.265 3389.110 2224.435 ;
        RECT 3383.500 2223.805 3383.670 2223.975 ;
        RECT 3388.940 2223.805 3389.110 2223.975 ;
        RECT 3383.500 2223.345 3383.670 2223.515 ;
        RECT 3388.940 2223.345 3389.110 2223.515 ;
        RECT 3383.500 2222.885 3383.670 2223.055 ;
        RECT 3388.940 2222.885 3389.110 2223.055 ;
        RECT 3383.500 2222.425 3383.670 2222.595 ;
        RECT 3388.940 2222.425 3389.110 2222.595 ;
        RECT 3383.500 2221.965 3383.670 2222.135 ;
        RECT 3388.940 2221.965 3389.110 2222.135 ;
        RECT 3383.500 2221.505 3383.670 2221.675 ;
        RECT 3388.940 2221.505 3389.110 2221.675 ;
        RECT 3383.500 2221.045 3383.670 2221.215 ;
        RECT 3388.940 2221.045 3389.110 2221.215 ;
        RECT 3383.500 2220.585 3383.670 2220.755 ;
        RECT 3388.940 2220.585 3389.110 2220.755 ;
        RECT 3383.500 2220.125 3383.670 2220.295 ;
        RECT 3388.940 2220.125 3389.110 2220.295 ;
        RECT 3383.500 2219.665 3383.670 2219.835 ;
        RECT 3388.940 2219.665 3389.110 2219.835 ;
        RECT 3383.500 2219.205 3383.670 2219.375 ;
        RECT 3388.940 2219.205 3389.110 2219.375 ;
        RECT 3383.500 2218.745 3383.670 2218.915 ;
        RECT 3388.940 2218.745 3389.110 2218.915 ;
        RECT 3383.500 2218.285 3383.670 2218.455 ;
        RECT 3388.940 2218.285 3389.110 2218.455 ;
        RECT 3383.500 2217.825 3383.670 2217.995 ;
        RECT 3388.940 2217.825 3389.110 2217.995 ;
        RECT 3383.500 2217.365 3383.670 2217.535 ;
        RECT 3388.940 2217.365 3389.110 2217.535 ;
        RECT 3383.500 2216.905 3383.670 2217.075 ;
        RECT 3388.940 2216.905 3389.110 2217.075 ;
        RECT 3383.500 2216.445 3383.670 2216.615 ;
        RECT 3388.940 2216.445 3389.110 2216.615 ;
        RECT 3383.500 2215.985 3383.670 2216.155 ;
        RECT 3388.940 2215.985 3389.110 2216.155 ;
        RECT 3383.500 2215.525 3383.670 2215.695 ;
        RECT 3388.940 2215.525 3389.110 2215.695 ;
        RECT 3383.500 2215.065 3383.670 2215.235 ;
        RECT 3388.940 2215.065 3389.110 2215.235 ;
        RECT 3383.500 2214.605 3383.670 2214.775 ;
        RECT 3388.940 2214.605 3389.110 2214.775 ;
        RECT 3383.500 2214.145 3383.670 2214.315 ;
        RECT 3388.940 2214.145 3389.110 2214.315 ;
        RECT 3383.500 2213.685 3383.670 2213.855 ;
        RECT 3388.940 2213.685 3389.110 2213.855 ;
        RECT 3383.500 2213.225 3383.670 2213.395 ;
        RECT 3388.940 2213.225 3389.110 2213.395 ;
        RECT 3383.500 2212.765 3383.670 2212.935 ;
        RECT 3388.940 2212.765 3389.110 2212.935 ;
        RECT 3383.500 2212.305 3383.670 2212.475 ;
        RECT 3388.940 2212.305 3389.110 2212.475 ;
        RECT 3383.500 2211.845 3383.670 2212.015 ;
        RECT 3388.940 2211.845 3389.110 2212.015 ;
        RECT 3383.500 2211.385 3383.670 2211.555 ;
        RECT 3388.940 2211.385 3389.110 2211.555 ;
        RECT 3383.500 2210.925 3383.670 2211.095 ;
        RECT 3388.940 2210.925 3389.110 2211.095 ;
        RECT 3383.500 2210.465 3383.670 2210.635 ;
        RECT 3388.940 2210.465 3389.110 2210.635 ;
        RECT 3383.500 2210.005 3383.670 2210.175 ;
        RECT 3388.940 2210.005 3389.110 2210.175 ;
        RECT 3383.500 2209.545 3383.670 2209.715 ;
        RECT 3388.940 2209.545 3389.110 2209.715 ;
        RECT 3383.500 2209.085 3383.670 2209.255 ;
        RECT 3388.940 2209.085 3389.110 2209.255 ;
        RECT 3383.500 2208.625 3383.670 2208.795 ;
        RECT 3388.940 2208.625 3389.110 2208.795 ;
        RECT 3383.500 2208.165 3383.670 2208.335 ;
        RECT 3388.940 2208.165 3389.110 2208.335 ;
        RECT 3383.500 2207.705 3383.670 2207.875 ;
        RECT 3388.940 2207.705 3389.110 2207.875 ;
        RECT 3383.500 2207.245 3383.670 2207.415 ;
        RECT 3388.940 2207.245 3389.110 2207.415 ;
        RECT 3383.500 2206.785 3383.670 2206.955 ;
        RECT 3388.940 2206.785 3389.110 2206.955 ;
        RECT 3383.500 2206.325 3383.670 2206.495 ;
        RECT 3388.940 2206.325 3389.110 2206.495 ;
        RECT 3383.500 2205.865 3383.670 2206.035 ;
        RECT 3388.940 2205.865 3389.110 2206.035 ;
        RECT 3383.500 2205.405 3383.670 2205.575 ;
        RECT 3388.940 2205.405 3389.110 2205.575 ;
        RECT 3383.500 2204.945 3383.670 2205.115 ;
        RECT 3388.940 2204.945 3389.110 2205.115 ;
        RECT 3383.500 2204.485 3383.670 2204.655 ;
        RECT 3388.940 2204.485 3389.110 2204.655 ;
        RECT 3383.500 2204.025 3383.670 2204.195 ;
        RECT 3388.940 2204.025 3389.110 2204.195 ;
        RECT 3383.500 2203.565 3383.670 2203.735 ;
        RECT 3388.940 2203.565 3389.110 2203.735 ;
        RECT 3383.500 2203.105 3383.670 2203.275 ;
        RECT 3388.940 2203.105 3389.110 2203.275 ;
        RECT 3383.500 2202.645 3383.670 2202.815 ;
        RECT 3388.940 2202.645 3389.110 2202.815 ;
        RECT 3383.500 2202.185 3383.670 2202.355 ;
        RECT 3388.940 2202.185 3389.110 2202.355 ;
        RECT 3383.500 2201.725 3383.670 2201.895 ;
        RECT 3388.940 2201.725 3389.110 2201.895 ;
        RECT 3383.500 2201.265 3383.670 2201.435 ;
        RECT 3388.940 2201.265 3389.110 2201.435 ;
        RECT 3383.500 2200.805 3383.670 2200.975 ;
        RECT 3388.940 2200.805 3389.110 2200.975 ;
        RECT 3383.500 2200.345 3383.670 2200.515 ;
        RECT 3388.940 2200.345 3389.110 2200.515 ;
        RECT 3383.500 2199.885 3383.670 2200.055 ;
        RECT 3388.940 2199.885 3389.110 2200.055 ;
        RECT 3383.500 2199.425 3383.670 2199.595 ;
        RECT 3388.940 2199.425 3389.110 2199.595 ;
        RECT 3383.500 2198.965 3383.670 2199.135 ;
        RECT 3388.940 2198.965 3389.110 2199.135 ;
        RECT 3383.500 2198.505 3383.670 2198.675 ;
        RECT 3388.940 2198.505 3389.110 2198.675 ;
        RECT 3383.500 2198.045 3383.670 2198.215 ;
        RECT 3388.940 2198.045 3389.110 2198.215 ;
        RECT 3383.500 2197.585 3383.670 2197.755 ;
        RECT 3388.940 2197.585 3389.110 2197.755 ;
        RECT 3383.500 2197.125 3383.670 2197.295 ;
        RECT 3388.940 2197.125 3389.110 2197.295 ;
        RECT 3383.500 2196.665 3383.670 2196.835 ;
        RECT 3388.940 2196.665 3389.110 2196.835 ;
        RECT 3383.500 2196.205 3383.670 2196.375 ;
        RECT 3388.940 2196.205 3389.110 2196.375 ;
      LAYER met1 ;
        RECT 3383.345 2196.060 3383.825 2268.280 ;
        RECT 3388.785 2196.060 3389.265 2268.280 ;
      LAYER via ;
        RECT 3383.425 2240.475 3383.725 2242.260 ;
        RECT 3388.835 2240.475 3389.135 2242.260 ;
      LAYER met2 ;
        RECT 3383.365 2240.435 3383.795 2242.300 ;
        RECT 3388.790 2240.435 3389.220 2242.300 ;
      LAYER via2 ;
        RECT 3383.425 2240.475 3383.725 2242.260 ;
        RECT 3388.835 2240.475 3389.135 2242.260 ;
      LAYER met3 ;
        RECT 3383.350 2240.440 3390.875 2242.305 ;
    END
  END vssd
  PIN vccd
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 3312.980 4984.485 3313.150 4984.655 ;
        RECT 3313.440 4984.485 3313.610 4984.655 ;
        RECT 3313.900 4984.485 3314.070 4984.655 ;
        RECT 3314.360 4984.485 3314.530 4984.655 ;
        RECT 3314.820 4984.485 3314.990 4984.655 ;
        RECT 3315.280 4984.485 3315.450 4984.655 ;
        RECT 3315.740 4984.485 3315.910 4984.655 ;
        RECT 3316.200 4984.485 3316.370 4984.655 ;
        RECT 3316.660 4984.485 3316.830 4984.655 ;
        RECT 3317.120 4984.485 3317.290 4984.655 ;
        RECT 3317.580 4984.485 3317.750 4984.655 ;
        RECT 3318.040 4984.485 3318.210 4984.655 ;
        RECT 3318.500 4984.485 3318.670 4984.655 ;
        RECT 3318.960 4984.485 3319.130 4984.655 ;
        RECT 3319.420 4984.485 3319.590 4984.655 ;
        RECT 3319.880 4984.485 3320.050 4984.655 ;
        RECT 3320.340 4984.485 3320.510 4984.655 ;
        RECT 3320.800 4984.485 3320.970 4984.655 ;
        RECT 3321.260 4984.485 3321.430 4984.655 ;
        RECT 3321.720 4984.485 3321.890 4984.655 ;
        RECT 3322.180 4984.485 3322.350 4984.655 ;
        RECT 3322.640 4984.485 3322.810 4984.655 ;
        RECT 3323.100 4984.485 3323.270 4984.655 ;
        RECT 3323.560 4984.485 3323.730 4984.655 ;
        RECT 3324.020 4984.485 3324.190 4984.655 ;
        RECT 3324.480 4984.485 3324.650 4984.655 ;
        RECT 3324.940 4984.485 3325.110 4984.655 ;
        RECT 3325.400 4984.485 3325.570 4984.655 ;
        RECT 3325.860 4984.485 3326.030 4984.655 ;
        RECT 3326.320 4984.485 3326.490 4984.655 ;
        RECT 3326.780 4984.485 3326.950 4984.655 ;
        RECT 3327.240 4984.485 3327.410 4984.655 ;
        RECT 3327.700 4984.485 3327.870 4984.655 ;
        RECT 3328.160 4984.485 3328.330 4984.655 ;
        RECT 3328.620 4984.485 3328.790 4984.655 ;
        RECT 3329.080 4984.485 3329.250 4984.655 ;
        RECT 3329.540 4984.485 3329.710 4984.655 ;
        RECT 3330.000 4984.485 3330.170 4984.655 ;
        RECT 3330.460 4984.485 3330.630 4984.655 ;
        RECT 3330.920 4984.485 3331.090 4984.655 ;
        RECT 3331.380 4984.485 3331.550 4984.655 ;
        RECT 3331.840 4984.485 3332.010 4984.655 ;
        RECT 3332.300 4984.485 3332.470 4984.655 ;
        RECT 3332.760 4984.485 3332.930 4984.655 ;
        RECT 3333.220 4984.485 3333.390 4984.655 ;
        RECT 3333.680 4984.485 3333.850 4984.655 ;
        RECT 3334.140 4984.485 3334.310 4984.655 ;
        RECT 3334.600 4984.485 3334.770 4984.655 ;
        RECT 3335.060 4984.485 3335.230 4984.655 ;
        RECT 3335.520 4984.485 3335.690 4984.655 ;
        RECT 3335.980 4984.485 3336.150 4984.655 ;
        RECT 3336.440 4984.485 3336.610 4984.655 ;
        RECT 3336.900 4984.485 3337.070 4984.655 ;
      LAYER met1 ;
        RECT 3312.835 4984.330 3337.215 4984.810 ;
      LAYER via ;
        RECT 3327.165 4984.420 3328.950 4984.720 ;
      LAYER met2 ;
        RECT 3327.125 4984.350 3328.990 4984.780 ;
      LAYER via2 ;
        RECT 3327.165 4984.420 3328.950 4984.720 ;
      LAYER met3 ;
        RECT 3327.130 4984.350 3328.980 4989.165 ;
    END
    PORT
      LAYER li1 ;
        RECT 2082.975 4984.895 2083.145 4985.065 ;
        RECT 2083.435 4984.895 2083.605 4985.065 ;
        RECT 2083.895 4984.895 2084.065 4985.065 ;
        RECT 2084.355 4984.895 2084.525 4985.065 ;
        RECT 2084.815 4984.895 2084.985 4985.065 ;
        RECT 2085.275 4984.895 2085.445 4985.065 ;
        RECT 2085.735 4984.895 2085.905 4985.065 ;
        RECT 2086.195 4984.895 2086.365 4985.065 ;
        RECT 2086.655 4984.895 2086.825 4985.065 ;
        RECT 2087.115 4984.895 2087.285 4985.065 ;
        RECT 2087.575 4984.895 2087.745 4985.065 ;
        RECT 2088.035 4984.895 2088.205 4985.065 ;
        RECT 2088.495 4984.895 2088.665 4985.065 ;
        RECT 2088.955 4984.895 2089.125 4985.065 ;
      LAYER met1 ;
        RECT 2082.830 4984.740 2092.990 4985.220 ;
      LAYER via ;
        RECT 2091.115 4984.830 2092.900 4985.130 ;
      LAYER met2 ;
        RECT 2091.075 4984.760 2092.940 4985.190 ;
      LAYER via2 ;
        RECT 2091.115 4984.830 2092.900 4985.130 ;
      LAYER met3 ;
        RECT 2091.080 4984.760 2092.930 4989.575 ;
    END
    PORT
      LAYER li1 ;
        RECT 834.795 4983.270 834.965 4983.440 ;
        RECT 835.255 4983.270 835.425 4983.440 ;
        RECT 835.715 4983.270 835.885 4983.440 ;
        RECT 836.175 4983.270 836.345 4983.440 ;
        RECT 836.635 4983.270 836.805 4983.440 ;
        RECT 837.095 4983.270 837.265 4983.440 ;
        RECT 837.555 4983.270 837.725 4983.440 ;
        RECT 838.015 4983.270 838.185 4983.440 ;
        RECT 838.475 4983.270 838.645 4983.440 ;
        RECT 838.935 4983.270 839.105 4983.440 ;
        RECT 839.395 4983.270 839.565 4983.440 ;
        RECT 839.855 4983.270 840.025 4983.440 ;
        RECT 840.315 4983.270 840.485 4983.440 ;
        RECT 840.775 4983.270 840.945 4983.440 ;
        RECT 841.235 4983.270 841.405 4983.440 ;
        RECT 841.695 4983.270 841.865 4983.440 ;
        RECT 842.155 4983.270 842.325 4983.440 ;
        RECT 842.615 4983.270 842.785 4983.440 ;
        RECT 843.075 4983.270 843.245 4983.440 ;
        RECT 843.535 4983.270 843.705 4983.440 ;
        RECT 843.995 4983.270 844.165 4983.440 ;
        RECT 844.455 4983.270 844.625 4983.440 ;
        RECT 844.915 4983.270 845.085 4983.440 ;
        RECT 845.375 4983.270 845.545 4983.440 ;
        RECT 845.835 4983.270 846.005 4983.440 ;
        RECT 846.295 4983.270 846.465 4983.440 ;
        RECT 846.755 4983.270 846.925 4983.440 ;
        RECT 847.215 4983.270 847.385 4983.440 ;
        RECT 847.675 4983.270 847.845 4983.440 ;
        RECT 848.135 4983.270 848.305 4983.440 ;
        RECT 848.595 4983.270 848.765 4983.440 ;
        RECT 849.055 4983.270 849.225 4983.440 ;
        RECT 849.515 4983.270 849.685 4983.440 ;
        RECT 849.975 4983.270 850.145 4983.440 ;
        RECT 850.435 4983.270 850.605 4983.440 ;
        RECT 850.895 4983.270 851.065 4983.440 ;
        RECT 851.355 4983.270 851.525 4983.440 ;
        RECT 851.815 4983.270 851.985 4983.440 ;
        RECT 852.275 4983.270 852.445 4983.440 ;
        RECT 852.735 4983.270 852.905 4983.440 ;
      LAYER met1 ;
        RECT 834.650 4983.115 853.050 4983.595 ;
      LAYER via ;
        RECT 848.930 4983.185 850.715 4983.485 ;
      LAYER met2 ;
        RECT 848.890 4983.115 850.755 4983.545 ;
      LAYER via2 ;
        RECT 848.930 4983.185 850.715 4983.485 ;
      LAYER met3 ;
        RECT 848.895 4983.115 850.745 4987.930 ;
    END
    PORT
      LAYER li1 ;
        RECT 669.145 1114.320 669.315 1114.490 ;
        RECT 669.605 1114.320 669.775 1114.490 ;
        RECT 670.065 1114.320 670.235 1114.490 ;
        RECT 670.525 1114.320 670.695 1114.490 ;
        RECT 670.985 1114.320 671.155 1114.490 ;
        RECT 671.445 1114.320 671.615 1114.490 ;
        RECT 671.905 1114.320 672.075 1114.490 ;
        RECT 672.365 1114.320 672.535 1114.490 ;
        RECT 672.825 1114.320 672.995 1114.490 ;
        RECT 673.285 1114.320 673.455 1114.490 ;
        RECT 673.745 1114.320 673.915 1114.490 ;
        RECT 674.205 1114.320 674.375 1114.490 ;
        RECT 674.665 1114.320 674.835 1114.490 ;
        RECT 675.125 1114.320 675.295 1114.490 ;
        RECT 675.585 1114.320 675.755 1114.490 ;
        RECT 676.045 1114.320 676.215 1114.490 ;
        RECT 676.505 1114.320 676.675 1114.490 ;
        RECT 676.965 1114.320 677.135 1114.490 ;
        RECT 677.425 1114.320 677.595 1114.490 ;
        RECT 677.885 1114.320 678.055 1114.490 ;
        RECT 678.345 1114.320 678.515 1114.490 ;
        RECT 678.805 1114.320 678.975 1114.490 ;
        RECT 679.265 1114.320 679.435 1114.490 ;
        RECT 679.725 1114.320 679.895 1114.490 ;
        RECT 680.185 1114.320 680.355 1114.490 ;
        RECT 680.645 1114.320 680.815 1114.490 ;
        RECT 681.105 1114.320 681.275 1114.490 ;
        RECT 681.565 1114.320 681.735 1114.490 ;
        RECT 682.025 1114.320 682.195 1114.490 ;
        RECT 682.485 1114.320 682.655 1114.490 ;
        RECT 682.945 1114.320 683.115 1114.490 ;
        RECT 683.405 1114.320 683.575 1114.490 ;
        RECT 683.865 1114.320 684.035 1114.490 ;
        RECT 684.325 1114.320 684.495 1114.490 ;
        RECT 684.785 1114.320 684.955 1114.490 ;
        RECT 685.245 1114.320 685.415 1114.490 ;
        RECT 685.705 1114.320 685.875 1114.490 ;
        RECT 686.165 1114.320 686.335 1114.490 ;
        RECT 686.625 1114.320 686.795 1114.490 ;
        RECT 687.085 1114.320 687.255 1114.490 ;
        RECT 687.545 1114.320 687.715 1114.490 ;
        RECT 688.005 1114.320 688.175 1114.490 ;
        RECT 688.465 1114.320 688.635 1114.490 ;
        RECT 688.925 1114.320 689.095 1114.490 ;
        RECT 689.385 1114.320 689.555 1114.490 ;
        RECT 689.845 1114.320 690.015 1114.490 ;
        RECT 690.305 1114.320 690.475 1114.490 ;
        RECT 690.765 1114.320 690.935 1114.490 ;
        RECT 691.225 1114.320 691.395 1114.490 ;
        RECT 691.685 1114.320 691.855 1114.490 ;
        RECT 692.145 1114.320 692.315 1114.490 ;
        RECT 692.605 1114.320 692.775 1114.490 ;
        RECT 693.065 1114.320 693.235 1114.490 ;
        RECT 693.525 1114.320 693.695 1114.490 ;
        RECT 693.985 1114.320 694.155 1114.490 ;
        RECT 694.445 1114.320 694.615 1114.490 ;
        RECT 694.905 1114.320 695.075 1114.490 ;
        RECT 695.365 1114.320 695.535 1114.490 ;
        RECT 695.825 1114.320 695.995 1114.490 ;
        RECT 696.285 1114.320 696.455 1114.490 ;
        RECT 696.745 1114.320 696.915 1114.490 ;
        RECT 697.205 1114.320 697.375 1114.490 ;
        RECT 697.665 1114.320 697.835 1114.490 ;
        RECT 698.125 1114.320 698.295 1114.490 ;
        RECT 698.585 1114.320 698.755 1114.490 ;
        RECT 699.045 1114.320 699.215 1114.490 ;
        RECT 699.505 1114.320 699.675 1114.490 ;
        RECT 699.965 1114.320 700.135 1114.490 ;
        RECT 700.425 1114.320 700.595 1114.490 ;
        RECT 700.885 1114.320 701.055 1114.490 ;
        RECT 701.345 1114.320 701.515 1114.490 ;
        RECT 701.805 1114.320 701.975 1114.490 ;
        RECT 702.265 1114.320 702.435 1114.490 ;
        RECT 702.725 1114.320 702.895 1114.490 ;
        RECT 703.185 1114.320 703.355 1114.490 ;
        RECT 703.645 1114.320 703.815 1114.490 ;
        RECT 704.105 1114.320 704.275 1114.490 ;
        RECT 704.565 1114.320 704.735 1114.490 ;
        RECT 705.025 1114.320 705.195 1114.490 ;
        RECT 705.485 1114.320 705.655 1114.490 ;
        RECT 705.945 1114.320 706.115 1114.490 ;
        RECT 706.405 1114.320 706.575 1114.490 ;
        RECT 706.865 1114.320 707.035 1114.490 ;
        RECT 707.325 1114.320 707.495 1114.490 ;
        RECT 707.785 1114.320 707.955 1114.490 ;
        RECT 708.245 1114.320 708.415 1114.490 ;
        RECT 708.705 1114.320 708.875 1114.490 ;
        RECT 709.165 1114.320 709.335 1114.490 ;
        RECT 709.625 1114.320 709.795 1114.490 ;
        RECT 710.085 1114.320 710.255 1114.490 ;
        RECT 710.545 1114.320 710.715 1114.490 ;
        RECT 711.005 1114.320 711.175 1114.490 ;
        RECT 711.465 1114.320 711.635 1114.490 ;
        RECT 711.925 1114.320 712.095 1114.490 ;
        RECT 712.385 1114.320 712.555 1114.490 ;
        RECT 712.845 1114.320 713.015 1114.490 ;
        RECT 713.305 1114.320 713.475 1114.490 ;
        RECT 713.765 1114.320 713.935 1114.490 ;
        RECT 714.225 1114.320 714.395 1114.490 ;
        RECT 714.685 1114.320 714.855 1114.490 ;
        RECT 715.145 1114.320 715.315 1114.490 ;
        RECT 715.605 1114.320 715.775 1114.490 ;
        RECT 716.065 1114.320 716.235 1114.490 ;
        RECT 716.525 1114.320 716.695 1114.490 ;
        RECT 716.985 1114.320 717.155 1114.490 ;
        RECT 717.445 1114.320 717.615 1114.490 ;
        RECT 717.905 1114.320 718.075 1114.490 ;
        RECT 718.365 1114.320 718.535 1114.490 ;
        RECT 718.825 1114.320 718.995 1114.490 ;
        RECT 719.285 1114.320 719.455 1114.490 ;
        RECT 719.745 1114.320 719.915 1114.490 ;
        RECT 720.205 1114.320 720.375 1114.490 ;
        RECT 720.665 1114.320 720.835 1114.490 ;
        RECT 721.125 1114.320 721.295 1114.490 ;
        RECT 721.585 1114.320 721.755 1114.490 ;
        RECT 722.045 1114.320 722.215 1114.490 ;
        RECT 722.505 1114.320 722.675 1114.490 ;
        RECT 722.965 1114.320 723.135 1114.490 ;
        RECT 723.425 1114.320 723.595 1114.490 ;
        RECT 723.885 1114.320 724.055 1114.490 ;
        RECT 724.345 1114.320 724.515 1114.490 ;
        RECT 724.805 1114.320 724.975 1114.490 ;
        RECT 725.265 1114.320 725.435 1114.490 ;
        RECT 725.725 1114.320 725.895 1114.490 ;
        RECT 726.185 1114.320 726.355 1114.490 ;
        RECT 726.645 1114.320 726.815 1114.490 ;
        RECT 727.105 1114.320 727.275 1114.490 ;
        RECT 727.565 1114.320 727.735 1114.490 ;
        RECT 728.025 1114.320 728.195 1114.490 ;
        RECT 728.485 1114.320 728.655 1114.490 ;
        RECT 728.945 1114.320 729.115 1114.490 ;
        RECT 729.405 1114.320 729.575 1114.490 ;
        RECT 729.865 1114.320 730.035 1114.490 ;
        RECT 730.325 1114.320 730.495 1114.490 ;
        RECT 730.785 1114.320 730.955 1114.490 ;
        RECT 731.245 1114.320 731.415 1114.490 ;
        RECT 731.705 1114.320 731.875 1114.490 ;
        RECT 732.165 1114.320 732.335 1114.490 ;
        RECT 732.625 1114.320 732.795 1114.490 ;
        RECT 733.085 1114.320 733.255 1114.490 ;
        RECT 733.545 1114.320 733.715 1114.490 ;
        RECT 734.005 1114.320 734.175 1114.490 ;
        RECT 734.465 1114.320 734.635 1114.490 ;
        RECT 734.925 1114.320 735.095 1114.490 ;
        RECT 735.385 1114.320 735.555 1114.490 ;
        RECT 735.845 1114.320 736.015 1114.490 ;
        RECT 736.305 1114.320 736.475 1114.490 ;
        RECT 736.765 1114.320 736.935 1114.490 ;
        RECT 737.225 1114.320 737.395 1114.490 ;
        RECT 737.685 1114.320 737.855 1114.490 ;
        RECT 738.145 1114.320 738.315 1114.490 ;
        RECT 738.605 1114.320 738.775 1114.490 ;
        RECT 739.065 1114.320 739.235 1114.490 ;
        RECT 739.525 1114.320 739.695 1114.490 ;
        RECT 739.985 1114.320 740.155 1114.490 ;
        RECT 740.445 1114.320 740.615 1114.490 ;
        RECT 740.905 1114.320 741.075 1114.490 ;
        RECT 741.365 1114.320 741.535 1114.490 ;
        RECT 741.825 1114.320 741.995 1114.490 ;
        RECT 742.285 1114.320 742.455 1114.490 ;
        RECT 742.745 1114.320 742.915 1114.490 ;
        RECT 743.205 1114.320 743.375 1114.490 ;
        RECT 743.665 1114.320 743.835 1114.490 ;
        RECT 744.125 1114.320 744.295 1114.490 ;
        RECT 744.585 1114.320 744.755 1114.490 ;
        RECT 745.045 1114.320 745.215 1114.490 ;
        RECT 745.505 1114.320 745.675 1114.490 ;
        RECT 745.965 1114.320 746.135 1114.490 ;
        RECT 746.425 1114.320 746.595 1114.490 ;
        RECT 746.885 1114.320 747.055 1114.490 ;
        RECT 747.345 1114.320 747.515 1114.490 ;
        RECT 747.805 1114.320 747.975 1114.490 ;
        RECT 748.265 1114.320 748.435 1114.490 ;
        RECT 748.725 1114.320 748.895 1114.490 ;
        RECT 749.185 1114.320 749.355 1114.490 ;
        RECT 749.645 1114.320 749.815 1114.490 ;
        RECT 750.105 1114.320 750.275 1114.490 ;
        RECT 750.565 1114.320 750.735 1114.490 ;
        RECT 751.025 1114.320 751.195 1114.490 ;
        RECT 751.485 1114.320 751.655 1114.490 ;
        RECT 751.945 1114.320 752.115 1114.490 ;
        RECT 752.405 1114.320 752.575 1114.490 ;
        RECT 752.865 1114.320 753.035 1114.490 ;
        RECT 753.325 1114.320 753.495 1114.490 ;
        RECT 753.785 1114.320 753.955 1114.490 ;
        RECT 754.245 1114.320 754.415 1114.490 ;
        RECT 754.705 1114.320 754.875 1114.490 ;
        RECT 755.165 1114.320 755.335 1114.490 ;
        RECT 755.625 1114.320 755.795 1114.490 ;
        RECT 756.085 1114.320 756.255 1114.490 ;
        RECT 756.545 1114.320 756.715 1114.490 ;
        RECT 757.005 1114.320 757.175 1114.490 ;
        RECT 757.465 1114.320 757.635 1114.490 ;
        RECT 757.925 1114.320 758.095 1114.490 ;
        RECT 758.385 1114.320 758.555 1114.490 ;
        RECT 758.845 1114.320 759.015 1114.490 ;
        RECT 759.305 1114.320 759.475 1114.490 ;
        RECT 759.765 1114.320 759.935 1114.490 ;
        RECT 760.225 1114.320 760.395 1114.490 ;
        RECT 760.685 1114.320 760.855 1114.490 ;
        RECT 761.145 1114.320 761.315 1114.490 ;
        RECT 761.605 1114.320 761.775 1114.490 ;
        RECT 762.065 1114.320 762.235 1114.490 ;
        RECT 762.525 1114.320 762.695 1114.490 ;
        RECT 762.985 1114.320 763.155 1114.490 ;
        RECT 763.445 1114.320 763.615 1114.490 ;
        RECT 763.905 1114.320 764.075 1114.490 ;
        RECT 764.365 1114.320 764.535 1114.490 ;
        RECT 764.825 1114.320 764.995 1114.490 ;
        RECT 765.285 1114.320 765.455 1114.490 ;
        RECT 765.745 1114.320 765.915 1114.490 ;
        RECT 766.205 1114.320 766.375 1114.490 ;
        RECT 766.665 1114.320 766.835 1114.490 ;
        RECT 767.125 1114.320 767.295 1114.490 ;
        RECT 767.585 1114.320 767.755 1114.490 ;
        RECT 768.045 1114.320 768.215 1114.490 ;
        RECT 768.505 1114.320 768.675 1114.490 ;
        RECT 768.965 1114.320 769.135 1114.490 ;
        RECT 769.425 1114.320 769.595 1114.490 ;
        RECT 769.885 1114.320 770.055 1114.490 ;
        RECT 770.345 1114.320 770.515 1114.490 ;
        RECT 770.805 1114.320 770.975 1114.490 ;
        RECT 771.265 1114.320 771.435 1114.490 ;
        RECT 771.725 1114.320 771.895 1114.490 ;
        RECT 772.185 1114.320 772.355 1114.490 ;
        RECT 772.645 1114.320 772.815 1114.490 ;
        RECT 773.105 1114.320 773.275 1114.490 ;
        RECT 773.565 1114.320 773.735 1114.490 ;
        RECT 774.025 1114.320 774.195 1114.490 ;
        RECT 774.485 1114.320 774.655 1114.490 ;
        RECT 774.945 1114.320 775.115 1114.490 ;
        RECT 775.405 1114.320 775.575 1114.490 ;
        RECT 775.865 1114.320 776.035 1114.490 ;
        RECT 776.325 1114.320 776.495 1114.490 ;
        RECT 776.785 1114.320 776.955 1114.490 ;
        RECT 777.245 1114.320 777.415 1114.490 ;
        RECT 777.705 1114.320 777.875 1114.490 ;
        RECT 778.165 1114.320 778.335 1114.490 ;
        RECT 778.625 1114.320 778.795 1114.490 ;
        RECT 779.085 1114.320 779.255 1114.490 ;
        RECT 779.545 1114.320 779.715 1114.490 ;
        RECT 780.005 1114.320 780.175 1114.490 ;
        RECT 780.465 1114.320 780.635 1114.490 ;
        RECT 780.925 1114.320 781.095 1114.490 ;
        RECT 781.385 1114.320 781.555 1114.490 ;
        RECT 781.845 1114.320 782.015 1114.490 ;
        RECT 782.305 1114.320 782.475 1114.490 ;
        RECT 782.765 1114.320 782.935 1114.490 ;
        RECT 783.225 1114.320 783.395 1114.490 ;
        RECT 783.685 1114.320 783.855 1114.490 ;
        RECT 784.145 1114.320 784.315 1114.490 ;
        RECT 784.605 1114.320 784.775 1114.490 ;
        RECT 785.065 1114.320 785.235 1114.490 ;
        RECT 785.525 1114.320 785.695 1114.490 ;
        RECT 785.985 1114.320 786.155 1114.490 ;
        RECT 786.445 1114.320 786.615 1114.490 ;
        RECT 786.905 1114.320 787.075 1114.490 ;
        RECT 787.365 1114.320 787.535 1114.490 ;
        RECT 787.825 1114.320 787.995 1114.490 ;
        RECT 788.285 1114.320 788.455 1114.490 ;
        RECT 788.745 1114.320 788.915 1114.490 ;
        RECT 789.205 1114.320 789.375 1114.490 ;
        RECT 789.665 1114.320 789.835 1114.490 ;
        RECT 790.125 1114.320 790.295 1114.490 ;
        RECT 790.585 1114.320 790.755 1114.490 ;
        RECT 791.045 1114.320 791.215 1114.490 ;
        RECT 791.505 1114.320 791.675 1114.490 ;
        RECT 791.965 1114.320 792.135 1114.490 ;
        RECT 792.425 1114.320 792.595 1114.490 ;
        RECT 792.885 1114.320 793.055 1114.490 ;
        RECT 793.345 1114.320 793.515 1114.490 ;
        RECT 793.805 1114.320 793.975 1114.490 ;
        RECT 794.265 1114.320 794.435 1114.490 ;
        RECT 794.725 1114.320 794.895 1114.490 ;
      LAYER met1 ;
        RECT 669.000 1114.165 795.040 1114.645 ;
      LAYER via ;
        RECT 730.995 1114.280 732.780 1114.580 ;
      LAYER met2 ;
        RECT 730.955 1114.220 732.820 1114.650 ;
      LAYER via2 ;
        RECT 730.995 1114.280 732.780 1114.580 ;
      LAYER met3 ;
        RECT 730.965 1109.835 732.815 1114.650 ;
    END
    PORT
      LAYER li1 ;
        RECT 1969.145 1114.320 1969.315 1114.490 ;
        RECT 1969.605 1114.320 1969.775 1114.490 ;
        RECT 1970.065 1114.320 1970.235 1114.490 ;
        RECT 1970.525 1114.320 1970.695 1114.490 ;
        RECT 1970.985 1114.320 1971.155 1114.490 ;
        RECT 1971.445 1114.320 1971.615 1114.490 ;
        RECT 1971.905 1114.320 1972.075 1114.490 ;
        RECT 1972.365 1114.320 1972.535 1114.490 ;
        RECT 1972.825 1114.320 1972.995 1114.490 ;
        RECT 1973.285 1114.320 1973.455 1114.490 ;
        RECT 1973.745 1114.320 1973.915 1114.490 ;
        RECT 1974.205 1114.320 1974.375 1114.490 ;
        RECT 1974.665 1114.320 1974.835 1114.490 ;
        RECT 1975.125 1114.320 1975.295 1114.490 ;
        RECT 1975.585 1114.320 1975.755 1114.490 ;
        RECT 1976.045 1114.320 1976.215 1114.490 ;
        RECT 1976.505 1114.320 1976.675 1114.490 ;
        RECT 1976.965 1114.320 1977.135 1114.490 ;
        RECT 1977.425 1114.320 1977.595 1114.490 ;
        RECT 1977.885 1114.320 1978.055 1114.490 ;
        RECT 1978.345 1114.320 1978.515 1114.490 ;
        RECT 1978.805 1114.320 1978.975 1114.490 ;
        RECT 1979.265 1114.320 1979.435 1114.490 ;
        RECT 1979.725 1114.320 1979.895 1114.490 ;
        RECT 1980.185 1114.320 1980.355 1114.490 ;
        RECT 1980.645 1114.320 1980.815 1114.490 ;
        RECT 1981.105 1114.320 1981.275 1114.490 ;
        RECT 1981.565 1114.320 1981.735 1114.490 ;
        RECT 1982.025 1114.320 1982.195 1114.490 ;
        RECT 1982.485 1114.320 1982.655 1114.490 ;
        RECT 1982.945 1114.320 1983.115 1114.490 ;
        RECT 1983.405 1114.320 1983.575 1114.490 ;
        RECT 1983.865 1114.320 1984.035 1114.490 ;
        RECT 1984.325 1114.320 1984.495 1114.490 ;
        RECT 1984.785 1114.320 1984.955 1114.490 ;
        RECT 1985.245 1114.320 1985.415 1114.490 ;
        RECT 1985.705 1114.320 1985.875 1114.490 ;
        RECT 1986.165 1114.320 1986.335 1114.490 ;
        RECT 1986.625 1114.320 1986.795 1114.490 ;
        RECT 1987.085 1114.320 1987.255 1114.490 ;
        RECT 1987.545 1114.320 1987.715 1114.490 ;
        RECT 1988.005 1114.320 1988.175 1114.490 ;
        RECT 1988.465 1114.320 1988.635 1114.490 ;
        RECT 1988.925 1114.320 1989.095 1114.490 ;
        RECT 1989.385 1114.320 1989.555 1114.490 ;
        RECT 1989.845 1114.320 1990.015 1114.490 ;
        RECT 1990.305 1114.320 1990.475 1114.490 ;
        RECT 1990.765 1114.320 1990.935 1114.490 ;
        RECT 1991.225 1114.320 1991.395 1114.490 ;
        RECT 1991.685 1114.320 1991.855 1114.490 ;
        RECT 1992.145 1114.320 1992.315 1114.490 ;
        RECT 1992.605 1114.320 1992.775 1114.490 ;
        RECT 1993.065 1114.320 1993.235 1114.490 ;
        RECT 1993.525 1114.320 1993.695 1114.490 ;
        RECT 1993.985 1114.320 1994.155 1114.490 ;
        RECT 1994.445 1114.320 1994.615 1114.490 ;
        RECT 1994.905 1114.320 1995.075 1114.490 ;
        RECT 1995.365 1114.320 1995.535 1114.490 ;
        RECT 1995.825 1114.320 1995.995 1114.490 ;
        RECT 1996.285 1114.320 1996.455 1114.490 ;
        RECT 1996.745 1114.320 1996.915 1114.490 ;
        RECT 1997.205 1114.320 1997.375 1114.490 ;
        RECT 1997.665 1114.320 1997.835 1114.490 ;
        RECT 1998.125 1114.320 1998.295 1114.490 ;
        RECT 1998.585 1114.320 1998.755 1114.490 ;
        RECT 1999.045 1114.320 1999.215 1114.490 ;
        RECT 1999.505 1114.320 1999.675 1114.490 ;
        RECT 1999.965 1114.320 2000.135 1114.490 ;
        RECT 2000.425 1114.320 2000.595 1114.490 ;
        RECT 2000.885 1114.320 2001.055 1114.490 ;
        RECT 2001.345 1114.320 2001.515 1114.490 ;
        RECT 2001.805 1114.320 2001.975 1114.490 ;
        RECT 2002.265 1114.320 2002.435 1114.490 ;
        RECT 2002.725 1114.320 2002.895 1114.490 ;
        RECT 2003.185 1114.320 2003.355 1114.490 ;
        RECT 2003.645 1114.320 2003.815 1114.490 ;
        RECT 2004.105 1114.320 2004.275 1114.490 ;
        RECT 2004.565 1114.320 2004.735 1114.490 ;
        RECT 2005.025 1114.320 2005.195 1114.490 ;
        RECT 2005.485 1114.320 2005.655 1114.490 ;
        RECT 2005.945 1114.320 2006.115 1114.490 ;
        RECT 2006.405 1114.320 2006.575 1114.490 ;
        RECT 2006.865 1114.320 2007.035 1114.490 ;
        RECT 2007.325 1114.320 2007.495 1114.490 ;
        RECT 2007.785 1114.320 2007.955 1114.490 ;
        RECT 2008.245 1114.320 2008.415 1114.490 ;
        RECT 2008.705 1114.320 2008.875 1114.490 ;
        RECT 2009.165 1114.320 2009.335 1114.490 ;
        RECT 2009.625 1114.320 2009.795 1114.490 ;
        RECT 2010.085 1114.320 2010.255 1114.490 ;
        RECT 2010.545 1114.320 2010.715 1114.490 ;
        RECT 2011.005 1114.320 2011.175 1114.490 ;
        RECT 2011.465 1114.320 2011.635 1114.490 ;
        RECT 2011.925 1114.320 2012.095 1114.490 ;
        RECT 2012.385 1114.320 2012.555 1114.490 ;
        RECT 2012.845 1114.320 2013.015 1114.490 ;
        RECT 2013.305 1114.320 2013.475 1114.490 ;
        RECT 2013.765 1114.320 2013.935 1114.490 ;
        RECT 2014.225 1114.320 2014.395 1114.490 ;
        RECT 2014.685 1114.320 2014.855 1114.490 ;
        RECT 2015.145 1114.320 2015.315 1114.490 ;
        RECT 2015.605 1114.320 2015.775 1114.490 ;
        RECT 2016.065 1114.320 2016.235 1114.490 ;
        RECT 2016.525 1114.320 2016.695 1114.490 ;
        RECT 2016.985 1114.320 2017.155 1114.490 ;
        RECT 2017.445 1114.320 2017.615 1114.490 ;
        RECT 2017.905 1114.320 2018.075 1114.490 ;
        RECT 2018.365 1114.320 2018.535 1114.490 ;
        RECT 2018.825 1114.320 2018.995 1114.490 ;
        RECT 2019.285 1114.320 2019.455 1114.490 ;
        RECT 2019.745 1114.320 2019.915 1114.490 ;
        RECT 2020.205 1114.320 2020.375 1114.490 ;
        RECT 2020.665 1114.320 2020.835 1114.490 ;
        RECT 2021.125 1114.320 2021.295 1114.490 ;
        RECT 2021.585 1114.320 2021.755 1114.490 ;
        RECT 2022.045 1114.320 2022.215 1114.490 ;
        RECT 2022.505 1114.320 2022.675 1114.490 ;
        RECT 2022.965 1114.320 2023.135 1114.490 ;
        RECT 2023.425 1114.320 2023.595 1114.490 ;
        RECT 2023.885 1114.320 2024.055 1114.490 ;
        RECT 2024.345 1114.320 2024.515 1114.490 ;
        RECT 2024.805 1114.320 2024.975 1114.490 ;
        RECT 2025.265 1114.320 2025.435 1114.490 ;
        RECT 2025.725 1114.320 2025.895 1114.490 ;
        RECT 2026.185 1114.320 2026.355 1114.490 ;
        RECT 2026.645 1114.320 2026.815 1114.490 ;
        RECT 2027.105 1114.320 2027.275 1114.490 ;
        RECT 2027.565 1114.320 2027.735 1114.490 ;
        RECT 2028.025 1114.320 2028.195 1114.490 ;
        RECT 2028.485 1114.320 2028.655 1114.490 ;
        RECT 2028.945 1114.320 2029.115 1114.490 ;
        RECT 2029.405 1114.320 2029.575 1114.490 ;
        RECT 2029.865 1114.320 2030.035 1114.490 ;
        RECT 2030.325 1114.320 2030.495 1114.490 ;
        RECT 2030.785 1114.320 2030.955 1114.490 ;
        RECT 2031.245 1114.320 2031.415 1114.490 ;
        RECT 2031.705 1114.320 2031.875 1114.490 ;
        RECT 2032.165 1114.320 2032.335 1114.490 ;
        RECT 2032.625 1114.320 2032.795 1114.490 ;
        RECT 2033.085 1114.320 2033.255 1114.490 ;
        RECT 2033.545 1114.320 2033.715 1114.490 ;
        RECT 2034.005 1114.320 2034.175 1114.490 ;
        RECT 2034.465 1114.320 2034.635 1114.490 ;
        RECT 2034.925 1114.320 2035.095 1114.490 ;
        RECT 2035.385 1114.320 2035.555 1114.490 ;
        RECT 2035.845 1114.320 2036.015 1114.490 ;
        RECT 2036.305 1114.320 2036.475 1114.490 ;
        RECT 2036.765 1114.320 2036.935 1114.490 ;
        RECT 2037.225 1114.320 2037.395 1114.490 ;
        RECT 2037.685 1114.320 2037.855 1114.490 ;
        RECT 2038.145 1114.320 2038.315 1114.490 ;
        RECT 2038.605 1114.320 2038.775 1114.490 ;
        RECT 2039.065 1114.320 2039.235 1114.490 ;
        RECT 2039.525 1114.320 2039.695 1114.490 ;
        RECT 2039.985 1114.320 2040.155 1114.490 ;
        RECT 2040.445 1114.320 2040.615 1114.490 ;
        RECT 2040.905 1114.320 2041.075 1114.490 ;
        RECT 2041.365 1114.320 2041.535 1114.490 ;
        RECT 2041.825 1114.320 2041.995 1114.490 ;
        RECT 2042.285 1114.320 2042.455 1114.490 ;
        RECT 2042.745 1114.320 2042.915 1114.490 ;
        RECT 2043.205 1114.320 2043.375 1114.490 ;
        RECT 2043.665 1114.320 2043.835 1114.490 ;
        RECT 2044.125 1114.320 2044.295 1114.490 ;
        RECT 2044.585 1114.320 2044.755 1114.490 ;
        RECT 2045.045 1114.320 2045.215 1114.490 ;
        RECT 2045.505 1114.320 2045.675 1114.490 ;
        RECT 2045.965 1114.320 2046.135 1114.490 ;
        RECT 2046.425 1114.320 2046.595 1114.490 ;
        RECT 2046.885 1114.320 2047.055 1114.490 ;
        RECT 2047.345 1114.320 2047.515 1114.490 ;
        RECT 2047.805 1114.320 2047.975 1114.490 ;
        RECT 2048.265 1114.320 2048.435 1114.490 ;
        RECT 2048.725 1114.320 2048.895 1114.490 ;
        RECT 2049.185 1114.320 2049.355 1114.490 ;
        RECT 2049.645 1114.320 2049.815 1114.490 ;
        RECT 2050.105 1114.320 2050.275 1114.490 ;
        RECT 2050.565 1114.320 2050.735 1114.490 ;
        RECT 2051.025 1114.320 2051.195 1114.490 ;
        RECT 2051.485 1114.320 2051.655 1114.490 ;
        RECT 2051.945 1114.320 2052.115 1114.490 ;
        RECT 2052.405 1114.320 2052.575 1114.490 ;
        RECT 2052.865 1114.320 2053.035 1114.490 ;
        RECT 2053.325 1114.320 2053.495 1114.490 ;
        RECT 2053.785 1114.320 2053.955 1114.490 ;
        RECT 2054.245 1114.320 2054.415 1114.490 ;
        RECT 2054.705 1114.320 2054.875 1114.490 ;
        RECT 2055.165 1114.320 2055.335 1114.490 ;
        RECT 2055.625 1114.320 2055.795 1114.490 ;
        RECT 2056.085 1114.320 2056.255 1114.490 ;
        RECT 2056.545 1114.320 2056.715 1114.490 ;
        RECT 2057.005 1114.320 2057.175 1114.490 ;
        RECT 2057.465 1114.320 2057.635 1114.490 ;
        RECT 2057.925 1114.320 2058.095 1114.490 ;
        RECT 2058.385 1114.320 2058.555 1114.490 ;
        RECT 2058.845 1114.320 2059.015 1114.490 ;
        RECT 2059.305 1114.320 2059.475 1114.490 ;
        RECT 2059.765 1114.320 2059.935 1114.490 ;
        RECT 2060.225 1114.320 2060.395 1114.490 ;
        RECT 2060.685 1114.320 2060.855 1114.490 ;
        RECT 2061.145 1114.320 2061.315 1114.490 ;
        RECT 2061.605 1114.320 2061.775 1114.490 ;
        RECT 2062.065 1114.320 2062.235 1114.490 ;
        RECT 2062.525 1114.320 2062.695 1114.490 ;
        RECT 2062.985 1114.320 2063.155 1114.490 ;
        RECT 2063.445 1114.320 2063.615 1114.490 ;
        RECT 2063.905 1114.320 2064.075 1114.490 ;
        RECT 2064.365 1114.320 2064.535 1114.490 ;
        RECT 2064.825 1114.320 2064.995 1114.490 ;
        RECT 2065.285 1114.320 2065.455 1114.490 ;
        RECT 2065.745 1114.320 2065.915 1114.490 ;
        RECT 2066.205 1114.320 2066.375 1114.490 ;
        RECT 2066.665 1114.320 2066.835 1114.490 ;
        RECT 2067.125 1114.320 2067.295 1114.490 ;
        RECT 2067.585 1114.320 2067.755 1114.490 ;
        RECT 2068.045 1114.320 2068.215 1114.490 ;
        RECT 2068.505 1114.320 2068.675 1114.490 ;
        RECT 2068.965 1114.320 2069.135 1114.490 ;
        RECT 2069.425 1114.320 2069.595 1114.490 ;
        RECT 2069.885 1114.320 2070.055 1114.490 ;
        RECT 2070.345 1114.320 2070.515 1114.490 ;
        RECT 2070.805 1114.320 2070.975 1114.490 ;
        RECT 2071.265 1114.320 2071.435 1114.490 ;
        RECT 2071.725 1114.320 2071.895 1114.490 ;
        RECT 2072.185 1114.320 2072.355 1114.490 ;
        RECT 2072.645 1114.320 2072.815 1114.490 ;
        RECT 2073.105 1114.320 2073.275 1114.490 ;
        RECT 2073.565 1114.320 2073.735 1114.490 ;
        RECT 2074.025 1114.320 2074.195 1114.490 ;
        RECT 2074.485 1114.320 2074.655 1114.490 ;
        RECT 2074.945 1114.320 2075.115 1114.490 ;
        RECT 2075.405 1114.320 2075.575 1114.490 ;
        RECT 2075.865 1114.320 2076.035 1114.490 ;
        RECT 2076.325 1114.320 2076.495 1114.490 ;
        RECT 2076.785 1114.320 2076.955 1114.490 ;
        RECT 2077.245 1114.320 2077.415 1114.490 ;
        RECT 2077.705 1114.320 2077.875 1114.490 ;
        RECT 2078.165 1114.320 2078.335 1114.490 ;
        RECT 2078.625 1114.320 2078.795 1114.490 ;
        RECT 2079.085 1114.320 2079.255 1114.490 ;
        RECT 2079.545 1114.320 2079.715 1114.490 ;
        RECT 2080.005 1114.320 2080.175 1114.490 ;
        RECT 2080.465 1114.320 2080.635 1114.490 ;
        RECT 2080.925 1114.320 2081.095 1114.490 ;
        RECT 2081.385 1114.320 2081.555 1114.490 ;
        RECT 2081.845 1114.320 2082.015 1114.490 ;
        RECT 2082.305 1114.320 2082.475 1114.490 ;
        RECT 2082.765 1114.320 2082.935 1114.490 ;
        RECT 2083.225 1114.320 2083.395 1114.490 ;
        RECT 2083.685 1114.320 2083.855 1114.490 ;
        RECT 2084.145 1114.320 2084.315 1114.490 ;
        RECT 2084.605 1114.320 2084.775 1114.490 ;
        RECT 2085.065 1114.320 2085.235 1114.490 ;
        RECT 2085.525 1114.320 2085.695 1114.490 ;
        RECT 2085.985 1114.320 2086.155 1114.490 ;
        RECT 2086.445 1114.320 2086.615 1114.490 ;
        RECT 2086.905 1114.320 2087.075 1114.490 ;
        RECT 2087.365 1114.320 2087.535 1114.490 ;
        RECT 2087.825 1114.320 2087.995 1114.490 ;
        RECT 2088.285 1114.320 2088.455 1114.490 ;
        RECT 2088.745 1114.320 2088.915 1114.490 ;
        RECT 2089.205 1114.320 2089.375 1114.490 ;
        RECT 2089.665 1114.320 2089.835 1114.490 ;
        RECT 2090.125 1114.320 2090.295 1114.490 ;
        RECT 2090.585 1114.320 2090.755 1114.490 ;
        RECT 2091.045 1114.320 2091.215 1114.490 ;
        RECT 2091.505 1114.320 2091.675 1114.490 ;
        RECT 2091.965 1114.320 2092.135 1114.490 ;
        RECT 2092.425 1114.320 2092.595 1114.490 ;
        RECT 2092.885 1114.320 2093.055 1114.490 ;
        RECT 2093.345 1114.320 2093.515 1114.490 ;
        RECT 2093.805 1114.320 2093.975 1114.490 ;
        RECT 2094.265 1114.320 2094.435 1114.490 ;
        RECT 2094.725 1114.320 2094.895 1114.490 ;
      LAYER met1 ;
        RECT 1969.000 1114.165 2095.040 1114.645 ;
      LAYER via ;
        RECT 2025.150 1114.245 2026.935 1114.545 ;
      LAYER met2 ;
        RECT 2025.110 1114.185 2026.975 1114.615 ;
      LAYER via2 ;
        RECT 2025.150 1114.245 2026.935 1114.545 ;
      LAYER met3 ;
        RECT 2025.120 1109.800 2026.970 1114.615 ;
    END
    PORT
      LAYER li1 ;
        RECT 201.515 1762.750 201.685 1762.920 ;
        RECT 201.515 1762.290 201.685 1762.460 ;
        RECT 201.515 1761.830 201.685 1762.000 ;
        RECT 201.515 1761.370 201.685 1761.540 ;
        RECT 201.515 1760.910 201.685 1761.080 ;
        RECT 201.515 1760.450 201.685 1760.620 ;
        RECT 201.515 1759.990 201.685 1760.160 ;
        RECT 201.515 1759.530 201.685 1759.700 ;
        RECT 201.515 1759.070 201.685 1759.240 ;
        RECT 201.515 1758.610 201.685 1758.780 ;
        RECT 201.515 1758.150 201.685 1758.320 ;
        RECT 201.515 1757.690 201.685 1757.860 ;
        RECT 201.515 1757.230 201.685 1757.400 ;
        RECT 201.515 1756.770 201.685 1756.940 ;
        RECT 201.515 1756.310 201.685 1756.480 ;
        RECT 201.515 1755.850 201.685 1756.020 ;
        RECT 201.515 1755.390 201.685 1755.560 ;
        RECT 201.515 1754.930 201.685 1755.100 ;
        RECT 201.515 1754.470 201.685 1754.640 ;
        RECT 201.515 1754.010 201.685 1754.180 ;
        RECT 201.515 1753.550 201.685 1753.720 ;
        RECT 201.515 1753.090 201.685 1753.260 ;
        RECT 201.515 1752.630 201.685 1752.800 ;
        RECT 201.515 1752.170 201.685 1752.340 ;
        RECT 201.515 1751.710 201.685 1751.880 ;
        RECT 201.515 1751.250 201.685 1751.420 ;
        RECT 201.515 1750.790 201.685 1750.960 ;
        RECT 201.515 1750.330 201.685 1750.500 ;
        RECT 201.515 1749.870 201.685 1750.040 ;
        RECT 201.515 1749.410 201.685 1749.580 ;
        RECT 201.515 1748.950 201.685 1749.120 ;
        RECT 201.515 1748.490 201.685 1748.660 ;
        RECT 201.515 1748.030 201.685 1748.200 ;
        RECT 201.515 1747.570 201.685 1747.740 ;
        RECT 201.515 1747.110 201.685 1747.280 ;
        RECT 201.515 1746.650 201.685 1746.820 ;
        RECT 201.515 1746.190 201.685 1746.360 ;
        RECT 201.515 1745.730 201.685 1745.900 ;
        RECT 201.515 1745.270 201.685 1745.440 ;
        RECT 201.515 1744.810 201.685 1744.980 ;
        RECT 201.515 1744.350 201.685 1744.520 ;
        RECT 201.515 1743.890 201.685 1744.060 ;
        RECT 201.515 1743.430 201.685 1743.600 ;
        RECT 201.515 1742.970 201.685 1743.140 ;
        RECT 201.515 1742.510 201.685 1742.680 ;
        RECT 201.515 1742.050 201.685 1742.220 ;
        RECT 201.515 1741.590 201.685 1741.760 ;
        RECT 201.515 1741.130 201.685 1741.300 ;
        RECT 201.515 1740.670 201.685 1740.840 ;
        RECT 201.515 1740.210 201.685 1740.380 ;
        RECT 201.515 1739.750 201.685 1739.920 ;
        RECT 201.515 1739.290 201.685 1739.460 ;
        RECT 201.515 1738.830 201.685 1739.000 ;
        RECT 201.515 1738.370 201.685 1738.540 ;
        RECT 201.515 1737.910 201.685 1738.080 ;
        RECT 201.515 1737.450 201.685 1737.620 ;
        RECT 201.515 1736.990 201.685 1737.160 ;
        RECT 201.515 1736.530 201.685 1736.700 ;
        RECT 201.515 1736.070 201.685 1736.240 ;
        RECT 201.515 1735.610 201.685 1735.780 ;
        RECT 201.515 1735.150 201.685 1735.320 ;
        RECT 201.515 1734.690 201.685 1734.860 ;
        RECT 201.515 1734.230 201.685 1734.400 ;
        RECT 201.515 1733.770 201.685 1733.940 ;
        RECT 201.515 1733.310 201.685 1733.480 ;
        RECT 201.515 1732.850 201.685 1733.020 ;
        RECT 201.515 1732.390 201.685 1732.560 ;
        RECT 201.515 1731.930 201.685 1732.100 ;
        RECT 201.515 1731.470 201.685 1731.640 ;
        RECT 201.515 1731.010 201.685 1731.180 ;
        RECT 201.515 1730.550 201.685 1730.720 ;
        RECT 201.515 1730.090 201.685 1730.260 ;
        RECT 201.515 1729.630 201.685 1729.800 ;
        RECT 201.515 1729.170 201.685 1729.340 ;
        RECT 201.515 1728.710 201.685 1728.880 ;
        RECT 201.515 1728.250 201.685 1728.420 ;
        RECT 201.515 1727.790 201.685 1727.960 ;
        RECT 201.515 1727.330 201.685 1727.500 ;
        RECT 201.515 1726.870 201.685 1727.040 ;
        RECT 201.515 1726.410 201.685 1726.580 ;
        RECT 201.515 1725.950 201.685 1726.120 ;
        RECT 201.515 1725.490 201.685 1725.660 ;
        RECT 201.515 1725.030 201.685 1725.200 ;
        RECT 201.515 1724.570 201.685 1724.740 ;
        RECT 201.515 1724.110 201.685 1724.280 ;
        RECT 201.515 1723.650 201.685 1723.820 ;
        RECT 201.515 1723.190 201.685 1723.360 ;
        RECT 201.515 1722.730 201.685 1722.900 ;
        RECT 201.515 1722.270 201.685 1722.440 ;
        RECT 201.515 1721.810 201.685 1721.980 ;
        RECT 201.515 1721.350 201.685 1721.520 ;
        RECT 201.515 1720.890 201.685 1721.060 ;
        RECT 201.515 1720.430 201.685 1720.600 ;
        RECT 201.515 1719.970 201.685 1720.140 ;
        RECT 201.515 1719.510 201.685 1719.680 ;
        RECT 201.515 1719.050 201.685 1719.220 ;
        RECT 201.515 1718.590 201.685 1718.760 ;
        RECT 201.515 1718.130 201.685 1718.300 ;
        RECT 201.515 1717.670 201.685 1717.840 ;
        RECT 201.515 1717.210 201.685 1717.380 ;
        RECT 201.515 1716.750 201.685 1716.920 ;
        RECT 201.515 1716.290 201.685 1716.460 ;
        RECT 201.515 1715.830 201.685 1716.000 ;
        RECT 201.515 1715.370 201.685 1715.540 ;
        RECT 201.515 1714.910 201.685 1715.080 ;
        RECT 201.515 1714.450 201.685 1714.620 ;
        RECT 201.515 1713.990 201.685 1714.160 ;
        RECT 201.515 1713.530 201.685 1713.700 ;
        RECT 201.515 1713.070 201.685 1713.240 ;
        RECT 201.515 1712.610 201.685 1712.780 ;
        RECT 201.515 1712.150 201.685 1712.320 ;
        RECT 201.515 1711.690 201.685 1711.860 ;
        RECT 201.515 1711.230 201.685 1711.400 ;
        RECT 201.515 1710.770 201.685 1710.940 ;
        RECT 201.515 1710.310 201.685 1710.480 ;
        RECT 201.515 1709.850 201.685 1710.020 ;
        RECT 201.515 1709.390 201.685 1709.560 ;
        RECT 201.515 1708.930 201.685 1709.100 ;
        RECT 201.515 1708.470 201.685 1708.640 ;
        RECT 201.515 1708.010 201.685 1708.180 ;
        RECT 201.515 1707.550 201.685 1707.720 ;
        RECT 201.515 1707.090 201.685 1707.260 ;
        RECT 201.515 1706.630 201.685 1706.800 ;
        RECT 201.515 1706.170 201.685 1706.340 ;
        RECT 201.515 1705.710 201.685 1705.880 ;
        RECT 201.515 1705.250 201.685 1705.420 ;
        RECT 201.515 1704.790 201.685 1704.960 ;
        RECT 201.515 1704.330 201.685 1704.500 ;
        RECT 201.515 1703.870 201.685 1704.040 ;
        RECT 201.515 1703.410 201.685 1703.580 ;
        RECT 201.515 1702.950 201.685 1703.120 ;
        RECT 201.515 1702.490 201.685 1702.660 ;
        RECT 201.515 1702.030 201.685 1702.200 ;
        RECT 201.515 1701.570 201.685 1701.740 ;
        RECT 201.515 1701.110 201.685 1701.280 ;
        RECT 201.515 1700.650 201.685 1700.820 ;
        RECT 201.515 1700.190 201.685 1700.360 ;
        RECT 201.515 1699.730 201.685 1699.900 ;
        RECT 201.515 1699.270 201.685 1699.440 ;
        RECT 201.515 1698.810 201.685 1698.980 ;
        RECT 201.515 1698.350 201.685 1698.520 ;
        RECT 201.515 1697.890 201.685 1698.060 ;
        RECT 201.515 1697.430 201.685 1697.600 ;
        RECT 201.515 1696.970 201.685 1697.140 ;
        RECT 201.515 1696.510 201.685 1696.680 ;
        RECT 201.515 1696.050 201.685 1696.220 ;
        RECT 201.515 1695.590 201.685 1695.760 ;
        RECT 201.515 1695.130 201.685 1695.300 ;
        RECT 201.515 1694.670 201.685 1694.840 ;
        RECT 201.515 1694.210 201.685 1694.380 ;
        RECT 201.515 1693.750 201.685 1693.920 ;
        RECT 201.515 1693.290 201.685 1693.460 ;
        RECT 201.515 1692.830 201.685 1693.000 ;
        RECT 201.515 1692.370 201.685 1692.540 ;
        RECT 201.515 1691.910 201.685 1692.080 ;
        RECT 201.515 1691.450 201.685 1691.620 ;
        RECT 201.515 1690.990 201.685 1691.160 ;
        RECT 201.515 1690.530 201.685 1690.700 ;
        RECT 201.515 1690.070 201.685 1690.240 ;
        RECT 201.515 1689.610 201.685 1689.780 ;
        RECT 201.515 1689.150 201.685 1689.320 ;
        RECT 201.515 1688.690 201.685 1688.860 ;
        RECT 201.515 1688.230 201.685 1688.400 ;
        RECT 201.515 1687.770 201.685 1687.940 ;
        RECT 201.515 1687.310 201.685 1687.480 ;
        RECT 201.515 1686.850 201.685 1687.020 ;
        RECT 201.515 1686.390 201.685 1686.560 ;
        RECT 201.515 1685.930 201.685 1686.100 ;
        RECT 201.515 1685.470 201.685 1685.640 ;
        RECT 201.515 1685.010 201.685 1685.180 ;
        RECT 201.515 1684.550 201.685 1684.720 ;
        RECT 201.515 1684.090 201.685 1684.260 ;
        RECT 201.515 1683.630 201.685 1683.800 ;
        RECT 201.515 1683.170 201.685 1683.340 ;
        RECT 201.515 1682.710 201.685 1682.880 ;
        RECT 201.515 1682.250 201.685 1682.420 ;
        RECT 201.515 1681.790 201.685 1681.960 ;
        RECT 201.515 1681.330 201.685 1681.500 ;
        RECT 201.515 1680.870 201.685 1681.040 ;
        RECT 201.515 1680.410 201.685 1680.580 ;
        RECT 201.515 1679.950 201.685 1680.120 ;
        RECT 201.515 1679.490 201.685 1679.660 ;
        RECT 201.515 1679.030 201.685 1679.200 ;
        RECT 201.515 1678.570 201.685 1678.740 ;
        RECT 201.515 1678.110 201.685 1678.280 ;
        RECT 201.515 1677.650 201.685 1677.820 ;
        RECT 201.515 1677.190 201.685 1677.360 ;
        RECT 201.515 1676.730 201.685 1676.900 ;
        RECT 201.515 1676.270 201.685 1676.440 ;
        RECT 201.515 1675.810 201.685 1675.980 ;
        RECT 201.515 1675.350 201.685 1675.520 ;
        RECT 201.515 1674.890 201.685 1675.060 ;
        RECT 201.515 1674.430 201.685 1674.600 ;
        RECT 201.515 1673.970 201.685 1674.140 ;
        RECT 201.515 1673.510 201.685 1673.680 ;
        RECT 201.515 1673.050 201.685 1673.220 ;
      LAYER met1 ;
        RECT 201.360 1672.905 201.840 1763.065 ;
      LAYER via ;
        RECT 201.455 1716.855 201.755 1718.640 ;
      LAYER met2 ;
        RECT 201.395 1716.815 201.825 1718.680 ;
      LAYER via2 ;
        RECT 201.455 1716.855 201.755 1718.640 ;
      LAYER met3 ;
        RECT 197.010 1716.820 201.825 1718.670 ;
    END
    PORT
      LAYER li1 ;
        RECT 201.405 3053.655 201.575 3053.825 ;
        RECT 201.405 3053.195 201.575 3053.365 ;
        RECT 201.405 3052.735 201.575 3052.905 ;
        RECT 201.405 3052.275 201.575 3052.445 ;
        RECT 201.405 3051.815 201.575 3051.985 ;
        RECT 201.405 3051.355 201.575 3051.525 ;
        RECT 201.405 3050.895 201.575 3051.065 ;
        RECT 201.405 3050.435 201.575 3050.605 ;
        RECT 201.405 3049.975 201.575 3050.145 ;
        RECT 201.405 3049.515 201.575 3049.685 ;
        RECT 201.405 3049.055 201.575 3049.225 ;
        RECT 201.405 3048.595 201.575 3048.765 ;
        RECT 201.405 3048.135 201.575 3048.305 ;
        RECT 201.405 3047.675 201.575 3047.845 ;
        RECT 201.405 3047.215 201.575 3047.385 ;
        RECT 201.405 3046.755 201.575 3046.925 ;
        RECT 201.405 3046.295 201.575 3046.465 ;
        RECT 201.405 3045.835 201.575 3046.005 ;
        RECT 201.405 3045.375 201.575 3045.545 ;
        RECT 201.405 3044.915 201.575 3045.085 ;
        RECT 201.405 3044.455 201.575 3044.625 ;
        RECT 201.405 3043.995 201.575 3044.165 ;
        RECT 201.405 3043.535 201.575 3043.705 ;
        RECT 201.405 3043.075 201.575 3043.245 ;
        RECT 201.405 3042.615 201.575 3042.785 ;
        RECT 201.405 3042.155 201.575 3042.325 ;
        RECT 201.405 3041.695 201.575 3041.865 ;
        RECT 201.405 3041.235 201.575 3041.405 ;
        RECT 201.405 3040.775 201.575 3040.945 ;
        RECT 201.405 3040.315 201.575 3040.485 ;
        RECT 201.405 3039.855 201.575 3040.025 ;
        RECT 201.405 3039.395 201.575 3039.565 ;
        RECT 201.405 3038.935 201.575 3039.105 ;
        RECT 201.405 3038.475 201.575 3038.645 ;
        RECT 201.405 3038.015 201.575 3038.185 ;
        RECT 201.405 3037.555 201.575 3037.725 ;
        RECT 201.405 3037.095 201.575 3037.265 ;
        RECT 201.405 3036.635 201.575 3036.805 ;
        RECT 201.405 3036.175 201.575 3036.345 ;
        RECT 201.405 3035.715 201.575 3035.885 ;
        RECT 201.405 3035.255 201.575 3035.425 ;
        RECT 201.405 3034.795 201.575 3034.965 ;
        RECT 201.405 3034.335 201.575 3034.505 ;
        RECT 201.405 3033.875 201.575 3034.045 ;
        RECT 201.405 3033.415 201.575 3033.585 ;
        RECT 201.405 3032.955 201.575 3033.125 ;
        RECT 201.405 3032.495 201.575 3032.665 ;
        RECT 201.405 3032.035 201.575 3032.205 ;
        RECT 201.405 3031.575 201.575 3031.745 ;
        RECT 201.405 3031.115 201.575 3031.285 ;
        RECT 201.405 3030.655 201.575 3030.825 ;
        RECT 201.405 3030.195 201.575 3030.365 ;
        RECT 201.405 3029.735 201.575 3029.905 ;
        RECT 201.405 3029.275 201.575 3029.445 ;
        RECT 201.405 3028.815 201.575 3028.985 ;
        RECT 201.405 3028.355 201.575 3028.525 ;
        RECT 201.405 3027.895 201.575 3028.065 ;
        RECT 201.405 3027.435 201.575 3027.605 ;
        RECT 201.405 3026.975 201.575 3027.145 ;
        RECT 201.405 3026.515 201.575 3026.685 ;
        RECT 201.405 3026.055 201.575 3026.225 ;
        RECT 201.405 3025.595 201.575 3025.765 ;
        RECT 201.405 3025.135 201.575 3025.305 ;
        RECT 201.405 3024.675 201.575 3024.845 ;
        RECT 201.405 3024.215 201.575 3024.385 ;
        RECT 201.405 3023.755 201.575 3023.925 ;
        RECT 201.405 3023.295 201.575 3023.465 ;
        RECT 201.405 3022.835 201.575 3023.005 ;
        RECT 201.405 3022.375 201.575 3022.545 ;
        RECT 201.405 3021.915 201.575 3022.085 ;
        RECT 201.405 3021.455 201.575 3021.625 ;
        RECT 201.405 3020.995 201.575 3021.165 ;
        RECT 201.405 3020.535 201.575 3020.705 ;
        RECT 201.405 3020.075 201.575 3020.245 ;
        RECT 201.405 3019.615 201.575 3019.785 ;
        RECT 201.405 3019.155 201.575 3019.325 ;
        RECT 201.405 3018.695 201.575 3018.865 ;
        RECT 201.405 3018.235 201.575 3018.405 ;
        RECT 201.405 3017.775 201.575 3017.945 ;
        RECT 201.405 3017.315 201.575 3017.485 ;
        RECT 201.405 3016.855 201.575 3017.025 ;
        RECT 201.405 3016.395 201.575 3016.565 ;
        RECT 201.405 3015.935 201.575 3016.105 ;
        RECT 201.405 3015.475 201.575 3015.645 ;
        RECT 201.405 3015.015 201.575 3015.185 ;
        RECT 201.405 3014.555 201.575 3014.725 ;
        RECT 201.405 3014.095 201.575 3014.265 ;
        RECT 201.405 3013.635 201.575 3013.805 ;
        RECT 201.405 3013.175 201.575 3013.345 ;
        RECT 201.405 3012.715 201.575 3012.885 ;
        RECT 201.405 3012.255 201.575 3012.425 ;
        RECT 201.405 3011.795 201.575 3011.965 ;
        RECT 201.405 3011.335 201.575 3011.505 ;
        RECT 201.405 3010.875 201.575 3011.045 ;
        RECT 201.405 3010.415 201.575 3010.585 ;
        RECT 201.405 3009.955 201.575 3010.125 ;
        RECT 201.405 3009.495 201.575 3009.665 ;
        RECT 201.405 3009.035 201.575 3009.205 ;
        RECT 201.405 3008.575 201.575 3008.745 ;
        RECT 201.405 3008.115 201.575 3008.285 ;
        RECT 201.405 3007.655 201.575 3007.825 ;
        RECT 201.405 3007.195 201.575 3007.365 ;
        RECT 201.405 3006.735 201.575 3006.905 ;
        RECT 201.405 3006.275 201.575 3006.445 ;
        RECT 201.405 3005.815 201.575 3005.985 ;
        RECT 201.405 3005.355 201.575 3005.525 ;
        RECT 201.405 3004.895 201.575 3005.065 ;
        RECT 201.405 3004.435 201.575 3004.605 ;
        RECT 201.405 3003.975 201.575 3004.145 ;
        RECT 201.405 3003.515 201.575 3003.685 ;
        RECT 201.405 3003.055 201.575 3003.225 ;
        RECT 201.405 3002.595 201.575 3002.765 ;
        RECT 201.405 3002.135 201.575 3002.305 ;
        RECT 201.405 3001.675 201.575 3001.845 ;
        RECT 201.405 3001.215 201.575 3001.385 ;
        RECT 201.405 3000.755 201.575 3000.925 ;
        RECT 201.405 3000.295 201.575 3000.465 ;
        RECT 201.405 2999.835 201.575 3000.005 ;
        RECT 201.405 2999.375 201.575 2999.545 ;
        RECT 201.405 2998.915 201.575 2999.085 ;
        RECT 201.405 2998.455 201.575 2998.625 ;
        RECT 201.405 2997.995 201.575 2998.165 ;
        RECT 201.405 2997.535 201.575 2997.705 ;
        RECT 201.405 2997.075 201.575 2997.245 ;
        RECT 201.405 2996.615 201.575 2996.785 ;
        RECT 201.405 2996.155 201.575 2996.325 ;
        RECT 201.405 2995.695 201.575 2995.865 ;
        RECT 201.405 2995.235 201.575 2995.405 ;
        RECT 201.405 2994.775 201.575 2994.945 ;
        RECT 201.405 2994.315 201.575 2994.485 ;
        RECT 201.405 2993.855 201.575 2994.025 ;
        RECT 201.405 2993.395 201.575 2993.565 ;
        RECT 201.405 2992.935 201.575 2993.105 ;
        RECT 201.405 2992.475 201.575 2992.645 ;
        RECT 201.405 2992.015 201.575 2992.185 ;
        RECT 201.405 2991.555 201.575 2991.725 ;
        RECT 201.405 2991.095 201.575 2991.265 ;
        RECT 201.405 2990.635 201.575 2990.805 ;
        RECT 201.405 2990.175 201.575 2990.345 ;
        RECT 201.405 2989.715 201.575 2989.885 ;
        RECT 201.405 2989.255 201.575 2989.425 ;
        RECT 201.405 2988.795 201.575 2988.965 ;
        RECT 201.405 2988.335 201.575 2988.505 ;
        RECT 201.405 2987.875 201.575 2988.045 ;
      LAYER met1 ;
        RECT 201.250 2987.730 201.730 3053.970 ;
      LAYER via ;
        RECT 201.360 3026.050 201.660 3027.835 ;
      LAYER met2 ;
        RECT 201.300 3026.010 201.730 3027.875 ;
      LAYER via2 ;
        RECT 201.360 3026.050 201.660 3027.835 ;
      LAYER met3 ;
        RECT 196.915 3026.015 201.730 3027.865 ;
    END
    PORT
      LAYER li1 ;
        RECT 201.280 4456.885 201.450 4457.055 ;
        RECT 201.280 4456.425 201.450 4456.595 ;
        RECT 201.280 4455.965 201.450 4456.135 ;
        RECT 201.280 4455.505 201.450 4455.675 ;
        RECT 201.280 4455.045 201.450 4455.215 ;
        RECT 201.280 4454.585 201.450 4454.755 ;
        RECT 201.280 4454.125 201.450 4454.295 ;
        RECT 201.280 4453.665 201.450 4453.835 ;
        RECT 201.280 4453.205 201.450 4453.375 ;
        RECT 201.280 4452.745 201.450 4452.915 ;
        RECT 201.280 4452.285 201.450 4452.455 ;
        RECT 201.280 4451.825 201.450 4451.995 ;
        RECT 201.280 4451.365 201.450 4451.535 ;
        RECT 201.280 4450.905 201.450 4451.075 ;
        RECT 201.280 4450.445 201.450 4450.615 ;
        RECT 201.280 4449.985 201.450 4450.155 ;
        RECT 201.280 4449.525 201.450 4449.695 ;
        RECT 201.280 4449.065 201.450 4449.235 ;
        RECT 201.280 4448.605 201.450 4448.775 ;
        RECT 201.280 4448.145 201.450 4448.315 ;
        RECT 201.280 4447.685 201.450 4447.855 ;
        RECT 201.280 4447.225 201.450 4447.395 ;
        RECT 201.280 4446.765 201.450 4446.935 ;
        RECT 201.280 4446.305 201.450 4446.475 ;
        RECT 201.280 4445.845 201.450 4446.015 ;
        RECT 201.280 4445.385 201.450 4445.555 ;
        RECT 201.280 4444.925 201.450 4445.095 ;
        RECT 201.280 4444.465 201.450 4444.635 ;
        RECT 201.280 4444.005 201.450 4444.175 ;
        RECT 201.280 4443.545 201.450 4443.715 ;
        RECT 201.280 4443.085 201.450 4443.255 ;
        RECT 201.280 4442.625 201.450 4442.795 ;
        RECT 201.280 4442.165 201.450 4442.335 ;
        RECT 201.280 4441.705 201.450 4441.875 ;
        RECT 201.280 4441.245 201.450 4441.415 ;
        RECT 201.280 4440.785 201.450 4440.955 ;
        RECT 201.280 4440.325 201.450 4440.495 ;
        RECT 201.280 4439.865 201.450 4440.035 ;
        RECT 201.280 4439.405 201.450 4439.575 ;
        RECT 201.280 4438.945 201.450 4439.115 ;
        RECT 201.280 4438.485 201.450 4438.655 ;
        RECT 201.280 4438.025 201.450 4438.195 ;
        RECT 201.280 4437.565 201.450 4437.735 ;
        RECT 201.280 4437.105 201.450 4437.275 ;
        RECT 201.280 4436.645 201.450 4436.815 ;
        RECT 201.280 4436.185 201.450 4436.355 ;
        RECT 201.280 4435.725 201.450 4435.895 ;
        RECT 201.280 4435.265 201.450 4435.435 ;
        RECT 201.280 4434.805 201.450 4434.975 ;
        RECT 201.280 4434.345 201.450 4434.515 ;
        RECT 201.280 4433.885 201.450 4434.055 ;
        RECT 201.280 4433.425 201.450 4433.595 ;
        RECT 201.280 4432.965 201.450 4433.135 ;
        RECT 201.280 4432.505 201.450 4432.675 ;
        RECT 201.280 4432.045 201.450 4432.215 ;
        RECT 201.280 4431.585 201.450 4431.755 ;
        RECT 201.280 4431.125 201.450 4431.295 ;
        RECT 201.280 4430.665 201.450 4430.835 ;
        RECT 201.280 4430.205 201.450 4430.375 ;
        RECT 201.280 4429.745 201.450 4429.915 ;
        RECT 201.280 4429.285 201.450 4429.455 ;
        RECT 201.280 4428.825 201.450 4428.995 ;
        RECT 201.280 4428.365 201.450 4428.535 ;
        RECT 201.280 4427.905 201.450 4428.075 ;
        RECT 201.280 4427.445 201.450 4427.615 ;
        RECT 201.280 4426.985 201.450 4427.155 ;
      LAYER met1 ;
        RECT 201.125 4426.840 201.605 4457.200 ;
      LAYER via ;
        RECT 201.205 4446.920 201.505 4448.705 ;
      LAYER met2 ;
        RECT 201.145 4446.880 201.575 4448.745 ;
      LAYER via2 ;
        RECT 201.205 4446.920 201.505 4448.705 ;
      LAYER met3 ;
        RECT 196.760 4446.885 201.575 4448.735 ;
    END
    PORT
      LAYER li1 ;
        RECT 3386.220 3572.085 3386.390 3572.255 ;
        RECT 3386.220 3571.625 3386.390 3571.795 ;
        RECT 3386.220 3571.165 3386.390 3571.335 ;
        RECT 3386.220 3570.705 3386.390 3570.875 ;
        RECT 3386.220 3570.245 3386.390 3570.415 ;
        RECT 3386.220 3569.785 3386.390 3569.955 ;
        RECT 3386.220 3569.325 3386.390 3569.495 ;
        RECT 3386.220 3568.865 3386.390 3569.035 ;
        RECT 3386.220 3568.405 3386.390 3568.575 ;
        RECT 3386.220 3567.945 3386.390 3568.115 ;
        RECT 3386.220 3567.485 3386.390 3567.655 ;
        RECT 3386.220 3567.025 3386.390 3567.195 ;
        RECT 3386.220 3566.565 3386.390 3566.735 ;
        RECT 3386.220 3566.105 3386.390 3566.275 ;
        RECT 3386.220 3565.645 3386.390 3565.815 ;
        RECT 3386.220 3565.185 3386.390 3565.355 ;
        RECT 3386.220 3564.725 3386.390 3564.895 ;
        RECT 3386.220 3564.265 3386.390 3564.435 ;
        RECT 3386.220 3563.805 3386.390 3563.975 ;
        RECT 3386.220 3563.345 3386.390 3563.515 ;
        RECT 3386.220 3562.885 3386.390 3563.055 ;
        RECT 3386.220 3562.425 3386.390 3562.595 ;
        RECT 3386.220 3561.965 3386.390 3562.135 ;
        RECT 3386.220 3561.505 3386.390 3561.675 ;
        RECT 3386.220 3561.045 3386.390 3561.215 ;
        RECT 3386.220 3560.585 3386.390 3560.755 ;
        RECT 3386.220 3560.125 3386.390 3560.295 ;
        RECT 3386.220 3559.665 3386.390 3559.835 ;
        RECT 3386.220 3559.205 3386.390 3559.375 ;
        RECT 3386.220 3558.745 3386.390 3558.915 ;
        RECT 3386.220 3558.285 3386.390 3558.455 ;
        RECT 3386.220 3557.825 3386.390 3557.995 ;
        RECT 3386.220 3557.365 3386.390 3557.535 ;
        RECT 3386.220 3556.905 3386.390 3557.075 ;
        RECT 3386.220 3556.445 3386.390 3556.615 ;
        RECT 3386.220 3555.985 3386.390 3556.155 ;
        RECT 3386.220 3555.525 3386.390 3555.695 ;
        RECT 3386.220 3555.065 3386.390 3555.235 ;
        RECT 3386.220 3554.605 3386.390 3554.775 ;
        RECT 3386.220 3554.145 3386.390 3554.315 ;
        RECT 3386.220 3553.685 3386.390 3553.855 ;
        RECT 3386.220 3553.225 3386.390 3553.395 ;
        RECT 3386.220 3552.765 3386.390 3552.935 ;
        RECT 3386.220 3552.305 3386.390 3552.475 ;
        RECT 3386.220 3551.845 3386.390 3552.015 ;
        RECT 3386.220 3551.385 3386.390 3551.555 ;
        RECT 3386.220 3550.925 3386.390 3551.095 ;
        RECT 3386.220 3550.465 3386.390 3550.635 ;
        RECT 3386.220 3550.005 3386.390 3550.175 ;
        RECT 3386.220 3549.545 3386.390 3549.715 ;
        RECT 3386.220 3549.085 3386.390 3549.255 ;
        RECT 3386.220 3548.625 3386.390 3548.795 ;
        RECT 3386.220 3548.165 3386.390 3548.335 ;
        RECT 3386.220 3547.705 3386.390 3547.875 ;
        RECT 3386.220 3547.245 3386.390 3547.415 ;
        RECT 3386.220 3546.785 3386.390 3546.955 ;
        RECT 3386.220 3546.325 3386.390 3546.495 ;
        RECT 3386.220 3545.865 3386.390 3546.035 ;
        RECT 3386.220 3545.405 3386.390 3545.575 ;
        RECT 3386.220 3544.945 3386.390 3545.115 ;
        RECT 3386.220 3544.485 3386.390 3544.655 ;
        RECT 3386.220 3544.025 3386.390 3544.195 ;
        RECT 3386.220 3543.565 3386.390 3543.735 ;
        RECT 3386.220 3543.105 3386.390 3543.275 ;
        RECT 3386.220 3542.645 3386.390 3542.815 ;
        RECT 3386.220 3542.185 3386.390 3542.355 ;
        RECT 3386.220 3541.725 3386.390 3541.895 ;
        RECT 3386.220 3541.265 3386.390 3541.435 ;
        RECT 3386.220 3540.805 3386.390 3540.975 ;
        RECT 3386.220 3540.345 3386.390 3540.515 ;
        RECT 3386.220 3539.885 3386.390 3540.055 ;
        RECT 3386.220 3539.425 3386.390 3539.595 ;
        RECT 3386.220 3538.965 3386.390 3539.135 ;
        RECT 3386.220 3538.505 3386.390 3538.675 ;
        RECT 3386.220 3538.045 3386.390 3538.215 ;
        RECT 3386.220 3537.585 3386.390 3537.755 ;
        RECT 3386.220 3537.125 3386.390 3537.295 ;
        RECT 3386.220 3536.665 3386.390 3536.835 ;
        RECT 3386.220 3536.205 3386.390 3536.375 ;
      LAYER met1 ;
        RECT 3386.065 3536.060 3386.545 3572.400 ;
      LAYER via ;
        RECT 3386.170 3550.500 3386.470 3552.285 ;
      LAYER met2 ;
        RECT 3386.100 3550.460 3386.530 3552.325 ;
      LAYER via2 ;
        RECT 3386.170 3550.500 3386.470 3552.285 ;
      LAYER met3 ;
        RECT 3386.100 3550.470 3390.915 3552.320 ;
    END
    PORT
      LAYER li1 ;
        RECT 3386.220 2267.965 3386.390 2268.135 ;
        RECT 3386.220 2267.505 3386.390 2267.675 ;
        RECT 3386.220 2267.045 3386.390 2267.215 ;
        RECT 3386.220 2266.585 3386.390 2266.755 ;
        RECT 3386.220 2266.125 3386.390 2266.295 ;
        RECT 3386.220 2265.665 3386.390 2265.835 ;
        RECT 3386.220 2265.205 3386.390 2265.375 ;
        RECT 3386.220 2264.745 3386.390 2264.915 ;
        RECT 3386.220 2264.285 3386.390 2264.455 ;
        RECT 3386.220 2263.825 3386.390 2263.995 ;
        RECT 3386.220 2263.365 3386.390 2263.535 ;
        RECT 3386.220 2262.905 3386.390 2263.075 ;
        RECT 3386.220 2262.445 3386.390 2262.615 ;
        RECT 3386.220 2261.985 3386.390 2262.155 ;
        RECT 3386.220 2261.525 3386.390 2261.695 ;
        RECT 3386.220 2261.065 3386.390 2261.235 ;
        RECT 3386.220 2260.605 3386.390 2260.775 ;
        RECT 3386.220 2260.145 3386.390 2260.315 ;
        RECT 3386.220 2259.685 3386.390 2259.855 ;
        RECT 3386.220 2259.225 3386.390 2259.395 ;
        RECT 3386.220 2258.765 3386.390 2258.935 ;
        RECT 3386.220 2258.305 3386.390 2258.475 ;
        RECT 3386.220 2257.845 3386.390 2258.015 ;
        RECT 3386.220 2257.385 3386.390 2257.555 ;
        RECT 3386.220 2256.925 3386.390 2257.095 ;
        RECT 3386.220 2256.465 3386.390 2256.635 ;
        RECT 3386.220 2256.005 3386.390 2256.175 ;
        RECT 3386.220 2255.545 3386.390 2255.715 ;
        RECT 3386.220 2255.085 3386.390 2255.255 ;
        RECT 3386.220 2254.625 3386.390 2254.795 ;
        RECT 3386.220 2254.165 3386.390 2254.335 ;
        RECT 3386.220 2253.705 3386.390 2253.875 ;
        RECT 3386.220 2253.245 3386.390 2253.415 ;
        RECT 3386.220 2252.785 3386.390 2252.955 ;
        RECT 3386.220 2252.325 3386.390 2252.495 ;
        RECT 3386.220 2251.865 3386.390 2252.035 ;
        RECT 3386.220 2251.405 3386.390 2251.575 ;
        RECT 3386.220 2250.945 3386.390 2251.115 ;
        RECT 3386.220 2250.485 3386.390 2250.655 ;
        RECT 3386.220 2250.025 3386.390 2250.195 ;
        RECT 3386.220 2249.565 3386.390 2249.735 ;
        RECT 3386.220 2249.105 3386.390 2249.275 ;
        RECT 3386.220 2248.645 3386.390 2248.815 ;
        RECT 3386.220 2248.185 3386.390 2248.355 ;
        RECT 3386.220 2247.725 3386.390 2247.895 ;
        RECT 3386.220 2247.265 3386.390 2247.435 ;
        RECT 3386.220 2246.805 3386.390 2246.975 ;
        RECT 3386.220 2246.345 3386.390 2246.515 ;
        RECT 3386.220 2245.885 3386.390 2246.055 ;
        RECT 3386.220 2245.425 3386.390 2245.595 ;
        RECT 3386.220 2244.965 3386.390 2245.135 ;
        RECT 3386.220 2244.505 3386.390 2244.675 ;
        RECT 3386.220 2244.045 3386.390 2244.215 ;
        RECT 3386.220 2243.585 3386.390 2243.755 ;
        RECT 3386.220 2243.125 3386.390 2243.295 ;
        RECT 3386.220 2242.665 3386.390 2242.835 ;
        RECT 3386.220 2242.205 3386.390 2242.375 ;
        RECT 3386.220 2241.745 3386.390 2241.915 ;
        RECT 3386.220 2241.285 3386.390 2241.455 ;
        RECT 3386.220 2240.825 3386.390 2240.995 ;
        RECT 3386.220 2240.365 3386.390 2240.535 ;
        RECT 3386.220 2239.905 3386.390 2240.075 ;
        RECT 3386.220 2239.445 3386.390 2239.615 ;
        RECT 3386.220 2238.985 3386.390 2239.155 ;
        RECT 3386.220 2238.525 3386.390 2238.695 ;
        RECT 3386.220 2238.065 3386.390 2238.235 ;
        RECT 3386.220 2237.605 3386.390 2237.775 ;
        RECT 3386.220 2237.145 3386.390 2237.315 ;
        RECT 3386.220 2236.685 3386.390 2236.855 ;
        RECT 3386.220 2236.225 3386.390 2236.395 ;
        RECT 3386.220 2235.765 3386.390 2235.935 ;
        RECT 3386.220 2235.305 3386.390 2235.475 ;
        RECT 3386.220 2234.845 3386.390 2235.015 ;
        RECT 3386.220 2234.385 3386.390 2234.555 ;
        RECT 3386.220 2233.925 3386.390 2234.095 ;
        RECT 3386.220 2233.465 3386.390 2233.635 ;
        RECT 3386.220 2233.005 3386.390 2233.175 ;
        RECT 3386.220 2232.545 3386.390 2232.715 ;
        RECT 3386.220 2232.085 3386.390 2232.255 ;
        RECT 3386.220 2231.625 3386.390 2231.795 ;
        RECT 3386.220 2231.165 3386.390 2231.335 ;
        RECT 3386.220 2230.705 3386.390 2230.875 ;
        RECT 3386.220 2230.245 3386.390 2230.415 ;
        RECT 3386.220 2229.785 3386.390 2229.955 ;
        RECT 3386.220 2229.325 3386.390 2229.495 ;
        RECT 3386.220 2228.865 3386.390 2229.035 ;
        RECT 3386.220 2228.405 3386.390 2228.575 ;
        RECT 3386.220 2227.945 3386.390 2228.115 ;
        RECT 3386.220 2227.485 3386.390 2227.655 ;
        RECT 3386.220 2227.025 3386.390 2227.195 ;
        RECT 3386.220 2226.565 3386.390 2226.735 ;
        RECT 3386.220 2226.105 3386.390 2226.275 ;
        RECT 3386.220 2225.645 3386.390 2225.815 ;
        RECT 3386.220 2225.185 3386.390 2225.355 ;
        RECT 3386.220 2224.725 3386.390 2224.895 ;
        RECT 3386.220 2224.265 3386.390 2224.435 ;
        RECT 3386.220 2223.805 3386.390 2223.975 ;
        RECT 3386.220 2223.345 3386.390 2223.515 ;
        RECT 3386.220 2222.885 3386.390 2223.055 ;
        RECT 3386.220 2222.425 3386.390 2222.595 ;
        RECT 3386.220 2221.965 3386.390 2222.135 ;
        RECT 3386.220 2221.505 3386.390 2221.675 ;
        RECT 3386.220 2221.045 3386.390 2221.215 ;
        RECT 3386.220 2220.585 3386.390 2220.755 ;
        RECT 3386.220 2220.125 3386.390 2220.295 ;
        RECT 3386.220 2219.665 3386.390 2219.835 ;
        RECT 3386.220 2219.205 3386.390 2219.375 ;
        RECT 3386.220 2218.745 3386.390 2218.915 ;
        RECT 3386.220 2218.285 3386.390 2218.455 ;
        RECT 3386.220 2217.825 3386.390 2217.995 ;
        RECT 3386.220 2217.365 3386.390 2217.535 ;
        RECT 3386.220 2216.905 3386.390 2217.075 ;
        RECT 3386.220 2216.445 3386.390 2216.615 ;
        RECT 3386.220 2215.985 3386.390 2216.155 ;
        RECT 3386.220 2215.525 3386.390 2215.695 ;
        RECT 3386.220 2215.065 3386.390 2215.235 ;
        RECT 3386.220 2214.605 3386.390 2214.775 ;
        RECT 3386.220 2214.145 3386.390 2214.315 ;
        RECT 3386.220 2213.685 3386.390 2213.855 ;
        RECT 3386.220 2213.225 3386.390 2213.395 ;
        RECT 3386.220 2212.765 3386.390 2212.935 ;
        RECT 3386.220 2212.305 3386.390 2212.475 ;
        RECT 3386.220 2211.845 3386.390 2212.015 ;
        RECT 3386.220 2211.385 3386.390 2211.555 ;
        RECT 3386.220 2210.925 3386.390 2211.095 ;
        RECT 3386.220 2210.465 3386.390 2210.635 ;
        RECT 3386.220 2210.005 3386.390 2210.175 ;
        RECT 3386.220 2209.545 3386.390 2209.715 ;
        RECT 3386.220 2209.085 3386.390 2209.255 ;
        RECT 3386.220 2208.625 3386.390 2208.795 ;
        RECT 3386.220 2208.165 3386.390 2208.335 ;
        RECT 3386.220 2207.705 3386.390 2207.875 ;
        RECT 3386.220 2207.245 3386.390 2207.415 ;
        RECT 3386.220 2206.785 3386.390 2206.955 ;
        RECT 3386.220 2206.325 3386.390 2206.495 ;
        RECT 3386.220 2205.865 3386.390 2206.035 ;
        RECT 3386.220 2205.405 3386.390 2205.575 ;
        RECT 3386.220 2204.945 3386.390 2205.115 ;
        RECT 3386.220 2204.485 3386.390 2204.655 ;
        RECT 3386.220 2204.025 3386.390 2204.195 ;
        RECT 3386.220 2203.565 3386.390 2203.735 ;
        RECT 3386.220 2203.105 3386.390 2203.275 ;
        RECT 3386.220 2202.645 3386.390 2202.815 ;
        RECT 3386.220 2202.185 3386.390 2202.355 ;
        RECT 3386.220 2201.725 3386.390 2201.895 ;
        RECT 3386.220 2201.265 3386.390 2201.435 ;
        RECT 3386.220 2200.805 3386.390 2200.975 ;
        RECT 3386.220 2200.345 3386.390 2200.515 ;
        RECT 3386.220 2199.885 3386.390 2200.055 ;
        RECT 3386.220 2199.425 3386.390 2199.595 ;
        RECT 3386.220 2198.965 3386.390 2199.135 ;
        RECT 3386.220 2198.505 3386.390 2198.675 ;
        RECT 3386.220 2198.045 3386.390 2198.215 ;
        RECT 3386.220 2197.585 3386.390 2197.755 ;
        RECT 3386.220 2197.125 3386.390 2197.295 ;
        RECT 3386.220 2196.665 3386.390 2196.835 ;
        RECT 3386.220 2196.205 3386.390 2196.375 ;
      LAYER met1 ;
        RECT 3386.065 2196.060 3386.545 2268.280 ;
      LAYER via ;
        RECT 3386.130 2234.495 3386.430 2236.280 ;
      LAYER met2 ;
        RECT 3386.060 2234.455 3386.490 2236.320 ;
      LAYER via2 ;
        RECT 3386.130 2234.495 3386.430 2236.280 ;
      LAYER met3 ;
        RECT 3386.060 2234.465 3390.875 2236.315 ;
    END
  END vccd
  OBS
      LAYER pwell ;
        RECT 2088.490 4987.595 2088.660 4987.785 ;
        RECT 2082.845 4986.725 2083.275 4987.510 ;
        RECT 2083.675 4986.685 2088.805 4987.595 ;
        RECT 2088.825 4986.725 2089.255 4987.510 ;
        RECT 3318.495 4987.185 3318.665 4987.375 ;
        RECT 3324.475 4987.185 3324.645 4987.375 ;
        RECT 3330.455 4987.185 3330.625 4987.375 ;
        RECT 3336.435 4987.185 3336.605 4987.375 ;
        RECT 835.260 4985.970 835.430 4986.160 ;
        RECT 841.240 4985.970 841.410 4986.160 ;
        RECT 847.220 4985.970 847.390 4986.160 ;
        RECT 834.665 4985.100 835.095 4985.885 ;
        RECT 835.115 4985.060 840.245 4985.970 ;
        RECT 840.645 4985.100 841.075 4985.885 ;
        RECT 841.095 4985.060 846.225 4985.970 ;
        RECT 846.625 4985.100 847.055 4985.885 ;
        RECT 847.075 4985.060 852.205 4985.970 ;
        RECT 852.605 4985.100 853.035 4985.885 ;
      LAYER nwell ;
        RECT 834.460 4981.940 853.240 4984.770 ;
        RECT 2082.640 4983.565 2089.460 4986.395 ;
      LAYER pwell ;
        RECT 3312.850 4986.315 3313.280 4987.100 ;
        RECT 3313.680 4986.275 3318.810 4987.185 ;
        RECT 3318.830 4986.315 3319.260 4987.100 ;
        RECT 3319.660 4986.275 3324.790 4987.185 ;
        RECT 3324.810 4986.315 3325.240 4987.100 ;
        RECT 3325.640 4986.275 3330.770 4987.185 ;
        RECT 3330.790 4986.315 3331.220 4987.100 ;
        RECT 3331.620 4986.275 3336.750 4987.185 ;
        RECT 3336.770 4986.315 3337.200 4987.100 ;
        RECT 2082.845 4982.450 2083.275 4983.235 ;
        RECT 2083.295 4982.365 2088.425 4983.275 ;
        RECT 2088.825 4982.450 2089.255 4983.235 ;
      LAYER nwell ;
        RECT 3312.645 4983.155 3337.405 4985.985 ;
      LAYER pwell ;
        RECT 2083.440 4982.175 2083.610 4982.365 ;
        RECT 3312.850 4982.040 3313.280 4982.825 ;
        RECT 3313.300 4981.955 3318.430 4982.865 ;
        RECT 3318.830 4982.040 3319.260 4982.825 ;
        RECT 3319.280 4981.955 3324.410 4982.865 ;
        RECT 3324.810 4982.040 3325.240 4982.825 ;
        RECT 3325.260 4981.955 3330.390 4982.865 ;
        RECT 3330.790 4982.040 3331.220 4982.825 ;
        RECT 3331.240 4981.955 3336.370 4982.865 ;
        RECT 3336.770 4982.040 3337.200 4982.825 ;
        RECT 3313.445 4981.765 3313.615 4981.955 ;
        RECT 3319.425 4981.765 3319.595 4981.955 ;
        RECT 3325.405 4981.765 3325.575 4981.955 ;
        RECT 3331.385 4981.765 3331.555 4981.955 ;
        RECT 834.665 4980.825 835.095 4981.610 ;
        RECT 835.495 4980.740 840.625 4981.650 ;
        RECT 840.645 4980.825 841.075 4981.610 ;
        RECT 841.475 4980.740 846.605 4981.650 ;
        RECT 846.625 4980.825 847.055 4981.610 ;
        RECT 847.455 4980.740 852.585 4981.650 ;
        RECT 852.605 4980.825 853.035 4981.610 ;
        RECT 840.310 4980.550 840.480 4980.740 ;
        RECT 846.290 4980.550 846.460 4980.740 ;
        RECT 852.270 4980.550 852.440 4980.740 ;
        RECT 198.835 4456.755 199.620 4457.185 ;
        RECT 198.750 4451.540 199.660 4456.355 ;
        RECT 198.560 4451.370 199.660 4451.540 ;
        RECT 198.750 4451.225 199.660 4451.370 ;
        RECT 198.835 4450.775 199.620 4451.205 ;
        RECT 198.750 4445.560 199.660 4450.375 ;
        RECT 198.560 4445.390 199.660 4445.560 ;
        RECT 198.750 4445.245 199.660 4445.390 ;
        RECT 198.835 4444.795 199.620 4445.225 ;
        RECT 198.750 4439.580 199.660 4444.395 ;
        RECT 198.560 4439.410 199.660 4439.580 ;
        RECT 198.750 4439.265 199.660 4439.410 ;
        RECT 198.835 4438.815 199.620 4439.245 ;
        RECT 198.750 4433.600 199.660 4438.415 ;
        RECT 198.560 4433.430 199.660 4433.600 ;
        RECT 198.750 4433.285 199.660 4433.430 ;
        RECT 198.835 4432.835 199.620 4433.265 ;
        RECT 198.750 4427.620 199.660 4432.435 ;
        RECT 198.560 4427.450 199.660 4427.620 ;
        RECT 198.750 4427.305 199.660 4427.450 ;
        RECT 198.835 4426.855 199.620 4427.285 ;
      LAYER nwell ;
        RECT 199.950 4426.650 202.780 4457.390 ;
      LAYER pwell ;
        RECT 203.110 4456.755 203.895 4457.185 ;
        RECT 203.070 4456.590 203.980 4456.735 ;
        RECT 203.070 4456.420 204.170 4456.590 ;
        RECT 203.070 4451.605 203.980 4456.420 ;
        RECT 203.110 4450.775 203.895 4451.205 ;
        RECT 203.070 4450.610 203.980 4450.755 ;
        RECT 203.070 4450.440 204.170 4450.610 ;
        RECT 203.070 4445.625 203.980 4450.440 ;
        RECT 203.110 4444.795 203.895 4445.225 ;
        RECT 203.070 4444.630 203.980 4444.775 ;
        RECT 203.070 4444.460 204.170 4444.630 ;
        RECT 203.070 4439.645 203.980 4444.460 ;
        RECT 203.110 4438.815 203.895 4439.245 ;
        RECT 203.070 4438.650 203.980 4438.795 ;
        RECT 203.070 4438.480 204.170 4438.650 ;
        RECT 203.070 4433.665 203.980 4438.480 ;
        RECT 203.110 4432.835 203.895 4433.265 ;
        RECT 203.070 4432.670 203.980 4432.815 ;
        RECT 203.070 4432.500 204.170 4432.670 ;
        RECT 203.070 4427.685 203.980 4432.500 ;
        RECT 203.110 4426.855 203.895 4427.285 ;
        RECT 3383.775 3571.955 3384.560 3572.385 ;
        RECT 3383.690 3571.790 3384.600 3571.935 ;
        RECT 3383.500 3571.620 3384.600 3571.790 ;
        RECT 3383.690 3566.805 3384.600 3571.620 ;
        RECT 3383.775 3565.975 3384.560 3566.405 ;
        RECT 3383.690 3565.810 3384.600 3565.955 ;
        RECT 3383.500 3565.640 3384.600 3565.810 ;
        RECT 3383.690 3560.825 3384.600 3565.640 ;
        RECT 3383.775 3559.995 3384.560 3560.425 ;
        RECT 3383.690 3559.830 3384.600 3559.975 ;
        RECT 3383.500 3559.660 3384.600 3559.830 ;
        RECT 3383.690 3554.845 3384.600 3559.660 ;
        RECT 3383.775 3554.015 3384.560 3554.445 ;
        RECT 3383.690 3553.850 3384.600 3553.995 ;
        RECT 3383.500 3553.680 3384.600 3553.850 ;
        RECT 3383.690 3548.865 3384.600 3553.680 ;
        RECT 3383.775 3548.035 3384.560 3548.465 ;
        RECT 3383.690 3547.870 3384.600 3548.015 ;
        RECT 3383.500 3547.700 3384.600 3547.870 ;
        RECT 3383.690 3542.885 3384.600 3547.700 ;
        RECT 3383.775 3542.055 3384.560 3542.485 ;
        RECT 3383.690 3541.890 3384.600 3542.035 ;
        RECT 3383.500 3541.720 3384.600 3541.890 ;
        RECT 3383.690 3536.905 3384.600 3541.720 ;
        RECT 3383.775 3536.075 3384.560 3536.505 ;
      LAYER nwell ;
        RECT 3384.890 3535.870 3387.720 3572.590 ;
      LAYER pwell ;
        RECT 3388.050 3571.955 3388.835 3572.385 ;
        RECT 3388.010 3566.740 3388.920 3571.555 ;
        RECT 3388.010 3566.570 3389.110 3566.740 ;
        RECT 3388.010 3566.425 3388.920 3566.570 ;
        RECT 3388.050 3565.975 3388.835 3566.405 ;
        RECT 3388.010 3560.760 3388.920 3565.575 ;
        RECT 3388.010 3560.590 3389.110 3560.760 ;
        RECT 3388.010 3560.445 3388.920 3560.590 ;
        RECT 3388.050 3559.995 3388.835 3560.425 ;
        RECT 3388.010 3554.780 3388.920 3559.595 ;
        RECT 3388.010 3554.610 3389.110 3554.780 ;
        RECT 3388.010 3554.465 3388.920 3554.610 ;
        RECT 3388.050 3554.015 3388.835 3554.445 ;
        RECT 3388.010 3548.800 3388.920 3553.615 ;
        RECT 3388.010 3548.630 3389.110 3548.800 ;
        RECT 3388.010 3548.485 3388.920 3548.630 ;
        RECT 3388.050 3548.035 3388.835 3548.465 ;
        RECT 3388.010 3542.820 3388.920 3547.635 ;
        RECT 3388.010 3542.650 3389.110 3542.820 ;
        RECT 3388.010 3542.505 3388.920 3542.650 ;
        RECT 3388.050 3542.055 3388.835 3542.485 ;
        RECT 3388.010 3536.840 3388.920 3541.655 ;
        RECT 3388.010 3536.670 3389.110 3536.840 ;
        RECT 3388.010 3536.525 3388.920 3536.670 ;
        RECT 3388.050 3536.075 3388.835 3536.505 ;
        RECT 198.960 3053.525 199.745 3053.955 ;
        RECT 198.875 3048.310 199.785 3053.125 ;
        RECT 198.685 3048.140 199.785 3048.310 ;
        RECT 198.875 3047.995 199.785 3048.140 ;
        RECT 198.960 3047.545 199.745 3047.975 ;
        RECT 198.875 3042.330 199.785 3047.145 ;
        RECT 198.685 3042.160 199.785 3042.330 ;
        RECT 198.875 3042.015 199.785 3042.160 ;
        RECT 198.960 3041.565 199.745 3041.995 ;
        RECT 198.875 3036.350 199.785 3041.165 ;
        RECT 198.685 3036.180 199.785 3036.350 ;
        RECT 198.875 3036.035 199.785 3036.180 ;
        RECT 198.960 3035.585 199.745 3036.015 ;
        RECT 198.875 3030.370 199.785 3035.185 ;
        RECT 198.685 3030.200 199.785 3030.370 ;
        RECT 198.875 3030.055 199.785 3030.200 ;
        RECT 198.960 3029.605 199.745 3030.035 ;
        RECT 198.875 3024.390 199.785 3029.205 ;
        RECT 198.685 3024.220 199.785 3024.390 ;
        RECT 198.875 3024.075 199.785 3024.220 ;
        RECT 198.960 3023.625 199.745 3024.055 ;
        RECT 198.875 3018.410 199.785 3023.225 ;
        RECT 198.685 3018.240 199.785 3018.410 ;
        RECT 198.875 3018.095 199.785 3018.240 ;
        RECT 198.960 3017.645 199.745 3018.075 ;
        RECT 198.875 3012.430 199.785 3017.245 ;
        RECT 198.685 3012.260 199.785 3012.430 ;
        RECT 198.875 3012.115 199.785 3012.260 ;
        RECT 198.960 3011.665 199.745 3012.095 ;
        RECT 198.875 3006.450 199.785 3011.265 ;
        RECT 198.685 3006.280 199.785 3006.450 ;
        RECT 198.875 3006.135 199.785 3006.280 ;
        RECT 198.960 3005.685 199.745 3006.115 ;
        RECT 198.875 3000.470 199.785 3005.285 ;
        RECT 198.685 3000.300 199.785 3000.470 ;
        RECT 198.875 3000.155 199.785 3000.300 ;
        RECT 198.960 2999.705 199.745 3000.135 ;
        RECT 198.875 2994.490 199.785 2999.305 ;
        RECT 198.685 2994.320 199.785 2994.490 ;
        RECT 198.875 2994.175 199.785 2994.320 ;
        RECT 198.960 2993.725 199.745 2994.155 ;
        RECT 198.875 2988.510 199.785 2993.325 ;
        RECT 198.685 2988.340 199.785 2988.510 ;
        RECT 198.875 2988.195 199.785 2988.340 ;
        RECT 198.960 2987.745 199.745 2988.175 ;
      LAYER nwell ;
        RECT 200.075 2987.540 202.905 3054.160 ;
      LAYER pwell ;
        RECT 203.235 3053.525 204.020 3053.955 ;
        RECT 203.195 3053.360 204.105 3053.505 ;
        RECT 203.195 3053.190 204.295 3053.360 ;
        RECT 203.195 3048.375 204.105 3053.190 ;
        RECT 203.235 3047.545 204.020 3047.975 ;
        RECT 203.195 3047.380 204.105 3047.525 ;
        RECT 203.195 3047.210 204.295 3047.380 ;
        RECT 203.195 3042.395 204.105 3047.210 ;
        RECT 203.235 3041.565 204.020 3041.995 ;
        RECT 203.195 3041.400 204.105 3041.545 ;
        RECT 203.195 3041.230 204.295 3041.400 ;
        RECT 203.195 3036.415 204.105 3041.230 ;
        RECT 203.235 3035.585 204.020 3036.015 ;
        RECT 203.195 3035.420 204.105 3035.565 ;
        RECT 203.195 3035.250 204.295 3035.420 ;
        RECT 203.195 3030.435 204.105 3035.250 ;
        RECT 203.235 3029.605 204.020 3030.035 ;
        RECT 203.195 3029.440 204.105 3029.585 ;
        RECT 203.195 3029.270 204.295 3029.440 ;
        RECT 203.195 3024.455 204.105 3029.270 ;
        RECT 203.235 3023.625 204.020 3024.055 ;
        RECT 203.195 3023.460 204.105 3023.605 ;
        RECT 203.195 3023.290 204.295 3023.460 ;
        RECT 203.195 3018.475 204.105 3023.290 ;
        RECT 203.235 3017.645 204.020 3018.075 ;
        RECT 203.195 3017.480 204.105 3017.625 ;
        RECT 203.195 3017.310 204.295 3017.480 ;
        RECT 203.195 3012.495 204.105 3017.310 ;
        RECT 203.235 3011.665 204.020 3012.095 ;
        RECT 203.195 3011.500 204.105 3011.645 ;
        RECT 203.195 3011.330 204.295 3011.500 ;
        RECT 203.195 3006.515 204.105 3011.330 ;
        RECT 203.235 3005.685 204.020 3006.115 ;
        RECT 203.195 3005.520 204.105 3005.665 ;
        RECT 203.195 3005.350 204.295 3005.520 ;
        RECT 203.195 3000.535 204.105 3005.350 ;
        RECT 203.235 2999.705 204.020 3000.135 ;
        RECT 203.195 2999.540 204.105 2999.685 ;
        RECT 203.195 2999.370 204.295 2999.540 ;
        RECT 203.195 2994.555 204.105 2999.370 ;
        RECT 203.235 2993.725 204.020 2994.155 ;
        RECT 203.195 2993.560 204.105 2993.705 ;
        RECT 203.195 2993.390 204.295 2993.560 ;
        RECT 203.195 2988.575 204.105 2993.390 ;
        RECT 203.235 2987.745 204.020 2988.175 ;
        RECT 3383.775 2267.835 3384.560 2268.265 ;
        RECT 3383.690 2267.670 3384.600 2267.815 ;
        RECT 3383.500 2267.500 3384.600 2267.670 ;
        RECT 3383.690 2262.685 3384.600 2267.500 ;
        RECT 3383.775 2261.855 3384.560 2262.285 ;
        RECT 3383.690 2261.690 3384.600 2261.835 ;
        RECT 3383.500 2261.520 3384.600 2261.690 ;
        RECT 3383.690 2256.705 3384.600 2261.520 ;
        RECT 3383.775 2255.875 3384.560 2256.305 ;
        RECT 3383.690 2255.710 3384.600 2255.855 ;
        RECT 3383.500 2255.540 3384.600 2255.710 ;
        RECT 3383.690 2250.725 3384.600 2255.540 ;
        RECT 3383.775 2249.895 3384.560 2250.325 ;
        RECT 3383.690 2249.730 3384.600 2249.875 ;
        RECT 3383.500 2249.560 3384.600 2249.730 ;
        RECT 3383.690 2244.745 3384.600 2249.560 ;
        RECT 3383.775 2243.915 3384.560 2244.345 ;
        RECT 3383.690 2243.750 3384.600 2243.895 ;
        RECT 3383.500 2243.580 3384.600 2243.750 ;
        RECT 3383.690 2238.765 3384.600 2243.580 ;
        RECT 3383.775 2237.935 3384.560 2238.365 ;
        RECT 3383.690 2237.770 3384.600 2237.915 ;
        RECT 3383.500 2237.600 3384.600 2237.770 ;
        RECT 3383.690 2232.785 3384.600 2237.600 ;
        RECT 3383.775 2231.955 3384.560 2232.385 ;
        RECT 3383.690 2231.790 3384.600 2231.935 ;
        RECT 3383.500 2231.620 3384.600 2231.790 ;
        RECT 3383.690 2226.805 3384.600 2231.620 ;
        RECT 3383.775 2225.975 3384.560 2226.405 ;
        RECT 3383.690 2225.810 3384.600 2225.955 ;
        RECT 3383.500 2225.640 3384.600 2225.810 ;
        RECT 3383.690 2220.825 3384.600 2225.640 ;
        RECT 3383.775 2219.995 3384.560 2220.425 ;
        RECT 3383.690 2219.830 3384.600 2219.975 ;
        RECT 3383.500 2219.660 3384.600 2219.830 ;
        RECT 3383.690 2214.845 3384.600 2219.660 ;
        RECT 3383.775 2214.015 3384.560 2214.445 ;
        RECT 3383.690 2213.850 3384.600 2213.995 ;
        RECT 3383.500 2213.680 3384.600 2213.850 ;
        RECT 3383.690 2208.865 3384.600 2213.680 ;
        RECT 3383.775 2208.035 3384.560 2208.465 ;
        RECT 3383.690 2207.870 3384.600 2208.015 ;
        RECT 3383.500 2207.700 3384.600 2207.870 ;
        RECT 3383.690 2202.885 3384.600 2207.700 ;
        RECT 3383.775 2202.055 3384.560 2202.485 ;
        RECT 3383.690 2201.890 3384.600 2202.035 ;
        RECT 3383.500 2201.720 3384.600 2201.890 ;
        RECT 3383.690 2196.905 3384.600 2201.720 ;
        RECT 3383.775 2196.075 3384.560 2196.505 ;
      LAYER nwell ;
        RECT 3384.890 2195.870 3387.720 2268.470 ;
      LAYER pwell ;
        RECT 3388.050 2267.835 3388.835 2268.265 ;
        RECT 3388.010 2262.620 3388.920 2267.435 ;
        RECT 3388.010 2262.450 3389.110 2262.620 ;
        RECT 3388.010 2262.305 3388.920 2262.450 ;
        RECT 3388.050 2261.855 3388.835 2262.285 ;
        RECT 3388.010 2256.640 3388.920 2261.455 ;
        RECT 3388.010 2256.470 3389.110 2256.640 ;
        RECT 3388.010 2256.325 3388.920 2256.470 ;
        RECT 3388.050 2255.875 3388.835 2256.305 ;
        RECT 3388.010 2250.660 3388.920 2255.475 ;
        RECT 3388.010 2250.490 3389.110 2250.660 ;
        RECT 3388.010 2250.345 3388.920 2250.490 ;
        RECT 3388.050 2249.895 3388.835 2250.325 ;
        RECT 3388.010 2244.680 3388.920 2249.495 ;
        RECT 3388.010 2244.510 3389.110 2244.680 ;
        RECT 3388.010 2244.365 3388.920 2244.510 ;
        RECT 3388.050 2243.915 3388.835 2244.345 ;
        RECT 3388.010 2238.700 3388.920 2243.515 ;
        RECT 3388.010 2238.530 3389.110 2238.700 ;
        RECT 3388.010 2238.385 3388.920 2238.530 ;
        RECT 3388.050 2237.935 3388.835 2238.365 ;
        RECT 3388.010 2232.720 3388.920 2237.535 ;
        RECT 3388.010 2232.550 3389.110 2232.720 ;
        RECT 3388.010 2232.405 3388.920 2232.550 ;
        RECT 3388.050 2231.955 3388.835 2232.385 ;
        RECT 3388.010 2226.740 3388.920 2231.555 ;
        RECT 3388.010 2226.570 3389.110 2226.740 ;
        RECT 3388.010 2226.425 3388.920 2226.570 ;
        RECT 3388.050 2225.975 3388.835 2226.405 ;
        RECT 3388.010 2220.760 3388.920 2225.575 ;
        RECT 3388.010 2220.590 3389.110 2220.760 ;
        RECT 3388.010 2220.445 3388.920 2220.590 ;
        RECT 3388.050 2219.995 3388.835 2220.425 ;
        RECT 3388.010 2214.780 3388.920 2219.595 ;
        RECT 3388.010 2214.610 3389.110 2214.780 ;
        RECT 3388.010 2214.465 3388.920 2214.610 ;
        RECT 3388.050 2214.015 3388.835 2214.445 ;
        RECT 3388.010 2208.800 3388.920 2213.615 ;
        RECT 3388.010 2208.630 3389.110 2208.800 ;
        RECT 3388.010 2208.485 3388.920 2208.630 ;
        RECT 3388.050 2208.035 3388.835 2208.465 ;
        RECT 3388.010 2202.820 3388.920 2207.635 ;
        RECT 3388.010 2202.650 3389.110 2202.820 ;
        RECT 3388.010 2202.505 3388.920 2202.650 ;
        RECT 3388.050 2202.055 3388.835 2202.485 ;
        RECT 3388.010 2196.840 3388.920 2201.655 ;
        RECT 3388.010 2196.670 3389.110 2196.840 ;
        RECT 3388.010 2196.525 3388.920 2196.670 ;
        RECT 3388.050 2196.075 3388.835 2196.505 ;
        RECT 199.070 1762.620 199.855 1763.050 ;
        RECT 198.985 1757.405 199.895 1762.220 ;
        RECT 198.795 1757.235 199.895 1757.405 ;
        RECT 198.985 1757.090 199.895 1757.235 ;
        RECT 199.070 1756.640 199.855 1757.070 ;
        RECT 198.985 1751.425 199.895 1756.240 ;
        RECT 198.795 1751.255 199.895 1751.425 ;
        RECT 198.985 1751.110 199.895 1751.255 ;
        RECT 199.070 1750.660 199.855 1751.090 ;
        RECT 198.985 1745.445 199.895 1750.260 ;
        RECT 198.795 1745.275 199.895 1745.445 ;
        RECT 198.985 1745.130 199.895 1745.275 ;
        RECT 199.070 1744.680 199.855 1745.110 ;
        RECT 198.985 1739.465 199.895 1744.280 ;
        RECT 198.795 1739.295 199.895 1739.465 ;
        RECT 198.985 1739.150 199.895 1739.295 ;
        RECT 199.070 1738.700 199.855 1739.130 ;
        RECT 198.985 1733.485 199.895 1738.300 ;
        RECT 198.795 1733.315 199.895 1733.485 ;
        RECT 198.985 1733.170 199.895 1733.315 ;
        RECT 199.070 1732.720 199.855 1733.150 ;
        RECT 198.985 1727.505 199.895 1732.320 ;
        RECT 198.795 1727.335 199.895 1727.505 ;
        RECT 198.985 1727.190 199.895 1727.335 ;
        RECT 199.070 1726.740 199.855 1727.170 ;
        RECT 198.985 1721.525 199.895 1726.340 ;
        RECT 198.795 1721.355 199.895 1721.525 ;
        RECT 198.985 1721.210 199.895 1721.355 ;
        RECT 199.070 1720.760 199.855 1721.190 ;
        RECT 198.985 1715.545 199.895 1720.360 ;
        RECT 198.795 1715.375 199.895 1715.545 ;
        RECT 198.985 1715.230 199.895 1715.375 ;
        RECT 199.070 1714.780 199.855 1715.210 ;
        RECT 198.985 1709.565 199.895 1714.380 ;
        RECT 198.795 1709.395 199.895 1709.565 ;
        RECT 198.985 1709.250 199.895 1709.395 ;
        RECT 199.070 1708.800 199.855 1709.230 ;
        RECT 198.985 1703.585 199.895 1708.400 ;
        RECT 198.795 1703.415 199.895 1703.585 ;
        RECT 198.985 1703.270 199.895 1703.415 ;
        RECT 199.070 1702.820 199.855 1703.250 ;
        RECT 198.985 1697.605 199.895 1702.420 ;
        RECT 198.795 1697.435 199.895 1697.605 ;
        RECT 198.985 1697.290 199.895 1697.435 ;
        RECT 199.070 1696.840 199.855 1697.270 ;
        RECT 198.985 1691.625 199.895 1696.440 ;
        RECT 198.795 1691.455 199.895 1691.625 ;
        RECT 198.985 1691.310 199.895 1691.455 ;
        RECT 199.070 1690.860 199.855 1691.290 ;
        RECT 198.985 1685.645 199.895 1690.460 ;
        RECT 198.795 1685.475 199.895 1685.645 ;
        RECT 198.985 1685.330 199.895 1685.475 ;
        RECT 199.070 1684.880 199.855 1685.310 ;
        RECT 198.985 1679.665 199.895 1684.480 ;
        RECT 198.795 1679.495 199.895 1679.665 ;
        RECT 198.985 1679.350 199.895 1679.495 ;
        RECT 199.070 1678.900 199.855 1679.330 ;
        RECT 198.985 1673.685 199.895 1678.500 ;
        RECT 198.795 1673.515 199.895 1673.685 ;
        RECT 198.985 1673.370 199.895 1673.515 ;
        RECT 199.070 1672.920 199.855 1673.350 ;
      LAYER nwell ;
        RECT 200.185 1672.715 203.015 1763.255 ;
      LAYER pwell ;
        RECT 203.345 1762.620 204.130 1763.050 ;
        RECT 203.305 1762.455 204.215 1762.600 ;
        RECT 203.305 1762.285 204.405 1762.455 ;
        RECT 203.305 1757.470 204.215 1762.285 ;
        RECT 203.345 1756.640 204.130 1757.070 ;
        RECT 203.305 1756.475 204.215 1756.620 ;
        RECT 203.305 1756.305 204.405 1756.475 ;
        RECT 203.305 1751.490 204.215 1756.305 ;
        RECT 203.345 1750.660 204.130 1751.090 ;
        RECT 203.305 1750.495 204.215 1750.640 ;
        RECT 203.305 1750.325 204.405 1750.495 ;
        RECT 203.305 1745.510 204.215 1750.325 ;
        RECT 203.345 1744.680 204.130 1745.110 ;
        RECT 203.305 1744.515 204.215 1744.660 ;
        RECT 203.305 1744.345 204.405 1744.515 ;
        RECT 203.305 1739.530 204.215 1744.345 ;
        RECT 203.345 1738.700 204.130 1739.130 ;
        RECT 203.305 1738.535 204.215 1738.680 ;
        RECT 203.305 1738.365 204.405 1738.535 ;
        RECT 203.305 1733.550 204.215 1738.365 ;
        RECT 203.345 1732.720 204.130 1733.150 ;
        RECT 203.305 1732.555 204.215 1732.700 ;
        RECT 203.305 1732.385 204.405 1732.555 ;
        RECT 203.305 1727.570 204.215 1732.385 ;
        RECT 203.345 1726.740 204.130 1727.170 ;
        RECT 203.305 1726.575 204.215 1726.720 ;
        RECT 203.305 1726.405 204.405 1726.575 ;
        RECT 203.305 1721.590 204.215 1726.405 ;
        RECT 203.345 1720.760 204.130 1721.190 ;
        RECT 203.305 1720.595 204.215 1720.740 ;
        RECT 203.305 1720.425 204.405 1720.595 ;
        RECT 203.305 1715.610 204.215 1720.425 ;
        RECT 203.345 1714.780 204.130 1715.210 ;
        RECT 203.305 1714.615 204.215 1714.760 ;
        RECT 203.305 1714.445 204.405 1714.615 ;
        RECT 203.305 1709.630 204.215 1714.445 ;
        RECT 203.345 1708.800 204.130 1709.230 ;
        RECT 203.305 1708.635 204.215 1708.780 ;
        RECT 203.305 1708.465 204.405 1708.635 ;
        RECT 203.305 1703.650 204.215 1708.465 ;
        RECT 203.345 1702.820 204.130 1703.250 ;
        RECT 203.305 1702.655 204.215 1702.800 ;
        RECT 203.305 1702.485 204.405 1702.655 ;
        RECT 203.305 1697.670 204.215 1702.485 ;
        RECT 203.345 1696.840 204.130 1697.270 ;
        RECT 203.305 1696.675 204.215 1696.820 ;
        RECT 203.305 1696.505 204.405 1696.675 ;
        RECT 203.305 1691.690 204.215 1696.505 ;
        RECT 203.345 1690.860 204.130 1691.290 ;
        RECT 203.305 1690.695 204.215 1690.840 ;
        RECT 203.305 1690.525 204.405 1690.695 ;
        RECT 203.305 1685.710 204.215 1690.525 ;
        RECT 203.345 1684.880 204.130 1685.310 ;
        RECT 203.305 1684.715 204.215 1684.860 ;
        RECT 203.305 1684.545 204.405 1684.715 ;
        RECT 203.305 1679.730 204.215 1684.545 ;
        RECT 203.345 1678.900 204.130 1679.330 ;
        RECT 203.305 1678.735 204.215 1678.880 ;
        RECT 203.305 1678.565 204.405 1678.735 ;
        RECT 203.305 1673.750 204.215 1678.565 ;
        RECT 203.345 1672.920 204.130 1673.350 ;
        RECT 674.660 1117.020 674.830 1117.210 ;
        RECT 680.640 1117.020 680.810 1117.210 ;
        RECT 686.620 1117.020 686.790 1117.210 ;
        RECT 692.600 1117.020 692.770 1117.210 ;
        RECT 698.580 1117.020 698.750 1117.210 ;
        RECT 704.560 1117.020 704.730 1117.210 ;
        RECT 710.540 1117.020 710.710 1117.210 ;
        RECT 716.520 1117.020 716.690 1117.210 ;
        RECT 722.500 1117.020 722.670 1117.210 ;
        RECT 728.480 1117.020 728.650 1117.210 ;
        RECT 734.460 1117.020 734.630 1117.210 ;
        RECT 740.440 1117.020 740.610 1117.210 ;
        RECT 746.420 1117.020 746.590 1117.210 ;
        RECT 752.400 1117.020 752.570 1117.210 ;
        RECT 758.380 1117.020 758.550 1117.210 ;
        RECT 764.360 1117.020 764.530 1117.210 ;
        RECT 770.340 1117.020 770.510 1117.210 ;
        RECT 776.320 1117.020 776.490 1117.210 ;
        RECT 782.300 1117.020 782.470 1117.210 ;
        RECT 788.280 1117.020 788.450 1117.210 ;
        RECT 794.260 1117.020 794.430 1117.210 ;
        RECT 1974.660 1117.020 1974.830 1117.210 ;
        RECT 1980.640 1117.020 1980.810 1117.210 ;
        RECT 1986.620 1117.020 1986.790 1117.210 ;
        RECT 1992.600 1117.020 1992.770 1117.210 ;
        RECT 1998.580 1117.020 1998.750 1117.210 ;
        RECT 2004.560 1117.020 2004.730 1117.210 ;
        RECT 2010.540 1117.020 2010.710 1117.210 ;
        RECT 2016.520 1117.020 2016.690 1117.210 ;
        RECT 2022.500 1117.020 2022.670 1117.210 ;
        RECT 2028.480 1117.020 2028.650 1117.210 ;
        RECT 2034.460 1117.020 2034.630 1117.210 ;
        RECT 2040.440 1117.020 2040.610 1117.210 ;
        RECT 2046.420 1117.020 2046.590 1117.210 ;
        RECT 2052.400 1117.020 2052.570 1117.210 ;
        RECT 2058.380 1117.020 2058.550 1117.210 ;
        RECT 2064.360 1117.020 2064.530 1117.210 ;
        RECT 2070.340 1117.020 2070.510 1117.210 ;
        RECT 2076.320 1117.020 2076.490 1117.210 ;
        RECT 2082.300 1117.020 2082.470 1117.210 ;
        RECT 2088.280 1117.020 2088.450 1117.210 ;
        RECT 2094.260 1117.020 2094.430 1117.210 ;
        RECT 669.015 1116.150 669.445 1116.935 ;
        RECT 669.845 1116.110 674.975 1117.020 ;
        RECT 674.995 1116.150 675.425 1116.935 ;
        RECT 675.825 1116.110 680.955 1117.020 ;
        RECT 680.975 1116.150 681.405 1116.935 ;
        RECT 681.805 1116.110 686.935 1117.020 ;
        RECT 686.955 1116.150 687.385 1116.935 ;
        RECT 687.785 1116.110 692.915 1117.020 ;
        RECT 692.935 1116.150 693.365 1116.935 ;
        RECT 693.765 1116.110 698.895 1117.020 ;
        RECT 698.915 1116.150 699.345 1116.935 ;
        RECT 699.745 1116.110 704.875 1117.020 ;
        RECT 704.895 1116.150 705.325 1116.935 ;
        RECT 705.725 1116.110 710.855 1117.020 ;
        RECT 710.875 1116.150 711.305 1116.935 ;
        RECT 711.705 1116.110 716.835 1117.020 ;
        RECT 716.855 1116.150 717.285 1116.935 ;
        RECT 717.685 1116.110 722.815 1117.020 ;
        RECT 722.835 1116.150 723.265 1116.935 ;
        RECT 723.665 1116.110 728.795 1117.020 ;
        RECT 728.815 1116.150 729.245 1116.935 ;
        RECT 729.645 1116.110 734.775 1117.020 ;
        RECT 734.795 1116.150 735.225 1116.935 ;
        RECT 735.625 1116.110 740.755 1117.020 ;
        RECT 740.775 1116.150 741.205 1116.935 ;
        RECT 741.605 1116.110 746.735 1117.020 ;
        RECT 746.755 1116.150 747.185 1116.935 ;
        RECT 747.585 1116.110 752.715 1117.020 ;
        RECT 752.735 1116.150 753.165 1116.935 ;
        RECT 753.565 1116.110 758.695 1117.020 ;
        RECT 758.715 1116.150 759.145 1116.935 ;
        RECT 759.545 1116.110 764.675 1117.020 ;
        RECT 764.695 1116.150 765.125 1116.935 ;
        RECT 765.525 1116.110 770.655 1117.020 ;
        RECT 770.675 1116.150 771.105 1116.935 ;
        RECT 771.505 1116.110 776.635 1117.020 ;
        RECT 776.655 1116.150 777.085 1116.935 ;
        RECT 777.485 1116.110 782.615 1117.020 ;
        RECT 782.635 1116.150 783.065 1116.935 ;
        RECT 783.465 1116.110 788.595 1117.020 ;
        RECT 788.615 1116.150 789.045 1116.935 ;
        RECT 789.445 1116.110 794.575 1117.020 ;
        RECT 794.595 1116.150 795.025 1116.935 ;
        RECT 1969.015 1116.150 1969.445 1116.935 ;
        RECT 1969.845 1116.110 1974.975 1117.020 ;
        RECT 1974.995 1116.150 1975.425 1116.935 ;
        RECT 1975.825 1116.110 1980.955 1117.020 ;
        RECT 1980.975 1116.150 1981.405 1116.935 ;
        RECT 1981.805 1116.110 1986.935 1117.020 ;
        RECT 1986.955 1116.150 1987.385 1116.935 ;
        RECT 1987.785 1116.110 1992.915 1117.020 ;
        RECT 1992.935 1116.150 1993.365 1116.935 ;
        RECT 1993.765 1116.110 1998.895 1117.020 ;
        RECT 1998.915 1116.150 1999.345 1116.935 ;
        RECT 1999.745 1116.110 2004.875 1117.020 ;
        RECT 2004.895 1116.150 2005.325 1116.935 ;
        RECT 2005.725 1116.110 2010.855 1117.020 ;
        RECT 2010.875 1116.150 2011.305 1116.935 ;
        RECT 2011.705 1116.110 2016.835 1117.020 ;
        RECT 2016.855 1116.150 2017.285 1116.935 ;
        RECT 2017.685 1116.110 2022.815 1117.020 ;
        RECT 2022.835 1116.150 2023.265 1116.935 ;
        RECT 2023.665 1116.110 2028.795 1117.020 ;
        RECT 2028.815 1116.150 2029.245 1116.935 ;
        RECT 2029.645 1116.110 2034.775 1117.020 ;
        RECT 2034.795 1116.150 2035.225 1116.935 ;
        RECT 2035.625 1116.110 2040.755 1117.020 ;
        RECT 2040.775 1116.150 2041.205 1116.935 ;
        RECT 2041.605 1116.110 2046.735 1117.020 ;
        RECT 2046.755 1116.150 2047.185 1116.935 ;
        RECT 2047.585 1116.110 2052.715 1117.020 ;
        RECT 2052.735 1116.150 2053.165 1116.935 ;
        RECT 2053.565 1116.110 2058.695 1117.020 ;
        RECT 2058.715 1116.150 2059.145 1116.935 ;
        RECT 2059.545 1116.110 2064.675 1117.020 ;
        RECT 2064.695 1116.150 2065.125 1116.935 ;
        RECT 2065.525 1116.110 2070.655 1117.020 ;
        RECT 2070.675 1116.150 2071.105 1116.935 ;
        RECT 2071.505 1116.110 2076.635 1117.020 ;
        RECT 2076.655 1116.150 2077.085 1116.935 ;
        RECT 2077.485 1116.110 2082.615 1117.020 ;
        RECT 2082.635 1116.150 2083.065 1116.935 ;
        RECT 2083.465 1116.110 2088.595 1117.020 ;
        RECT 2088.615 1116.150 2089.045 1116.935 ;
        RECT 2089.445 1116.110 2094.575 1117.020 ;
        RECT 2094.595 1116.150 2095.025 1116.935 ;
      LAYER nwell ;
        RECT 668.810 1114.215 795.230 1115.820 ;
        RECT 1968.810 1114.215 2095.230 1115.820 ;
        RECT 674.790 1112.990 795.230 1114.215 ;
        RECT 1974.790 1112.990 2095.230 1114.215 ;
      LAYER pwell ;
        RECT 674.995 1111.875 675.425 1112.660 ;
        RECT 675.445 1111.790 680.575 1112.700 ;
        RECT 680.975 1111.875 681.405 1112.660 ;
        RECT 681.425 1111.790 686.555 1112.700 ;
        RECT 686.955 1111.875 687.385 1112.660 ;
        RECT 687.405 1111.790 692.535 1112.700 ;
        RECT 692.935 1111.875 693.365 1112.660 ;
        RECT 693.385 1111.790 698.515 1112.700 ;
        RECT 698.915 1111.875 699.345 1112.660 ;
        RECT 699.365 1111.790 704.495 1112.700 ;
        RECT 704.895 1111.875 705.325 1112.660 ;
        RECT 705.345 1111.790 710.475 1112.700 ;
        RECT 710.875 1111.875 711.305 1112.660 ;
        RECT 711.325 1111.790 716.455 1112.700 ;
        RECT 716.855 1111.875 717.285 1112.660 ;
        RECT 717.305 1111.790 722.435 1112.700 ;
        RECT 722.835 1111.875 723.265 1112.660 ;
        RECT 723.285 1111.790 728.415 1112.700 ;
        RECT 728.815 1111.875 729.245 1112.660 ;
        RECT 729.265 1111.790 734.395 1112.700 ;
        RECT 734.795 1111.875 735.225 1112.660 ;
        RECT 735.245 1111.790 740.375 1112.700 ;
        RECT 740.775 1111.875 741.205 1112.660 ;
        RECT 741.225 1111.790 746.355 1112.700 ;
        RECT 746.755 1111.875 747.185 1112.660 ;
        RECT 747.205 1111.790 752.335 1112.700 ;
        RECT 752.735 1111.875 753.165 1112.660 ;
        RECT 753.185 1111.790 758.315 1112.700 ;
        RECT 758.715 1111.875 759.145 1112.660 ;
        RECT 759.165 1111.790 764.295 1112.700 ;
        RECT 764.695 1111.875 765.125 1112.660 ;
        RECT 765.145 1111.790 770.275 1112.700 ;
        RECT 770.675 1111.875 771.105 1112.660 ;
        RECT 771.125 1111.790 776.255 1112.700 ;
        RECT 776.655 1111.875 777.085 1112.660 ;
        RECT 777.105 1111.790 782.235 1112.700 ;
        RECT 782.635 1111.875 783.065 1112.660 ;
        RECT 783.085 1111.790 788.215 1112.700 ;
        RECT 788.615 1111.875 789.045 1112.660 ;
        RECT 789.445 1111.790 794.575 1112.700 ;
        RECT 794.595 1111.875 795.025 1112.660 ;
        RECT 1974.995 1111.875 1975.425 1112.660 ;
        RECT 1975.445 1111.790 1980.575 1112.700 ;
        RECT 1980.975 1111.875 1981.405 1112.660 ;
        RECT 1981.425 1111.790 1986.555 1112.700 ;
        RECT 1986.955 1111.875 1987.385 1112.660 ;
        RECT 1987.405 1111.790 1992.535 1112.700 ;
        RECT 1992.935 1111.875 1993.365 1112.660 ;
        RECT 1993.385 1111.790 1998.515 1112.700 ;
        RECT 1998.915 1111.875 1999.345 1112.660 ;
        RECT 1999.365 1111.790 2004.495 1112.700 ;
        RECT 2004.895 1111.875 2005.325 1112.660 ;
        RECT 2005.345 1111.790 2010.475 1112.700 ;
        RECT 2010.875 1111.875 2011.305 1112.660 ;
        RECT 2011.325 1111.790 2016.455 1112.700 ;
        RECT 2016.855 1111.875 2017.285 1112.660 ;
        RECT 2017.305 1111.790 2022.435 1112.700 ;
        RECT 2022.835 1111.875 2023.265 1112.660 ;
        RECT 2023.285 1111.790 2028.415 1112.700 ;
        RECT 2028.815 1111.875 2029.245 1112.660 ;
        RECT 2029.265 1111.790 2034.395 1112.700 ;
        RECT 2034.795 1111.875 2035.225 1112.660 ;
        RECT 2035.245 1111.790 2040.375 1112.700 ;
        RECT 2040.775 1111.875 2041.205 1112.660 ;
        RECT 2041.225 1111.790 2046.355 1112.700 ;
        RECT 2046.755 1111.875 2047.185 1112.660 ;
        RECT 2047.205 1111.790 2052.335 1112.700 ;
        RECT 2052.735 1111.875 2053.165 1112.660 ;
        RECT 2053.185 1111.790 2058.315 1112.700 ;
        RECT 2058.715 1111.875 2059.145 1112.660 ;
        RECT 2059.165 1111.790 2064.295 1112.700 ;
        RECT 2064.695 1111.875 2065.125 1112.660 ;
        RECT 2065.145 1111.790 2070.275 1112.700 ;
        RECT 2070.675 1111.875 2071.105 1112.660 ;
        RECT 2071.125 1111.790 2076.255 1112.700 ;
        RECT 2076.655 1111.875 2077.085 1112.660 ;
        RECT 2077.105 1111.790 2082.235 1112.700 ;
        RECT 2082.635 1111.875 2083.065 1112.660 ;
        RECT 2083.085 1111.790 2088.215 1112.700 ;
        RECT 2088.615 1111.875 2089.045 1112.660 ;
        RECT 2089.445 1111.790 2094.575 1112.700 ;
        RECT 2094.595 1111.875 2095.025 1112.660 ;
        RECT 675.590 1111.600 675.760 1111.790 ;
        RECT 681.570 1111.600 681.740 1111.790 ;
        RECT 687.550 1111.600 687.720 1111.790 ;
        RECT 693.530 1111.600 693.700 1111.790 ;
        RECT 699.510 1111.600 699.680 1111.790 ;
        RECT 705.490 1111.600 705.660 1111.790 ;
        RECT 711.470 1111.600 711.640 1111.790 ;
        RECT 717.450 1111.600 717.620 1111.790 ;
        RECT 723.430 1111.600 723.600 1111.790 ;
        RECT 729.410 1111.600 729.580 1111.790 ;
        RECT 735.390 1111.600 735.560 1111.790 ;
        RECT 741.370 1111.600 741.540 1111.790 ;
        RECT 747.350 1111.600 747.520 1111.790 ;
        RECT 753.330 1111.600 753.500 1111.790 ;
        RECT 759.310 1111.600 759.480 1111.790 ;
        RECT 765.290 1111.600 765.460 1111.790 ;
        RECT 771.270 1111.600 771.440 1111.790 ;
        RECT 777.250 1111.600 777.420 1111.790 ;
        RECT 783.230 1111.600 783.400 1111.790 ;
        RECT 794.260 1111.600 794.430 1111.790 ;
        RECT 1975.590 1111.600 1975.760 1111.790 ;
        RECT 1981.570 1111.600 1981.740 1111.790 ;
        RECT 1987.550 1111.600 1987.720 1111.790 ;
        RECT 1993.530 1111.600 1993.700 1111.790 ;
        RECT 1999.510 1111.600 1999.680 1111.790 ;
        RECT 2005.490 1111.600 2005.660 1111.790 ;
        RECT 2011.470 1111.600 2011.640 1111.790 ;
        RECT 2017.450 1111.600 2017.620 1111.790 ;
        RECT 2023.430 1111.600 2023.600 1111.790 ;
        RECT 2029.410 1111.600 2029.580 1111.790 ;
        RECT 2035.390 1111.600 2035.560 1111.790 ;
        RECT 2041.370 1111.600 2041.540 1111.790 ;
        RECT 2047.350 1111.600 2047.520 1111.790 ;
        RECT 2053.330 1111.600 2053.500 1111.790 ;
        RECT 2059.310 1111.600 2059.480 1111.790 ;
        RECT 2065.290 1111.600 2065.460 1111.790 ;
        RECT 2071.270 1111.600 2071.440 1111.790 ;
        RECT 2077.250 1111.600 2077.420 1111.790 ;
        RECT 2083.230 1111.600 2083.400 1111.790 ;
        RECT 2094.260 1111.600 2094.430 1111.790 ;
      LAYER li1 ;
        RECT 2082.830 4987.615 2082.975 4987.785 ;
        RECT 2083.145 4987.615 2083.435 4987.785 ;
        RECT 2083.605 4987.615 2083.895 4987.785 ;
        RECT 2084.065 4987.615 2084.355 4987.785 ;
        RECT 2084.525 4987.615 2084.815 4987.785 ;
        RECT 2084.985 4987.615 2085.275 4987.785 ;
        RECT 2085.445 4987.615 2085.735 4987.785 ;
        RECT 2085.905 4987.615 2086.195 4987.785 ;
        RECT 2086.365 4987.615 2086.655 4987.785 ;
        RECT 2086.825 4987.615 2087.115 4987.785 ;
        RECT 2087.285 4987.615 2087.575 4987.785 ;
        RECT 2087.745 4987.615 2088.035 4987.785 ;
        RECT 2088.205 4987.615 2088.495 4987.785 ;
        RECT 2088.665 4987.615 2088.955 4987.785 ;
        RECT 2089.125 4987.615 2089.270 4987.785 ;
        RECT 2082.915 4986.890 2083.205 4987.615 ;
        RECT 2083.765 4986.815 2084.095 4987.615 ;
        RECT 2084.605 4987.135 2084.935 4987.615 ;
        RECT 2085.445 4987.135 2085.775 4987.615 ;
        RECT 2086.285 4987.135 2086.615 4987.615 ;
        RECT 2087.125 4987.135 2087.455 4987.615 ;
        RECT 2087.625 4986.965 2087.795 4987.440 ;
        RECT 2087.965 4987.135 2088.295 4987.615 ;
        RECT 2088.465 4986.965 2088.635 4987.445 ;
        RECT 2087.215 4986.795 2088.635 4986.965 ;
        RECT 2088.895 4986.890 2089.185 4987.615 ;
        RECT 3312.835 4987.205 3312.980 4987.375 ;
        RECT 3313.150 4987.205 3313.440 4987.375 ;
        RECT 3313.610 4987.205 3313.900 4987.375 ;
        RECT 3314.070 4987.205 3314.360 4987.375 ;
        RECT 3314.530 4987.205 3314.820 4987.375 ;
        RECT 3314.990 4987.205 3315.280 4987.375 ;
        RECT 3315.450 4987.205 3315.740 4987.375 ;
        RECT 3315.910 4987.205 3316.200 4987.375 ;
        RECT 3316.370 4987.205 3316.660 4987.375 ;
        RECT 3316.830 4987.205 3317.120 4987.375 ;
        RECT 3317.290 4987.205 3317.580 4987.375 ;
        RECT 3317.750 4987.205 3318.040 4987.375 ;
        RECT 3318.210 4987.205 3318.500 4987.375 ;
        RECT 3318.670 4987.205 3318.960 4987.375 ;
        RECT 3319.130 4987.205 3319.420 4987.375 ;
        RECT 3319.590 4987.205 3319.880 4987.375 ;
        RECT 3320.050 4987.205 3320.340 4987.375 ;
        RECT 3320.510 4987.205 3320.800 4987.375 ;
        RECT 3320.970 4987.205 3321.260 4987.375 ;
        RECT 3321.430 4987.205 3321.720 4987.375 ;
        RECT 3321.890 4987.205 3322.180 4987.375 ;
        RECT 3322.350 4987.205 3322.640 4987.375 ;
        RECT 3322.810 4987.205 3323.100 4987.375 ;
        RECT 3323.270 4987.205 3323.560 4987.375 ;
        RECT 3323.730 4987.205 3324.020 4987.375 ;
        RECT 3324.190 4987.205 3324.480 4987.375 ;
        RECT 3324.650 4987.205 3324.940 4987.375 ;
        RECT 3325.110 4987.205 3325.400 4987.375 ;
        RECT 3325.570 4987.205 3325.860 4987.375 ;
        RECT 3326.030 4987.205 3326.320 4987.375 ;
        RECT 3326.490 4987.205 3326.780 4987.375 ;
        RECT 3326.950 4987.205 3327.240 4987.375 ;
        RECT 3327.410 4987.205 3327.700 4987.375 ;
        RECT 3327.870 4987.205 3328.160 4987.375 ;
        RECT 3328.330 4987.205 3328.620 4987.375 ;
        RECT 3328.790 4987.205 3329.080 4987.375 ;
        RECT 3329.250 4987.205 3329.540 4987.375 ;
        RECT 3329.710 4987.205 3330.000 4987.375 ;
        RECT 3330.170 4987.205 3330.460 4987.375 ;
        RECT 3330.630 4987.205 3330.920 4987.375 ;
        RECT 3331.090 4987.205 3331.380 4987.375 ;
        RECT 3331.550 4987.205 3331.840 4987.375 ;
        RECT 3332.010 4987.205 3332.300 4987.375 ;
        RECT 3332.470 4987.205 3332.760 4987.375 ;
        RECT 3332.930 4987.205 3333.220 4987.375 ;
        RECT 3333.390 4987.205 3333.680 4987.375 ;
        RECT 3333.850 4987.205 3334.140 4987.375 ;
        RECT 3334.310 4987.205 3334.600 4987.375 ;
        RECT 3334.770 4987.205 3335.060 4987.375 ;
        RECT 3335.230 4987.205 3335.520 4987.375 ;
        RECT 3335.690 4987.205 3335.980 4987.375 ;
        RECT 3336.150 4987.205 3336.440 4987.375 ;
        RECT 3336.610 4987.205 3336.900 4987.375 ;
        RECT 3337.070 4987.205 3337.215 4987.375 ;
        RECT 2087.215 4986.625 2087.390 4986.795 ;
        RECT 2084.765 4986.455 2087.390 4986.625 ;
        RECT 2087.215 4986.255 2087.390 4986.455 ;
      LAYER li1 ;
        RECT 2087.570 4986.425 2088.670 4986.625 ;
      LAYER li1 ;
        RECT 3312.920 4986.480 3313.210 4987.205 ;
        RECT 3313.770 4986.405 3314.100 4987.205 ;
      LAYER li1 ;
        RECT 3314.270 4986.555 3314.440 4987.035 ;
      LAYER li1 ;
        RECT 3314.610 4986.725 3314.940 4987.205 ;
      LAYER li1 ;
        RECT 3315.110 4986.555 3315.280 4987.035 ;
      LAYER li1 ;
        RECT 3315.450 4986.725 3315.780 4987.205 ;
      LAYER li1 ;
        RECT 3315.950 4986.555 3316.120 4987.035 ;
      LAYER li1 ;
        RECT 3316.290 4986.725 3316.620 4987.205 ;
      LAYER li1 ;
        RECT 3316.790 4986.555 3316.960 4987.035 ;
      LAYER li1 ;
        RECT 3317.130 4986.725 3317.460 4987.205 ;
        RECT 3317.630 4986.555 3317.800 4987.030 ;
        RECT 3317.970 4986.725 3318.300 4987.205 ;
        RECT 3318.470 4986.555 3318.640 4987.035 ;
      LAYER li1 ;
        RECT 3314.270 4986.385 3316.960 4986.555 ;
      LAYER li1 ;
        RECT 3317.220 4986.385 3318.640 4986.555 ;
        RECT 3318.900 4986.480 3319.190 4987.205 ;
        RECT 3319.750 4986.405 3320.080 4987.205 ;
        RECT 3320.590 4986.725 3320.920 4987.205 ;
        RECT 3321.430 4986.725 3321.760 4987.205 ;
        RECT 3322.270 4986.725 3322.600 4987.205 ;
        RECT 3323.110 4986.725 3323.440 4987.205 ;
        RECT 3323.610 4986.555 3323.780 4987.030 ;
        RECT 3323.950 4986.725 3324.280 4987.205 ;
        RECT 3324.450 4986.555 3324.620 4987.035 ;
        RECT 3323.200 4986.385 3324.620 4986.555 ;
        RECT 3324.880 4986.480 3325.170 4987.205 ;
        RECT 3325.730 4986.405 3326.060 4987.205 ;
        RECT 3326.570 4986.725 3326.900 4987.205 ;
        RECT 3327.410 4986.725 3327.740 4987.205 ;
        RECT 3328.250 4986.725 3328.580 4987.205 ;
        RECT 3329.090 4986.725 3329.420 4987.205 ;
        RECT 3329.590 4986.555 3329.760 4987.030 ;
        RECT 3329.930 4986.725 3330.260 4987.205 ;
        RECT 3330.430 4986.555 3330.600 4987.035 ;
        RECT 3329.180 4986.385 3330.600 4986.555 ;
        RECT 3330.860 4986.480 3331.150 4987.205 ;
        RECT 3331.710 4986.405 3332.040 4987.205 ;
        RECT 3332.550 4986.725 3332.880 4987.205 ;
        RECT 3333.390 4986.725 3333.720 4987.205 ;
        RECT 3334.230 4986.725 3334.560 4987.205 ;
        RECT 3335.070 4986.725 3335.400 4987.205 ;
        RECT 3335.570 4986.555 3335.740 4987.030 ;
        RECT 3335.910 4986.725 3336.240 4987.205 ;
        RECT 3336.410 4986.555 3336.580 4987.035 ;
        RECT 3335.160 4986.385 3336.580 4986.555 ;
        RECT 3336.840 4986.480 3337.130 4987.205 ;
        RECT 834.650 4985.990 834.795 4986.160 ;
        RECT 834.965 4985.990 835.255 4986.160 ;
        RECT 835.425 4985.990 835.715 4986.160 ;
        RECT 835.885 4985.990 836.175 4986.160 ;
        RECT 836.345 4985.990 836.635 4986.160 ;
        RECT 836.805 4985.990 837.095 4986.160 ;
        RECT 837.265 4985.990 837.555 4986.160 ;
        RECT 837.725 4985.990 838.015 4986.160 ;
        RECT 838.185 4985.990 838.475 4986.160 ;
        RECT 838.645 4985.990 838.935 4986.160 ;
        RECT 839.105 4985.990 839.395 4986.160 ;
        RECT 839.565 4985.990 839.855 4986.160 ;
        RECT 840.025 4985.990 840.315 4986.160 ;
        RECT 840.485 4985.990 840.775 4986.160 ;
        RECT 840.945 4985.990 841.235 4986.160 ;
        RECT 841.405 4985.990 841.695 4986.160 ;
        RECT 841.865 4985.990 842.155 4986.160 ;
        RECT 842.325 4985.990 842.615 4986.160 ;
        RECT 842.785 4985.990 843.075 4986.160 ;
        RECT 843.245 4985.990 843.535 4986.160 ;
        RECT 843.705 4985.990 843.995 4986.160 ;
        RECT 844.165 4985.990 844.455 4986.160 ;
        RECT 844.625 4985.990 844.915 4986.160 ;
        RECT 845.085 4985.990 845.375 4986.160 ;
        RECT 845.545 4985.990 845.835 4986.160 ;
        RECT 846.005 4985.990 846.295 4986.160 ;
        RECT 846.465 4985.990 846.755 4986.160 ;
        RECT 846.925 4985.990 847.215 4986.160 ;
        RECT 847.385 4985.990 847.675 4986.160 ;
        RECT 847.845 4985.990 848.135 4986.160 ;
        RECT 848.305 4985.990 848.595 4986.160 ;
        RECT 848.765 4985.990 849.055 4986.160 ;
        RECT 849.225 4985.990 849.515 4986.160 ;
        RECT 849.685 4985.990 849.975 4986.160 ;
        RECT 850.145 4985.990 850.435 4986.160 ;
        RECT 850.605 4985.990 850.895 4986.160 ;
        RECT 851.065 4985.990 851.355 4986.160 ;
        RECT 851.525 4985.990 851.815 4986.160 ;
        RECT 851.985 4985.990 852.275 4986.160 ;
        RECT 852.445 4985.990 852.735 4986.160 ;
        RECT 852.905 4985.990 853.050 4986.160 ;
        RECT 834.735 4985.265 835.025 4985.990 ;
        RECT 835.285 4985.340 835.455 4985.820 ;
        RECT 835.625 4985.510 835.955 4985.990 ;
        RECT 836.125 4985.340 836.295 4985.815 ;
        RECT 836.465 4985.510 836.795 4985.990 ;
        RECT 837.305 4985.510 837.635 4985.990 ;
        RECT 838.145 4985.510 838.475 4985.990 ;
        RECT 838.985 4985.510 839.315 4985.990 ;
        RECT 835.285 4985.170 836.705 4985.340 ;
        RECT 839.825 4985.190 840.155 4985.990 ;
        RECT 840.715 4985.265 841.005 4985.990 ;
        RECT 841.265 4985.340 841.435 4985.820 ;
        RECT 841.605 4985.510 841.935 4985.990 ;
        RECT 842.105 4985.340 842.275 4985.815 ;
        RECT 842.445 4985.510 842.775 4985.990 ;
        RECT 843.285 4985.510 843.615 4985.990 ;
        RECT 844.125 4985.510 844.455 4985.990 ;
        RECT 844.965 4985.510 845.295 4985.990 ;
        RECT 841.265 4985.170 842.685 4985.340 ;
        RECT 845.805 4985.190 846.135 4985.990 ;
        RECT 846.695 4985.265 846.985 4985.990 ;
        RECT 847.245 4985.340 847.415 4985.820 ;
        RECT 847.585 4985.510 847.915 4985.990 ;
        RECT 848.085 4985.340 848.255 4985.815 ;
        RECT 848.425 4985.510 848.755 4985.990 ;
        RECT 849.265 4985.510 849.595 4985.990 ;
        RECT 850.105 4985.510 850.435 4985.990 ;
        RECT 850.945 4985.510 851.275 4985.990 ;
        RECT 847.245 4985.170 848.665 4985.340 ;
        RECT 851.785 4985.190 852.115 4985.990 ;
        RECT 852.675 4985.265 852.965 4985.990 ;
        RECT 836.530 4985.000 836.705 4985.170 ;
        RECT 842.510 4985.000 842.685 4985.170 ;
        RECT 848.490 4985.000 848.665 4985.170 ;
        RECT 2082.915 4985.065 2083.205 4986.230 ;
        RECT 2083.765 4985.065 2084.095 4986.215 ;
        RECT 2087.215 4986.085 2088.715 4986.255 ;
        RECT 2084.605 4985.065 2084.935 4985.865 ;
        RECT 2085.445 4985.065 2085.775 4985.865 ;
        RECT 2086.285 4985.065 2086.615 4985.865 ;
        RECT 2087.205 4985.065 2087.375 4985.865 ;
        RECT 2087.545 4985.235 2087.875 4986.085 ;
        RECT 2088.045 4985.065 2088.215 4985.865 ;
        RECT 2088.385 4985.235 2088.715 4986.085 ;
        RECT 2088.895 4985.065 2089.185 4986.230 ;
      LAYER li1 ;
        RECT 3314.270 4985.845 3314.525 4986.385 ;
      LAYER li1 ;
        RECT 3317.220 4986.215 3317.395 4986.385 ;
        RECT 3323.200 4986.215 3323.375 4986.385 ;
        RECT 3329.180 4986.215 3329.355 4986.385 ;
        RECT 3335.160 4986.215 3335.335 4986.385 ;
        RECT 3314.770 4986.045 3317.395 4986.215 ;
        RECT 3317.220 4985.845 3317.395 4986.045 ;
      LAYER li1 ;
        RECT 3317.575 4986.015 3318.675 4986.215 ;
      LAYER li1 ;
        RECT 3320.750 4986.045 3323.375 4986.215 ;
        RECT 3323.200 4985.845 3323.375 4986.045 ;
      LAYER li1 ;
        RECT 3323.555 4986.015 3324.655 4986.215 ;
      LAYER li1 ;
        RECT 3326.730 4986.045 3329.355 4986.215 ;
        RECT 3329.180 4985.845 3329.355 4986.045 ;
      LAYER li1 ;
        RECT 3329.535 4986.015 3330.635 4986.215 ;
      LAYER li1 ;
        RECT 3332.710 4986.045 3335.335 4986.215 ;
        RECT 3335.160 4985.845 3335.335 4986.045 ;
      LAYER li1 ;
        RECT 3335.515 4986.015 3336.615 4986.215 ;
        RECT 835.250 4984.800 836.350 4985.000 ;
      LAYER li1 ;
        RECT 836.530 4984.830 839.155 4985.000 ;
        RECT 836.530 4984.630 836.705 4984.830 ;
      LAYER li1 ;
        RECT 841.230 4984.800 842.330 4985.000 ;
      LAYER li1 ;
        RECT 842.510 4984.830 845.135 4985.000 ;
        RECT 842.510 4984.630 842.685 4984.830 ;
      LAYER li1 ;
        RECT 847.210 4984.800 848.310 4985.000 ;
      LAYER li1 ;
        RECT 848.490 4984.830 851.115 4985.000 ;
        RECT 2082.830 4984.895 2082.975 4985.065 ;
        RECT 2083.145 4984.895 2083.435 4985.065 ;
        RECT 2083.605 4984.895 2083.895 4985.065 ;
        RECT 2084.065 4984.895 2084.355 4985.065 ;
        RECT 2084.525 4984.895 2084.815 4985.065 ;
        RECT 2084.985 4984.895 2085.275 4985.065 ;
        RECT 2085.445 4984.895 2085.735 4985.065 ;
        RECT 2085.905 4984.895 2086.195 4985.065 ;
        RECT 2086.365 4984.895 2086.655 4985.065 ;
        RECT 2086.825 4984.895 2087.115 4985.065 ;
        RECT 2087.285 4984.895 2087.575 4985.065 ;
        RECT 2087.745 4984.895 2088.035 4985.065 ;
        RECT 2088.205 4984.895 2088.495 4985.065 ;
        RECT 2088.665 4984.895 2088.955 4985.065 ;
        RECT 2089.125 4984.895 2089.270 4985.065 ;
        RECT 848.490 4984.630 848.665 4984.830 ;
        RECT 834.735 4983.440 835.025 4984.605 ;
        RECT 835.205 4984.460 836.705 4984.630 ;
        RECT 835.205 4983.610 835.535 4984.460 ;
        RECT 835.705 4983.440 835.875 4984.240 ;
        RECT 836.045 4983.610 836.375 4984.460 ;
        RECT 836.545 4983.440 836.715 4984.240 ;
        RECT 837.305 4983.440 837.635 4984.240 ;
        RECT 838.145 4983.440 838.475 4984.240 ;
        RECT 838.985 4983.440 839.315 4984.240 ;
        RECT 839.825 4983.440 840.155 4984.590 ;
        RECT 840.715 4983.440 841.005 4984.605 ;
        RECT 841.185 4984.460 842.685 4984.630 ;
        RECT 841.185 4983.610 841.515 4984.460 ;
        RECT 841.685 4983.440 841.855 4984.240 ;
        RECT 842.025 4983.610 842.355 4984.460 ;
        RECT 842.525 4983.440 842.695 4984.240 ;
        RECT 843.285 4983.440 843.615 4984.240 ;
        RECT 844.125 4983.440 844.455 4984.240 ;
        RECT 844.965 4983.440 845.295 4984.240 ;
        RECT 845.805 4983.440 846.135 4984.590 ;
        RECT 846.695 4983.440 846.985 4984.605 ;
        RECT 847.165 4984.460 848.665 4984.630 ;
        RECT 847.165 4983.610 847.495 4984.460 ;
        RECT 847.665 4983.440 847.835 4984.240 ;
        RECT 848.005 4983.610 848.335 4984.460 ;
        RECT 848.505 4983.440 848.675 4984.240 ;
        RECT 849.265 4983.440 849.595 4984.240 ;
        RECT 850.105 4983.440 850.435 4984.240 ;
        RECT 850.945 4983.440 851.275 4984.240 ;
        RECT 851.785 4983.440 852.115 4984.590 ;
        RECT 852.675 4983.440 852.965 4984.605 ;
        RECT 2082.915 4983.730 2083.205 4984.895 ;
        RECT 2083.385 4983.875 2083.715 4984.725 ;
        RECT 2083.885 4984.095 2084.055 4984.895 ;
        RECT 2084.225 4983.875 2084.555 4984.725 ;
        RECT 2084.725 4984.095 2084.895 4984.895 ;
      LAYER li1 ;
        RECT 2085.145 4983.875 2085.315 4984.725 ;
      LAYER li1 ;
        RECT 2085.485 4984.095 2085.815 4984.895 ;
      LAYER li1 ;
        RECT 2085.985 4983.875 2086.155 4984.725 ;
      LAYER li1 ;
        RECT 2086.325 4984.095 2086.655 4984.895 ;
      LAYER li1 ;
        RECT 2086.825 4983.875 2086.995 4984.725 ;
      LAYER li1 ;
        RECT 2087.165 4984.095 2087.495 4984.895 ;
      LAYER li1 ;
        RECT 2087.665 4983.875 2087.835 4984.725 ;
      LAYER li1 ;
        RECT 2083.385 4983.705 2084.885 4983.875 ;
      LAYER li1 ;
        RECT 2085.145 4983.705 2087.835 4983.875 ;
      LAYER li1 ;
        RECT 2088.005 4983.745 2088.335 4984.895 ;
        RECT 2088.895 4983.730 2089.185 4984.895 ;
        RECT 3312.920 4984.655 3313.210 4985.820 ;
        RECT 3313.770 4984.655 3314.100 4985.805 ;
      LAYER li1 ;
        RECT 3314.270 4985.675 3316.960 4985.845 ;
      LAYER li1 ;
        RECT 3317.220 4985.675 3318.720 4985.845 ;
      LAYER li1 ;
        RECT 3314.270 4984.825 3314.440 4985.675 ;
      LAYER li1 ;
        RECT 3314.610 4984.655 3314.940 4985.455 ;
      LAYER li1 ;
        RECT 3315.110 4984.825 3315.280 4985.675 ;
      LAYER li1 ;
        RECT 3315.450 4984.655 3315.780 4985.455 ;
      LAYER li1 ;
        RECT 3315.950 4984.825 3316.120 4985.675 ;
      LAYER li1 ;
        RECT 3316.290 4984.655 3316.620 4985.455 ;
      LAYER li1 ;
        RECT 3316.790 4984.825 3316.960 4985.675 ;
      LAYER li1 ;
        RECT 3317.210 4984.655 3317.380 4985.455 ;
        RECT 3317.550 4984.825 3317.880 4985.675 ;
        RECT 3318.050 4984.655 3318.220 4985.455 ;
        RECT 3318.390 4984.825 3318.720 4985.675 ;
        RECT 3318.900 4984.655 3319.190 4985.820 ;
        RECT 3319.750 4984.655 3320.080 4985.805 ;
        RECT 3323.200 4985.675 3324.700 4985.845 ;
        RECT 3320.590 4984.655 3320.920 4985.455 ;
        RECT 3321.430 4984.655 3321.760 4985.455 ;
        RECT 3322.270 4984.655 3322.600 4985.455 ;
        RECT 3323.190 4984.655 3323.360 4985.455 ;
        RECT 3323.530 4984.825 3323.860 4985.675 ;
        RECT 3324.030 4984.655 3324.200 4985.455 ;
        RECT 3324.370 4984.825 3324.700 4985.675 ;
        RECT 3324.880 4984.655 3325.170 4985.820 ;
        RECT 3325.730 4984.655 3326.060 4985.805 ;
        RECT 3329.180 4985.675 3330.680 4985.845 ;
        RECT 3326.570 4984.655 3326.900 4985.455 ;
        RECT 3327.410 4984.655 3327.740 4985.455 ;
        RECT 3328.250 4984.655 3328.580 4985.455 ;
        RECT 3329.170 4984.655 3329.340 4985.455 ;
        RECT 3329.510 4984.825 3329.840 4985.675 ;
        RECT 3330.010 4984.655 3330.180 4985.455 ;
        RECT 3330.350 4984.825 3330.680 4985.675 ;
        RECT 3330.860 4984.655 3331.150 4985.820 ;
        RECT 3331.710 4984.655 3332.040 4985.805 ;
        RECT 3335.160 4985.675 3336.660 4985.845 ;
        RECT 3332.550 4984.655 3332.880 4985.455 ;
        RECT 3333.390 4984.655 3333.720 4985.455 ;
        RECT 3334.230 4984.655 3334.560 4985.455 ;
        RECT 3335.150 4984.655 3335.320 4985.455 ;
        RECT 3335.490 4984.825 3335.820 4985.675 ;
        RECT 3335.990 4984.655 3336.160 4985.455 ;
        RECT 3336.330 4984.825 3336.660 4985.675 ;
        RECT 3336.840 4984.655 3337.130 4985.820 ;
        RECT 3312.835 4984.485 3312.980 4984.655 ;
        RECT 3313.150 4984.485 3313.440 4984.655 ;
        RECT 3313.610 4984.485 3313.900 4984.655 ;
        RECT 3314.070 4984.485 3314.360 4984.655 ;
        RECT 3314.530 4984.485 3314.820 4984.655 ;
        RECT 3314.990 4984.485 3315.280 4984.655 ;
        RECT 3315.450 4984.485 3315.740 4984.655 ;
        RECT 3315.910 4984.485 3316.200 4984.655 ;
        RECT 3316.370 4984.485 3316.660 4984.655 ;
        RECT 3316.830 4984.485 3317.120 4984.655 ;
        RECT 3317.290 4984.485 3317.580 4984.655 ;
        RECT 3317.750 4984.485 3318.040 4984.655 ;
        RECT 3318.210 4984.485 3318.500 4984.655 ;
        RECT 3318.670 4984.485 3318.960 4984.655 ;
        RECT 3319.130 4984.485 3319.420 4984.655 ;
        RECT 3319.590 4984.485 3319.880 4984.655 ;
        RECT 3320.050 4984.485 3320.340 4984.655 ;
        RECT 3320.510 4984.485 3320.800 4984.655 ;
        RECT 3320.970 4984.485 3321.260 4984.655 ;
        RECT 3321.430 4984.485 3321.720 4984.655 ;
        RECT 3321.890 4984.485 3322.180 4984.655 ;
        RECT 3322.350 4984.485 3322.640 4984.655 ;
        RECT 3322.810 4984.485 3323.100 4984.655 ;
        RECT 3323.270 4984.485 3323.560 4984.655 ;
        RECT 3323.730 4984.485 3324.020 4984.655 ;
        RECT 3324.190 4984.485 3324.480 4984.655 ;
        RECT 3324.650 4984.485 3324.940 4984.655 ;
        RECT 3325.110 4984.485 3325.400 4984.655 ;
        RECT 3325.570 4984.485 3325.860 4984.655 ;
        RECT 3326.030 4984.485 3326.320 4984.655 ;
        RECT 3326.490 4984.485 3326.780 4984.655 ;
        RECT 3326.950 4984.485 3327.240 4984.655 ;
        RECT 3327.410 4984.485 3327.700 4984.655 ;
        RECT 3327.870 4984.485 3328.160 4984.655 ;
        RECT 3328.330 4984.485 3328.620 4984.655 ;
        RECT 3328.790 4984.485 3329.080 4984.655 ;
        RECT 3329.250 4984.485 3329.540 4984.655 ;
        RECT 3329.710 4984.485 3330.000 4984.655 ;
        RECT 3330.170 4984.485 3330.460 4984.655 ;
        RECT 3330.630 4984.485 3330.920 4984.655 ;
        RECT 3331.090 4984.485 3331.380 4984.655 ;
        RECT 3331.550 4984.485 3331.840 4984.655 ;
        RECT 3332.010 4984.485 3332.300 4984.655 ;
        RECT 3332.470 4984.485 3332.760 4984.655 ;
        RECT 3332.930 4984.485 3333.220 4984.655 ;
        RECT 3333.390 4984.485 3333.680 4984.655 ;
        RECT 3333.850 4984.485 3334.140 4984.655 ;
        RECT 3334.310 4984.485 3334.600 4984.655 ;
        RECT 3334.770 4984.485 3335.060 4984.655 ;
        RECT 3335.230 4984.485 3335.520 4984.655 ;
        RECT 3335.690 4984.485 3335.980 4984.655 ;
        RECT 3336.150 4984.485 3336.440 4984.655 ;
        RECT 3336.610 4984.485 3336.900 4984.655 ;
        RECT 3337.070 4984.485 3337.215 4984.655 ;
        RECT 2084.710 4983.505 2084.885 4983.705 ;
        RECT 834.650 4983.270 834.795 4983.440 ;
        RECT 834.965 4983.270 835.255 4983.440 ;
        RECT 835.425 4983.270 835.715 4983.440 ;
        RECT 835.885 4983.270 836.175 4983.440 ;
        RECT 836.345 4983.270 836.635 4983.440 ;
        RECT 836.805 4983.270 837.095 4983.440 ;
        RECT 837.265 4983.270 837.555 4983.440 ;
        RECT 837.725 4983.270 838.015 4983.440 ;
        RECT 838.185 4983.270 838.475 4983.440 ;
        RECT 838.645 4983.270 838.935 4983.440 ;
        RECT 839.105 4983.270 839.395 4983.440 ;
        RECT 839.565 4983.270 839.855 4983.440 ;
        RECT 840.025 4983.270 840.315 4983.440 ;
        RECT 840.485 4983.270 840.775 4983.440 ;
        RECT 840.945 4983.270 841.235 4983.440 ;
        RECT 841.405 4983.270 841.695 4983.440 ;
        RECT 841.865 4983.270 842.155 4983.440 ;
        RECT 842.325 4983.270 842.615 4983.440 ;
        RECT 842.785 4983.270 843.075 4983.440 ;
        RECT 843.245 4983.270 843.535 4983.440 ;
        RECT 843.705 4983.270 843.995 4983.440 ;
        RECT 844.165 4983.270 844.455 4983.440 ;
        RECT 844.625 4983.270 844.915 4983.440 ;
        RECT 845.085 4983.270 845.375 4983.440 ;
        RECT 845.545 4983.270 845.835 4983.440 ;
        RECT 846.005 4983.270 846.295 4983.440 ;
        RECT 846.465 4983.270 846.755 4983.440 ;
        RECT 846.925 4983.270 847.215 4983.440 ;
        RECT 847.385 4983.270 847.675 4983.440 ;
        RECT 847.845 4983.270 848.135 4983.440 ;
        RECT 848.305 4983.270 848.595 4983.440 ;
        RECT 848.765 4983.270 849.055 4983.440 ;
        RECT 849.225 4983.270 849.515 4983.440 ;
        RECT 849.685 4983.270 849.975 4983.440 ;
        RECT 850.145 4983.270 850.435 4983.440 ;
        RECT 850.605 4983.270 850.895 4983.440 ;
        RECT 851.065 4983.270 851.355 4983.440 ;
        RECT 851.525 4983.270 851.815 4983.440 ;
        RECT 851.985 4983.270 852.275 4983.440 ;
        RECT 852.445 4983.270 852.735 4983.440 ;
        RECT 852.905 4983.270 853.050 4983.440 ;
        RECT 2084.710 4983.335 2087.335 4983.505 ;
        RECT 834.735 4982.105 835.025 4983.270 ;
        RECT 835.585 4982.120 835.915 4983.270 ;
      LAYER li1 ;
        RECT 836.085 4982.250 836.255 4983.100 ;
      LAYER li1 ;
        RECT 836.425 4982.470 836.755 4983.270 ;
      LAYER li1 ;
        RECT 836.925 4982.250 837.095 4983.100 ;
      LAYER li1 ;
        RECT 837.265 4982.470 837.595 4983.270 ;
      LAYER li1 ;
        RECT 837.765 4982.250 837.935 4983.100 ;
      LAYER li1 ;
        RECT 838.105 4982.470 838.435 4983.270 ;
      LAYER li1 ;
        RECT 838.605 4982.250 838.775 4983.100 ;
      LAYER li1 ;
        RECT 839.025 4982.470 839.195 4983.270 ;
        RECT 839.365 4982.250 839.695 4983.100 ;
        RECT 839.865 4982.470 840.035 4983.270 ;
        RECT 840.205 4982.250 840.535 4983.100 ;
      LAYER li1 ;
        RECT 836.085 4982.080 838.775 4982.250 ;
      LAYER li1 ;
        RECT 839.035 4982.080 840.535 4982.250 ;
        RECT 840.715 4982.105 841.005 4983.270 ;
        RECT 841.565 4982.120 841.895 4983.270 ;
      LAYER li1 ;
        RECT 842.065 4982.250 842.235 4983.100 ;
      LAYER li1 ;
        RECT 842.405 4982.470 842.735 4983.270 ;
      LAYER li1 ;
        RECT 842.905 4982.250 843.075 4983.100 ;
      LAYER li1 ;
        RECT 843.245 4982.470 843.575 4983.270 ;
      LAYER li1 ;
        RECT 843.745 4982.250 843.915 4983.100 ;
      LAYER li1 ;
        RECT 844.085 4982.470 844.415 4983.270 ;
      LAYER li1 ;
        RECT 844.585 4982.250 844.755 4983.100 ;
      LAYER li1 ;
        RECT 845.005 4982.470 845.175 4983.270 ;
        RECT 845.345 4982.250 845.675 4983.100 ;
        RECT 845.845 4982.470 846.015 4983.270 ;
        RECT 846.185 4982.250 846.515 4983.100 ;
      LAYER li1 ;
        RECT 842.065 4982.080 844.755 4982.250 ;
      LAYER li1 ;
        RECT 845.015 4982.080 846.515 4982.250 ;
        RECT 846.695 4982.105 846.985 4983.270 ;
        RECT 847.545 4982.120 847.875 4983.270 ;
      LAYER li1 ;
        RECT 848.045 4982.250 848.215 4983.100 ;
      LAYER li1 ;
        RECT 848.385 4982.470 848.715 4983.270 ;
      LAYER li1 ;
        RECT 848.885 4982.250 849.055 4983.100 ;
      LAYER li1 ;
        RECT 849.225 4982.470 849.555 4983.270 ;
      LAYER li1 ;
        RECT 849.725 4982.250 849.895 4983.100 ;
      LAYER li1 ;
        RECT 850.065 4982.470 850.395 4983.270 ;
      LAYER li1 ;
        RECT 850.565 4982.250 850.735 4983.100 ;
      LAYER li1 ;
        RECT 850.985 4982.470 851.155 4983.270 ;
        RECT 851.325 4982.250 851.655 4983.100 ;
        RECT 851.825 4982.470 851.995 4983.270 ;
        RECT 852.165 4982.250 852.495 4983.100 ;
      LAYER li1 ;
        RECT 848.045 4982.080 850.735 4982.250 ;
      LAYER li1 ;
        RECT 850.995 4982.080 852.495 4982.250 ;
        RECT 852.675 4982.105 852.965 4983.270 ;
        RECT 2084.710 4983.165 2084.885 4983.335 ;
      LAYER li1 ;
        RECT 2087.580 4983.165 2087.835 4983.705 ;
      LAYER li1 ;
        RECT 3312.920 4983.320 3313.210 4984.485 ;
        RECT 3313.390 4983.465 3313.720 4984.315 ;
        RECT 3313.890 4983.685 3314.060 4984.485 ;
        RECT 3314.230 4983.465 3314.560 4984.315 ;
        RECT 3314.730 4983.685 3314.900 4984.485 ;
      LAYER li1 ;
        RECT 3315.150 4983.465 3315.320 4984.315 ;
      LAYER li1 ;
        RECT 3315.490 4983.685 3315.820 4984.485 ;
      LAYER li1 ;
        RECT 3315.990 4983.465 3316.160 4984.315 ;
      LAYER li1 ;
        RECT 3316.330 4983.685 3316.660 4984.485 ;
      LAYER li1 ;
        RECT 3316.830 4983.465 3317.000 4984.315 ;
      LAYER li1 ;
        RECT 3317.170 4983.685 3317.500 4984.485 ;
      LAYER li1 ;
        RECT 3317.670 4983.465 3317.840 4984.315 ;
      LAYER li1 ;
        RECT 3313.390 4983.295 3314.890 4983.465 ;
      LAYER li1 ;
        RECT 3315.150 4983.295 3317.840 4983.465 ;
      LAYER li1 ;
        RECT 3318.010 4983.335 3318.340 4984.485 ;
        RECT 3318.900 4983.320 3319.190 4984.485 ;
        RECT 3319.370 4983.465 3319.700 4984.315 ;
        RECT 3319.870 4983.685 3320.040 4984.485 ;
        RECT 3320.210 4983.465 3320.540 4984.315 ;
        RECT 3320.710 4983.685 3320.880 4984.485 ;
      LAYER li1 ;
        RECT 3321.130 4983.465 3321.300 4984.315 ;
      LAYER li1 ;
        RECT 3321.470 4983.685 3321.800 4984.485 ;
      LAYER li1 ;
        RECT 3321.970 4983.465 3322.140 4984.315 ;
      LAYER li1 ;
        RECT 3322.310 4983.685 3322.640 4984.485 ;
      LAYER li1 ;
        RECT 3322.810 4983.465 3322.980 4984.315 ;
      LAYER li1 ;
        RECT 3323.150 4983.685 3323.480 4984.485 ;
      LAYER li1 ;
        RECT 3323.650 4983.465 3323.820 4984.315 ;
      LAYER li1 ;
        RECT 3319.370 4983.295 3320.870 4983.465 ;
      LAYER li1 ;
        RECT 3321.130 4983.295 3323.820 4983.465 ;
      LAYER li1 ;
        RECT 3323.990 4983.335 3324.320 4984.485 ;
        RECT 3324.880 4983.320 3325.170 4984.485 ;
        RECT 3325.350 4983.465 3325.680 4984.315 ;
        RECT 3325.850 4983.685 3326.020 4984.485 ;
        RECT 3326.190 4983.465 3326.520 4984.315 ;
        RECT 3326.690 4983.685 3326.860 4984.485 ;
      LAYER li1 ;
        RECT 3327.110 4983.465 3327.280 4984.315 ;
      LAYER li1 ;
        RECT 3327.450 4983.685 3327.780 4984.485 ;
      LAYER li1 ;
        RECT 3327.950 4983.465 3328.120 4984.315 ;
      LAYER li1 ;
        RECT 3328.290 4983.685 3328.620 4984.485 ;
      LAYER li1 ;
        RECT 3328.790 4983.465 3328.960 4984.315 ;
      LAYER li1 ;
        RECT 3329.130 4983.685 3329.460 4984.485 ;
      LAYER li1 ;
        RECT 3329.630 4983.465 3329.800 4984.315 ;
      LAYER li1 ;
        RECT 3325.350 4983.295 3326.850 4983.465 ;
      LAYER li1 ;
        RECT 3327.110 4983.295 3329.800 4983.465 ;
      LAYER li1 ;
        RECT 3329.970 4983.335 3330.300 4984.485 ;
        RECT 3330.860 4983.320 3331.150 4984.485 ;
        RECT 3331.330 4983.465 3331.660 4984.315 ;
        RECT 3331.830 4983.685 3332.000 4984.485 ;
        RECT 3332.170 4983.465 3332.500 4984.315 ;
        RECT 3332.670 4983.685 3332.840 4984.485 ;
      LAYER li1 ;
        RECT 3333.090 4983.465 3333.260 4984.315 ;
      LAYER li1 ;
        RECT 3333.430 4983.685 3333.760 4984.485 ;
      LAYER li1 ;
        RECT 3333.930 4983.465 3334.100 4984.315 ;
      LAYER li1 ;
        RECT 3334.270 4983.685 3334.600 4984.485 ;
      LAYER li1 ;
        RECT 3334.770 4983.465 3334.940 4984.315 ;
      LAYER li1 ;
        RECT 3335.110 4983.685 3335.440 4984.485 ;
      LAYER li1 ;
        RECT 3335.610 4983.465 3335.780 4984.315 ;
      LAYER li1 ;
        RECT 3331.330 4983.295 3332.830 4983.465 ;
      LAYER li1 ;
        RECT 3333.090 4983.295 3335.780 4983.465 ;
      LAYER li1 ;
        RECT 3335.950 4983.335 3336.280 4984.485 ;
        RECT 3336.840 4983.320 3337.130 4984.485 ;
        RECT 2082.915 4982.345 2083.205 4983.070 ;
        RECT 2083.465 4982.995 2084.885 4983.165 ;
      LAYER li1 ;
        RECT 2085.145 4982.995 2087.835 4983.165 ;
      LAYER li1 ;
        RECT 2083.465 4982.515 2083.635 4982.995 ;
        RECT 2083.805 4982.345 2084.135 4982.825 ;
        RECT 2084.305 4982.520 2084.475 4982.995 ;
        RECT 2084.645 4982.345 2084.975 4982.825 ;
      LAYER li1 ;
        RECT 2085.145 4982.515 2085.315 4982.995 ;
      LAYER li1 ;
        RECT 2085.485 4982.345 2085.815 4982.825 ;
      LAYER li1 ;
        RECT 2085.985 4982.515 2086.155 4982.995 ;
      LAYER li1 ;
        RECT 2086.325 4982.345 2086.655 4982.825 ;
      LAYER li1 ;
        RECT 2086.825 4982.515 2086.995 4982.995 ;
      LAYER li1 ;
        RECT 2087.165 4982.345 2087.495 4982.825 ;
      LAYER li1 ;
        RECT 2087.665 4982.515 2087.835 4982.995 ;
      LAYER li1 ;
        RECT 2088.005 4982.345 2088.335 4983.145 ;
        RECT 2088.895 4982.345 2089.185 4983.070 ;
      LAYER li1 ;
        RECT 3312.945 4982.925 3314.535 4983.125 ;
      LAYER li1 ;
        RECT 3314.715 4983.095 3314.890 4983.295 ;
        RECT 3314.715 4982.925 3317.340 4983.095 ;
        RECT 3314.715 4982.755 3314.890 4982.925 ;
      LAYER li1 ;
        RECT 3317.585 4982.755 3317.840 4983.295 ;
      LAYER li1 ;
        RECT 3320.695 4983.095 3320.870 4983.295 ;
        RECT 3320.695 4982.925 3323.320 4983.095 ;
        RECT 3320.695 4982.755 3320.870 4982.925 ;
      LAYER li1 ;
        RECT 3323.565 4982.755 3323.820 4983.295 ;
      LAYER li1 ;
        RECT 3326.675 4983.095 3326.850 4983.295 ;
        RECT 3326.675 4982.925 3329.300 4983.095 ;
        RECT 3326.675 4982.755 3326.850 4982.925 ;
      LAYER li1 ;
        RECT 3329.545 4982.755 3329.800 4983.295 ;
      LAYER li1 ;
        RECT 3332.655 4983.095 3332.830 4983.295 ;
        RECT 3332.655 4982.925 3335.280 4983.095 ;
        RECT 3332.655 4982.755 3332.830 4982.925 ;
      LAYER li1 ;
        RECT 3335.525 4982.755 3335.780 4983.295 ;
      LAYER li1 ;
        RECT 2082.830 4982.175 2082.975 4982.345 ;
        RECT 2083.145 4982.175 2083.435 4982.345 ;
        RECT 2083.605 4982.175 2083.895 4982.345 ;
        RECT 2084.065 4982.175 2084.355 4982.345 ;
        RECT 2084.525 4982.175 2084.815 4982.345 ;
        RECT 2084.985 4982.175 2085.275 4982.345 ;
        RECT 2085.445 4982.175 2085.735 4982.345 ;
        RECT 2085.905 4982.175 2086.195 4982.345 ;
        RECT 2086.365 4982.175 2086.655 4982.345 ;
        RECT 2086.825 4982.175 2087.115 4982.345 ;
        RECT 2087.285 4982.175 2087.575 4982.345 ;
        RECT 2087.745 4982.175 2088.035 4982.345 ;
        RECT 2088.205 4982.175 2088.495 4982.345 ;
        RECT 2088.665 4982.175 2088.955 4982.345 ;
        RECT 2089.125 4982.175 2089.270 4982.345 ;
      LAYER li1 ;
        RECT 836.085 4981.540 836.340 4982.080 ;
      LAYER li1 ;
        RECT 839.035 4981.880 839.210 4982.080 ;
        RECT 836.585 4981.710 839.210 4981.880 ;
        RECT 839.035 4981.540 839.210 4981.710 ;
      LAYER li1 ;
        RECT 842.065 4981.540 842.320 4982.080 ;
      LAYER li1 ;
        RECT 845.015 4981.880 845.190 4982.080 ;
        RECT 842.565 4981.710 845.190 4981.880 ;
        RECT 845.015 4981.540 845.190 4981.710 ;
      LAYER li1 ;
        RECT 848.045 4981.540 848.300 4982.080 ;
      LAYER li1 ;
        RECT 850.995 4981.880 851.170 4982.080 ;
        RECT 3312.920 4981.935 3313.210 4982.660 ;
        RECT 3313.470 4982.585 3314.890 4982.755 ;
      LAYER li1 ;
        RECT 3315.150 4982.585 3317.840 4982.755 ;
      LAYER li1 ;
        RECT 3313.470 4982.105 3313.640 4982.585 ;
        RECT 3313.810 4981.935 3314.140 4982.415 ;
        RECT 3314.310 4982.110 3314.480 4982.585 ;
        RECT 3314.650 4981.935 3314.980 4982.415 ;
      LAYER li1 ;
        RECT 3315.150 4982.105 3315.320 4982.585 ;
      LAYER li1 ;
        RECT 3315.490 4981.935 3315.820 4982.415 ;
      LAYER li1 ;
        RECT 3315.990 4982.105 3316.160 4982.585 ;
      LAYER li1 ;
        RECT 3316.330 4981.935 3316.660 4982.415 ;
      LAYER li1 ;
        RECT 3316.830 4982.105 3317.000 4982.585 ;
      LAYER li1 ;
        RECT 3317.170 4981.935 3317.500 4982.415 ;
      LAYER li1 ;
        RECT 3317.670 4982.105 3317.840 4982.585 ;
      LAYER li1 ;
        RECT 3318.010 4981.935 3318.340 4982.735 ;
        RECT 3318.900 4981.935 3319.190 4982.660 ;
        RECT 3319.450 4982.585 3320.870 4982.755 ;
      LAYER li1 ;
        RECT 3321.130 4982.585 3323.820 4982.755 ;
      LAYER li1 ;
        RECT 3319.450 4982.105 3319.620 4982.585 ;
        RECT 3319.790 4981.935 3320.120 4982.415 ;
        RECT 3320.290 4982.110 3320.460 4982.585 ;
        RECT 3320.630 4981.935 3320.960 4982.415 ;
      LAYER li1 ;
        RECT 3321.130 4982.105 3321.300 4982.585 ;
      LAYER li1 ;
        RECT 3321.470 4981.935 3321.800 4982.415 ;
      LAYER li1 ;
        RECT 3321.970 4982.105 3322.140 4982.585 ;
      LAYER li1 ;
        RECT 3322.310 4981.935 3322.640 4982.415 ;
      LAYER li1 ;
        RECT 3322.810 4982.105 3322.980 4982.585 ;
      LAYER li1 ;
        RECT 3323.150 4981.935 3323.480 4982.415 ;
      LAYER li1 ;
        RECT 3323.650 4982.105 3323.820 4982.585 ;
      LAYER li1 ;
        RECT 3323.990 4981.935 3324.320 4982.735 ;
        RECT 3324.880 4981.935 3325.170 4982.660 ;
        RECT 3325.430 4982.585 3326.850 4982.755 ;
      LAYER li1 ;
        RECT 3327.110 4982.585 3329.800 4982.755 ;
      LAYER li1 ;
        RECT 3325.430 4982.105 3325.600 4982.585 ;
        RECT 3325.770 4981.935 3326.100 4982.415 ;
        RECT 3326.270 4982.110 3326.440 4982.585 ;
        RECT 3326.610 4981.935 3326.940 4982.415 ;
      LAYER li1 ;
        RECT 3327.110 4982.105 3327.280 4982.585 ;
      LAYER li1 ;
        RECT 3327.450 4981.935 3327.780 4982.415 ;
      LAYER li1 ;
        RECT 3327.950 4982.105 3328.120 4982.585 ;
      LAYER li1 ;
        RECT 3328.290 4981.935 3328.620 4982.415 ;
      LAYER li1 ;
        RECT 3328.790 4982.105 3328.960 4982.585 ;
      LAYER li1 ;
        RECT 3329.130 4981.935 3329.460 4982.415 ;
      LAYER li1 ;
        RECT 3329.630 4982.105 3329.800 4982.585 ;
      LAYER li1 ;
        RECT 3329.970 4981.935 3330.300 4982.735 ;
        RECT 3330.860 4981.935 3331.150 4982.660 ;
        RECT 3331.410 4982.585 3332.830 4982.755 ;
      LAYER li1 ;
        RECT 3333.090 4982.585 3335.780 4982.755 ;
      LAYER li1 ;
        RECT 3331.410 4982.105 3331.580 4982.585 ;
        RECT 3331.750 4981.935 3332.080 4982.415 ;
        RECT 3332.250 4982.110 3332.420 4982.585 ;
        RECT 3332.590 4981.935 3332.920 4982.415 ;
      LAYER li1 ;
        RECT 3333.090 4982.105 3333.260 4982.585 ;
      LAYER li1 ;
        RECT 3333.430 4981.935 3333.760 4982.415 ;
      LAYER li1 ;
        RECT 3333.930 4982.105 3334.100 4982.585 ;
      LAYER li1 ;
        RECT 3334.270 4981.935 3334.600 4982.415 ;
      LAYER li1 ;
        RECT 3334.770 4982.105 3334.940 4982.585 ;
      LAYER li1 ;
        RECT 3335.110 4981.935 3335.440 4982.415 ;
      LAYER li1 ;
        RECT 3335.610 4982.105 3335.780 4982.585 ;
      LAYER li1 ;
        RECT 3335.950 4981.935 3336.280 4982.735 ;
        RECT 3336.840 4981.935 3337.130 4982.660 ;
        RECT 848.545 4981.710 851.170 4981.880 ;
        RECT 3312.835 4981.765 3312.980 4981.935 ;
        RECT 3313.150 4981.765 3313.440 4981.935 ;
        RECT 3313.610 4981.765 3313.900 4981.935 ;
        RECT 3314.070 4981.765 3314.360 4981.935 ;
        RECT 3314.530 4981.765 3314.820 4981.935 ;
        RECT 3314.990 4981.765 3315.280 4981.935 ;
        RECT 3315.450 4981.765 3315.740 4981.935 ;
        RECT 3315.910 4981.765 3316.200 4981.935 ;
        RECT 3316.370 4981.765 3316.660 4981.935 ;
        RECT 3316.830 4981.765 3317.120 4981.935 ;
        RECT 3317.290 4981.765 3317.580 4981.935 ;
        RECT 3317.750 4981.765 3318.040 4981.935 ;
        RECT 3318.210 4981.765 3318.500 4981.935 ;
        RECT 3318.670 4981.765 3318.960 4981.935 ;
        RECT 3319.130 4981.765 3319.420 4981.935 ;
        RECT 3319.590 4981.765 3319.880 4981.935 ;
        RECT 3320.050 4981.765 3320.340 4981.935 ;
        RECT 3320.510 4981.765 3320.800 4981.935 ;
        RECT 3320.970 4981.765 3321.260 4981.935 ;
        RECT 3321.430 4981.765 3321.720 4981.935 ;
        RECT 3321.890 4981.765 3322.180 4981.935 ;
        RECT 3322.350 4981.765 3322.640 4981.935 ;
        RECT 3322.810 4981.765 3323.100 4981.935 ;
        RECT 3323.270 4981.765 3323.560 4981.935 ;
        RECT 3323.730 4981.765 3324.020 4981.935 ;
        RECT 3324.190 4981.765 3324.480 4981.935 ;
        RECT 3324.650 4981.765 3324.940 4981.935 ;
        RECT 3325.110 4981.765 3325.400 4981.935 ;
        RECT 3325.570 4981.765 3325.860 4981.935 ;
        RECT 3326.030 4981.765 3326.320 4981.935 ;
        RECT 3326.490 4981.765 3326.780 4981.935 ;
        RECT 3326.950 4981.765 3327.240 4981.935 ;
        RECT 3327.410 4981.765 3327.700 4981.935 ;
        RECT 3327.870 4981.765 3328.160 4981.935 ;
        RECT 3328.330 4981.765 3328.620 4981.935 ;
        RECT 3328.790 4981.765 3329.080 4981.935 ;
        RECT 3329.250 4981.765 3329.540 4981.935 ;
        RECT 3329.710 4981.765 3330.000 4981.935 ;
        RECT 3330.170 4981.765 3330.460 4981.935 ;
        RECT 3330.630 4981.765 3330.920 4981.935 ;
        RECT 3331.090 4981.765 3331.380 4981.935 ;
        RECT 3331.550 4981.765 3331.840 4981.935 ;
        RECT 3332.010 4981.765 3332.300 4981.935 ;
        RECT 3332.470 4981.765 3332.760 4981.935 ;
        RECT 3332.930 4981.765 3333.220 4981.935 ;
        RECT 3333.390 4981.765 3333.680 4981.935 ;
        RECT 3333.850 4981.765 3334.140 4981.935 ;
        RECT 3334.310 4981.765 3334.600 4981.935 ;
        RECT 3334.770 4981.765 3335.060 4981.935 ;
        RECT 3335.230 4981.765 3335.520 4981.935 ;
        RECT 3335.690 4981.765 3335.980 4981.935 ;
        RECT 3336.150 4981.765 3336.440 4981.935 ;
        RECT 3336.610 4981.765 3336.900 4981.935 ;
        RECT 3337.070 4981.765 3337.215 4981.935 ;
        RECT 850.995 4981.540 851.170 4981.710 ;
        RECT 834.735 4980.720 835.025 4981.445 ;
        RECT 835.585 4980.720 835.915 4981.520 ;
      LAYER li1 ;
        RECT 836.085 4981.370 838.775 4981.540 ;
      LAYER li1 ;
        RECT 839.035 4981.370 840.455 4981.540 ;
      LAYER li1 ;
        RECT 836.085 4980.890 836.255 4981.370 ;
      LAYER li1 ;
        RECT 836.425 4980.720 836.755 4981.200 ;
      LAYER li1 ;
        RECT 836.925 4980.890 837.095 4981.370 ;
      LAYER li1 ;
        RECT 837.265 4980.720 837.595 4981.200 ;
      LAYER li1 ;
        RECT 837.765 4980.890 837.935 4981.370 ;
      LAYER li1 ;
        RECT 838.105 4980.720 838.435 4981.200 ;
      LAYER li1 ;
        RECT 838.605 4980.890 838.775 4981.370 ;
      LAYER li1 ;
        RECT 838.945 4980.720 839.275 4981.200 ;
        RECT 839.445 4980.895 839.615 4981.370 ;
        RECT 839.785 4980.720 840.115 4981.200 ;
        RECT 840.285 4980.890 840.455 4981.370 ;
        RECT 840.715 4980.720 841.005 4981.445 ;
        RECT 841.565 4980.720 841.895 4981.520 ;
      LAYER li1 ;
        RECT 842.065 4981.370 844.755 4981.540 ;
      LAYER li1 ;
        RECT 845.015 4981.370 846.435 4981.540 ;
      LAYER li1 ;
        RECT 842.065 4980.890 842.235 4981.370 ;
      LAYER li1 ;
        RECT 842.405 4980.720 842.735 4981.200 ;
      LAYER li1 ;
        RECT 842.905 4980.890 843.075 4981.370 ;
      LAYER li1 ;
        RECT 843.245 4980.720 843.575 4981.200 ;
      LAYER li1 ;
        RECT 843.745 4980.890 843.915 4981.370 ;
      LAYER li1 ;
        RECT 844.085 4980.720 844.415 4981.200 ;
      LAYER li1 ;
        RECT 844.585 4980.890 844.755 4981.370 ;
      LAYER li1 ;
        RECT 844.925 4980.720 845.255 4981.200 ;
        RECT 845.425 4980.895 845.595 4981.370 ;
        RECT 845.765 4980.720 846.095 4981.200 ;
        RECT 846.265 4980.890 846.435 4981.370 ;
        RECT 846.695 4980.720 846.985 4981.445 ;
        RECT 847.545 4980.720 847.875 4981.520 ;
      LAYER li1 ;
        RECT 848.045 4981.370 850.735 4981.540 ;
      LAYER li1 ;
        RECT 850.995 4981.370 852.415 4981.540 ;
      LAYER li1 ;
        RECT 848.045 4980.890 848.215 4981.370 ;
      LAYER li1 ;
        RECT 848.385 4980.720 848.715 4981.200 ;
      LAYER li1 ;
        RECT 848.885 4980.890 849.055 4981.370 ;
      LAYER li1 ;
        RECT 849.225 4980.720 849.555 4981.200 ;
      LAYER li1 ;
        RECT 849.725 4980.890 849.895 4981.370 ;
      LAYER li1 ;
        RECT 850.065 4980.720 850.395 4981.200 ;
      LAYER li1 ;
        RECT 850.565 4980.890 850.735 4981.370 ;
      LAYER li1 ;
        RECT 850.905 4980.720 851.235 4981.200 ;
        RECT 851.405 4980.895 851.575 4981.370 ;
        RECT 851.745 4980.720 852.075 4981.200 ;
        RECT 852.245 4980.890 852.415 4981.370 ;
        RECT 852.675 4980.720 852.965 4981.445 ;
        RECT 834.650 4980.550 834.795 4980.720 ;
        RECT 834.965 4980.550 835.255 4980.720 ;
        RECT 835.425 4980.550 835.715 4980.720 ;
        RECT 835.885 4980.550 836.175 4980.720 ;
        RECT 836.345 4980.550 836.635 4980.720 ;
        RECT 836.805 4980.550 837.095 4980.720 ;
        RECT 837.265 4980.550 837.555 4980.720 ;
        RECT 837.725 4980.550 838.015 4980.720 ;
        RECT 838.185 4980.550 838.475 4980.720 ;
        RECT 838.645 4980.550 838.935 4980.720 ;
        RECT 839.105 4980.550 839.395 4980.720 ;
        RECT 839.565 4980.550 839.855 4980.720 ;
        RECT 840.025 4980.550 840.315 4980.720 ;
        RECT 840.485 4980.550 840.775 4980.720 ;
        RECT 840.945 4980.550 841.235 4980.720 ;
        RECT 841.405 4980.550 841.695 4980.720 ;
        RECT 841.865 4980.550 842.155 4980.720 ;
        RECT 842.325 4980.550 842.615 4980.720 ;
        RECT 842.785 4980.550 843.075 4980.720 ;
        RECT 843.245 4980.550 843.535 4980.720 ;
        RECT 843.705 4980.550 843.995 4980.720 ;
        RECT 844.165 4980.550 844.455 4980.720 ;
        RECT 844.625 4980.550 844.915 4980.720 ;
        RECT 845.085 4980.550 845.375 4980.720 ;
        RECT 845.545 4980.550 845.835 4980.720 ;
        RECT 846.005 4980.550 846.295 4980.720 ;
        RECT 846.465 4980.550 846.755 4980.720 ;
        RECT 846.925 4980.550 847.215 4980.720 ;
        RECT 847.385 4980.550 847.675 4980.720 ;
        RECT 847.845 4980.550 848.135 4980.720 ;
        RECT 848.305 4980.550 848.595 4980.720 ;
        RECT 848.765 4980.550 849.055 4980.720 ;
        RECT 849.225 4980.550 849.515 4980.720 ;
        RECT 849.685 4980.550 849.975 4980.720 ;
        RECT 850.145 4980.550 850.435 4980.720 ;
        RECT 850.605 4980.550 850.895 4980.720 ;
        RECT 851.065 4980.550 851.355 4980.720 ;
        RECT 851.525 4980.550 851.815 4980.720 ;
        RECT 851.985 4980.550 852.275 4980.720 ;
        RECT 852.445 4980.550 852.735 4980.720 ;
        RECT 852.905 4980.550 853.050 4980.720 ;
        RECT 198.560 4457.115 198.730 4457.200 ;
        RECT 201.280 4457.115 201.450 4457.200 ;
        RECT 204.000 4457.115 204.170 4457.200 ;
        RECT 198.560 4457.055 199.455 4457.115 ;
        RECT 198.730 4456.885 199.455 4457.055 ;
        RECT 198.560 4456.825 199.455 4456.885 ;
        RECT 200.115 4457.055 202.615 4457.115 ;
        RECT 200.115 4456.885 201.280 4457.055 ;
        RECT 201.450 4456.885 202.615 4457.055 ;
        RECT 200.115 4456.825 202.615 4456.885 ;
        RECT 198.560 4456.595 198.730 4456.825 ;
        RECT 201.280 4456.595 201.450 4456.825 ;
        RECT 198.560 4456.265 198.730 4456.425 ;
        RECT 201.280 4456.265 201.450 4456.425 ;
        RECT 201.620 4456.315 202.640 4456.645 ;
        RECT 198.560 4456.135 199.530 4456.265 ;
        RECT 198.730 4455.965 199.530 4456.135 ;
        RECT 198.560 4455.935 199.530 4455.965 ;
        RECT 200.130 4456.145 201.450 4456.265 ;
        RECT 200.130 4456.135 202.250 4456.145 ;
        RECT 200.130 4455.965 201.280 4456.135 ;
        RECT 201.450 4455.975 202.250 4456.135 ;
        RECT 200.130 4455.935 201.450 4455.965 ;
        RECT 198.560 4455.675 198.730 4455.935 ;
      LAYER li1 ;
        RECT 198.900 4455.595 201.110 4455.765 ;
      LAYER li1 ;
        RECT 201.280 4455.675 201.450 4455.935 ;
        RECT 202.470 4455.805 202.640 4456.315 ;
      LAYER li1 ;
        RECT 199.380 4455.510 200.260 4455.595 ;
      LAYER li1 ;
        RECT 198.560 4455.425 198.730 4455.505 ;
        RECT 198.560 4455.215 199.210 4455.425 ;
        RECT 198.730 4455.095 199.210 4455.215 ;
        RECT 198.560 4454.755 198.730 4455.045 ;
      LAYER li1 ;
        RECT 199.380 4454.925 199.550 4455.510 ;
        RECT 198.900 4454.755 199.550 4454.925 ;
      LAYER li1 ;
        RECT 198.560 4454.295 199.210 4454.585 ;
        RECT 198.730 4454.255 199.210 4454.295 ;
        RECT 198.560 4453.835 198.730 4454.125 ;
      LAYER li1 ;
        RECT 199.380 4454.085 199.550 4454.755 ;
        RECT 198.900 4453.915 199.550 4454.085 ;
      LAYER li1 ;
        RECT 198.730 4453.665 199.210 4453.745 ;
        RECT 198.560 4453.415 199.210 4453.665 ;
        RECT 198.560 4453.375 198.730 4453.415 ;
      LAYER li1 ;
        RECT 199.380 4453.245 199.550 4453.915 ;
      LAYER li1 ;
        RECT 198.560 4452.915 198.730 4453.205 ;
      LAYER li1 ;
        RECT 198.900 4453.075 199.550 4453.245 ;
      LAYER li1 ;
        RECT 198.730 4452.745 199.210 4452.905 ;
        RECT 199.720 4452.815 199.890 4455.265 ;
      LAYER li1 ;
        RECT 200.090 4454.925 200.260 4455.510 ;
      LAYER li1 ;
        RECT 201.280 4455.425 201.450 4455.505 ;
        RECT 201.620 4455.475 202.640 4455.805 ;
      LAYER li1 ;
        RECT 202.810 4455.500 203.010 4457.090 ;
      LAYER li1 ;
        RECT 203.275 4457.055 204.170 4457.115 ;
        RECT 203.275 4456.885 204.000 4457.055 ;
        RECT 203.275 4456.825 204.170 4456.885 ;
        RECT 204.000 4456.595 204.170 4456.825 ;
        RECT 203.180 4456.395 203.830 4456.565 ;
        RECT 203.180 4455.725 203.350 4456.395 ;
        RECT 204.000 4456.225 204.170 4456.425 ;
        RECT 203.520 4456.135 204.170 4456.225 ;
        RECT 203.520 4455.965 204.000 4456.135 ;
        RECT 203.520 4455.895 204.170 4455.965 ;
        RECT 203.180 4455.555 203.825 4455.725 ;
        RECT 204.000 4455.675 204.170 4455.895 ;
        RECT 200.480 4455.305 201.450 4455.425 ;
        RECT 202.470 4455.320 202.640 4455.475 ;
        RECT 203.180 4455.320 203.350 4455.555 ;
        RECT 204.000 4455.385 204.170 4455.505 ;
        RECT 200.480 4455.215 202.250 4455.305 ;
        RECT 200.480 4455.095 201.280 4455.215 ;
        RECT 201.450 4455.135 202.250 4455.215 ;
        RECT 202.470 4455.145 203.350 4455.320 ;
        RECT 203.520 4455.215 204.170 4455.385 ;
      LAYER li1 ;
        RECT 200.090 4454.755 201.110 4454.925 ;
      LAYER li1 ;
        RECT 201.280 4454.755 201.450 4455.045 ;
      LAYER li1 ;
        RECT 200.090 4454.085 200.260 4454.755 ;
        RECT 201.620 4454.715 202.640 4454.885 ;
      LAYER li1 ;
        RECT 200.480 4454.545 201.450 4454.585 ;
        RECT 200.480 4454.295 202.250 4454.545 ;
        RECT 200.480 4454.255 201.280 4454.295 ;
        RECT 201.450 4454.215 202.250 4454.295 ;
      LAYER li1 ;
        RECT 200.090 4453.915 201.110 4454.085 ;
        RECT 200.090 4453.245 200.260 4453.915 ;
      LAYER li1 ;
        RECT 201.280 4453.835 201.450 4454.125 ;
      LAYER li1 ;
        RECT 202.470 4454.045 202.640 4454.715 ;
        RECT 201.620 4453.875 202.640 4454.045 ;
      LAYER li1 ;
        RECT 200.480 4453.665 201.280 4453.745 ;
        RECT 201.450 4453.665 202.250 4453.705 ;
        RECT 200.480 4453.415 202.250 4453.665 ;
        RECT 201.280 4453.375 202.250 4453.415 ;
      LAYER li1 ;
        RECT 200.090 4453.075 201.110 4453.245 ;
        RECT 202.470 4453.205 202.640 4453.875 ;
      LAYER li1 ;
        RECT 201.280 4452.915 201.450 4453.205 ;
      LAYER li1 ;
        RECT 201.620 4453.035 202.640 4453.205 ;
      LAYER li1 ;
        RECT 198.560 4452.575 199.210 4452.745 ;
        RECT 199.380 4452.640 200.260 4452.815 ;
        RECT 200.480 4452.745 201.280 4452.825 ;
        RECT 201.450 4452.745 202.250 4452.865 ;
        RECT 200.480 4452.655 202.250 4452.745 ;
        RECT 198.560 4452.455 198.730 4452.575 ;
        RECT 199.380 4452.405 199.550 4452.640 ;
        RECT 200.090 4452.485 200.260 4452.640 ;
        RECT 201.280 4452.535 202.250 4452.655 ;
        RECT 198.560 4452.065 198.730 4452.285 ;
        RECT 198.905 4452.235 199.550 4452.405 ;
        RECT 198.560 4451.995 199.210 4452.065 ;
        RECT 198.730 4451.825 199.210 4451.995 ;
        RECT 198.560 4451.735 199.210 4451.825 ;
        RECT 198.560 4451.535 198.730 4451.735 ;
        RECT 199.380 4451.565 199.550 4452.235 ;
        RECT 198.900 4451.395 199.550 4451.565 ;
        RECT 198.560 4451.135 198.730 4451.365 ;
      LAYER li1 ;
        RECT 199.720 4451.360 199.920 4452.460 ;
      LAYER li1 ;
        RECT 200.090 4452.155 201.110 4452.485 ;
        RECT 201.280 4452.455 201.450 4452.535 ;
      LAYER li1 ;
        RECT 202.470 4452.450 202.640 4453.035 ;
      LAYER li1 ;
        RECT 202.840 4452.695 203.010 4455.145 ;
        RECT 203.520 4455.055 204.000 4455.215 ;
      LAYER li1 ;
        RECT 203.180 4454.715 203.830 4454.885 ;
      LAYER li1 ;
        RECT 204.000 4454.755 204.170 4455.045 ;
      LAYER li1 ;
        RECT 203.180 4454.045 203.350 4454.715 ;
      LAYER li1 ;
        RECT 204.000 4454.545 204.170 4454.585 ;
        RECT 203.520 4454.295 204.170 4454.545 ;
        RECT 203.520 4454.215 204.000 4454.295 ;
      LAYER li1 ;
        RECT 203.180 4453.875 203.830 4454.045 ;
        RECT 203.180 4453.205 203.350 4453.875 ;
      LAYER li1 ;
        RECT 204.000 4453.835 204.170 4454.125 ;
        RECT 203.520 4453.665 204.000 4453.705 ;
        RECT 203.520 4453.375 204.170 4453.665 ;
      LAYER li1 ;
        RECT 203.180 4453.035 203.830 4453.205 ;
        RECT 203.180 4452.450 203.350 4453.035 ;
      LAYER li1 ;
        RECT 204.000 4452.915 204.170 4453.205 ;
        RECT 203.520 4452.745 204.000 4452.865 ;
        RECT 203.520 4452.535 204.170 4452.745 ;
        RECT 204.000 4452.455 204.170 4452.535 ;
      LAYER li1 ;
        RECT 202.470 4452.365 203.350 4452.450 ;
      LAYER li1 ;
        RECT 200.090 4451.645 200.260 4452.155 ;
        RECT 201.280 4452.025 201.450 4452.285 ;
      LAYER li1 ;
        RECT 201.620 4452.195 203.830 4452.365 ;
      LAYER li1 ;
        RECT 204.000 4452.025 204.170 4452.285 ;
        RECT 201.280 4451.995 202.600 4452.025 ;
        RECT 200.480 4451.825 201.280 4451.985 ;
        RECT 201.450 4451.825 202.600 4451.995 ;
        RECT 200.480 4451.815 202.600 4451.825 ;
        RECT 201.280 4451.695 202.600 4451.815 ;
        RECT 203.200 4451.995 204.170 4452.025 ;
        RECT 203.200 4451.825 204.000 4451.995 ;
        RECT 203.200 4451.695 204.170 4451.825 ;
        RECT 200.090 4451.315 201.110 4451.645 ;
        RECT 201.280 4451.535 201.450 4451.695 ;
        RECT 204.000 4451.535 204.170 4451.695 ;
        RECT 201.280 4451.135 201.450 4451.365 ;
        RECT 204.000 4451.135 204.170 4451.365 ;
        RECT 198.560 4451.075 199.455 4451.135 ;
        RECT 198.730 4450.905 199.455 4451.075 ;
        RECT 198.560 4450.845 199.455 4450.905 ;
        RECT 200.115 4451.075 202.615 4451.135 ;
        RECT 200.115 4450.905 201.280 4451.075 ;
        RECT 201.450 4450.905 202.615 4451.075 ;
        RECT 200.115 4450.845 202.615 4450.905 ;
        RECT 198.560 4450.615 198.730 4450.845 ;
        RECT 201.280 4450.615 201.450 4450.845 ;
        RECT 198.560 4450.285 198.730 4450.445 ;
        RECT 201.280 4450.285 201.450 4450.445 ;
        RECT 201.620 4450.335 202.640 4450.665 ;
        RECT 198.560 4450.155 199.530 4450.285 ;
        RECT 198.730 4449.985 199.530 4450.155 ;
        RECT 198.560 4449.955 199.530 4449.985 ;
        RECT 200.130 4450.165 201.450 4450.285 ;
        RECT 200.130 4450.155 202.250 4450.165 ;
        RECT 200.130 4449.985 201.280 4450.155 ;
        RECT 201.450 4449.995 202.250 4450.155 ;
        RECT 200.130 4449.955 201.450 4449.985 ;
        RECT 198.560 4449.695 198.730 4449.955 ;
      LAYER li1 ;
        RECT 198.900 4449.615 201.110 4449.785 ;
      LAYER li1 ;
        RECT 201.280 4449.695 201.450 4449.955 ;
        RECT 202.470 4449.825 202.640 4450.335 ;
      LAYER li1 ;
        RECT 199.380 4449.530 200.260 4449.615 ;
      LAYER li1 ;
        RECT 198.560 4449.445 198.730 4449.525 ;
        RECT 198.560 4449.235 199.210 4449.445 ;
        RECT 198.730 4449.115 199.210 4449.235 ;
        RECT 198.560 4448.775 198.730 4449.065 ;
      LAYER li1 ;
        RECT 199.380 4448.945 199.550 4449.530 ;
        RECT 198.900 4448.775 199.550 4448.945 ;
      LAYER li1 ;
        RECT 198.560 4448.315 199.210 4448.605 ;
        RECT 198.730 4448.275 199.210 4448.315 ;
        RECT 198.560 4447.855 198.730 4448.145 ;
      LAYER li1 ;
        RECT 199.380 4448.105 199.550 4448.775 ;
        RECT 198.900 4447.935 199.550 4448.105 ;
      LAYER li1 ;
        RECT 198.730 4447.685 199.210 4447.765 ;
        RECT 198.560 4447.435 199.210 4447.685 ;
        RECT 198.560 4447.395 198.730 4447.435 ;
      LAYER li1 ;
        RECT 199.380 4447.265 199.550 4447.935 ;
      LAYER li1 ;
        RECT 198.560 4446.935 198.730 4447.225 ;
      LAYER li1 ;
        RECT 198.900 4447.095 199.550 4447.265 ;
      LAYER li1 ;
        RECT 198.730 4446.765 199.210 4446.925 ;
        RECT 199.720 4446.835 199.890 4449.285 ;
      LAYER li1 ;
        RECT 200.090 4448.945 200.260 4449.530 ;
      LAYER li1 ;
        RECT 201.280 4449.445 201.450 4449.525 ;
        RECT 201.620 4449.495 202.640 4449.825 ;
      LAYER li1 ;
        RECT 202.810 4449.520 203.010 4451.110 ;
      LAYER li1 ;
        RECT 203.275 4451.075 204.170 4451.135 ;
        RECT 203.275 4450.905 204.000 4451.075 ;
        RECT 203.275 4450.845 204.170 4450.905 ;
        RECT 204.000 4450.615 204.170 4450.845 ;
        RECT 203.180 4450.415 203.830 4450.585 ;
        RECT 203.180 4449.745 203.350 4450.415 ;
        RECT 204.000 4450.245 204.170 4450.445 ;
        RECT 203.520 4450.155 204.170 4450.245 ;
        RECT 203.520 4449.985 204.000 4450.155 ;
        RECT 203.520 4449.915 204.170 4449.985 ;
        RECT 203.180 4449.575 203.825 4449.745 ;
        RECT 204.000 4449.695 204.170 4449.915 ;
        RECT 200.480 4449.325 201.450 4449.445 ;
        RECT 202.470 4449.340 202.640 4449.495 ;
        RECT 203.180 4449.340 203.350 4449.575 ;
        RECT 204.000 4449.405 204.170 4449.525 ;
        RECT 200.480 4449.235 202.250 4449.325 ;
        RECT 200.480 4449.115 201.280 4449.235 ;
        RECT 201.450 4449.155 202.250 4449.235 ;
        RECT 202.470 4449.165 203.350 4449.340 ;
        RECT 203.520 4449.235 204.170 4449.405 ;
      LAYER li1 ;
        RECT 200.090 4448.775 201.110 4448.945 ;
      LAYER li1 ;
        RECT 201.280 4448.775 201.450 4449.065 ;
      LAYER li1 ;
        RECT 200.090 4448.105 200.260 4448.775 ;
        RECT 201.620 4448.735 202.640 4448.905 ;
      LAYER li1 ;
        RECT 200.480 4448.565 201.450 4448.605 ;
        RECT 200.480 4448.315 202.250 4448.565 ;
        RECT 200.480 4448.275 201.280 4448.315 ;
        RECT 201.450 4448.235 202.250 4448.315 ;
      LAYER li1 ;
        RECT 200.090 4447.935 201.110 4448.105 ;
        RECT 200.090 4447.265 200.260 4447.935 ;
      LAYER li1 ;
        RECT 201.280 4447.855 201.450 4448.145 ;
      LAYER li1 ;
        RECT 202.470 4448.065 202.640 4448.735 ;
        RECT 201.620 4447.895 202.640 4448.065 ;
      LAYER li1 ;
        RECT 200.480 4447.685 201.280 4447.765 ;
        RECT 201.450 4447.685 202.250 4447.725 ;
        RECT 200.480 4447.435 202.250 4447.685 ;
        RECT 201.280 4447.395 202.250 4447.435 ;
      LAYER li1 ;
        RECT 200.090 4447.095 201.110 4447.265 ;
        RECT 202.470 4447.225 202.640 4447.895 ;
      LAYER li1 ;
        RECT 201.280 4446.935 201.450 4447.225 ;
      LAYER li1 ;
        RECT 201.620 4447.055 202.640 4447.225 ;
      LAYER li1 ;
        RECT 198.560 4446.595 199.210 4446.765 ;
        RECT 199.380 4446.660 200.260 4446.835 ;
        RECT 200.480 4446.765 201.280 4446.845 ;
        RECT 201.450 4446.765 202.250 4446.885 ;
        RECT 200.480 4446.675 202.250 4446.765 ;
        RECT 198.560 4446.475 198.730 4446.595 ;
        RECT 199.380 4446.425 199.550 4446.660 ;
        RECT 200.090 4446.505 200.260 4446.660 ;
        RECT 201.280 4446.555 202.250 4446.675 ;
        RECT 198.560 4446.085 198.730 4446.305 ;
        RECT 198.905 4446.255 199.550 4446.425 ;
        RECT 198.560 4446.015 199.210 4446.085 ;
        RECT 198.730 4445.845 199.210 4446.015 ;
        RECT 198.560 4445.755 199.210 4445.845 ;
        RECT 198.560 4445.555 198.730 4445.755 ;
        RECT 199.380 4445.585 199.550 4446.255 ;
        RECT 198.900 4445.415 199.550 4445.585 ;
        RECT 198.560 4445.155 198.730 4445.385 ;
      LAYER li1 ;
        RECT 199.720 4445.380 199.920 4446.480 ;
      LAYER li1 ;
        RECT 200.090 4446.175 201.110 4446.505 ;
        RECT 201.280 4446.475 201.450 4446.555 ;
      LAYER li1 ;
        RECT 202.470 4446.470 202.640 4447.055 ;
      LAYER li1 ;
        RECT 202.840 4446.715 203.010 4449.165 ;
        RECT 203.520 4449.075 204.000 4449.235 ;
      LAYER li1 ;
        RECT 203.180 4448.735 203.830 4448.905 ;
      LAYER li1 ;
        RECT 204.000 4448.775 204.170 4449.065 ;
      LAYER li1 ;
        RECT 203.180 4448.065 203.350 4448.735 ;
      LAYER li1 ;
        RECT 204.000 4448.565 204.170 4448.605 ;
        RECT 203.520 4448.315 204.170 4448.565 ;
        RECT 203.520 4448.235 204.000 4448.315 ;
      LAYER li1 ;
        RECT 203.180 4447.895 203.830 4448.065 ;
        RECT 203.180 4447.225 203.350 4447.895 ;
      LAYER li1 ;
        RECT 204.000 4447.855 204.170 4448.145 ;
        RECT 203.520 4447.685 204.000 4447.725 ;
        RECT 203.520 4447.395 204.170 4447.685 ;
      LAYER li1 ;
        RECT 203.180 4447.055 203.830 4447.225 ;
        RECT 203.180 4446.470 203.350 4447.055 ;
      LAYER li1 ;
        RECT 204.000 4446.935 204.170 4447.225 ;
        RECT 203.520 4446.765 204.000 4446.885 ;
        RECT 203.520 4446.555 204.170 4446.765 ;
        RECT 204.000 4446.475 204.170 4446.555 ;
      LAYER li1 ;
        RECT 202.470 4446.385 203.350 4446.470 ;
      LAYER li1 ;
        RECT 200.090 4445.665 200.260 4446.175 ;
        RECT 201.280 4446.045 201.450 4446.305 ;
      LAYER li1 ;
        RECT 201.620 4446.215 203.830 4446.385 ;
      LAYER li1 ;
        RECT 204.000 4446.045 204.170 4446.305 ;
        RECT 201.280 4446.015 202.600 4446.045 ;
        RECT 200.480 4445.845 201.280 4446.005 ;
        RECT 201.450 4445.845 202.600 4446.015 ;
        RECT 200.480 4445.835 202.600 4445.845 ;
        RECT 201.280 4445.715 202.600 4445.835 ;
        RECT 203.200 4446.015 204.170 4446.045 ;
        RECT 203.200 4445.845 204.000 4446.015 ;
        RECT 203.200 4445.715 204.170 4445.845 ;
        RECT 200.090 4445.335 201.110 4445.665 ;
        RECT 201.280 4445.555 201.450 4445.715 ;
        RECT 204.000 4445.555 204.170 4445.715 ;
        RECT 201.280 4445.155 201.450 4445.385 ;
        RECT 204.000 4445.155 204.170 4445.385 ;
        RECT 198.560 4445.095 199.455 4445.155 ;
        RECT 198.730 4444.925 199.455 4445.095 ;
        RECT 198.560 4444.865 199.455 4444.925 ;
        RECT 200.115 4445.095 202.615 4445.155 ;
        RECT 200.115 4444.925 201.280 4445.095 ;
        RECT 201.450 4444.925 202.615 4445.095 ;
        RECT 200.115 4444.865 202.615 4444.925 ;
        RECT 198.560 4444.635 198.730 4444.865 ;
        RECT 201.280 4444.635 201.450 4444.865 ;
        RECT 198.560 4444.305 198.730 4444.465 ;
        RECT 201.280 4444.305 201.450 4444.465 ;
        RECT 201.620 4444.355 202.640 4444.685 ;
        RECT 198.560 4444.175 199.530 4444.305 ;
        RECT 198.730 4444.005 199.530 4444.175 ;
        RECT 198.560 4443.975 199.530 4444.005 ;
        RECT 200.130 4444.185 201.450 4444.305 ;
        RECT 200.130 4444.175 202.250 4444.185 ;
        RECT 200.130 4444.005 201.280 4444.175 ;
        RECT 201.450 4444.015 202.250 4444.175 ;
        RECT 200.130 4443.975 201.450 4444.005 ;
        RECT 198.560 4443.715 198.730 4443.975 ;
      LAYER li1 ;
        RECT 198.900 4443.635 201.110 4443.805 ;
      LAYER li1 ;
        RECT 201.280 4443.715 201.450 4443.975 ;
        RECT 202.470 4443.845 202.640 4444.355 ;
      LAYER li1 ;
        RECT 199.380 4443.550 200.260 4443.635 ;
      LAYER li1 ;
        RECT 198.560 4443.465 198.730 4443.545 ;
        RECT 198.560 4443.255 199.210 4443.465 ;
        RECT 198.730 4443.135 199.210 4443.255 ;
        RECT 198.560 4442.795 198.730 4443.085 ;
      LAYER li1 ;
        RECT 199.380 4442.965 199.550 4443.550 ;
        RECT 198.900 4442.795 199.550 4442.965 ;
      LAYER li1 ;
        RECT 198.560 4442.335 199.210 4442.625 ;
        RECT 198.730 4442.295 199.210 4442.335 ;
        RECT 198.560 4441.875 198.730 4442.165 ;
      LAYER li1 ;
        RECT 199.380 4442.125 199.550 4442.795 ;
        RECT 198.900 4441.955 199.550 4442.125 ;
      LAYER li1 ;
        RECT 198.730 4441.705 199.210 4441.785 ;
        RECT 198.560 4441.455 199.210 4441.705 ;
        RECT 198.560 4441.415 198.730 4441.455 ;
      LAYER li1 ;
        RECT 199.380 4441.285 199.550 4441.955 ;
      LAYER li1 ;
        RECT 198.560 4440.955 198.730 4441.245 ;
      LAYER li1 ;
        RECT 198.900 4441.115 199.550 4441.285 ;
      LAYER li1 ;
        RECT 198.730 4440.785 199.210 4440.945 ;
        RECT 199.720 4440.855 199.890 4443.305 ;
      LAYER li1 ;
        RECT 200.090 4442.965 200.260 4443.550 ;
      LAYER li1 ;
        RECT 201.280 4443.465 201.450 4443.545 ;
        RECT 201.620 4443.515 202.640 4443.845 ;
      LAYER li1 ;
        RECT 202.810 4443.540 203.010 4445.130 ;
      LAYER li1 ;
        RECT 203.275 4445.095 204.170 4445.155 ;
        RECT 203.275 4444.925 204.000 4445.095 ;
        RECT 203.275 4444.865 204.170 4444.925 ;
        RECT 204.000 4444.635 204.170 4444.865 ;
        RECT 203.180 4444.435 203.830 4444.605 ;
        RECT 203.180 4443.765 203.350 4444.435 ;
        RECT 204.000 4444.265 204.170 4444.465 ;
        RECT 203.520 4444.175 204.170 4444.265 ;
        RECT 203.520 4444.005 204.000 4444.175 ;
        RECT 203.520 4443.935 204.170 4444.005 ;
        RECT 203.180 4443.595 203.825 4443.765 ;
        RECT 204.000 4443.715 204.170 4443.935 ;
        RECT 200.480 4443.345 201.450 4443.465 ;
        RECT 202.470 4443.360 202.640 4443.515 ;
        RECT 203.180 4443.360 203.350 4443.595 ;
        RECT 204.000 4443.425 204.170 4443.545 ;
        RECT 200.480 4443.255 202.250 4443.345 ;
        RECT 200.480 4443.135 201.280 4443.255 ;
        RECT 201.450 4443.175 202.250 4443.255 ;
        RECT 202.470 4443.185 203.350 4443.360 ;
        RECT 203.520 4443.255 204.170 4443.425 ;
      LAYER li1 ;
        RECT 200.090 4442.795 201.110 4442.965 ;
      LAYER li1 ;
        RECT 201.280 4442.795 201.450 4443.085 ;
      LAYER li1 ;
        RECT 200.090 4442.125 200.260 4442.795 ;
        RECT 201.620 4442.755 202.640 4442.925 ;
      LAYER li1 ;
        RECT 200.480 4442.585 201.450 4442.625 ;
        RECT 200.480 4442.335 202.250 4442.585 ;
        RECT 200.480 4442.295 201.280 4442.335 ;
        RECT 201.450 4442.255 202.250 4442.335 ;
      LAYER li1 ;
        RECT 200.090 4441.955 201.110 4442.125 ;
        RECT 200.090 4441.285 200.260 4441.955 ;
      LAYER li1 ;
        RECT 201.280 4441.875 201.450 4442.165 ;
      LAYER li1 ;
        RECT 202.470 4442.085 202.640 4442.755 ;
        RECT 201.620 4441.915 202.640 4442.085 ;
      LAYER li1 ;
        RECT 200.480 4441.705 201.280 4441.785 ;
        RECT 201.450 4441.705 202.250 4441.745 ;
        RECT 200.480 4441.455 202.250 4441.705 ;
        RECT 201.280 4441.415 202.250 4441.455 ;
      LAYER li1 ;
        RECT 200.090 4441.115 201.110 4441.285 ;
        RECT 202.470 4441.245 202.640 4441.915 ;
      LAYER li1 ;
        RECT 201.280 4440.955 201.450 4441.245 ;
      LAYER li1 ;
        RECT 201.620 4441.075 202.640 4441.245 ;
      LAYER li1 ;
        RECT 198.560 4440.615 199.210 4440.785 ;
        RECT 199.380 4440.680 200.260 4440.855 ;
        RECT 200.480 4440.785 201.280 4440.865 ;
        RECT 201.450 4440.785 202.250 4440.905 ;
        RECT 200.480 4440.695 202.250 4440.785 ;
        RECT 198.560 4440.495 198.730 4440.615 ;
        RECT 199.380 4440.445 199.550 4440.680 ;
        RECT 200.090 4440.525 200.260 4440.680 ;
        RECT 201.280 4440.575 202.250 4440.695 ;
        RECT 198.560 4440.105 198.730 4440.325 ;
        RECT 198.905 4440.275 199.550 4440.445 ;
        RECT 198.560 4440.035 199.210 4440.105 ;
        RECT 198.730 4439.865 199.210 4440.035 ;
        RECT 198.560 4439.775 199.210 4439.865 ;
        RECT 198.560 4439.575 198.730 4439.775 ;
        RECT 199.380 4439.605 199.550 4440.275 ;
        RECT 198.900 4439.435 199.550 4439.605 ;
        RECT 198.560 4439.175 198.730 4439.405 ;
      LAYER li1 ;
        RECT 199.720 4439.400 199.920 4440.500 ;
      LAYER li1 ;
        RECT 200.090 4440.195 201.110 4440.525 ;
        RECT 201.280 4440.495 201.450 4440.575 ;
      LAYER li1 ;
        RECT 202.470 4440.490 202.640 4441.075 ;
      LAYER li1 ;
        RECT 202.840 4440.735 203.010 4443.185 ;
        RECT 203.520 4443.095 204.000 4443.255 ;
      LAYER li1 ;
        RECT 203.180 4442.755 203.830 4442.925 ;
      LAYER li1 ;
        RECT 204.000 4442.795 204.170 4443.085 ;
      LAYER li1 ;
        RECT 203.180 4442.085 203.350 4442.755 ;
      LAYER li1 ;
        RECT 204.000 4442.585 204.170 4442.625 ;
        RECT 203.520 4442.335 204.170 4442.585 ;
        RECT 203.520 4442.255 204.000 4442.335 ;
      LAYER li1 ;
        RECT 203.180 4441.915 203.830 4442.085 ;
        RECT 203.180 4441.245 203.350 4441.915 ;
      LAYER li1 ;
        RECT 204.000 4441.875 204.170 4442.165 ;
        RECT 203.520 4441.705 204.000 4441.745 ;
        RECT 203.520 4441.415 204.170 4441.705 ;
      LAYER li1 ;
        RECT 203.180 4441.075 203.830 4441.245 ;
        RECT 203.180 4440.490 203.350 4441.075 ;
      LAYER li1 ;
        RECT 204.000 4440.955 204.170 4441.245 ;
        RECT 203.520 4440.785 204.000 4440.905 ;
        RECT 203.520 4440.575 204.170 4440.785 ;
        RECT 204.000 4440.495 204.170 4440.575 ;
      LAYER li1 ;
        RECT 202.470 4440.405 203.350 4440.490 ;
      LAYER li1 ;
        RECT 200.090 4439.685 200.260 4440.195 ;
        RECT 201.280 4440.065 201.450 4440.325 ;
      LAYER li1 ;
        RECT 201.620 4440.235 203.830 4440.405 ;
      LAYER li1 ;
        RECT 204.000 4440.065 204.170 4440.325 ;
        RECT 201.280 4440.035 202.600 4440.065 ;
        RECT 200.480 4439.865 201.280 4440.025 ;
        RECT 201.450 4439.865 202.600 4440.035 ;
        RECT 200.480 4439.855 202.600 4439.865 ;
        RECT 201.280 4439.735 202.600 4439.855 ;
        RECT 203.200 4440.035 204.170 4440.065 ;
        RECT 203.200 4439.865 204.000 4440.035 ;
        RECT 203.200 4439.735 204.170 4439.865 ;
        RECT 200.090 4439.355 201.110 4439.685 ;
        RECT 201.280 4439.575 201.450 4439.735 ;
        RECT 204.000 4439.575 204.170 4439.735 ;
        RECT 201.280 4439.175 201.450 4439.405 ;
        RECT 204.000 4439.175 204.170 4439.405 ;
        RECT 198.560 4439.115 199.455 4439.175 ;
        RECT 198.730 4438.945 199.455 4439.115 ;
        RECT 198.560 4438.885 199.455 4438.945 ;
        RECT 200.115 4439.115 202.615 4439.175 ;
        RECT 200.115 4438.945 201.280 4439.115 ;
        RECT 201.450 4438.945 202.615 4439.115 ;
        RECT 200.115 4438.885 202.615 4438.945 ;
        RECT 203.275 4439.115 204.170 4439.175 ;
        RECT 203.275 4438.945 204.000 4439.115 ;
        RECT 203.275 4438.885 204.170 4438.945 ;
        RECT 198.560 4438.655 198.730 4438.885 ;
        RECT 201.280 4438.655 201.450 4438.885 ;
        RECT 198.560 4438.325 198.730 4438.485 ;
        RECT 201.280 4438.325 201.450 4438.485 ;
        RECT 201.620 4438.375 202.640 4438.705 ;
        RECT 204.000 4438.655 204.170 4438.885 ;
        RECT 198.560 4438.195 199.530 4438.325 ;
        RECT 198.730 4438.025 199.530 4438.195 ;
        RECT 198.560 4437.995 199.530 4438.025 ;
        RECT 200.130 4438.205 201.450 4438.325 ;
        RECT 200.130 4438.195 202.250 4438.205 ;
        RECT 200.130 4438.025 201.280 4438.195 ;
        RECT 201.450 4438.035 202.250 4438.195 ;
        RECT 200.130 4437.995 201.450 4438.025 ;
        RECT 198.560 4437.735 198.730 4437.995 ;
        RECT 201.280 4437.735 201.450 4437.995 ;
        RECT 202.470 4437.865 202.640 4438.375 ;
        RECT 198.560 4437.485 198.730 4437.565 ;
        RECT 201.280 4437.485 201.450 4437.565 ;
        RECT 201.620 4437.535 202.640 4437.865 ;
        RECT 198.560 4437.275 199.210 4437.485 ;
        RECT 200.480 4437.365 201.450 4437.485 ;
        RECT 202.470 4437.380 202.640 4437.535 ;
        RECT 203.180 4438.455 203.830 4438.625 ;
        RECT 203.180 4437.785 203.350 4438.455 ;
        RECT 204.000 4438.285 204.170 4438.485 ;
        RECT 203.520 4438.195 204.170 4438.285 ;
        RECT 203.520 4438.025 204.000 4438.195 ;
        RECT 203.520 4437.955 204.170 4438.025 ;
        RECT 203.180 4437.615 203.825 4437.785 ;
        RECT 204.000 4437.735 204.170 4437.955 ;
        RECT 203.180 4437.380 203.350 4437.615 ;
        RECT 204.000 4437.445 204.170 4437.565 ;
        RECT 198.730 4437.155 199.210 4437.275 ;
        RECT 198.560 4436.815 198.730 4437.105 ;
        RECT 198.560 4436.355 199.210 4436.645 ;
        RECT 198.730 4436.315 199.210 4436.355 ;
        RECT 198.560 4435.895 198.730 4436.185 ;
        RECT 198.730 4435.725 199.210 4435.805 ;
        RECT 198.560 4435.475 199.210 4435.725 ;
        RECT 198.560 4435.435 198.730 4435.475 ;
        RECT 198.560 4434.975 198.730 4435.265 ;
        RECT 198.730 4434.805 199.210 4434.965 ;
        RECT 199.720 4434.875 199.890 4437.325 ;
        RECT 200.480 4437.275 202.250 4437.365 ;
        RECT 200.480 4437.155 201.280 4437.275 ;
        RECT 201.450 4437.195 202.250 4437.275 ;
        RECT 202.470 4437.205 203.350 4437.380 ;
        RECT 203.520 4437.275 204.170 4437.445 ;
        RECT 201.280 4436.815 201.450 4437.105 ;
      LAYER li1 ;
        RECT 201.620 4436.775 202.640 4436.945 ;
      LAYER li1 ;
        RECT 200.480 4436.605 201.450 4436.645 ;
        RECT 200.480 4436.355 202.250 4436.605 ;
        RECT 200.480 4436.315 201.280 4436.355 ;
        RECT 201.450 4436.275 202.250 4436.355 ;
        RECT 201.280 4435.895 201.450 4436.185 ;
      LAYER li1 ;
        RECT 202.470 4436.105 202.640 4436.775 ;
        RECT 201.620 4435.935 202.640 4436.105 ;
      LAYER li1 ;
        RECT 200.480 4435.725 201.280 4435.805 ;
        RECT 201.450 4435.725 202.250 4435.765 ;
        RECT 200.480 4435.475 202.250 4435.725 ;
        RECT 201.280 4435.435 202.250 4435.475 ;
      LAYER li1 ;
        RECT 202.470 4435.265 202.640 4435.935 ;
      LAYER li1 ;
        RECT 201.280 4434.975 201.450 4435.265 ;
      LAYER li1 ;
        RECT 201.620 4435.095 202.640 4435.265 ;
      LAYER li1 ;
        RECT 198.560 4434.635 199.210 4434.805 ;
        RECT 199.380 4434.700 200.260 4434.875 ;
        RECT 200.480 4434.805 201.280 4434.885 ;
        RECT 201.450 4434.805 202.250 4434.925 ;
        RECT 200.480 4434.715 202.250 4434.805 ;
        RECT 198.560 4434.515 198.730 4434.635 ;
        RECT 199.380 4434.465 199.550 4434.700 ;
        RECT 200.090 4434.545 200.260 4434.700 ;
        RECT 201.280 4434.595 202.250 4434.715 ;
        RECT 198.560 4434.125 198.730 4434.345 ;
        RECT 198.905 4434.295 199.550 4434.465 ;
        RECT 198.560 4434.055 199.210 4434.125 ;
        RECT 198.730 4433.885 199.210 4434.055 ;
        RECT 198.560 4433.795 199.210 4433.885 ;
        RECT 198.560 4433.595 198.730 4433.795 ;
        RECT 199.380 4433.625 199.550 4434.295 ;
        RECT 198.900 4433.455 199.550 4433.625 ;
        RECT 198.560 4433.195 198.730 4433.425 ;
      LAYER li1 ;
        RECT 199.720 4433.420 199.920 4434.520 ;
      LAYER li1 ;
        RECT 200.090 4434.215 201.110 4434.545 ;
        RECT 201.280 4434.515 201.450 4434.595 ;
      LAYER li1 ;
        RECT 202.470 4434.510 202.640 4435.095 ;
      LAYER li1 ;
        RECT 202.840 4434.755 203.010 4437.205 ;
        RECT 203.520 4437.115 204.000 4437.275 ;
      LAYER li1 ;
        RECT 203.180 4436.775 203.830 4436.945 ;
      LAYER li1 ;
        RECT 204.000 4436.815 204.170 4437.105 ;
      LAYER li1 ;
        RECT 203.180 4436.105 203.350 4436.775 ;
      LAYER li1 ;
        RECT 204.000 4436.605 204.170 4436.645 ;
        RECT 203.520 4436.355 204.170 4436.605 ;
        RECT 203.520 4436.275 204.000 4436.355 ;
      LAYER li1 ;
        RECT 203.180 4435.935 203.830 4436.105 ;
        RECT 203.180 4435.265 203.350 4435.935 ;
      LAYER li1 ;
        RECT 204.000 4435.895 204.170 4436.185 ;
        RECT 203.520 4435.725 204.000 4435.765 ;
        RECT 203.520 4435.435 204.170 4435.725 ;
      LAYER li1 ;
        RECT 203.180 4435.095 203.830 4435.265 ;
        RECT 203.180 4434.510 203.350 4435.095 ;
      LAYER li1 ;
        RECT 204.000 4434.975 204.170 4435.265 ;
        RECT 203.520 4434.805 204.000 4434.925 ;
        RECT 203.520 4434.595 204.170 4434.805 ;
        RECT 204.000 4434.515 204.170 4434.595 ;
      LAYER li1 ;
        RECT 202.470 4434.425 203.350 4434.510 ;
      LAYER li1 ;
        RECT 200.090 4433.705 200.260 4434.215 ;
        RECT 201.280 4434.085 201.450 4434.345 ;
      LAYER li1 ;
        RECT 201.620 4434.255 203.830 4434.425 ;
      LAYER li1 ;
        RECT 204.000 4434.085 204.170 4434.345 ;
        RECT 201.280 4434.055 202.600 4434.085 ;
        RECT 200.480 4433.885 201.280 4434.045 ;
        RECT 201.450 4433.885 202.600 4434.055 ;
        RECT 200.480 4433.875 202.600 4433.885 ;
        RECT 201.280 4433.755 202.600 4433.875 ;
        RECT 203.200 4434.055 204.170 4434.085 ;
        RECT 203.200 4433.885 204.000 4434.055 ;
        RECT 203.200 4433.755 204.170 4433.885 ;
        RECT 200.090 4433.375 201.110 4433.705 ;
        RECT 201.280 4433.595 201.450 4433.755 ;
        RECT 204.000 4433.595 204.170 4433.755 ;
        RECT 201.280 4433.195 201.450 4433.425 ;
        RECT 204.000 4433.195 204.170 4433.425 ;
        RECT 198.560 4433.135 199.455 4433.195 ;
        RECT 198.730 4432.965 199.455 4433.135 ;
        RECT 198.560 4432.905 199.455 4432.965 ;
        RECT 200.115 4433.135 202.615 4433.195 ;
        RECT 200.115 4432.965 201.280 4433.135 ;
        RECT 201.450 4432.965 202.615 4433.135 ;
        RECT 200.115 4432.905 202.615 4432.965 ;
        RECT 203.275 4433.135 204.170 4433.195 ;
        RECT 203.275 4432.965 204.000 4433.135 ;
        RECT 203.275 4432.905 204.170 4432.965 ;
        RECT 198.560 4432.675 198.730 4432.905 ;
        RECT 201.280 4432.675 201.450 4432.905 ;
        RECT 198.560 4432.345 198.730 4432.505 ;
        RECT 201.280 4432.345 201.450 4432.505 ;
        RECT 201.620 4432.395 202.640 4432.725 ;
        RECT 204.000 4432.675 204.170 4432.905 ;
        RECT 198.560 4432.215 199.530 4432.345 ;
        RECT 198.730 4432.045 199.530 4432.215 ;
        RECT 198.560 4432.015 199.530 4432.045 ;
        RECT 200.130 4432.225 201.450 4432.345 ;
        RECT 200.130 4432.215 202.250 4432.225 ;
        RECT 200.130 4432.045 201.280 4432.215 ;
        RECT 201.450 4432.055 202.250 4432.215 ;
        RECT 200.130 4432.015 201.450 4432.045 ;
        RECT 198.560 4431.755 198.730 4432.015 ;
        RECT 201.280 4431.755 201.450 4432.015 ;
        RECT 202.470 4431.885 202.640 4432.395 ;
        RECT 198.560 4431.505 198.730 4431.585 ;
        RECT 201.280 4431.505 201.450 4431.585 ;
        RECT 201.620 4431.555 202.640 4431.885 ;
        RECT 198.560 4431.295 199.210 4431.505 ;
        RECT 200.480 4431.385 201.450 4431.505 ;
        RECT 202.470 4431.400 202.640 4431.555 ;
        RECT 203.180 4432.475 203.830 4432.645 ;
        RECT 203.180 4431.805 203.350 4432.475 ;
        RECT 204.000 4432.305 204.170 4432.505 ;
        RECT 203.520 4432.215 204.170 4432.305 ;
        RECT 203.520 4432.045 204.000 4432.215 ;
        RECT 203.520 4431.975 204.170 4432.045 ;
        RECT 203.180 4431.635 203.825 4431.805 ;
        RECT 204.000 4431.755 204.170 4431.975 ;
        RECT 203.180 4431.400 203.350 4431.635 ;
        RECT 204.000 4431.465 204.170 4431.585 ;
        RECT 198.730 4431.175 199.210 4431.295 ;
        RECT 198.560 4430.835 198.730 4431.125 ;
        RECT 198.560 4430.375 199.210 4430.665 ;
        RECT 198.730 4430.335 199.210 4430.375 ;
        RECT 198.560 4429.915 198.730 4430.205 ;
        RECT 198.730 4429.745 199.210 4429.825 ;
        RECT 198.560 4429.495 199.210 4429.745 ;
        RECT 198.560 4429.455 198.730 4429.495 ;
        RECT 198.560 4428.995 198.730 4429.285 ;
        RECT 198.730 4428.825 199.210 4428.985 ;
        RECT 199.720 4428.895 199.890 4431.345 ;
        RECT 200.480 4431.295 202.250 4431.385 ;
        RECT 200.480 4431.175 201.280 4431.295 ;
        RECT 201.450 4431.215 202.250 4431.295 ;
        RECT 202.470 4431.225 203.350 4431.400 ;
        RECT 203.520 4431.295 204.170 4431.465 ;
        RECT 201.280 4430.835 201.450 4431.125 ;
      LAYER li1 ;
        RECT 201.620 4430.795 202.640 4430.965 ;
      LAYER li1 ;
        RECT 200.480 4430.625 201.450 4430.665 ;
        RECT 200.480 4430.375 202.250 4430.625 ;
        RECT 200.480 4430.335 201.280 4430.375 ;
        RECT 201.450 4430.295 202.250 4430.375 ;
        RECT 201.280 4429.915 201.450 4430.205 ;
      LAYER li1 ;
        RECT 202.470 4430.125 202.640 4430.795 ;
        RECT 201.620 4429.955 202.640 4430.125 ;
      LAYER li1 ;
        RECT 200.480 4429.745 201.280 4429.825 ;
        RECT 201.450 4429.745 202.250 4429.785 ;
        RECT 200.480 4429.495 202.250 4429.745 ;
        RECT 201.280 4429.455 202.250 4429.495 ;
      LAYER li1 ;
        RECT 202.470 4429.285 202.640 4429.955 ;
      LAYER li1 ;
        RECT 201.280 4428.995 201.450 4429.285 ;
      LAYER li1 ;
        RECT 201.620 4429.115 202.640 4429.285 ;
      LAYER li1 ;
        RECT 198.560 4428.655 199.210 4428.825 ;
        RECT 199.380 4428.720 200.260 4428.895 ;
        RECT 200.480 4428.825 201.280 4428.905 ;
        RECT 201.450 4428.825 202.250 4428.945 ;
        RECT 200.480 4428.735 202.250 4428.825 ;
        RECT 198.560 4428.535 198.730 4428.655 ;
        RECT 199.380 4428.485 199.550 4428.720 ;
        RECT 200.090 4428.565 200.260 4428.720 ;
        RECT 201.280 4428.615 202.250 4428.735 ;
        RECT 198.560 4428.145 198.730 4428.365 ;
        RECT 198.905 4428.315 199.550 4428.485 ;
        RECT 198.560 4428.075 199.210 4428.145 ;
        RECT 198.730 4427.905 199.210 4428.075 ;
        RECT 198.560 4427.815 199.210 4427.905 ;
        RECT 198.560 4427.615 198.730 4427.815 ;
        RECT 199.380 4427.645 199.550 4428.315 ;
        RECT 198.900 4427.475 199.550 4427.645 ;
        RECT 198.560 4427.215 198.730 4427.445 ;
      LAYER li1 ;
        RECT 199.720 4427.440 199.920 4428.540 ;
      LAYER li1 ;
        RECT 200.090 4428.235 201.110 4428.565 ;
        RECT 201.280 4428.535 201.450 4428.615 ;
      LAYER li1 ;
        RECT 202.470 4428.530 202.640 4429.115 ;
      LAYER li1 ;
        RECT 202.840 4428.775 203.010 4431.225 ;
        RECT 203.520 4431.135 204.000 4431.295 ;
      LAYER li1 ;
        RECT 203.180 4430.795 203.830 4430.965 ;
      LAYER li1 ;
        RECT 204.000 4430.835 204.170 4431.125 ;
      LAYER li1 ;
        RECT 203.180 4430.125 203.350 4430.795 ;
      LAYER li1 ;
        RECT 204.000 4430.625 204.170 4430.665 ;
        RECT 203.520 4430.375 204.170 4430.625 ;
        RECT 203.520 4430.295 204.000 4430.375 ;
      LAYER li1 ;
        RECT 203.180 4429.955 203.830 4430.125 ;
        RECT 203.180 4429.285 203.350 4429.955 ;
      LAYER li1 ;
        RECT 204.000 4429.915 204.170 4430.205 ;
        RECT 203.520 4429.745 204.000 4429.785 ;
        RECT 203.520 4429.455 204.170 4429.745 ;
      LAYER li1 ;
        RECT 203.180 4429.115 203.830 4429.285 ;
        RECT 203.180 4428.530 203.350 4429.115 ;
      LAYER li1 ;
        RECT 204.000 4428.995 204.170 4429.285 ;
        RECT 203.520 4428.825 204.000 4428.945 ;
        RECT 203.520 4428.615 204.170 4428.825 ;
        RECT 204.000 4428.535 204.170 4428.615 ;
      LAYER li1 ;
        RECT 202.470 4428.445 203.350 4428.530 ;
      LAYER li1 ;
        RECT 200.090 4427.725 200.260 4428.235 ;
        RECT 201.280 4428.105 201.450 4428.365 ;
      LAYER li1 ;
        RECT 201.620 4428.275 203.830 4428.445 ;
      LAYER li1 ;
        RECT 204.000 4428.105 204.170 4428.365 ;
        RECT 201.280 4428.075 202.600 4428.105 ;
        RECT 200.480 4427.905 201.280 4428.065 ;
        RECT 201.450 4427.905 202.600 4428.075 ;
        RECT 200.480 4427.895 202.600 4427.905 ;
        RECT 201.280 4427.775 202.600 4427.895 ;
        RECT 203.200 4428.075 204.170 4428.105 ;
        RECT 203.200 4427.905 204.000 4428.075 ;
        RECT 203.200 4427.775 204.170 4427.905 ;
        RECT 200.090 4427.395 201.110 4427.725 ;
        RECT 201.280 4427.615 201.450 4427.775 ;
        RECT 204.000 4427.615 204.170 4427.775 ;
        RECT 201.280 4427.215 201.450 4427.445 ;
        RECT 204.000 4427.215 204.170 4427.445 ;
        RECT 198.560 4427.155 199.455 4427.215 ;
        RECT 198.730 4426.985 199.455 4427.155 ;
        RECT 198.560 4426.925 199.455 4426.985 ;
        RECT 200.115 4427.155 202.615 4427.215 ;
        RECT 200.115 4426.985 201.280 4427.155 ;
        RECT 201.450 4426.985 202.615 4427.155 ;
        RECT 200.115 4426.925 202.615 4426.985 ;
        RECT 203.275 4427.155 204.170 4427.215 ;
        RECT 203.275 4426.985 204.000 4427.155 ;
        RECT 203.275 4426.925 204.170 4426.985 ;
        RECT 198.560 4426.840 198.730 4426.925 ;
        RECT 201.280 4426.840 201.450 4426.925 ;
        RECT 204.000 4426.840 204.170 4426.925 ;
        RECT 3383.500 3572.315 3383.670 3572.400 ;
        RECT 3386.220 3572.315 3386.390 3572.400 ;
        RECT 3388.940 3572.315 3389.110 3572.400 ;
        RECT 3383.500 3572.255 3384.395 3572.315 ;
        RECT 3383.670 3572.085 3384.395 3572.255 ;
        RECT 3383.500 3572.025 3384.395 3572.085 ;
        RECT 3383.500 3571.795 3383.670 3572.025 ;
        RECT 3383.500 3571.425 3383.670 3571.625 ;
        RECT 3383.840 3571.595 3384.490 3571.765 ;
        RECT 3383.500 3571.335 3384.150 3571.425 ;
        RECT 3383.670 3571.165 3384.150 3571.335 ;
        RECT 3383.500 3571.095 3384.150 3571.165 ;
        RECT 3383.500 3570.875 3383.670 3571.095 ;
        RECT 3384.320 3570.925 3384.490 3571.595 ;
        RECT 3383.845 3570.755 3384.490 3570.925 ;
        RECT 3383.500 3570.585 3383.670 3570.705 ;
        RECT 3383.500 3570.415 3384.150 3570.585 ;
        RECT 3383.670 3570.255 3384.150 3570.415 ;
        RECT 3384.320 3570.520 3384.490 3570.755 ;
      LAYER li1 ;
        RECT 3384.660 3570.700 3384.860 3572.290 ;
      LAYER li1 ;
        RECT 3385.055 3572.255 3387.555 3572.315 ;
        RECT 3385.055 3572.085 3386.220 3572.255 ;
        RECT 3386.390 3572.085 3387.555 3572.255 ;
        RECT 3385.055 3572.025 3387.555 3572.085 ;
        RECT 3388.215 3572.255 3389.110 3572.315 ;
        RECT 3388.215 3572.085 3388.940 3572.255 ;
        RECT 3388.215 3572.025 3389.110 3572.085 ;
        RECT 3385.030 3571.515 3386.050 3571.845 ;
        RECT 3386.220 3571.795 3386.390 3572.025 ;
        RECT 3388.940 3571.795 3389.110 3572.025 ;
        RECT 3385.030 3571.005 3385.200 3571.515 ;
        RECT 3386.220 3571.465 3386.390 3571.625 ;
        RECT 3388.940 3571.465 3389.110 3571.625 ;
        RECT 3386.220 3571.345 3387.540 3571.465 ;
        RECT 3385.420 3571.335 3387.540 3571.345 ;
        RECT 3385.420 3571.175 3386.220 3571.335 ;
        RECT 3386.390 3571.165 3387.540 3571.335 ;
        RECT 3386.220 3571.135 3387.540 3571.165 ;
        RECT 3388.140 3571.335 3389.110 3571.465 ;
        RECT 3388.140 3571.165 3388.940 3571.335 ;
        RECT 3388.140 3571.135 3389.110 3571.165 ;
        RECT 3385.030 3570.675 3386.050 3571.005 ;
        RECT 3386.220 3570.875 3386.390 3571.135 ;
      LAYER li1 ;
        RECT 3386.560 3570.795 3388.770 3570.965 ;
      LAYER li1 ;
        RECT 3388.940 3570.875 3389.110 3571.135 ;
      LAYER li1 ;
        RECT 3387.410 3570.710 3388.290 3570.795 ;
      LAYER li1 ;
        RECT 3385.030 3570.520 3385.200 3570.675 ;
        RECT 3384.320 3570.345 3385.200 3570.520 ;
        RECT 3386.220 3570.625 3386.390 3570.705 ;
        RECT 3386.220 3570.505 3387.190 3570.625 ;
        RECT 3385.420 3570.415 3387.190 3570.505 ;
        RECT 3383.500 3569.955 3383.670 3570.245 ;
      LAYER li1 ;
        RECT 3383.840 3569.915 3384.490 3570.085 ;
      LAYER li1 ;
        RECT 3383.500 3569.745 3383.670 3569.785 ;
        RECT 3383.500 3569.495 3384.150 3569.745 ;
        RECT 3383.670 3569.415 3384.150 3569.495 ;
        RECT 3383.500 3569.035 3383.670 3569.325 ;
      LAYER li1 ;
        RECT 3384.320 3569.245 3384.490 3569.915 ;
        RECT 3383.840 3569.075 3384.490 3569.245 ;
      LAYER li1 ;
        RECT 3383.670 3568.865 3384.150 3568.905 ;
        RECT 3383.500 3568.575 3384.150 3568.865 ;
      LAYER li1 ;
        RECT 3384.320 3568.405 3384.490 3569.075 ;
      LAYER li1 ;
        RECT 3383.500 3568.115 3383.670 3568.405 ;
      LAYER li1 ;
        RECT 3383.840 3568.235 3384.490 3568.405 ;
      LAYER li1 ;
        RECT 3383.670 3567.945 3384.150 3568.065 ;
        RECT 3383.500 3567.735 3384.150 3567.945 ;
        RECT 3383.500 3567.655 3383.670 3567.735 ;
      LAYER li1 ;
        RECT 3384.320 3567.650 3384.490 3568.235 ;
      LAYER li1 ;
        RECT 3384.660 3567.895 3384.830 3570.345 ;
        RECT 3385.420 3570.335 3386.220 3570.415 ;
        RECT 3386.390 3570.295 3387.190 3570.415 ;
      LAYER li1 ;
        RECT 3385.030 3569.915 3386.050 3570.085 ;
      LAYER li1 ;
        RECT 3386.220 3569.955 3386.390 3570.245 ;
      LAYER li1 ;
        RECT 3387.410 3570.125 3387.580 3570.710 ;
        RECT 3386.560 3569.955 3387.580 3570.125 ;
        RECT 3385.030 3569.245 3385.200 3569.915 ;
      LAYER li1 ;
        RECT 3386.220 3569.745 3387.190 3569.785 ;
        RECT 3385.420 3569.495 3387.190 3569.745 ;
        RECT 3385.420 3569.415 3386.220 3569.495 ;
        RECT 3386.390 3569.455 3387.190 3569.495 ;
      LAYER li1 ;
        RECT 3385.030 3569.075 3386.050 3569.245 ;
        RECT 3385.030 3568.405 3385.200 3569.075 ;
      LAYER li1 ;
        RECT 3386.220 3569.035 3386.390 3569.325 ;
      LAYER li1 ;
        RECT 3387.410 3569.285 3387.580 3569.955 ;
        RECT 3386.560 3569.115 3387.580 3569.285 ;
      LAYER li1 ;
        RECT 3385.420 3568.865 3386.220 3568.905 ;
        RECT 3386.390 3568.865 3387.190 3568.945 ;
        RECT 3385.420 3568.615 3387.190 3568.865 ;
        RECT 3385.420 3568.575 3386.390 3568.615 ;
      LAYER li1 ;
        RECT 3387.410 3568.445 3387.580 3569.115 ;
        RECT 3385.030 3568.235 3386.050 3568.405 ;
        RECT 3385.030 3567.650 3385.200 3568.235 ;
      LAYER li1 ;
        RECT 3386.220 3568.115 3386.390 3568.405 ;
      LAYER li1 ;
        RECT 3386.560 3568.275 3387.580 3568.445 ;
      LAYER li1 ;
        RECT 3385.420 3567.945 3386.220 3568.065 ;
        RECT 3386.390 3567.945 3387.190 3568.025 ;
        RECT 3387.780 3568.015 3387.950 3570.465 ;
      LAYER li1 ;
        RECT 3388.120 3570.125 3388.290 3570.710 ;
      LAYER li1 ;
        RECT 3388.940 3570.625 3389.110 3570.705 ;
        RECT 3388.460 3570.415 3389.110 3570.625 ;
        RECT 3388.460 3570.295 3388.940 3570.415 ;
      LAYER li1 ;
        RECT 3388.120 3569.955 3388.770 3570.125 ;
      LAYER li1 ;
        RECT 3388.940 3569.955 3389.110 3570.245 ;
      LAYER li1 ;
        RECT 3388.120 3569.285 3388.290 3569.955 ;
      LAYER li1 ;
        RECT 3388.460 3569.495 3389.110 3569.785 ;
        RECT 3388.460 3569.455 3388.940 3569.495 ;
      LAYER li1 ;
        RECT 3388.120 3569.115 3388.770 3569.285 ;
        RECT 3388.120 3568.445 3388.290 3569.115 ;
      LAYER li1 ;
        RECT 3388.940 3569.035 3389.110 3569.325 ;
        RECT 3388.460 3568.865 3388.940 3568.945 ;
        RECT 3388.460 3568.615 3389.110 3568.865 ;
        RECT 3388.940 3568.575 3389.110 3568.615 ;
      LAYER li1 ;
        RECT 3388.120 3568.275 3388.770 3568.445 ;
      LAYER li1 ;
        RECT 3388.940 3568.115 3389.110 3568.405 ;
        RECT 3385.420 3567.855 3387.190 3567.945 ;
        RECT 3385.420 3567.735 3386.390 3567.855 ;
        RECT 3386.220 3567.655 3386.390 3567.735 ;
        RECT 3387.410 3567.840 3388.290 3568.015 ;
        RECT 3387.410 3567.685 3387.580 3567.840 ;
      LAYER li1 ;
        RECT 3384.320 3567.565 3385.200 3567.650 ;
      LAYER li1 ;
        RECT 3383.500 3567.225 3383.670 3567.485 ;
      LAYER li1 ;
        RECT 3383.840 3567.395 3386.050 3567.565 ;
      LAYER li1 ;
        RECT 3386.220 3567.225 3386.390 3567.485 ;
        RECT 3386.560 3567.355 3387.580 3567.685 ;
        RECT 3383.500 3567.195 3384.470 3567.225 ;
        RECT 3383.670 3567.025 3384.470 3567.195 ;
        RECT 3383.500 3566.895 3384.470 3567.025 ;
        RECT 3385.070 3567.195 3386.390 3567.225 ;
        RECT 3385.070 3567.025 3386.220 3567.195 ;
        RECT 3386.390 3567.025 3387.190 3567.185 ;
        RECT 3385.070 3567.015 3387.190 3567.025 ;
        RECT 3385.070 3566.895 3386.390 3567.015 ;
        RECT 3383.500 3566.735 3383.670 3566.895 ;
        RECT 3386.220 3566.735 3386.390 3566.895 ;
        RECT 3387.410 3566.845 3387.580 3567.355 ;
        RECT 3383.500 3566.335 3383.670 3566.565 ;
        RECT 3386.220 3566.335 3386.390 3566.565 ;
        RECT 3386.560 3566.515 3387.580 3566.845 ;
      LAYER li1 ;
        RECT 3387.750 3566.560 3387.950 3567.660 ;
      LAYER li1 ;
        RECT 3388.120 3567.605 3388.290 3567.840 ;
        RECT 3388.460 3567.945 3388.940 3568.105 ;
        RECT 3388.460 3567.775 3389.110 3567.945 ;
        RECT 3388.940 3567.655 3389.110 3567.775 ;
        RECT 3388.120 3567.435 3388.765 3567.605 ;
        RECT 3388.120 3566.765 3388.290 3567.435 ;
        RECT 3388.940 3567.265 3389.110 3567.485 ;
        RECT 3388.460 3567.195 3389.110 3567.265 ;
        RECT 3388.460 3567.025 3388.940 3567.195 ;
        RECT 3388.460 3566.935 3389.110 3567.025 ;
        RECT 3388.120 3566.595 3388.770 3566.765 ;
        RECT 3388.940 3566.735 3389.110 3566.935 ;
        RECT 3388.940 3566.335 3389.110 3566.565 ;
        RECT 3383.500 3566.275 3384.395 3566.335 ;
        RECT 3383.670 3566.105 3384.395 3566.275 ;
        RECT 3383.500 3566.045 3384.395 3566.105 ;
        RECT 3383.500 3565.815 3383.670 3566.045 ;
        RECT 3383.500 3565.445 3383.670 3565.645 ;
        RECT 3383.840 3565.615 3384.490 3565.785 ;
        RECT 3383.500 3565.355 3384.150 3565.445 ;
        RECT 3383.670 3565.185 3384.150 3565.355 ;
        RECT 3383.500 3565.115 3384.150 3565.185 ;
        RECT 3383.500 3564.895 3383.670 3565.115 ;
        RECT 3384.320 3564.945 3384.490 3565.615 ;
        RECT 3383.845 3564.775 3384.490 3564.945 ;
        RECT 3383.500 3564.605 3383.670 3564.725 ;
        RECT 3383.500 3564.435 3384.150 3564.605 ;
        RECT 3383.670 3564.275 3384.150 3564.435 ;
        RECT 3384.320 3564.540 3384.490 3564.775 ;
      LAYER li1 ;
        RECT 3384.660 3564.720 3384.860 3566.310 ;
      LAYER li1 ;
        RECT 3385.055 3566.275 3387.555 3566.335 ;
        RECT 3385.055 3566.105 3386.220 3566.275 ;
        RECT 3386.390 3566.105 3387.555 3566.275 ;
        RECT 3385.055 3566.045 3387.555 3566.105 ;
        RECT 3388.215 3566.275 3389.110 3566.335 ;
        RECT 3388.215 3566.105 3388.940 3566.275 ;
        RECT 3388.215 3566.045 3389.110 3566.105 ;
        RECT 3385.030 3565.535 3386.050 3565.865 ;
        RECT 3386.220 3565.815 3386.390 3566.045 ;
        RECT 3388.940 3565.815 3389.110 3566.045 ;
        RECT 3385.030 3565.025 3385.200 3565.535 ;
        RECT 3386.220 3565.485 3386.390 3565.645 ;
        RECT 3388.940 3565.485 3389.110 3565.645 ;
        RECT 3386.220 3565.365 3387.540 3565.485 ;
        RECT 3385.420 3565.355 3387.540 3565.365 ;
        RECT 3385.420 3565.195 3386.220 3565.355 ;
        RECT 3386.390 3565.185 3387.540 3565.355 ;
        RECT 3386.220 3565.155 3387.540 3565.185 ;
        RECT 3388.140 3565.355 3389.110 3565.485 ;
        RECT 3388.140 3565.185 3388.940 3565.355 ;
        RECT 3388.140 3565.155 3389.110 3565.185 ;
        RECT 3385.030 3564.695 3386.050 3565.025 ;
        RECT 3386.220 3564.895 3386.390 3565.155 ;
      LAYER li1 ;
        RECT 3386.560 3564.815 3388.770 3564.985 ;
      LAYER li1 ;
        RECT 3388.940 3564.895 3389.110 3565.155 ;
      LAYER li1 ;
        RECT 3387.410 3564.730 3388.290 3564.815 ;
      LAYER li1 ;
        RECT 3385.030 3564.540 3385.200 3564.695 ;
        RECT 3384.320 3564.365 3385.200 3564.540 ;
        RECT 3386.220 3564.645 3386.390 3564.725 ;
        RECT 3386.220 3564.525 3387.190 3564.645 ;
        RECT 3385.420 3564.435 3387.190 3564.525 ;
        RECT 3383.500 3563.975 3383.670 3564.265 ;
      LAYER li1 ;
        RECT 3383.840 3563.935 3384.490 3564.105 ;
      LAYER li1 ;
        RECT 3383.500 3563.765 3383.670 3563.805 ;
        RECT 3383.500 3563.515 3384.150 3563.765 ;
        RECT 3383.670 3563.435 3384.150 3563.515 ;
        RECT 3383.500 3563.055 3383.670 3563.345 ;
      LAYER li1 ;
        RECT 3384.320 3563.265 3384.490 3563.935 ;
        RECT 3383.840 3563.095 3384.490 3563.265 ;
      LAYER li1 ;
        RECT 3383.670 3562.885 3384.150 3562.925 ;
        RECT 3383.500 3562.595 3384.150 3562.885 ;
      LAYER li1 ;
        RECT 3384.320 3562.425 3384.490 3563.095 ;
      LAYER li1 ;
        RECT 3383.500 3562.135 3383.670 3562.425 ;
      LAYER li1 ;
        RECT 3383.840 3562.255 3384.490 3562.425 ;
      LAYER li1 ;
        RECT 3383.670 3561.965 3384.150 3562.085 ;
        RECT 3383.500 3561.755 3384.150 3561.965 ;
        RECT 3383.500 3561.675 3383.670 3561.755 ;
      LAYER li1 ;
        RECT 3384.320 3561.670 3384.490 3562.255 ;
      LAYER li1 ;
        RECT 3384.660 3561.915 3384.830 3564.365 ;
        RECT 3385.420 3564.355 3386.220 3564.435 ;
        RECT 3386.390 3564.315 3387.190 3564.435 ;
      LAYER li1 ;
        RECT 3385.030 3563.935 3386.050 3564.105 ;
      LAYER li1 ;
        RECT 3386.220 3563.975 3386.390 3564.265 ;
      LAYER li1 ;
        RECT 3387.410 3564.145 3387.580 3564.730 ;
        RECT 3386.560 3563.975 3387.580 3564.145 ;
        RECT 3385.030 3563.265 3385.200 3563.935 ;
      LAYER li1 ;
        RECT 3386.220 3563.765 3387.190 3563.805 ;
        RECT 3385.420 3563.515 3387.190 3563.765 ;
        RECT 3385.420 3563.435 3386.220 3563.515 ;
        RECT 3386.390 3563.475 3387.190 3563.515 ;
      LAYER li1 ;
        RECT 3385.030 3563.095 3386.050 3563.265 ;
        RECT 3385.030 3562.425 3385.200 3563.095 ;
      LAYER li1 ;
        RECT 3386.220 3563.055 3386.390 3563.345 ;
      LAYER li1 ;
        RECT 3387.410 3563.305 3387.580 3563.975 ;
        RECT 3386.560 3563.135 3387.580 3563.305 ;
      LAYER li1 ;
        RECT 3385.420 3562.885 3386.220 3562.925 ;
        RECT 3386.390 3562.885 3387.190 3562.965 ;
        RECT 3385.420 3562.635 3387.190 3562.885 ;
        RECT 3385.420 3562.595 3386.390 3562.635 ;
      LAYER li1 ;
        RECT 3387.410 3562.465 3387.580 3563.135 ;
        RECT 3385.030 3562.255 3386.050 3562.425 ;
        RECT 3385.030 3561.670 3385.200 3562.255 ;
      LAYER li1 ;
        RECT 3386.220 3562.135 3386.390 3562.425 ;
      LAYER li1 ;
        RECT 3386.560 3562.295 3387.580 3562.465 ;
      LAYER li1 ;
        RECT 3385.420 3561.965 3386.220 3562.085 ;
        RECT 3386.390 3561.965 3387.190 3562.045 ;
        RECT 3387.780 3562.035 3387.950 3564.485 ;
      LAYER li1 ;
        RECT 3388.120 3564.145 3388.290 3564.730 ;
      LAYER li1 ;
        RECT 3388.940 3564.645 3389.110 3564.725 ;
        RECT 3388.460 3564.435 3389.110 3564.645 ;
        RECT 3388.460 3564.315 3388.940 3564.435 ;
      LAYER li1 ;
        RECT 3388.120 3563.975 3388.770 3564.145 ;
      LAYER li1 ;
        RECT 3388.940 3563.975 3389.110 3564.265 ;
      LAYER li1 ;
        RECT 3388.120 3563.305 3388.290 3563.975 ;
      LAYER li1 ;
        RECT 3388.460 3563.515 3389.110 3563.805 ;
        RECT 3388.460 3563.475 3388.940 3563.515 ;
      LAYER li1 ;
        RECT 3388.120 3563.135 3388.770 3563.305 ;
        RECT 3388.120 3562.465 3388.290 3563.135 ;
      LAYER li1 ;
        RECT 3388.940 3563.055 3389.110 3563.345 ;
        RECT 3388.460 3562.885 3388.940 3562.965 ;
        RECT 3388.460 3562.635 3389.110 3562.885 ;
        RECT 3388.940 3562.595 3389.110 3562.635 ;
      LAYER li1 ;
        RECT 3388.120 3562.295 3388.770 3562.465 ;
      LAYER li1 ;
        RECT 3388.940 3562.135 3389.110 3562.425 ;
        RECT 3385.420 3561.875 3387.190 3561.965 ;
        RECT 3385.420 3561.755 3386.390 3561.875 ;
        RECT 3386.220 3561.675 3386.390 3561.755 ;
        RECT 3387.410 3561.860 3388.290 3562.035 ;
        RECT 3387.410 3561.705 3387.580 3561.860 ;
      LAYER li1 ;
        RECT 3384.320 3561.585 3385.200 3561.670 ;
      LAYER li1 ;
        RECT 3383.500 3561.245 3383.670 3561.505 ;
      LAYER li1 ;
        RECT 3383.840 3561.415 3386.050 3561.585 ;
      LAYER li1 ;
        RECT 3386.220 3561.245 3386.390 3561.505 ;
        RECT 3386.560 3561.375 3387.580 3561.705 ;
        RECT 3383.500 3561.215 3384.470 3561.245 ;
        RECT 3383.670 3561.045 3384.470 3561.215 ;
        RECT 3383.500 3560.915 3384.470 3561.045 ;
        RECT 3385.070 3561.215 3386.390 3561.245 ;
        RECT 3385.070 3561.045 3386.220 3561.215 ;
        RECT 3386.390 3561.045 3387.190 3561.205 ;
        RECT 3385.070 3561.035 3387.190 3561.045 ;
        RECT 3385.070 3560.915 3386.390 3561.035 ;
        RECT 3383.500 3560.755 3383.670 3560.915 ;
        RECT 3386.220 3560.755 3386.390 3560.915 ;
        RECT 3387.410 3560.865 3387.580 3561.375 ;
        RECT 3383.500 3560.355 3383.670 3560.585 ;
        RECT 3386.220 3560.355 3386.390 3560.585 ;
        RECT 3386.560 3560.535 3387.580 3560.865 ;
      LAYER li1 ;
        RECT 3387.750 3560.580 3387.950 3561.680 ;
      LAYER li1 ;
        RECT 3388.120 3561.625 3388.290 3561.860 ;
        RECT 3388.460 3561.965 3388.940 3562.125 ;
        RECT 3388.460 3561.795 3389.110 3561.965 ;
        RECT 3388.940 3561.675 3389.110 3561.795 ;
        RECT 3388.120 3561.455 3388.765 3561.625 ;
        RECT 3388.120 3560.785 3388.290 3561.455 ;
        RECT 3388.940 3561.285 3389.110 3561.505 ;
        RECT 3388.460 3561.215 3389.110 3561.285 ;
        RECT 3388.460 3561.045 3388.940 3561.215 ;
        RECT 3388.460 3560.955 3389.110 3561.045 ;
        RECT 3388.120 3560.615 3388.770 3560.785 ;
        RECT 3388.940 3560.755 3389.110 3560.955 ;
        RECT 3388.940 3560.355 3389.110 3560.585 ;
        RECT 3383.500 3560.295 3384.395 3560.355 ;
        RECT 3383.670 3560.125 3384.395 3560.295 ;
        RECT 3383.500 3560.065 3384.395 3560.125 ;
        RECT 3383.500 3559.835 3383.670 3560.065 ;
        RECT 3383.500 3559.465 3383.670 3559.665 ;
        RECT 3383.840 3559.635 3384.490 3559.805 ;
        RECT 3383.500 3559.375 3384.150 3559.465 ;
        RECT 3383.670 3559.205 3384.150 3559.375 ;
        RECT 3383.500 3559.135 3384.150 3559.205 ;
        RECT 3383.500 3558.915 3383.670 3559.135 ;
        RECT 3384.320 3558.965 3384.490 3559.635 ;
        RECT 3383.845 3558.795 3384.490 3558.965 ;
        RECT 3383.500 3558.625 3383.670 3558.745 ;
        RECT 3383.500 3558.455 3384.150 3558.625 ;
        RECT 3383.670 3558.295 3384.150 3558.455 ;
        RECT 3384.320 3558.560 3384.490 3558.795 ;
      LAYER li1 ;
        RECT 3384.660 3558.740 3384.860 3560.330 ;
      LAYER li1 ;
        RECT 3385.055 3560.295 3387.555 3560.355 ;
        RECT 3385.055 3560.125 3386.220 3560.295 ;
        RECT 3386.390 3560.125 3387.555 3560.295 ;
        RECT 3385.055 3560.065 3387.555 3560.125 ;
        RECT 3388.215 3560.295 3389.110 3560.355 ;
        RECT 3388.215 3560.125 3388.940 3560.295 ;
        RECT 3388.215 3560.065 3389.110 3560.125 ;
        RECT 3385.030 3559.555 3386.050 3559.885 ;
        RECT 3386.220 3559.835 3386.390 3560.065 ;
        RECT 3388.940 3559.835 3389.110 3560.065 ;
        RECT 3385.030 3559.045 3385.200 3559.555 ;
        RECT 3386.220 3559.505 3386.390 3559.665 ;
        RECT 3388.940 3559.505 3389.110 3559.665 ;
        RECT 3386.220 3559.385 3387.540 3559.505 ;
        RECT 3385.420 3559.375 3387.540 3559.385 ;
        RECT 3385.420 3559.215 3386.220 3559.375 ;
        RECT 3386.390 3559.205 3387.540 3559.375 ;
        RECT 3386.220 3559.175 3387.540 3559.205 ;
        RECT 3388.140 3559.375 3389.110 3559.505 ;
        RECT 3388.140 3559.205 3388.940 3559.375 ;
        RECT 3388.140 3559.175 3389.110 3559.205 ;
        RECT 3385.030 3558.715 3386.050 3559.045 ;
        RECT 3386.220 3558.915 3386.390 3559.175 ;
      LAYER li1 ;
        RECT 3386.560 3558.835 3388.770 3559.005 ;
      LAYER li1 ;
        RECT 3388.940 3558.915 3389.110 3559.175 ;
      LAYER li1 ;
        RECT 3387.410 3558.750 3388.290 3558.835 ;
      LAYER li1 ;
        RECT 3385.030 3558.560 3385.200 3558.715 ;
        RECT 3384.320 3558.385 3385.200 3558.560 ;
        RECT 3386.220 3558.665 3386.390 3558.745 ;
        RECT 3386.220 3558.545 3387.190 3558.665 ;
        RECT 3385.420 3558.455 3387.190 3558.545 ;
        RECT 3383.500 3557.995 3383.670 3558.285 ;
      LAYER li1 ;
        RECT 3383.840 3557.955 3384.490 3558.125 ;
      LAYER li1 ;
        RECT 3383.500 3557.785 3383.670 3557.825 ;
        RECT 3383.500 3557.535 3384.150 3557.785 ;
        RECT 3383.670 3557.455 3384.150 3557.535 ;
        RECT 3383.500 3557.075 3383.670 3557.365 ;
      LAYER li1 ;
        RECT 3384.320 3557.285 3384.490 3557.955 ;
        RECT 3383.840 3557.115 3384.490 3557.285 ;
      LAYER li1 ;
        RECT 3383.670 3556.905 3384.150 3556.945 ;
        RECT 3383.500 3556.615 3384.150 3556.905 ;
      LAYER li1 ;
        RECT 3384.320 3556.445 3384.490 3557.115 ;
      LAYER li1 ;
        RECT 3383.500 3556.155 3383.670 3556.445 ;
      LAYER li1 ;
        RECT 3383.840 3556.275 3384.490 3556.445 ;
      LAYER li1 ;
        RECT 3383.670 3555.985 3384.150 3556.105 ;
        RECT 3383.500 3555.775 3384.150 3555.985 ;
        RECT 3383.500 3555.695 3383.670 3555.775 ;
      LAYER li1 ;
        RECT 3384.320 3555.690 3384.490 3556.275 ;
      LAYER li1 ;
        RECT 3384.660 3555.935 3384.830 3558.385 ;
        RECT 3385.420 3558.375 3386.220 3558.455 ;
        RECT 3386.390 3558.335 3387.190 3558.455 ;
      LAYER li1 ;
        RECT 3385.030 3557.955 3386.050 3558.125 ;
      LAYER li1 ;
        RECT 3386.220 3557.995 3386.390 3558.285 ;
      LAYER li1 ;
        RECT 3387.410 3558.165 3387.580 3558.750 ;
        RECT 3386.560 3557.995 3387.580 3558.165 ;
        RECT 3385.030 3557.285 3385.200 3557.955 ;
      LAYER li1 ;
        RECT 3386.220 3557.785 3387.190 3557.825 ;
        RECT 3385.420 3557.535 3387.190 3557.785 ;
        RECT 3385.420 3557.455 3386.220 3557.535 ;
        RECT 3386.390 3557.495 3387.190 3557.535 ;
      LAYER li1 ;
        RECT 3385.030 3557.115 3386.050 3557.285 ;
        RECT 3385.030 3556.445 3385.200 3557.115 ;
      LAYER li1 ;
        RECT 3386.220 3557.075 3386.390 3557.365 ;
      LAYER li1 ;
        RECT 3387.410 3557.325 3387.580 3557.995 ;
        RECT 3386.560 3557.155 3387.580 3557.325 ;
      LAYER li1 ;
        RECT 3385.420 3556.905 3386.220 3556.945 ;
        RECT 3386.390 3556.905 3387.190 3556.985 ;
        RECT 3385.420 3556.655 3387.190 3556.905 ;
        RECT 3385.420 3556.615 3386.390 3556.655 ;
      LAYER li1 ;
        RECT 3387.410 3556.485 3387.580 3557.155 ;
        RECT 3385.030 3556.275 3386.050 3556.445 ;
        RECT 3385.030 3555.690 3385.200 3556.275 ;
      LAYER li1 ;
        RECT 3386.220 3556.155 3386.390 3556.445 ;
      LAYER li1 ;
        RECT 3386.560 3556.315 3387.580 3556.485 ;
      LAYER li1 ;
        RECT 3385.420 3555.985 3386.220 3556.105 ;
        RECT 3386.390 3555.985 3387.190 3556.065 ;
        RECT 3387.780 3556.055 3387.950 3558.505 ;
      LAYER li1 ;
        RECT 3388.120 3558.165 3388.290 3558.750 ;
      LAYER li1 ;
        RECT 3388.940 3558.665 3389.110 3558.745 ;
        RECT 3388.460 3558.455 3389.110 3558.665 ;
        RECT 3388.460 3558.335 3388.940 3558.455 ;
      LAYER li1 ;
        RECT 3388.120 3557.995 3388.770 3558.165 ;
      LAYER li1 ;
        RECT 3388.940 3557.995 3389.110 3558.285 ;
      LAYER li1 ;
        RECT 3388.120 3557.325 3388.290 3557.995 ;
      LAYER li1 ;
        RECT 3388.460 3557.535 3389.110 3557.825 ;
        RECT 3388.460 3557.495 3388.940 3557.535 ;
      LAYER li1 ;
        RECT 3388.120 3557.155 3388.770 3557.325 ;
        RECT 3388.120 3556.485 3388.290 3557.155 ;
      LAYER li1 ;
        RECT 3388.940 3557.075 3389.110 3557.365 ;
        RECT 3388.460 3556.905 3388.940 3556.985 ;
        RECT 3388.460 3556.655 3389.110 3556.905 ;
        RECT 3388.940 3556.615 3389.110 3556.655 ;
      LAYER li1 ;
        RECT 3388.120 3556.315 3388.770 3556.485 ;
      LAYER li1 ;
        RECT 3388.940 3556.155 3389.110 3556.445 ;
        RECT 3385.420 3555.895 3387.190 3555.985 ;
        RECT 3385.420 3555.775 3386.390 3555.895 ;
        RECT 3386.220 3555.695 3386.390 3555.775 ;
        RECT 3387.410 3555.880 3388.290 3556.055 ;
        RECT 3387.410 3555.725 3387.580 3555.880 ;
      LAYER li1 ;
        RECT 3384.320 3555.605 3385.200 3555.690 ;
      LAYER li1 ;
        RECT 3383.500 3555.265 3383.670 3555.525 ;
      LAYER li1 ;
        RECT 3383.840 3555.435 3386.050 3555.605 ;
      LAYER li1 ;
        RECT 3386.220 3555.265 3386.390 3555.525 ;
        RECT 3386.560 3555.395 3387.580 3555.725 ;
        RECT 3383.500 3555.235 3384.470 3555.265 ;
        RECT 3383.670 3555.065 3384.470 3555.235 ;
        RECT 3383.500 3554.935 3384.470 3555.065 ;
        RECT 3385.070 3555.235 3386.390 3555.265 ;
        RECT 3385.070 3555.065 3386.220 3555.235 ;
        RECT 3386.390 3555.065 3387.190 3555.225 ;
        RECT 3385.070 3555.055 3387.190 3555.065 ;
        RECT 3385.070 3554.935 3386.390 3555.055 ;
        RECT 3383.500 3554.775 3383.670 3554.935 ;
        RECT 3386.220 3554.775 3386.390 3554.935 ;
        RECT 3387.410 3554.885 3387.580 3555.395 ;
        RECT 3383.500 3554.375 3383.670 3554.605 ;
        RECT 3386.220 3554.375 3386.390 3554.605 ;
        RECT 3386.560 3554.555 3387.580 3554.885 ;
      LAYER li1 ;
        RECT 3387.750 3554.600 3387.950 3555.700 ;
      LAYER li1 ;
        RECT 3388.120 3555.645 3388.290 3555.880 ;
        RECT 3388.460 3555.985 3388.940 3556.145 ;
        RECT 3388.460 3555.815 3389.110 3555.985 ;
        RECT 3388.940 3555.695 3389.110 3555.815 ;
        RECT 3388.120 3555.475 3388.765 3555.645 ;
        RECT 3388.120 3554.805 3388.290 3555.475 ;
        RECT 3388.940 3555.305 3389.110 3555.525 ;
        RECT 3388.460 3555.235 3389.110 3555.305 ;
        RECT 3388.460 3555.065 3388.940 3555.235 ;
        RECT 3388.460 3554.975 3389.110 3555.065 ;
        RECT 3388.120 3554.635 3388.770 3554.805 ;
        RECT 3388.940 3554.775 3389.110 3554.975 ;
        RECT 3388.940 3554.375 3389.110 3554.605 ;
        RECT 3383.500 3554.315 3384.395 3554.375 ;
        RECT 3383.670 3554.145 3384.395 3554.315 ;
        RECT 3383.500 3554.085 3384.395 3554.145 ;
        RECT 3383.500 3553.855 3383.670 3554.085 ;
        RECT 3383.500 3553.485 3383.670 3553.685 ;
        RECT 3383.840 3553.655 3384.490 3553.825 ;
        RECT 3383.500 3553.395 3384.150 3553.485 ;
        RECT 3383.670 3553.225 3384.150 3553.395 ;
        RECT 3383.500 3553.155 3384.150 3553.225 ;
        RECT 3383.500 3552.935 3383.670 3553.155 ;
        RECT 3384.320 3552.985 3384.490 3553.655 ;
        RECT 3383.845 3552.815 3384.490 3552.985 ;
        RECT 3383.500 3552.645 3383.670 3552.765 ;
        RECT 3383.500 3552.475 3384.150 3552.645 ;
        RECT 3383.670 3552.315 3384.150 3552.475 ;
        RECT 3384.320 3552.580 3384.490 3552.815 ;
      LAYER li1 ;
        RECT 3384.660 3552.760 3384.860 3554.350 ;
      LAYER li1 ;
        RECT 3385.055 3554.315 3387.555 3554.375 ;
        RECT 3385.055 3554.145 3386.220 3554.315 ;
        RECT 3386.390 3554.145 3387.555 3554.315 ;
        RECT 3385.055 3554.085 3387.555 3554.145 ;
        RECT 3388.215 3554.315 3389.110 3554.375 ;
        RECT 3388.215 3554.145 3388.940 3554.315 ;
        RECT 3388.215 3554.085 3389.110 3554.145 ;
        RECT 3385.030 3553.575 3386.050 3553.905 ;
        RECT 3386.220 3553.855 3386.390 3554.085 ;
        RECT 3388.940 3553.855 3389.110 3554.085 ;
        RECT 3385.030 3553.065 3385.200 3553.575 ;
        RECT 3386.220 3553.525 3386.390 3553.685 ;
        RECT 3388.940 3553.525 3389.110 3553.685 ;
        RECT 3386.220 3553.405 3387.540 3553.525 ;
        RECT 3385.420 3553.395 3387.540 3553.405 ;
        RECT 3385.420 3553.235 3386.220 3553.395 ;
        RECT 3386.390 3553.225 3387.540 3553.395 ;
        RECT 3386.220 3553.195 3387.540 3553.225 ;
        RECT 3388.140 3553.395 3389.110 3553.525 ;
        RECT 3388.140 3553.225 3388.940 3553.395 ;
        RECT 3388.140 3553.195 3389.110 3553.225 ;
        RECT 3385.030 3552.735 3386.050 3553.065 ;
        RECT 3386.220 3552.935 3386.390 3553.195 ;
      LAYER li1 ;
        RECT 3386.560 3552.855 3388.770 3553.025 ;
      LAYER li1 ;
        RECT 3388.940 3552.935 3389.110 3553.195 ;
      LAYER li1 ;
        RECT 3387.410 3552.770 3388.290 3552.855 ;
      LAYER li1 ;
        RECT 3385.030 3552.580 3385.200 3552.735 ;
        RECT 3384.320 3552.405 3385.200 3552.580 ;
        RECT 3386.220 3552.685 3386.390 3552.765 ;
        RECT 3386.220 3552.565 3387.190 3552.685 ;
        RECT 3385.420 3552.475 3387.190 3552.565 ;
        RECT 3383.500 3552.015 3383.670 3552.305 ;
      LAYER li1 ;
        RECT 3383.840 3551.975 3384.490 3552.145 ;
      LAYER li1 ;
        RECT 3383.500 3551.805 3383.670 3551.845 ;
        RECT 3383.500 3551.555 3384.150 3551.805 ;
        RECT 3383.670 3551.475 3384.150 3551.555 ;
        RECT 3383.500 3551.095 3383.670 3551.385 ;
      LAYER li1 ;
        RECT 3384.320 3551.305 3384.490 3551.975 ;
        RECT 3383.840 3551.135 3384.490 3551.305 ;
      LAYER li1 ;
        RECT 3383.670 3550.925 3384.150 3550.965 ;
        RECT 3383.500 3550.635 3384.150 3550.925 ;
      LAYER li1 ;
        RECT 3384.320 3550.465 3384.490 3551.135 ;
      LAYER li1 ;
        RECT 3383.500 3550.175 3383.670 3550.465 ;
      LAYER li1 ;
        RECT 3383.840 3550.295 3384.490 3550.465 ;
      LAYER li1 ;
        RECT 3383.670 3550.005 3384.150 3550.125 ;
        RECT 3383.500 3549.795 3384.150 3550.005 ;
        RECT 3383.500 3549.715 3383.670 3549.795 ;
      LAYER li1 ;
        RECT 3384.320 3549.710 3384.490 3550.295 ;
      LAYER li1 ;
        RECT 3384.660 3549.955 3384.830 3552.405 ;
        RECT 3385.420 3552.395 3386.220 3552.475 ;
        RECT 3386.390 3552.355 3387.190 3552.475 ;
      LAYER li1 ;
        RECT 3385.030 3551.975 3386.050 3552.145 ;
      LAYER li1 ;
        RECT 3386.220 3552.015 3386.390 3552.305 ;
      LAYER li1 ;
        RECT 3387.410 3552.185 3387.580 3552.770 ;
        RECT 3386.560 3552.015 3387.580 3552.185 ;
        RECT 3385.030 3551.305 3385.200 3551.975 ;
      LAYER li1 ;
        RECT 3386.220 3551.805 3387.190 3551.845 ;
        RECT 3385.420 3551.555 3387.190 3551.805 ;
        RECT 3385.420 3551.475 3386.220 3551.555 ;
        RECT 3386.390 3551.515 3387.190 3551.555 ;
      LAYER li1 ;
        RECT 3385.030 3551.135 3386.050 3551.305 ;
        RECT 3385.030 3550.465 3385.200 3551.135 ;
      LAYER li1 ;
        RECT 3386.220 3551.095 3386.390 3551.385 ;
      LAYER li1 ;
        RECT 3387.410 3551.345 3387.580 3552.015 ;
        RECT 3386.560 3551.175 3387.580 3551.345 ;
      LAYER li1 ;
        RECT 3385.420 3550.925 3386.220 3550.965 ;
        RECT 3386.390 3550.925 3387.190 3551.005 ;
        RECT 3385.420 3550.675 3387.190 3550.925 ;
        RECT 3385.420 3550.635 3386.390 3550.675 ;
      LAYER li1 ;
        RECT 3387.410 3550.505 3387.580 3551.175 ;
        RECT 3385.030 3550.295 3386.050 3550.465 ;
        RECT 3385.030 3549.710 3385.200 3550.295 ;
      LAYER li1 ;
        RECT 3386.220 3550.175 3386.390 3550.465 ;
      LAYER li1 ;
        RECT 3386.560 3550.335 3387.580 3550.505 ;
      LAYER li1 ;
        RECT 3385.420 3550.005 3386.220 3550.125 ;
        RECT 3386.390 3550.005 3387.190 3550.085 ;
        RECT 3387.780 3550.075 3387.950 3552.525 ;
      LAYER li1 ;
        RECT 3388.120 3552.185 3388.290 3552.770 ;
      LAYER li1 ;
        RECT 3388.940 3552.685 3389.110 3552.765 ;
        RECT 3388.460 3552.475 3389.110 3552.685 ;
        RECT 3388.460 3552.355 3388.940 3552.475 ;
      LAYER li1 ;
        RECT 3388.120 3552.015 3388.770 3552.185 ;
      LAYER li1 ;
        RECT 3388.940 3552.015 3389.110 3552.305 ;
      LAYER li1 ;
        RECT 3388.120 3551.345 3388.290 3552.015 ;
      LAYER li1 ;
        RECT 3388.460 3551.555 3389.110 3551.845 ;
        RECT 3388.460 3551.515 3388.940 3551.555 ;
      LAYER li1 ;
        RECT 3388.120 3551.175 3388.770 3551.345 ;
        RECT 3388.120 3550.505 3388.290 3551.175 ;
      LAYER li1 ;
        RECT 3388.940 3551.095 3389.110 3551.385 ;
        RECT 3388.460 3550.925 3388.940 3551.005 ;
        RECT 3388.460 3550.675 3389.110 3550.925 ;
        RECT 3388.940 3550.635 3389.110 3550.675 ;
      LAYER li1 ;
        RECT 3388.120 3550.335 3388.770 3550.505 ;
      LAYER li1 ;
        RECT 3388.940 3550.175 3389.110 3550.465 ;
        RECT 3385.420 3549.915 3387.190 3550.005 ;
        RECT 3385.420 3549.795 3386.390 3549.915 ;
        RECT 3386.220 3549.715 3386.390 3549.795 ;
        RECT 3387.410 3549.900 3388.290 3550.075 ;
        RECT 3387.410 3549.745 3387.580 3549.900 ;
      LAYER li1 ;
        RECT 3384.320 3549.625 3385.200 3549.710 ;
      LAYER li1 ;
        RECT 3383.500 3549.285 3383.670 3549.545 ;
      LAYER li1 ;
        RECT 3383.840 3549.455 3386.050 3549.625 ;
      LAYER li1 ;
        RECT 3386.220 3549.285 3386.390 3549.545 ;
        RECT 3386.560 3549.415 3387.580 3549.745 ;
        RECT 3383.500 3549.255 3384.470 3549.285 ;
        RECT 3383.670 3549.085 3384.470 3549.255 ;
        RECT 3383.500 3548.955 3384.470 3549.085 ;
        RECT 3385.070 3549.255 3386.390 3549.285 ;
        RECT 3385.070 3549.085 3386.220 3549.255 ;
        RECT 3386.390 3549.085 3387.190 3549.245 ;
        RECT 3385.070 3549.075 3387.190 3549.085 ;
        RECT 3385.070 3548.955 3386.390 3549.075 ;
        RECT 3383.500 3548.795 3383.670 3548.955 ;
        RECT 3386.220 3548.795 3386.390 3548.955 ;
        RECT 3387.410 3548.905 3387.580 3549.415 ;
        RECT 3383.500 3548.395 3383.670 3548.625 ;
        RECT 3386.220 3548.395 3386.390 3548.625 ;
        RECT 3386.560 3548.575 3387.580 3548.905 ;
      LAYER li1 ;
        RECT 3387.750 3548.620 3387.950 3549.720 ;
      LAYER li1 ;
        RECT 3388.120 3549.665 3388.290 3549.900 ;
        RECT 3388.460 3550.005 3388.940 3550.165 ;
        RECT 3388.460 3549.835 3389.110 3550.005 ;
        RECT 3388.940 3549.715 3389.110 3549.835 ;
        RECT 3388.120 3549.495 3388.765 3549.665 ;
        RECT 3388.120 3548.825 3388.290 3549.495 ;
        RECT 3388.940 3549.325 3389.110 3549.545 ;
        RECT 3388.460 3549.255 3389.110 3549.325 ;
        RECT 3388.460 3549.085 3388.940 3549.255 ;
        RECT 3388.460 3548.995 3389.110 3549.085 ;
        RECT 3388.120 3548.655 3388.770 3548.825 ;
        RECT 3388.940 3548.795 3389.110 3548.995 ;
        RECT 3388.940 3548.395 3389.110 3548.625 ;
        RECT 3383.500 3548.335 3384.395 3548.395 ;
        RECT 3383.670 3548.165 3384.395 3548.335 ;
        RECT 3383.500 3548.105 3384.395 3548.165 ;
        RECT 3385.055 3548.335 3387.555 3548.395 ;
        RECT 3385.055 3548.165 3386.220 3548.335 ;
        RECT 3386.390 3548.165 3387.555 3548.335 ;
        RECT 3385.055 3548.105 3387.555 3548.165 ;
        RECT 3388.215 3548.335 3389.110 3548.395 ;
        RECT 3388.215 3548.165 3388.940 3548.335 ;
        RECT 3388.215 3548.105 3389.110 3548.165 ;
        RECT 3383.500 3547.875 3383.670 3548.105 ;
        RECT 3383.500 3547.505 3383.670 3547.705 ;
        RECT 3383.840 3547.675 3384.490 3547.845 ;
        RECT 3383.500 3547.415 3384.150 3547.505 ;
        RECT 3383.670 3547.245 3384.150 3547.415 ;
        RECT 3383.500 3547.175 3384.150 3547.245 ;
        RECT 3383.500 3546.955 3383.670 3547.175 ;
        RECT 3384.320 3547.005 3384.490 3547.675 ;
        RECT 3383.845 3546.835 3384.490 3547.005 ;
        RECT 3383.500 3546.665 3383.670 3546.785 ;
        RECT 3383.500 3546.495 3384.150 3546.665 ;
        RECT 3383.670 3546.335 3384.150 3546.495 ;
        RECT 3384.320 3546.600 3384.490 3546.835 ;
        RECT 3385.030 3547.595 3386.050 3547.925 ;
        RECT 3386.220 3547.875 3386.390 3548.105 ;
        RECT 3388.940 3547.875 3389.110 3548.105 ;
        RECT 3385.030 3547.085 3385.200 3547.595 ;
        RECT 3386.220 3547.545 3386.390 3547.705 ;
        RECT 3388.940 3547.545 3389.110 3547.705 ;
        RECT 3386.220 3547.425 3387.540 3547.545 ;
        RECT 3385.420 3547.415 3387.540 3547.425 ;
        RECT 3385.420 3547.255 3386.220 3547.415 ;
        RECT 3386.390 3547.245 3387.540 3547.415 ;
        RECT 3386.220 3547.215 3387.540 3547.245 ;
        RECT 3388.140 3547.415 3389.110 3547.545 ;
        RECT 3388.140 3547.245 3388.940 3547.415 ;
        RECT 3388.140 3547.215 3389.110 3547.245 ;
        RECT 3385.030 3546.755 3386.050 3547.085 ;
        RECT 3386.220 3546.955 3386.390 3547.215 ;
        RECT 3388.940 3546.955 3389.110 3547.215 ;
        RECT 3385.030 3546.600 3385.200 3546.755 ;
        RECT 3384.320 3546.425 3385.200 3546.600 ;
        RECT 3386.220 3546.705 3386.390 3546.785 ;
        RECT 3388.940 3546.705 3389.110 3546.785 ;
        RECT 3386.220 3546.585 3387.190 3546.705 ;
        RECT 3385.420 3546.495 3387.190 3546.585 ;
        RECT 3383.500 3546.035 3383.670 3546.325 ;
      LAYER li1 ;
        RECT 3383.840 3545.995 3384.490 3546.165 ;
      LAYER li1 ;
        RECT 3383.500 3545.825 3383.670 3545.865 ;
        RECT 3383.500 3545.575 3384.150 3545.825 ;
        RECT 3383.670 3545.495 3384.150 3545.575 ;
        RECT 3383.500 3545.115 3383.670 3545.405 ;
      LAYER li1 ;
        RECT 3384.320 3545.325 3384.490 3545.995 ;
        RECT 3383.840 3545.155 3384.490 3545.325 ;
      LAYER li1 ;
        RECT 3383.670 3544.945 3384.150 3544.985 ;
        RECT 3383.500 3544.655 3384.150 3544.945 ;
      LAYER li1 ;
        RECT 3384.320 3544.485 3384.490 3545.155 ;
      LAYER li1 ;
        RECT 3383.500 3544.195 3383.670 3544.485 ;
      LAYER li1 ;
        RECT 3383.840 3544.315 3384.490 3544.485 ;
      LAYER li1 ;
        RECT 3383.670 3544.025 3384.150 3544.145 ;
        RECT 3383.500 3543.815 3384.150 3544.025 ;
        RECT 3383.500 3543.735 3383.670 3543.815 ;
      LAYER li1 ;
        RECT 3384.320 3543.730 3384.490 3544.315 ;
      LAYER li1 ;
        RECT 3384.660 3543.975 3384.830 3546.425 ;
        RECT 3385.420 3546.415 3386.220 3546.495 ;
        RECT 3386.390 3546.375 3387.190 3546.495 ;
      LAYER li1 ;
        RECT 3385.030 3545.995 3386.050 3546.165 ;
      LAYER li1 ;
        RECT 3386.220 3546.035 3386.390 3546.325 ;
      LAYER li1 ;
        RECT 3385.030 3545.325 3385.200 3545.995 ;
      LAYER li1 ;
        RECT 3386.220 3545.825 3387.190 3545.865 ;
        RECT 3385.420 3545.575 3387.190 3545.825 ;
        RECT 3385.420 3545.495 3386.220 3545.575 ;
        RECT 3386.390 3545.535 3387.190 3545.575 ;
      LAYER li1 ;
        RECT 3385.030 3545.155 3386.050 3545.325 ;
        RECT 3385.030 3544.485 3385.200 3545.155 ;
      LAYER li1 ;
        RECT 3386.220 3545.115 3386.390 3545.405 ;
        RECT 3385.420 3544.945 3386.220 3544.985 ;
        RECT 3386.390 3544.945 3387.190 3545.025 ;
        RECT 3385.420 3544.695 3387.190 3544.945 ;
        RECT 3385.420 3544.655 3386.390 3544.695 ;
      LAYER li1 ;
        RECT 3385.030 3544.315 3386.050 3544.485 ;
        RECT 3385.030 3543.730 3385.200 3544.315 ;
      LAYER li1 ;
        RECT 3386.220 3544.195 3386.390 3544.485 ;
        RECT 3385.420 3544.025 3386.220 3544.145 ;
        RECT 3386.390 3544.025 3387.190 3544.105 ;
        RECT 3387.780 3544.095 3387.950 3546.545 ;
        RECT 3388.460 3546.495 3389.110 3546.705 ;
        RECT 3388.460 3546.375 3388.940 3546.495 ;
        RECT 3388.940 3546.035 3389.110 3546.325 ;
        RECT 3388.460 3545.575 3389.110 3545.865 ;
        RECT 3388.460 3545.535 3388.940 3545.575 ;
        RECT 3388.940 3545.115 3389.110 3545.405 ;
        RECT 3388.460 3544.945 3388.940 3545.025 ;
        RECT 3388.460 3544.695 3389.110 3544.945 ;
        RECT 3388.940 3544.655 3389.110 3544.695 ;
        RECT 3388.940 3544.195 3389.110 3544.485 ;
        RECT 3385.420 3543.935 3387.190 3544.025 ;
        RECT 3385.420 3543.815 3386.390 3543.935 ;
        RECT 3386.220 3543.735 3386.390 3543.815 ;
        RECT 3387.410 3543.920 3388.290 3544.095 ;
        RECT 3387.410 3543.765 3387.580 3543.920 ;
      LAYER li1 ;
        RECT 3384.320 3543.645 3385.200 3543.730 ;
      LAYER li1 ;
        RECT 3383.500 3543.305 3383.670 3543.565 ;
      LAYER li1 ;
        RECT 3383.840 3543.475 3386.050 3543.645 ;
      LAYER li1 ;
        RECT 3386.220 3543.305 3386.390 3543.565 ;
        RECT 3386.560 3543.435 3387.580 3543.765 ;
        RECT 3383.500 3543.275 3384.470 3543.305 ;
        RECT 3383.670 3543.105 3384.470 3543.275 ;
        RECT 3383.500 3542.975 3384.470 3543.105 ;
        RECT 3385.070 3543.275 3386.390 3543.305 ;
        RECT 3385.070 3543.105 3386.220 3543.275 ;
        RECT 3386.390 3543.105 3387.190 3543.265 ;
        RECT 3385.070 3543.095 3387.190 3543.105 ;
        RECT 3385.070 3542.975 3386.390 3543.095 ;
        RECT 3383.500 3542.815 3383.670 3542.975 ;
        RECT 3386.220 3542.815 3386.390 3542.975 ;
        RECT 3387.410 3542.925 3387.580 3543.435 ;
        RECT 3383.500 3542.415 3383.670 3542.645 ;
        RECT 3386.220 3542.415 3386.390 3542.645 ;
        RECT 3386.560 3542.595 3387.580 3542.925 ;
      LAYER li1 ;
        RECT 3387.750 3542.640 3387.950 3543.740 ;
      LAYER li1 ;
        RECT 3388.120 3543.685 3388.290 3543.920 ;
        RECT 3388.460 3544.025 3388.940 3544.185 ;
        RECT 3388.460 3543.855 3389.110 3544.025 ;
        RECT 3388.940 3543.735 3389.110 3543.855 ;
        RECT 3388.120 3543.515 3388.765 3543.685 ;
        RECT 3388.120 3542.845 3388.290 3543.515 ;
        RECT 3388.940 3543.345 3389.110 3543.565 ;
        RECT 3388.460 3543.275 3389.110 3543.345 ;
        RECT 3388.460 3543.105 3388.940 3543.275 ;
        RECT 3388.460 3543.015 3389.110 3543.105 ;
        RECT 3388.120 3542.675 3388.770 3542.845 ;
        RECT 3388.940 3542.815 3389.110 3543.015 ;
        RECT 3388.940 3542.415 3389.110 3542.645 ;
        RECT 3383.500 3542.355 3384.395 3542.415 ;
        RECT 3383.670 3542.185 3384.395 3542.355 ;
        RECT 3383.500 3542.125 3384.395 3542.185 ;
        RECT 3385.055 3542.355 3387.555 3542.415 ;
        RECT 3385.055 3542.185 3386.220 3542.355 ;
        RECT 3386.390 3542.185 3387.555 3542.355 ;
        RECT 3385.055 3542.125 3387.555 3542.185 ;
        RECT 3388.215 3542.355 3389.110 3542.415 ;
        RECT 3388.215 3542.185 3388.940 3542.355 ;
        RECT 3388.215 3542.125 3389.110 3542.185 ;
        RECT 3383.500 3541.895 3383.670 3542.125 ;
        RECT 3383.500 3541.525 3383.670 3541.725 ;
        RECT 3383.840 3541.695 3384.490 3541.865 ;
        RECT 3383.500 3541.435 3384.150 3541.525 ;
        RECT 3383.670 3541.265 3384.150 3541.435 ;
        RECT 3383.500 3541.195 3384.150 3541.265 ;
        RECT 3383.500 3540.975 3383.670 3541.195 ;
        RECT 3384.320 3541.025 3384.490 3541.695 ;
        RECT 3383.845 3540.855 3384.490 3541.025 ;
        RECT 3383.500 3540.685 3383.670 3540.805 ;
        RECT 3383.500 3540.515 3384.150 3540.685 ;
        RECT 3383.670 3540.355 3384.150 3540.515 ;
        RECT 3384.320 3540.620 3384.490 3540.855 ;
        RECT 3385.030 3541.615 3386.050 3541.945 ;
        RECT 3386.220 3541.895 3386.390 3542.125 ;
        RECT 3388.940 3541.895 3389.110 3542.125 ;
        RECT 3385.030 3541.105 3385.200 3541.615 ;
        RECT 3386.220 3541.565 3386.390 3541.725 ;
        RECT 3388.940 3541.565 3389.110 3541.725 ;
        RECT 3386.220 3541.445 3387.540 3541.565 ;
        RECT 3385.420 3541.435 3387.540 3541.445 ;
        RECT 3385.420 3541.275 3386.220 3541.435 ;
        RECT 3386.390 3541.265 3387.540 3541.435 ;
        RECT 3386.220 3541.235 3387.540 3541.265 ;
        RECT 3388.140 3541.435 3389.110 3541.565 ;
        RECT 3388.140 3541.265 3388.940 3541.435 ;
        RECT 3388.140 3541.235 3389.110 3541.265 ;
        RECT 3385.030 3540.775 3386.050 3541.105 ;
        RECT 3386.220 3540.975 3386.390 3541.235 ;
        RECT 3388.940 3540.975 3389.110 3541.235 ;
        RECT 3385.030 3540.620 3385.200 3540.775 ;
        RECT 3384.320 3540.445 3385.200 3540.620 ;
        RECT 3386.220 3540.725 3386.390 3540.805 ;
        RECT 3388.940 3540.725 3389.110 3540.805 ;
        RECT 3386.220 3540.605 3387.190 3540.725 ;
        RECT 3385.420 3540.515 3387.190 3540.605 ;
        RECT 3383.500 3540.055 3383.670 3540.345 ;
      LAYER li1 ;
        RECT 3383.840 3540.015 3384.490 3540.185 ;
      LAYER li1 ;
        RECT 3383.500 3539.845 3383.670 3539.885 ;
        RECT 3383.500 3539.595 3384.150 3539.845 ;
        RECT 3383.670 3539.515 3384.150 3539.595 ;
        RECT 3383.500 3539.135 3383.670 3539.425 ;
      LAYER li1 ;
        RECT 3384.320 3539.345 3384.490 3540.015 ;
        RECT 3383.840 3539.175 3384.490 3539.345 ;
      LAYER li1 ;
        RECT 3383.670 3538.965 3384.150 3539.005 ;
        RECT 3383.500 3538.675 3384.150 3538.965 ;
      LAYER li1 ;
        RECT 3384.320 3538.505 3384.490 3539.175 ;
      LAYER li1 ;
        RECT 3383.500 3538.215 3383.670 3538.505 ;
      LAYER li1 ;
        RECT 3383.840 3538.335 3384.490 3538.505 ;
      LAYER li1 ;
        RECT 3383.670 3538.045 3384.150 3538.165 ;
        RECT 3383.500 3537.835 3384.150 3538.045 ;
        RECT 3383.500 3537.755 3383.670 3537.835 ;
      LAYER li1 ;
        RECT 3384.320 3537.750 3384.490 3538.335 ;
      LAYER li1 ;
        RECT 3384.660 3537.995 3384.830 3540.445 ;
        RECT 3385.420 3540.435 3386.220 3540.515 ;
        RECT 3386.390 3540.395 3387.190 3540.515 ;
      LAYER li1 ;
        RECT 3385.030 3540.015 3386.050 3540.185 ;
      LAYER li1 ;
        RECT 3386.220 3540.055 3386.390 3540.345 ;
      LAYER li1 ;
        RECT 3385.030 3539.345 3385.200 3540.015 ;
      LAYER li1 ;
        RECT 3386.220 3539.845 3387.190 3539.885 ;
        RECT 3385.420 3539.595 3387.190 3539.845 ;
        RECT 3385.420 3539.515 3386.220 3539.595 ;
        RECT 3386.390 3539.555 3387.190 3539.595 ;
      LAYER li1 ;
        RECT 3385.030 3539.175 3386.050 3539.345 ;
        RECT 3385.030 3538.505 3385.200 3539.175 ;
      LAYER li1 ;
        RECT 3386.220 3539.135 3386.390 3539.425 ;
        RECT 3385.420 3538.965 3386.220 3539.005 ;
        RECT 3386.390 3538.965 3387.190 3539.045 ;
        RECT 3385.420 3538.715 3387.190 3538.965 ;
        RECT 3385.420 3538.675 3386.390 3538.715 ;
      LAYER li1 ;
        RECT 3385.030 3538.335 3386.050 3538.505 ;
        RECT 3385.030 3537.750 3385.200 3538.335 ;
      LAYER li1 ;
        RECT 3386.220 3538.215 3386.390 3538.505 ;
        RECT 3385.420 3538.045 3386.220 3538.165 ;
        RECT 3386.390 3538.045 3387.190 3538.125 ;
        RECT 3387.780 3538.115 3387.950 3540.565 ;
        RECT 3388.460 3540.515 3389.110 3540.725 ;
        RECT 3388.460 3540.395 3388.940 3540.515 ;
        RECT 3388.940 3540.055 3389.110 3540.345 ;
        RECT 3388.460 3539.595 3389.110 3539.885 ;
        RECT 3388.460 3539.555 3388.940 3539.595 ;
        RECT 3388.940 3539.135 3389.110 3539.425 ;
        RECT 3388.460 3538.965 3388.940 3539.045 ;
        RECT 3388.460 3538.715 3389.110 3538.965 ;
        RECT 3388.940 3538.675 3389.110 3538.715 ;
        RECT 3388.940 3538.215 3389.110 3538.505 ;
        RECT 3385.420 3537.955 3387.190 3538.045 ;
        RECT 3385.420 3537.835 3386.390 3537.955 ;
        RECT 3386.220 3537.755 3386.390 3537.835 ;
        RECT 3387.410 3537.940 3388.290 3538.115 ;
        RECT 3387.410 3537.785 3387.580 3537.940 ;
      LAYER li1 ;
        RECT 3384.320 3537.665 3385.200 3537.750 ;
      LAYER li1 ;
        RECT 3383.500 3537.325 3383.670 3537.585 ;
      LAYER li1 ;
        RECT 3383.840 3537.495 3386.050 3537.665 ;
      LAYER li1 ;
        RECT 3386.220 3537.325 3386.390 3537.585 ;
        RECT 3386.560 3537.455 3387.580 3537.785 ;
        RECT 3383.500 3537.295 3384.470 3537.325 ;
        RECT 3383.670 3537.125 3384.470 3537.295 ;
        RECT 3383.500 3536.995 3384.470 3537.125 ;
        RECT 3385.070 3537.295 3386.390 3537.325 ;
        RECT 3385.070 3537.125 3386.220 3537.295 ;
        RECT 3386.390 3537.125 3387.190 3537.285 ;
        RECT 3385.070 3537.115 3387.190 3537.125 ;
        RECT 3385.070 3536.995 3386.390 3537.115 ;
        RECT 3383.500 3536.835 3383.670 3536.995 ;
        RECT 3386.220 3536.835 3386.390 3536.995 ;
        RECT 3387.410 3536.945 3387.580 3537.455 ;
        RECT 3383.500 3536.435 3383.670 3536.665 ;
        RECT 3386.220 3536.435 3386.390 3536.665 ;
        RECT 3386.560 3536.615 3387.580 3536.945 ;
      LAYER li1 ;
        RECT 3387.750 3536.660 3387.950 3537.760 ;
      LAYER li1 ;
        RECT 3388.120 3537.705 3388.290 3537.940 ;
        RECT 3388.460 3538.045 3388.940 3538.205 ;
        RECT 3388.460 3537.875 3389.110 3538.045 ;
        RECT 3388.940 3537.755 3389.110 3537.875 ;
        RECT 3388.120 3537.535 3388.765 3537.705 ;
        RECT 3388.120 3536.865 3388.290 3537.535 ;
        RECT 3388.940 3537.365 3389.110 3537.585 ;
        RECT 3388.460 3537.295 3389.110 3537.365 ;
        RECT 3388.460 3537.125 3388.940 3537.295 ;
        RECT 3388.460 3537.035 3389.110 3537.125 ;
        RECT 3388.120 3536.695 3388.770 3536.865 ;
        RECT 3388.940 3536.835 3389.110 3537.035 ;
        RECT 3388.940 3536.435 3389.110 3536.665 ;
        RECT 3383.500 3536.375 3384.395 3536.435 ;
        RECT 3383.670 3536.205 3384.395 3536.375 ;
        RECT 3383.500 3536.145 3384.395 3536.205 ;
        RECT 3385.055 3536.375 3387.555 3536.435 ;
        RECT 3385.055 3536.205 3386.220 3536.375 ;
        RECT 3386.390 3536.205 3387.555 3536.375 ;
        RECT 3385.055 3536.145 3387.555 3536.205 ;
        RECT 3388.215 3536.375 3389.110 3536.435 ;
        RECT 3388.215 3536.205 3388.940 3536.375 ;
        RECT 3388.215 3536.145 3389.110 3536.205 ;
        RECT 3383.500 3536.060 3383.670 3536.145 ;
        RECT 3386.220 3536.060 3386.390 3536.145 ;
        RECT 3388.940 3536.060 3389.110 3536.145 ;
        RECT 198.685 3053.885 198.855 3053.970 ;
        RECT 201.405 3053.885 201.575 3053.970 ;
        RECT 204.125 3053.885 204.295 3053.970 ;
        RECT 198.685 3053.825 199.580 3053.885 ;
        RECT 198.855 3053.655 199.580 3053.825 ;
        RECT 198.685 3053.595 199.580 3053.655 ;
        RECT 200.240 3053.825 202.740 3053.885 ;
        RECT 200.240 3053.655 201.405 3053.825 ;
        RECT 201.575 3053.655 202.740 3053.825 ;
        RECT 200.240 3053.595 202.740 3053.655 ;
        RECT 198.685 3053.365 198.855 3053.595 ;
        RECT 201.405 3053.365 201.575 3053.595 ;
        RECT 198.685 3053.035 198.855 3053.195 ;
        RECT 201.405 3053.035 201.575 3053.195 ;
        RECT 201.745 3053.085 202.765 3053.415 ;
        RECT 198.685 3052.905 199.655 3053.035 ;
        RECT 198.855 3052.735 199.655 3052.905 ;
        RECT 198.685 3052.705 199.655 3052.735 ;
        RECT 200.255 3052.915 201.575 3053.035 ;
        RECT 200.255 3052.905 202.375 3052.915 ;
        RECT 200.255 3052.735 201.405 3052.905 ;
        RECT 201.575 3052.745 202.375 3052.905 ;
        RECT 200.255 3052.705 201.575 3052.735 ;
        RECT 198.685 3052.445 198.855 3052.705 ;
      LAYER li1 ;
        RECT 199.025 3052.365 201.235 3052.535 ;
      LAYER li1 ;
        RECT 201.405 3052.445 201.575 3052.705 ;
        RECT 202.595 3052.575 202.765 3053.085 ;
      LAYER li1 ;
        RECT 199.505 3052.280 200.385 3052.365 ;
      LAYER li1 ;
        RECT 198.685 3052.195 198.855 3052.275 ;
        RECT 198.685 3051.985 199.335 3052.195 ;
        RECT 198.855 3051.865 199.335 3051.985 ;
        RECT 198.685 3051.525 198.855 3051.815 ;
      LAYER li1 ;
        RECT 199.505 3051.695 199.675 3052.280 ;
        RECT 199.025 3051.525 199.675 3051.695 ;
      LAYER li1 ;
        RECT 198.685 3051.065 199.335 3051.355 ;
        RECT 198.855 3051.025 199.335 3051.065 ;
        RECT 198.685 3050.605 198.855 3050.895 ;
      LAYER li1 ;
        RECT 199.505 3050.855 199.675 3051.525 ;
        RECT 199.025 3050.685 199.675 3050.855 ;
      LAYER li1 ;
        RECT 198.855 3050.435 199.335 3050.515 ;
        RECT 198.685 3050.185 199.335 3050.435 ;
        RECT 198.685 3050.145 198.855 3050.185 ;
      LAYER li1 ;
        RECT 199.505 3050.015 199.675 3050.685 ;
      LAYER li1 ;
        RECT 198.685 3049.685 198.855 3049.975 ;
      LAYER li1 ;
        RECT 199.025 3049.845 199.675 3050.015 ;
      LAYER li1 ;
        RECT 198.855 3049.515 199.335 3049.675 ;
        RECT 199.845 3049.585 200.015 3052.035 ;
      LAYER li1 ;
        RECT 200.215 3051.695 200.385 3052.280 ;
      LAYER li1 ;
        RECT 201.405 3052.195 201.575 3052.275 ;
        RECT 201.745 3052.245 202.765 3052.575 ;
      LAYER li1 ;
        RECT 202.935 3052.270 203.135 3053.860 ;
      LAYER li1 ;
        RECT 203.400 3053.825 204.295 3053.885 ;
        RECT 203.400 3053.655 204.125 3053.825 ;
        RECT 203.400 3053.595 204.295 3053.655 ;
        RECT 204.125 3053.365 204.295 3053.595 ;
        RECT 203.305 3053.165 203.955 3053.335 ;
        RECT 203.305 3052.495 203.475 3053.165 ;
        RECT 204.125 3052.995 204.295 3053.195 ;
        RECT 203.645 3052.905 204.295 3052.995 ;
        RECT 203.645 3052.735 204.125 3052.905 ;
        RECT 203.645 3052.665 204.295 3052.735 ;
        RECT 203.305 3052.325 203.950 3052.495 ;
        RECT 204.125 3052.445 204.295 3052.665 ;
        RECT 200.605 3052.075 201.575 3052.195 ;
        RECT 202.595 3052.090 202.765 3052.245 ;
        RECT 203.305 3052.090 203.475 3052.325 ;
        RECT 204.125 3052.155 204.295 3052.275 ;
        RECT 200.605 3051.985 202.375 3052.075 ;
        RECT 200.605 3051.865 201.405 3051.985 ;
        RECT 201.575 3051.905 202.375 3051.985 ;
        RECT 202.595 3051.915 203.475 3052.090 ;
        RECT 203.645 3051.985 204.295 3052.155 ;
      LAYER li1 ;
        RECT 200.215 3051.525 201.235 3051.695 ;
      LAYER li1 ;
        RECT 201.405 3051.525 201.575 3051.815 ;
      LAYER li1 ;
        RECT 200.215 3050.855 200.385 3051.525 ;
        RECT 201.745 3051.485 202.765 3051.655 ;
      LAYER li1 ;
        RECT 200.605 3051.315 201.575 3051.355 ;
        RECT 200.605 3051.065 202.375 3051.315 ;
        RECT 200.605 3051.025 201.405 3051.065 ;
        RECT 201.575 3050.985 202.375 3051.065 ;
      LAYER li1 ;
        RECT 200.215 3050.685 201.235 3050.855 ;
        RECT 200.215 3050.015 200.385 3050.685 ;
      LAYER li1 ;
        RECT 201.405 3050.605 201.575 3050.895 ;
      LAYER li1 ;
        RECT 202.595 3050.815 202.765 3051.485 ;
        RECT 201.745 3050.645 202.765 3050.815 ;
      LAYER li1 ;
        RECT 200.605 3050.435 201.405 3050.515 ;
        RECT 201.575 3050.435 202.375 3050.475 ;
        RECT 200.605 3050.185 202.375 3050.435 ;
        RECT 201.405 3050.145 202.375 3050.185 ;
      LAYER li1 ;
        RECT 200.215 3049.845 201.235 3050.015 ;
        RECT 202.595 3049.975 202.765 3050.645 ;
      LAYER li1 ;
        RECT 201.405 3049.685 201.575 3049.975 ;
      LAYER li1 ;
        RECT 201.745 3049.805 202.765 3049.975 ;
      LAYER li1 ;
        RECT 198.685 3049.345 199.335 3049.515 ;
        RECT 199.505 3049.410 200.385 3049.585 ;
        RECT 200.605 3049.515 201.405 3049.595 ;
        RECT 201.575 3049.515 202.375 3049.635 ;
        RECT 200.605 3049.425 202.375 3049.515 ;
        RECT 198.685 3049.225 198.855 3049.345 ;
        RECT 199.505 3049.175 199.675 3049.410 ;
        RECT 200.215 3049.255 200.385 3049.410 ;
        RECT 201.405 3049.305 202.375 3049.425 ;
        RECT 198.685 3048.835 198.855 3049.055 ;
        RECT 199.030 3049.005 199.675 3049.175 ;
        RECT 198.685 3048.765 199.335 3048.835 ;
        RECT 198.855 3048.595 199.335 3048.765 ;
        RECT 198.685 3048.505 199.335 3048.595 ;
        RECT 198.685 3048.305 198.855 3048.505 ;
        RECT 199.505 3048.335 199.675 3049.005 ;
        RECT 199.025 3048.165 199.675 3048.335 ;
        RECT 198.685 3047.905 198.855 3048.135 ;
      LAYER li1 ;
        RECT 199.845 3048.130 200.045 3049.230 ;
      LAYER li1 ;
        RECT 200.215 3048.925 201.235 3049.255 ;
        RECT 201.405 3049.225 201.575 3049.305 ;
      LAYER li1 ;
        RECT 202.595 3049.220 202.765 3049.805 ;
      LAYER li1 ;
        RECT 202.965 3049.465 203.135 3051.915 ;
        RECT 203.645 3051.825 204.125 3051.985 ;
      LAYER li1 ;
        RECT 203.305 3051.485 203.955 3051.655 ;
      LAYER li1 ;
        RECT 204.125 3051.525 204.295 3051.815 ;
      LAYER li1 ;
        RECT 203.305 3050.815 203.475 3051.485 ;
      LAYER li1 ;
        RECT 204.125 3051.315 204.295 3051.355 ;
        RECT 203.645 3051.065 204.295 3051.315 ;
        RECT 203.645 3050.985 204.125 3051.065 ;
      LAYER li1 ;
        RECT 203.305 3050.645 203.955 3050.815 ;
        RECT 203.305 3049.975 203.475 3050.645 ;
      LAYER li1 ;
        RECT 204.125 3050.605 204.295 3050.895 ;
        RECT 203.645 3050.435 204.125 3050.475 ;
        RECT 203.645 3050.145 204.295 3050.435 ;
      LAYER li1 ;
        RECT 203.305 3049.805 203.955 3049.975 ;
        RECT 203.305 3049.220 203.475 3049.805 ;
      LAYER li1 ;
        RECT 204.125 3049.685 204.295 3049.975 ;
        RECT 203.645 3049.515 204.125 3049.635 ;
        RECT 203.645 3049.305 204.295 3049.515 ;
        RECT 204.125 3049.225 204.295 3049.305 ;
      LAYER li1 ;
        RECT 202.595 3049.135 203.475 3049.220 ;
      LAYER li1 ;
        RECT 200.215 3048.415 200.385 3048.925 ;
        RECT 201.405 3048.795 201.575 3049.055 ;
      LAYER li1 ;
        RECT 201.745 3048.965 203.955 3049.135 ;
      LAYER li1 ;
        RECT 204.125 3048.795 204.295 3049.055 ;
        RECT 201.405 3048.765 202.725 3048.795 ;
        RECT 200.605 3048.595 201.405 3048.755 ;
        RECT 201.575 3048.595 202.725 3048.765 ;
        RECT 200.605 3048.585 202.725 3048.595 ;
        RECT 201.405 3048.465 202.725 3048.585 ;
        RECT 203.325 3048.765 204.295 3048.795 ;
        RECT 203.325 3048.595 204.125 3048.765 ;
        RECT 203.325 3048.465 204.295 3048.595 ;
        RECT 200.215 3048.085 201.235 3048.415 ;
        RECT 201.405 3048.305 201.575 3048.465 ;
        RECT 204.125 3048.305 204.295 3048.465 ;
        RECT 201.405 3047.905 201.575 3048.135 ;
        RECT 204.125 3047.905 204.295 3048.135 ;
        RECT 198.685 3047.845 199.580 3047.905 ;
        RECT 198.855 3047.675 199.580 3047.845 ;
        RECT 198.685 3047.615 199.580 3047.675 ;
        RECT 200.240 3047.845 202.740 3047.905 ;
        RECT 200.240 3047.675 201.405 3047.845 ;
        RECT 201.575 3047.675 202.740 3047.845 ;
        RECT 200.240 3047.615 202.740 3047.675 ;
        RECT 198.685 3047.385 198.855 3047.615 ;
        RECT 201.405 3047.385 201.575 3047.615 ;
        RECT 198.685 3047.055 198.855 3047.215 ;
        RECT 201.405 3047.055 201.575 3047.215 ;
        RECT 201.745 3047.105 202.765 3047.435 ;
        RECT 198.685 3046.925 199.655 3047.055 ;
        RECT 198.855 3046.755 199.655 3046.925 ;
        RECT 198.685 3046.725 199.655 3046.755 ;
        RECT 200.255 3046.935 201.575 3047.055 ;
        RECT 200.255 3046.925 202.375 3046.935 ;
        RECT 200.255 3046.755 201.405 3046.925 ;
        RECT 201.575 3046.765 202.375 3046.925 ;
        RECT 200.255 3046.725 201.575 3046.755 ;
        RECT 198.685 3046.465 198.855 3046.725 ;
      LAYER li1 ;
        RECT 199.025 3046.385 201.235 3046.555 ;
      LAYER li1 ;
        RECT 201.405 3046.465 201.575 3046.725 ;
        RECT 202.595 3046.595 202.765 3047.105 ;
      LAYER li1 ;
        RECT 199.505 3046.300 200.385 3046.385 ;
      LAYER li1 ;
        RECT 198.685 3046.215 198.855 3046.295 ;
        RECT 198.685 3046.005 199.335 3046.215 ;
        RECT 198.855 3045.885 199.335 3046.005 ;
        RECT 198.685 3045.545 198.855 3045.835 ;
      LAYER li1 ;
        RECT 199.505 3045.715 199.675 3046.300 ;
        RECT 199.025 3045.545 199.675 3045.715 ;
      LAYER li1 ;
        RECT 198.685 3045.085 199.335 3045.375 ;
        RECT 198.855 3045.045 199.335 3045.085 ;
        RECT 198.685 3044.625 198.855 3044.915 ;
      LAYER li1 ;
        RECT 199.505 3044.875 199.675 3045.545 ;
        RECT 199.025 3044.705 199.675 3044.875 ;
      LAYER li1 ;
        RECT 198.855 3044.455 199.335 3044.535 ;
        RECT 198.685 3044.205 199.335 3044.455 ;
        RECT 198.685 3044.165 198.855 3044.205 ;
      LAYER li1 ;
        RECT 199.505 3044.035 199.675 3044.705 ;
      LAYER li1 ;
        RECT 198.685 3043.705 198.855 3043.995 ;
      LAYER li1 ;
        RECT 199.025 3043.865 199.675 3044.035 ;
      LAYER li1 ;
        RECT 198.855 3043.535 199.335 3043.695 ;
        RECT 199.845 3043.605 200.015 3046.055 ;
      LAYER li1 ;
        RECT 200.215 3045.715 200.385 3046.300 ;
      LAYER li1 ;
        RECT 201.405 3046.215 201.575 3046.295 ;
        RECT 201.745 3046.265 202.765 3046.595 ;
      LAYER li1 ;
        RECT 202.935 3046.290 203.135 3047.880 ;
      LAYER li1 ;
        RECT 203.400 3047.845 204.295 3047.905 ;
        RECT 203.400 3047.675 204.125 3047.845 ;
        RECT 203.400 3047.615 204.295 3047.675 ;
        RECT 204.125 3047.385 204.295 3047.615 ;
        RECT 203.305 3047.185 203.955 3047.355 ;
        RECT 203.305 3046.515 203.475 3047.185 ;
        RECT 204.125 3047.015 204.295 3047.215 ;
        RECT 203.645 3046.925 204.295 3047.015 ;
        RECT 203.645 3046.755 204.125 3046.925 ;
        RECT 203.645 3046.685 204.295 3046.755 ;
        RECT 203.305 3046.345 203.950 3046.515 ;
        RECT 204.125 3046.465 204.295 3046.685 ;
        RECT 200.605 3046.095 201.575 3046.215 ;
        RECT 202.595 3046.110 202.765 3046.265 ;
        RECT 203.305 3046.110 203.475 3046.345 ;
        RECT 204.125 3046.175 204.295 3046.295 ;
        RECT 200.605 3046.005 202.375 3046.095 ;
        RECT 200.605 3045.885 201.405 3046.005 ;
        RECT 201.575 3045.925 202.375 3046.005 ;
        RECT 202.595 3045.935 203.475 3046.110 ;
        RECT 203.645 3046.005 204.295 3046.175 ;
      LAYER li1 ;
        RECT 200.215 3045.545 201.235 3045.715 ;
      LAYER li1 ;
        RECT 201.405 3045.545 201.575 3045.835 ;
      LAYER li1 ;
        RECT 200.215 3044.875 200.385 3045.545 ;
        RECT 201.745 3045.505 202.765 3045.675 ;
      LAYER li1 ;
        RECT 200.605 3045.335 201.575 3045.375 ;
        RECT 200.605 3045.085 202.375 3045.335 ;
        RECT 200.605 3045.045 201.405 3045.085 ;
        RECT 201.575 3045.005 202.375 3045.085 ;
      LAYER li1 ;
        RECT 200.215 3044.705 201.235 3044.875 ;
        RECT 200.215 3044.035 200.385 3044.705 ;
      LAYER li1 ;
        RECT 201.405 3044.625 201.575 3044.915 ;
      LAYER li1 ;
        RECT 202.595 3044.835 202.765 3045.505 ;
        RECT 201.745 3044.665 202.765 3044.835 ;
      LAYER li1 ;
        RECT 200.605 3044.455 201.405 3044.535 ;
        RECT 201.575 3044.455 202.375 3044.495 ;
        RECT 200.605 3044.205 202.375 3044.455 ;
        RECT 201.405 3044.165 202.375 3044.205 ;
      LAYER li1 ;
        RECT 200.215 3043.865 201.235 3044.035 ;
        RECT 202.595 3043.995 202.765 3044.665 ;
      LAYER li1 ;
        RECT 201.405 3043.705 201.575 3043.995 ;
      LAYER li1 ;
        RECT 201.745 3043.825 202.765 3043.995 ;
      LAYER li1 ;
        RECT 198.685 3043.365 199.335 3043.535 ;
        RECT 199.505 3043.430 200.385 3043.605 ;
        RECT 200.605 3043.535 201.405 3043.615 ;
        RECT 201.575 3043.535 202.375 3043.655 ;
        RECT 200.605 3043.445 202.375 3043.535 ;
        RECT 198.685 3043.245 198.855 3043.365 ;
        RECT 199.505 3043.195 199.675 3043.430 ;
        RECT 200.215 3043.275 200.385 3043.430 ;
        RECT 201.405 3043.325 202.375 3043.445 ;
        RECT 198.685 3042.855 198.855 3043.075 ;
        RECT 199.030 3043.025 199.675 3043.195 ;
        RECT 198.685 3042.785 199.335 3042.855 ;
        RECT 198.855 3042.615 199.335 3042.785 ;
        RECT 198.685 3042.525 199.335 3042.615 ;
        RECT 198.685 3042.325 198.855 3042.525 ;
        RECT 199.505 3042.355 199.675 3043.025 ;
        RECT 199.025 3042.185 199.675 3042.355 ;
        RECT 198.685 3041.925 198.855 3042.155 ;
      LAYER li1 ;
        RECT 199.845 3042.150 200.045 3043.250 ;
      LAYER li1 ;
        RECT 200.215 3042.945 201.235 3043.275 ;
        RECT 201.405 3043.245 201.575 3043.325 ;
      LAYER li1 ;
        RECT 202.595 3043.240 202.765 3043.825 ;
      LAYER li1 ;
        RECT 202.965 3043.485 203.135 3045.935 ;
        RECT 203.645 3045.845 204.125 3046.005 ;
      LAYER li1 ;
        RECT 203.305 3045.505 203.955 3045.675 ;
      LAYER li1 ;
        RECT 204.125 3045.545 204.295 3045.835 ;
      LAYER li1 ;
        RECT 203.305 3044.835 203.475 3045.505 ;
      LAYER li1 ;
        RECT 204.125 3045.335 204.295 3045.375 ;
        RECT 203.645 3045.085 204.295 3045.335 ;
        RECT 203.645 3045.005 204.125 3045.085 ;
      LAYER li1 ;
        RECT 203.305 3044.665 203.955 3044.835 ;
        RECT 203.305 3043.995 203.475 3044.665 ;
      LAYER li1 ;
        RECT 204.125 3044.625 204.295 3044.915 ;
        RECT 203.645 3044.455 204.125 3044.495 ;
        RECT 203.645 3044.165 204.295 3044.455 ;
      LAYER li1 ;
        RECT 203.305 3043.825 203.955 3043.995 ;
        RECT 203.305 3043.240 203.475 3043.825 ;
      LAYER li1 ;
        RECT 204.125 3043.705 204.295 3043.995 ;
        RECT 203.645 3043.535 204.125 3043.655 ;
        RECT 203.645 3043.325 204.295 3043.535 ;
        RECT 204.125 3043.245 204.295 3043.325 ;
      LAYER li1 ;
        RECT 202.595 3043.155 203.475 3043.240 ;
      LAYER li1 ;
        RECT 200.215 3042.435 200.385 3042.945 ;
        RECT 201.405 3042.815 201.575 3043.075 ;
      LAYER li1 ;
        RECT 201.745 3042.985 203.955 3043.155 ;
      LAYER li1 ;
        RECT 204.125 3042.815 204.295 3043.075 ;
        RECT 201.405 3042.785 202.725 3042.815 ;
        RECT 200.605 3042.615 201.405 3042.775 ;
        RECT 201.575 3042.615 202.725 3042.785 ;
        RECT 200.605 3042.605 202.725 3042.615 ;
        RECT 201.405 3042.485 202.725 3042.605 ;
        RECT 203.325 3042.785 204.295 3042.815 ;
        RECT 203.325 3042.615 204.125 3042.785 ;
        RECT 203.325 3042.485 204.295 3042.615 ;
        RECT 200.215 3042.105 201.235 3042.435 ;
        RECT 201.405 3042.325 201.575 3042.485 ;
        RECT 204.125 3042.325 204.295 3042.485 ;
        RECT 201.405 3041.925 201.575 3042.155 ;
        RECT 204.125 3041.925 204.295 3042.155 ;
        RECT 198.685 3041.865 199.580 3041.925 ;
        RECT 198.855 3041.695 199.580 3041.865 ;
        RECT 198.685 3041.635 199.580 3041.695 ;
        RECT 200.240 3041.865 202.740 3041.925 ;
        RECT 200.240 3041.695 201.405 3041.865 ;
        RECT 201.575 3041.695 202.740 3041.865 ;
        RECT 200.240 3041.635 202.740 3041.695 ;
        RECT 198.685 3041.405 198.855 3041.635 ;
        RECT 201.405 3041.405 201.575 3041.635 ;
        RECT 198.685 3041.075 198.855 3041.235 ;
        RECT 201.405 3041.075 201.575 3041.235 ;
        RECT 201.745 3041.125 202.765 3041.455 ;
        RECT 198.685 3040.945 199.655 3041.075 ;
        RECT 198.855 3040.775 199.655 3040.945 ;
        RECT 198.685 3040.745 199.655 3040.775 ;
        RECT 200.255 3040.955 201.575 3041.075 ;
        RECT 200.255 3040.945 202.375 3040.955 ;
        RECT 200.255 3040.775 201.405 3040.945 ;
        RECT 201.575 3040.785 202.375 3040.945 ;
        RECT 200.255 3040.745 201.575 3040.775 ;
        RECT 198.685 3040.485 198.855 3040.745 ;
      LAYER li1 ;
        RECT 199.025 3040.405 201.235 3040.575 ;
      LAYER li1 ;
        RECT 201.405 3040.485 201.575 3040.745 ;
        RECT 202.595 3040.615 202.765 3041.125 ;
      LAYER li1 ;
        RECT 199.505 3040.320 200.385 3040.405 ;
      LAYER li1 ;
        RECT 198.685 3040.235 198.855 3040.315 ;
        RECT 198.685 3040.025 199.335 3040.235 ;
        RECT 198.855 3039.905 199.335 3040.025 ;
        RECT 198.685 3039.565 198.855 3039.855 ;
      LAYER li1 ;
        RECT 199.505 3039.735 199.675 3040.320 ;
        RECT 199.025 3039.565 199.675 3039.735 ;
      LAYER li1 ;
        RECT 198.685 3039.105 199.335 3039.395 ;
        RECT 198.855 3039.065 199.335 3039.105 ;
        RECT 198.685 3038.645 198.855 3038.935 ;
      LAYER li1 ;
        RECT 199.505 3038.895 199.675 3039.565 ;
        RECT 199.025 3038.725 199.675 3038.895 ;
      LAYER li1 ;
        RECT 198.855 3038.475 199.335 3038.555 ;
        RECT 198.685 3038.225 199.335 3038.475 ;
        RECT 198.685 3038.185 198.855 3038.225 ;
      LAYER li1 ;
        RECT 199.505 3038.055 199.675 3038.725 ;
      LAYER li1 ;
        RECT 198.685 3037.725 198.855 3038.015 ;
      LAYER li1 ;
        RECT 199.025 3037.885 199.675 3038.055 ;
      LAYER li1 ;
        RECT 198.855 3037.555 199.335 3037.715 ;
        RECT 199.845 3037.625 200.015 3040.075 ;
      LAYER li1 ;
        RECT 200.215 3039.735 200.385 3040.320 ;
      LAYER li1 ;
        RECT 201.405 3040.235 201.575 3040.315 ;
        RECT 201.745 3040.285 202.765 3040.615 ;
      LAYER li1 ;
        RECT 202.935 3040.310 203.135 3041.900 ;
      LAYER li1 ;
        RECT 203.400 3041.865 204.295 3041.925 ;
        RECT 203.400 3041.695 204.125 3041.865 ;
        RECT 203.400 3041.635 204.295 3041.695 ;
        RECT 204.125 3041.405 204.295 3041.635 ;
        RECT 203.305 3041.205 203.955 3041.375 ;
        RECT 203.305 3040.535 203.475 3041.205 ;
        RECT 204.125 3041.035 204.295 3041.235 ;
        RECT 203.645 3040.945 204.295 3041.035 ;
        RECT 203.645 3040.775 204.125 3040.945 ;
        RECT 203.645 3040.705 204.295 3040.775 ;
        RECT 203.305 3040.365 203.950 3040.535 ;
        RECT 204.125 3040.485 204.295 3040.705 ;
        RECT 200.605 3040.115 201.575 3040.235 ;
        RECT 202.595 3040.130 202.765 3040.285 ;
        RECT 203.305 3040.130 203.475 3040.365 ;
        RECT 204.125 3040.195 204.295 3040.315 ;
        RECT 200.605 3040.025 202.375 3040.115 ;
        RECT 200.605 3039.905 201.405 3040.025 ;
        RECT 201.575 3039.945 202.375 3040.025 ;
        RECT 202.595 3039.955 203.475 3040.130 ;
        RECT 203.645 3040.025 204.295 3040.195 ;
      LAYER li1 ;
        RECT 200.215 3039.565 201.235 3039.735 ;
      LAYER li1 ;
        RECT 201.405 3039.565 201.575 3039.855 ;
      LAYER li1 ;
        RECT 200.215 3038.895 200.385 3039.565 ;
        RECT 201.745 3039.525 202.765 3039.695 ;
      LAYER li1 ;
        RECT 200.605 3039.355 201.575 3039.395 ;
        RECT 200.605 3039.105 202.375 3039.355 ;
        RECT 200.605 3039.065 201.405 3039.105 ;
        RECT 201.575 3039.025 202.375 3039.105 ;
      LAYER li1 ;
        RECT 200.215 3038.725 201.235 3038.895 ;
        RECT 200.215 3038.055 200.385 3038.725 ;
      LAYER li1 ;
        RECT 201.405 3038.645 201.575 3038.935 ;
      LAYER li1 ;
        RECT 202.595 3038.855 202.765 3039.525 ;
        RECT 201.745 3038.685 202.765 3038.855 ;
      LAYER li1 ;
        RECT 200.605 3038.475 201.405 3038.555 ;
        RECT 201.575 3038.475 202.375 3038.515 ;
        RECT 200.605 3038.225 202.375 3038.475 ;
        RECT 201.405 3038.185 202.375 3038.225 ;
      LAYER li1 ;
        RECT 200.215 3037.885 201.235 3038.055 ;
        RECT 202.595 3038.015 202.765 3038.685 ;
      LAYER li1 ;
        RECT 201.405 3037.725 201.575 3038.015 ;
      LAYER li1 ;
        RECT 201.745 3037.845 202.765 3038.015 ;
      LAYER li1 ;
        RECT 198.685 3037.385 199.335 3037.555 ;
        RECT 199.505 3037.450 200.385 3037.625 ;
        RECT 200.605 3037.555 201.405 3037.635 ;
        RECT 201.575 3037.555 202.375 3037.675 ;
        RECT 200.605 3037.465 202.375 3037.555 ;
        RECT 198.685 3037.265 198.855 3037.385 ;
        RECT 199.505 3037.215 199.675 3037.450 ;
        RECT 200.215 3037.295 200.385 3037.450 ;
        RECT 201.405 3037.345 202.375 3037.465 ;
        RECT 198.685 3036.875 198.855 3037.095 ;
        RECT 199.030 3037.045 199.675 3037.215 ;
        RECT 198.685 3036.805 199.335 3036.875 ;
        RECT 198.855 3036.635 199.335 3036.805 ;
        RECT 198.685 3036.545 199.335 3036.635 ;
        RECT 198.685 3036.345 198.855 3036.545 ;
        RECT 199.505 3036.375 199.675 3037.045 ;
        RECT 199.025 3036.205 199.675 3036.375 ;
        RECT 198.685 3035.945 198.855 3036.175 ;
      LAYER li1 ;
        RECT 199.845 3036.170 200.045 3037.270 ;
      LAYER li1 ;
        RECT 200.215 3036.965 201.235 3037.295 ;
        RECT 201.405 3037.265 201.575 3037.345 ;
      LAYER li1 ;
        RECT 202.595 3037.260 202.765 3037.845 ;
      LAYER li1 ;
        RECT 202.965 3037.505 203.135 3039.955 ;
        RECT 203.645 3039.865 204.125 3040.025 ;
      LAYER li1 ;
        RECT 203.305 3039.525 203.955 3039.695 ;
      LAYER li1 ;
        RECT 204.125 3039.565 204.295 3039.855 ;
      LAYER li1 ;
        RECT 203.305 3038.855 203.475 3039.525 ;
      LAYER li1 ;
        RECT 204.125 3039.355 204.295 3039.395 ;
        RECT 203.645 3039.105 204.295 3039.355 ;
        RECT 203.645 3039.025 204.125 3039.105 ;
      LAYER li1 ;
        RECT 203.305 3038.685 203.955 3038.855 ;
        RECT 203.305 3038.015 203.475 3038.685 ;
      LAYER li1 ;
        RECT 204.125 3038.645 204.295 3038.935 ;
        RECT 203.645 3038.475 204.125 3038.515 ;
        RECT 203.645 3038.185 204.295 3038.475 ;
      LAYER li1 ;
        RECT 203.305 3037.845 203.955 3038.015 ;
        RECT 203.305 3037.260 203.475 3037.845 ;
      LAYER li1 ;
        RECT 204.125 3037.725 204.295 3038.015 ;
        RECT 203.645 3037.555 204.125 3037.675 ;
        RECT 203.645 3037.345 204.295 3037.555 ;
        RECT 204.125 3037.265 204.295 3037.345 ;
      LAYER li1 ;
        RECT 202.595 3037.175 203.475 3037.260 ;
      LAYER li1 ;
        RECT 200.215 3036.455 200.385 3036.965 ;
        RECT 201.405 3036.835 201.575 3037.095 ;
      LAYER li1 ;
        RECT 201.745 3037.005 203.955 3037.175 ;
      LAYER li1 ;
        RECT 204.125 3036.835 204.295 3037.095 ;
        RECT 201.405 3036.805 202.725 3036.835 ;
        RECT 200.605 3036.635 201.405 3036.795 ;
        RECT 201.575 3036.635 202.725 3036.805 ;
        RECT 200.605 3036.625 202.725 3036.635 ;
        RECT 201.405 3036.505 202.725 3036.625 ;
        RECT 203.325 3036.805 204.295 3036.835 ;
        RECT 203.325 3036.635 204.125 3036.805 ;
        RECT 203.325 3036.505 204.295 3036.635 ;
        RECT 200.215 3036.125 201.235 3036.455 ;
        RECT 201.405 3036.345 201.575 3036.505 ;
        RECT 204.125 3036.345 204.295 3036.505 ;
        RECT 201.405 3035.945 201.575 3036.175 ;
        RECT 204.125 3035.945 204.295 3036.175 ;
        RECT 198.685 3035.885 199.580 3035.945 ;
        RECT 198.855 3035.715 199.580 3035.885 ;
        RECT 198.685 3035.655 199.580 3035.715 ;
        RECT 200.240 3035.885 202.740 3035.945 ;
        RECT 200.240 3035.715 201.405 3035.885 ;
        RECT 201.575 3035.715 202.740 3035.885 ;
        RECT 200.240 3035.655 202.740 3035.715 ;
        RECT 198.685 3035.425 198.855 3035.655 ;
        RECT 201.405 3035.425 201.575 3035.655 ;
        RECT 198.685 3035.095 198.855 3035.255 ;
        RECT 201.405 3035.095 201.575 3035.255 ;
        RECT 201.745 3035.145 202.765 3035.475 ;
        RECT 198.685 3034.965 199.655 3035.095 ;
        RECT 198.855 3034.795 199.655 3034.965 ;
        RECT 198.685 3034.765 199.655 3034.795 ;
        RECT 200.255 3034.975 201.575 3035.095 ;
        RECT 200.255 3034.965 202.375 3034.975 ;
        RECT 200.255 3034.795 201.405 3034.965 ;
        RECT 201.575 3034.805 202.375 3034.965 ;
        RECT 200.255 3034.765 201.575 3034.795 ;
        RECT 198.685 3034.505 198.855 3034.765 ;
      LAYER li1 ;
        RECT 199.025 3034.425 201.235 3034.595 ;
      LAYER li1 ;
        RECT 201.405 3034.505 201.575 3034.765 ;
        RECT 202.595 3034.635 202.765 3035.145 ;
      LAYER li1 ;
        RECT 199.505 3034.340 200.385 3034.425 ;
      LAYER li1 ;
        RECT 198.685 3034.255 198.855 3034.335 ;
        RECT 198.685 3034.045 199.335 3034.255 ;
        RECT 198.855 3033.925 199.335 3034.045 ;
        RECT 198.685 3033.585 198.855 3033.875 ;
      LAYER li1 ;
        RECT 199.505 3033.755 199.675 3034.340 ;
        RECT 199.025 3033.585 199.675 3033.755 ;
      LAYER li1 ;
        RECT 198.685 3033.125 199.335 3033.415 ;
        RECT 198.855 3033.085 199.335 3033.125 ;
        RECT 198.685 3032.665 198.855 3032.955 ;
      LAYER li1 ;
        RECT 199.505 3032.915 199.675 3033.585 ;
        RECT 199.025 3032.745 199.675 3032.915 ;
      LAYER li1 ;
        RECT 198.855 3032.495 199.335 3032.575 ;
        RECT 198.685 3032.245 199.335 3032.495 ;
        RECT 198.685 3032.205 198.855 3032.245 ;
      LAYER li1 ;
        RECT 199.505 3032.075 199.675 3032.745 ;
      LAYER li1 ;
        RECT 198.685 3031.745 198.855 3032.035 ;
      LAYER li1 ;
        RECT 199.025 3031.905 199.675 3032.075 ;
      LAYER li1 ;
        RECT 198.855 3031.575 199.335 3031.735 ;
        RECT 199.845 3031.645 200.015 3034.095 ;
      LAYER li1 ;
        RECT 200.215 3033.755 200.385 3034.340 ;
      LAYER li1 ;
        RECT 201.405 3034.255 201.575 3034.335 ;
        RECT 201.745 3034.305 202.765 3034.635 ;
      LAYER li1 ;
        RECT 202.935 3034.330 203.135 3035.920 ;
      LAYER li1 ;
        RECT 203.400 3035.885 204.295 3035.945 ;
        RECT 203.400 3035.715 204.125 3035.885 ;
        RECT 203.400 3035.655 204.295 3035.715 ;
        RECT 204.125 3035.425 204.295 3035.655 ;
        RECT 203.305 3035.225 203.955 3035.395 ;
        RECT 203.305 3034.555 203.475 3035.225 ;
        RECT 204.125 3035.055 204.295 3035.255 ;
        RECT 203.645 3034.965 204.295 3035.055 ;
        RECT 203.645 3034.795 204.125 3034.965 ;
        RECT 203.645 3034.725 204.295 3034.795 ;
        RECT 203.305 3034.385 203.950 3034.555 ;
        RECT 204.125 3034.505 204.295 3034.725 ;
        RECT 200.605 3034.135 201.575 3034.255 ;
        RECT 202.595 3034.150 202.765 3034.305 ;
        RECT 203.305 3034.150 203.475 3034.385 ;
        RECT 204.125 3034.215 204.295 3034.335 ;
        RECT 200.605 3034.045 202.375 3034.135 ;
        RECT 200.605 3033.925 201.405 3034.045 ;
        RECT 201.575 3033.965 202.375 3034.045 ;
        RECT 202.595 3033.975 203.475 3034.150 ;
        RECT 203.645 3034.045 204.295 3034.215 ;
      LAYER li1 ;
        RECT 200.215 3033.585 201.235 3033.755 ;
      LAYER li1 ;
        RECT 201.405 3033.585 201.575 3033.875 ;
      LAYER li1 ;
        RECT 200.215 3032.915 200.385 3033.585 ;
        RECT 201.745 3033.545 202.765 3033.715 ;
      LAYER li1 ;
        RECT 200.605 3033.375 201.575 3033.415 ;
        RECT 200.605 3033.125 202.375 3033.375 ;
        RECT 200.605 3033.085 201.405 3033.125 ;
        RECT 201.575 3033.045 202.375 3033.125 ;
      LAYER li1 ;
        RECT 200.215 3032.745 201.235 3032.915 ;
        RECT 200.215 3032.075 200.385 3032.745 ;
      LAYER li1 ;
        RECT 201.405 3032.665 201.575 3032.955 ;
      LAYER li1 ;
        RECT 202.595 3032.875 202.765 3033.545 ;
        RECT 201.745 3032.705 202.765 3032.875 ;
      LAYER li1 ;
        RECT 200.605 3032.495 201.405 3032.575 ;
        RECT 201.575 3032.495 202.375 3032.535 ;
        RECT 200.605 3032.245 202.375 3032.495 ;
        RECT 201.405 3032.205 202.375 3032.245 ;
      LAYER li1 ;
        RECT 200.215 3031.905 201.235 3032.075 ;
        RECT 202.595 3032.035 202.765 3032.705 ;
      LAYER li1 ;
        RECT 201.405 3031.745 201.575 3032.035 ;
      LAYER li1 ;
        RECT 201.745 3031.865 202.765 3032.035 ;
      LAYER li1 ;
        RECT 198.685 3031.405 199.335 3031.575 ;
        RECT 199.505 3031.470 200.385 3031.645 ;
        RECT 200.605 3031.575 201.405 3031.655 ;
        RECT 201.575 3031.575 202.375 3031.695 ;
        RECT 200.605 3031.485 202.375 3031.575 ;
        RECT 198.685 3031.285 198.855 3031.405 ;
        RECT 199.505 3031.235 199.675 3031.470 ;
        RECT 200.215 3031.315 200.385 3031.470 ;
        RECT 201.405 3031.365 202.375 3031.485 ;
        RECT 198.685 3030.895 198.855 3031.115 ;
        RECT 199.030 3031.065 199.675 3031.235 ;
        RECT 198.685 3030.825 199.335 3030.895 ;
        RECT 198.855 3030.655 199.335 3030.825 ;
        RECT 198.685 3030.565 199.335 3030.655 ;
        RECT 198.685 3030.365 198.855 3030.565 ;
        RECT 199.505 3030.395 199.675 3031.065 ;
        RECT 199.025 3030.225 199.675 3030.395 ;
        RECT 198.685 3029.965 198.855 3030.195 ;
      LAYER li1 ;
        RECT 199.845 3030.190 200.045 3031.290 ;
      LAYER li1 ;
        RECT 200.215 3030.985 201.235 3031.315 ;
        RECT 201.405 3031.285 201.575 3031.365 ;
      LAYER li1 ;
        RECT 202.595 3031.280 202.765 3031.865 ;
      LAYER li1 ;
        RECT 202.965 3031.525 203.135 3033.975 ;
        RECT 203.645 3033.885 204.125 3034.045 ;
      LAYER li1 ;
        RECT 203.305 3033.545 203.955 3033.715 ;
      LAYER li1 ;
        RECT 204.125 3033.585 204.295 3033.875 ;
      LAYER li1 ;
        RECT 203.305 3032.875 203.475 3033.545 ;
      LAYER li1 ;
        RECT 204.125 3033.375 204.295 3033.415 ;
        RECT 203.645 3033.125 204.295 3033.375 ;
        RECT 203.645 3033.045 204.125 3033.125 ;
      LAYER li1 ;
        RECT 203.305 3032.705 203.955 3032.875 ;
        RECT 203.305 3032.035 203.475 3032.705 ;
      LAYER li1 ;
        RECT 204.125 3032.665 204.295 3032.955 ;
        RECT 203.645 3032.495 204.125 3032.535 ;
        RECT 203.645 3032.205 204.295 3032.495 ;
      LAYER li1 ;
        RECT 203.305 3031.865 203.955 3032.035 ;
        RECT 203.305 3031.280 203.475 3031.865 ;
      LAYER li1 ;
        RECT 204.125 3031.745 204.295 3032.035 ;
        RECT 203.645 3031.575 204.125 3031.695 ;
        RECT 203.645 3031.365 204.295 3031.575 ;
        RECT 204.125 3031.285 204.295 3031.365 ;
      LAYER li1 ;
        RECT 202.595 3031.195 203.475 3031.280 ;
      LAYER li1 ;
        RECT 200.215 3030.475 200.385 3030.985 ;
        RECT 201.405 3030.855 201.575 3031.115 ;
      LAYER li1 ;
        RECT 201.745 3031.025 203.955 3031.195 ;
      LAYER li1 ;
        RECT 204.125 3030.855 204.295 3031.115 ;
        RECT 201.405 3030.825 202.725 3030.855 ;
        RECT 200.605 3030.655 201.405 3030.815 ;
        RECT 201.575 3030.655 202.725 3030.825 ;
        RECT 200.605 3030.645 202.725 3030.655 ;
        RECT 201.405 3030.525 202.725 3030.645 ;
        RECT 203.325 3030.825 204.295 3030.855 ;
        RECT 203.325 3030.655 204.125 3030.825 ;
        RECT 203.325 3030.525 204.295 3030.655 ;
        RECT 200.215 3030.145 201.235 3030.475 ;
        RECT 201.405 3030.365 201.575 3030.525 ;
        RECT 204.125 3030.365 204.295 3030.525 ;
        RECT 201.405 3029.965 201.575 3030.195 ;
        RECT 204.125 3029.965 204.295 3030.195 ;
        RECT 198.685 3029.905 199.580 3029.965 ;
        RECT 198.855 3029.735 199.580 3029.905 ;
        RECT 198.685 3029.675 199.580 3029.735 ;
        RECT 200.240 3029.905 202.740 3029.965 ;
        RECT 200.240 3029.735 201.405 3029.905 ;
        RECT 201.575 3029.735 202.740 3029.905 ;
        RECT 200.240 3029.675 202.740 3029.735 ;
        RECT 198.685 3029.445 198.855 3029.675 ;
        RECT 201.405 3029.445 201.575 3029.675 ;
        RECT 198.685 3029.115 198.855 3029.275 ;
        RECT 201.405 3029.115 201.575 3029.275 ;
        RECT 201.745 3029.165 202.765 3029.495 ;
        RECT 198.685 3028.985 199.655 3029.115 ;
        RECT 198.855 3028.815 199.655 3028.985 ;
        RECT 198.685 3028.785 199.655 3028.815 ;
        RECT 200.255 3028.995 201.575 3029.115 ;
        RECT 200.255 3028.985 202.375 3028.995 ;
        RECT 200.255 3028.815 201.405 3028.985 ;
        RECT 201.575 3028.825 202.375 3028.985 ;
        RECT 200.255 3028.785 201.575 3028.815 ;
        RECT 198.685 3028.525 198.855 3028.785 ;
      LAYER li1 ;
        RECT 199.025 3028.445 201.235 3028.615 ;
      LAYER li1 ;
        RECT 201.405 3028.525 201.575 3028.785 ;
        RECT 202.595 3028.655 202.765 3029.165 ;
      LAYER li1 ;
        RECT 199.505 3028.360 200.385 3028.445 ;
      LAYER li1 ;
        RECT 198.685 3028.275 198.855 3028.355 ;
        RECT 198.685 3028.065 199.335 3028.275 ;
        RECT 198.855 3027.945 199.335 3028.065 ;
        RECT 198.685 3027.605 198.855 3027.895 ;
      LAYER li1 ;
        RECT 199.505 3027.775 199.675 3028.360 ;
        RECT 199.025 3027.605 199.675 3027.775 ;
      LAYER li1 ;
        RECT 198.685 3027.145 199.335 3027.435 ;
        RECT 198.855 3027.105 199.335 3027.145 ;
        RECT 198.685 3026.685 198.855 3026.975 ;
      LAYER li1 ;
        RECT 199.505 3026.935 199.675 3027.605 ;
        RECT 199.025 3026.765 199.675 3026.935 ;
      LAYER li1 ;
        RECT 198.855 3026.515 199.335 3026.595 ;
        RECT 198.685 3026.265 199.335 3026.515 ;
        RECT 198.685 3026.225 198.855 3026.265 ;
      LAYER li1 ;
        RECT 199.505 3026.095 199.675 3026.765 ;
      LAYER li1 ;
        RECT 198.685 3025.765 198.855 3026.055 ;
      LAYER li1 ;
        RECT 199.025 3025.925 199.675 3026.095 ;
      LAYER li1 ;
        RECT 198.855 3025.595 199.335 3025.755 ;
        RECT 199.845 3025.665 200.015 3028.115 ;
      LAYER li1 ;
        RECT 200.215 3027.775 200.385 3028.360 ;
      LAYER li1 ;
        RECT 201.405 3028.275 201.575 3028.355 ;
        RECT 201.745 3028.325 202.765 3028.655 ;
      LAYER li1 ;
        RECT 202.935 3028.350 203.135 3029.940 ;
      LAYER li1 ;
        RECT 203.400 3029.905 204.295 3029.965 ;
        RECT 203.400 3029.735 204.125 3029.905 ;
        RECT 203.400 3029.675 204.295 3029.735 ;
        RECT 204.125 3029.445 204.295 3029.675 ;
        RECT 203.305 3029.245 203.955 3029.415 ;
        RECT 203.305 3028.575 203.475 3029.245 ;
        RECT 204.125 3029.075 204.295 3029.275 ;
        RECT 203.645 3028.985 204.295 3029.075 ;
        RECT 203.645 3028.815 204.125 3028.985 ;
        RECT 203.645 3028.745 204.295 3028.815 ;
        RECT 203.305 3028.405 203.950 3028.575 ;
        RECT 204.125 3028.525 204.295 3028.745 ;
        RECT 200.605 3028.155 201.575 3028.275 ;
        RECT 202.595 3028.170 202.765 3028.325 ;
        RECT 203.305 3028.170 203.475 3028.405 ;
        RECT 204.125 3028.235 204.295 3028.355 ;
        RECT 200.605 3028.065 202.375 3028.155 ;
        RECT 200.605 3027.945 201.405 3028.065 ;
        RECT 201.575 3027.985 202.375 3028.065 ;
        RECT 202.595 3027.995 203.475 3028.170 ;
        RECT 203.645 3028.065 204.295 3028.235 ;
      LAYER li1 ;
        RECT 200.215 3027.605 201.235 3027.775 ;
      LAYER li1 ;
        RECT 201.405 3027.605 201.575 3027.895 ;
      LAYER li1 ;
        RECT 200.215 3026.935 200.385 3027.605 ;
        RECT 201.745 3027.565 202.765 3027.735 ;
      LAYER li1 ;
        RECT 200.605 3027.395 201.575 3027.435 ;
        RECT 200.605 3027.145 202.375 3027.395 ;
        RECT 200.605 3027.105 201.405 3027.145 ;
        RECT 201.575 3027.065 202.375 3027.145 ;
      LAYER li1 ;
        RECT 200.215 3026.765 201.235 3026.935 ;
        RECT 200.215 3026.095 200.385 3026.765 ;
      LAYER li1 ;
        RECT 201.405 3026.685 201.575 3026.975 ;
      LAYER li1 ;
        RECT 202.595 3026.895 202.765 3027.565 ;
        RECT 201.745 3026.725 202.765 3026.895 ;
      LAYER li1 ;
        RECT 200.605 3026.515 201.405 3026.595 ;
        RECT 201.575 3026.515 202.375 3026.555 ;
        RECT 200.605 3026.265 202.375 3026.515 ;
        RECT 201.405 3026.225 202.375 3026.265 ;
      LAYER li1 ;
        RECT 200.215 3025.925 201.235 3026.095 ;
        RECT 202.595 3026.055 202.765 3026.725 ;
      LAYER li1 ;
        RECT 201.405 3025.765 201.575 3026.055 ;
      LAYER li1 ;
        RECT 201.745 3025.885 202.765 3026.055 ;
      LAYER li1 ;
        RECT 198.685 3025.425 199.335 3025.595 ;
        RECT 199.505 3025.490 200.385 3025.665 ;
        RECT 200.605 3025.595 201.405 3025.675 ;
        RECT 201.575 3025.595 202.375 3025.715 ;
        RECT 200.605 3025.505 202.375 3025.595 ;
        RECT 198.685 3025.305 198.855 3025.425 ;
        RECT 199.505 3025.255 199.675 3025.490 ;
        RECT 200.215 3025.335 200.385 3025.490 ;
        RECT 201.405 3025.385 202.375 3025.505 ;
        RECT 198.685 3024.915 198.855 3025.135 ;
        RECT 199.030 3025.085 199.675 3025.255 ;
        RECT 198.685 3024.845 199.335 3024.915 ;
        RECT 198.855 3024.675 199.335 3024.845 ;
        RECT 198.685 3024.585 199.335 3024.675 ;
        RECT 198.685 3024.385 198.855 3024.585 ;
        RECT 199.505 3024.415 199.675 3025.085 ;
        RECT 199.025 3024.245 199.675 3024.415 ;
        RECT 198.685 3023.985 198.855 3024.215 ;
      LAYER li1 ;
        RECT 199.845 3024.210 200.045 3025.310 ;
      LAYER li1 ;
        RECT 200.215 3025.005 201.235 3025.335 ;
        RECT 201.405 3025.305 201.575 3025.385 ;
      LAYER li1 ;
        RECT 202.595 3025.300 202.765 3025.885 ;
      LAYER li1 ;
        RECT 202.965 3025.545 203.135 3027.995 ;
        RECT 203.645 3027.905 204.125 3028.065 ;
      LAYER li1 ;
        RECT 203.305 3027.565 203.955 3027.735 ;
      LAYER li1 ;
        RECT 204.125 3027.605 204.295 3027.895 ;
      LAYER li1 ;
        RECT 203.305 3026.895 203.475 3027.565 ;
      LAYER li1 ;
        RECT 204.125 3027.395 204.295 3027.435 ;
        RECT 203.645 3027.145 204.295 3027.395 ;
        RECT 203.645 3027.065 204.125 3027.145 ;
      LAYER li1 ;
        RECT 203.305 3026.725 203.955 3026.895 ;
        RECT 203.305 3026.055 203.475 3026.725 ;
      LAYER li1 ;
        RECT 204.125 3026.685 204.295 3026.975 ;
        RECT 203.645 3026.515 204.125 3026.555 ;
        RECT 203.645 3026.225 204.295 3026.515 ;
      LAYER li1 ;
        RECT 203.305 3025.885 203.955 3026.055 ;
        RECT 203.305 3025.300 203.475 3025.885 ;
      LAYER li1 ;
        RECT 204.125 3025.765 204.295 3026.055 ;
        RECT 203.645 3025.595 204.125 3025.715 ;
        RECT 203.645 3025.385 204.295 3025.595 ;
        RECT 204.125 3025.305 204.295 3025.385 ;
      LAYER li1 ;
        RECT 202.595 3025.215 203.475 3025.300 ;
      LAYER li1 ;
        RECT 200.215 3024.495 200.385 3025.005 ;
        RECT 201.405 3024.875 201.575 3025.135 ;
      LAYER li1 ;
        RECT 201.745 3025.045 203.955 3025.215 ;
      LAYER li1 ;
        RECT 204.125 3024.875 204.295 3025.135 ;
        RECT 201.405 3024.845 202.725 3024.875 ;
        RECT 200.605 3024.675 201.405 3024.835 ;
        RECT 201.575 3024.675 202.725 3024.845 ;
        RECT 200.605 3024.665 202.725 3024.675 ;
        RECT 201.405 3024.545 202.725 3024.665 ;
        RECT 203.325 3024.845 204.295 3024.875 ;
        RECT 203.325 3024.675 204.125 3024.845 ;
        RECT 203.325 3024.545 204.295 3024.675 ;
        RECT 200.215 3024.165 201.235 3024.495 ;
        RECT 201.405 3024.385 201.575 3024.545 ;
        RECT 204.125 3024.385 204.295 3024.545 ;
        RECT 201.405 3023.985 201.575 3024.215 ;
        RECT 204.125 3023.985 204.295 3024.215 ;
        RECT 198.685 3023.925 199.580 3023.985 ;
        RECT 198.855 3023.755 199.580 3023.925 ;
        RECT 198.685 3023.695 199.580 3023.755 ;
        RECT 200.240 3023.925 202.740 3023.985 ;
        RECT 200.240 3023.755 201.405 3023.925 ;
        RECT 201.575 3023.755 202.740 3023.925 ;
        RECT 200.240 3023.695 202.740 3023.755 ;
        RECT 203.400 3023.925 204.295 3023.985 ;
        RECT 203.400 3023.755 204.125 3023.925 ;
        RECT 203.400 3023.695 204.295 3023.755 ;
        RECT 198.685 3023.465 198.855 3023.695 ;
        RECT 201.405 3023.465 201.575 3023.695 ;
        RECT 198.685 3023.135 198.855 3023.295 ;
        RECT 201.405 3023.135 201.575 3023.295 ;
        RECT 201.745 3023.185 202.765 3023.515 ;
        RECT 204.125 3023.465 204.295 3023.695 ;
        RECT 198.685 3023.005 199.655 3023.135 ;
        RECT 198.855 3022.835 199.655 3023.005 ;
        RECT 198.685 3022.805 199.655 3022.835 ;
        RECT 200.255 3023.015 201.575 3023.135 ;
        RECT 200.255 3023.005 202.375 3023.015 ;
        RECT 200.255 3022.835 201.405 3023.005 ;
        RECT 201.575 3022.845 202.375 3023.005 ;
        RECT 200.255 3022.805 201.575 3022.835 ;
        RECT 198.685 3022.545 198.855 3022.805 ;
        RECT 201.405 3022.545 201.575 3022.805 ;
        RECT 202.595 3022.675 202.765 3023.185 ;
        RECT 198.685 3022.295 198.855 3022.375 ;
        RECT 201.405 3022.295 201.575 3022.375 ;
        RECT 201.745 3022.345 202.765 3022.675 ;
        RECT 198.685 3022.085 199.335 3022.295 ;
        RECT 200.605 3022.175 201.575 3022.295 ;
        RECT 202.595 3022.190 202.765 3022.345 ;
        RECT 203.305 3023.265 203.955 3023.435 ;
        RECT 203.305 3022.595 203.475 3023.265 ;
        RECT 204.125 3023.095 204.295 3023.295 ;
        RECT 203.645 3023.005 204.295 3023.095 ;
        RECT 203.645 3022.835 204.125 3023.005 ;
        RECT 203.645 3022.765 204.295 3022.835 ;
        RECT 203.305 3022.425 203.950 3022.595 ;
        RECT 204.125 3022.545 204.295 3022.765 ;
        RECT 203.305 3022.190 203.475 3022.425 ;
        RECT 204.125 3022.255 204.295 3022.375 ;
        RECT 198.855 3021.965 199.335 3022.085 ;
        RECT 198.685 3021.625 198.855 3021.915 ;
        RECT 198.685 3021.165 199.335 3021.455 ;
        RECT 198.855 3021.125 199.335 3021.165 ;
        RECT 198.685 3020.705 198.855 3020.995 ;
        RECT 198.855 3020.535 199.335 3020.615 ;
        RECT 198.685 3020.285 199.335 3020.535 ;
        RECT 198.685 3020.245 198.855 3020.285 ;
        RECT 198.685 3019.785 198.855 3020.075 ;
        RECT 198.855 3019.615 199.335 3019.775 ;
        RECT 199.845 3019.685 200.015 3022.135 ;
        RECT 200.605 3022.085 202.375 3022.175 ;
        RECT 200.605 3021.965 201.405 3022.085 ;
        RECT 201.575 3022.005 202.375 3022.085 ;
        RECT 202.595 3022.015 203.475 3022.190 ;
        RECT 203.645 3022.085 204.295 3022.255 ;
        RECT 201.405 3021.625 201.575 3021.915 ;
      LAYER li1 ;
        RECT 201.745 3021.585 202.765 3021.755 ;
      LAYER li1 ;
        RECT 200.605 3021.415 201.575 3021.455 ;
        RECT 200.605 3021.165 202.375 3021.415 ;
        RECT 200.605 3021.125 201.405 3021.165 ;
        RECT 201.575 3021.085 202.375 3021.165 ;
        RECT 201.405 3020.705 201.575 3020.995 ;
      LAYER li1 ;
        RECT 202.595 3020.915 202.765 3021.585 ;
        RECT 201.745 3020.745 202.765 3020.915 ;
      LAYER li1 ;
        RECT 200.605 3020.535 201.405 3020.615 ;
        RECT 201.575 3020.535 202.375 3020.575 ;
        RECT 200.605 3020.285 202.375 3020.535 ;
        RECT 201.405 3020.245 202.375 3020.285 ;
      LAYER li1 ;
        RECT 202.595 3020.075 202.765 3020.745 ;
      LAYER li1 ;
        RECT 201.405 3019.785 201.575 3020.075 ;
      LAYER li1 ;
        RECT 201.745 3019.905 202.765 3020.075 ;
      LAYER li1 ;
        RECT 198.685 3019.445 199.335 3019.615 ;
        RECT 199.505 3019.510 200.385 3019.685 ;
        RECT 200.605 3019.615 201.405 3019.695 ;
        RECT 201.575 3019.615 202.375 3019.735 ;
        RECT 200.605 3019.525 202.375 3019.615 ;
        RECT 198.685 3019.325 198.855 3019.445 ;
        RECT 199.505 3019.275 199.675 3019.510 ;
        RECT 200.215 3019.355 200.385 3019.510 ;
        RECT 201.405 3019.405 202.375 3019.525 ;
        RECT 198.685 3018.935 198.855 3019.155 ;
        RECT 199.030 3019.105 199.675 3019.275 ;
        RECT 198.685 3018.865 199.335 3018.935 ;
        RECT 198.855 3018.695 199.335 3018.865 ;
        RECT 198.685 3018.605 199.335 3018.695 ;
        RECT 198.685 3018.405 198.855 3018.605 ;
        RECT 199.505 3018.435 199.675 3019.105 ;
        RECT 199.025 3018.265 199.675 3018.435 ;
        RECT 198.685 3018.005 198.855 3018.235 ;
      LAYER li1 ;
        RECT 199.845 3018.230 200.045 3019.330 ;
      LAYER li1 ;
        RECT 200.215 3019.025 201.235 3019.355 ;
        RECT 201.405 3019.325 201.575 3019.405 ;
      LAYER li1 ;
        RECT 202.595 3019.320 202.765 3019.905 ;
      LAYER li1 ;
        RECT 202.965 3019.565 203.135 3022.015 ;
        RECT 203.645 3021.925 204.125 3022.085 ;
      LAYER li1 ;
        RECT 203.305 3021.585 203.955 3021.755 ;
      LAYER li1 ;
        RECT 204.125 3021.625 204.295 3021.915 ;
      LAYER li1 ;
        RECT 203.305 3020.915 203.475 3021.585 ;
      LAYER li1 ;
        RECT 204.125 3021.415 204.295 3021.455 ;
        RECT 203.645 3021.165 204.295 3021.415 ;
        RECT 203.645 3021.085 204.125 3021.165 ;
      LAYER li1 ;
        RECT 203.305 3020.745 203.955 3020.915 ;
        RECT 203.305 3020.075 203.475 3020.745 ;
      LAYER li1 ;
        RECT 204.125 3020.705 204.295 3020.995 ;
        RECT 203.645 3020.535 204.125 3020.575 ;
        RECT 203.645 3020.245 204.295 3020.535 ;
      LAYER li1 ;
        RECT 203.305 3019.905 203.955 3020.075 ;
        RECT 203.305 3019.320 203.475 3019.905 ;
      LAYER li1 ;
        RECT 204.125 3019.785 204.295 3020.075 ;
        RECT 203.645 3019.615 204.125 3019.735 ;
        RECT 203.645 3019.405 204.295 3019.615 ;
        RECT 204.125 3019.325 204.295 3019.405 ;
      LAYER li1 ;
        RECT 202.595 3019.235 203.475 3019.320 ;
      LAYER li1 ;
        RECT 200.215 3018.515 200.385 3019.025 ;
        RECT 201.405 3018.895 201.575 3019.155 ;
      LAYER li1 ;
        RECT 201.745 3019.065 203.955 3019.235 ;
      LAYER li1 ;
        RECT 204.125 3018.895 204.295 3019.155 ;
        RECT 201.405 3018.865 202.725 3018.895 ;
        RECT 200.605 3018.695 201.405 3018.855 ;
        RECT 201.575 3018.695 202.725 3018.865 ;
        RECT 200.605 3018.685 202.725 3018.695 ;
        RECT 201.405 3018.565 202.725 3018.685 ;
        RECT 203.325 3018.865 204.295 3018.895 ;
        RECT 203.325 3018.695 204.125 3018.865 ;
        RECT 203.325 3018.565 204.295 3018.695 ;
        RECT 200.215 3018.185 201.235 3018.515 ;
        RECT 201.405 3018.405 201.575 3018.565 ;
        RECT 204.125 3018.405 204.295 3018.565 ;
        RECT 201.405 3018.005 201.575 3018.235 ;
        RECT 204.125 3018.005 204.295 3018.235 ;
        RECT 198.685 3017.945 199.580 3018.005 ;
        RECT 198.855 3017.775 199.580 3017.945 ;
        RECT 198.685 3017.715 199.580 3017.775 ;
        RECT 200.240 3017.945 202.740 3018.005 ;
        RECT 200.240 3017.775 201.405 3017.945 ;
        RECT 201.575 3017.775 202.740 3017.945 ;
        RECT 200.240 3017.715 202.740 3017.775 ;
        RECT 203.400 3017.945 204.295 3018.005 ;
        RECT 203.400 3017.775 204.125 3017.945 ;
        RECT 203.400 3017.715 204.295 3017.775 ;
        RECT 198.685 3017.485 198.855 3017.715 ;
        RECT 201.405 3017.485 201.575 3017.715 ;
        RECT 198.685 3017.155 198.855 3017.315 ;
        RECT 201.405 3017.155 201.575 3017.315 ;
        RECT 201.745 3017.205 202.765 3017.535 ;
        RECT 204.125 3017.485 204.295 3017.715 ;
        RECT 198.685 3017.025 199.655 3017.155 ;
        RECT 198.855 3016.855 199.655 3017.025 ;
        RECT 198.685 3016.825 199.655 3016.855 ;
        RECT 200.255 3017.035 201.575 3017.155 ;
        RECT 200.255 3017.025 202.375 3017.035 ;
        RECT 200.255 3016.855 201.405 3017.025 ;
        RECT 201.575 3016.865 202.375 3017.025 ;
        RECT 200.255 3016.825 201.575 3016.855 ;
        RECT 198.685 3016.565 198.855 3016.825 ;
        RECT 201.405 3016.565 201.575 3016.825 ;
        RECT 202.595 3016.695 202.765 3017.205 ;
        RECT 198.685 3016.315 198.855 3016.395 ;
        RECT 201.405 3016.315 201.575 3016.395 ;
        RECT 201.745 3016.365 202.765 3016.695 ;
        RECT 198.685 3016.105 199.335 3016.315 ;
        RECT 200.605 3016.195 201.575 3016.315 ;
        RECT 202.595 3016.210 202.765 3016.365 ;
        RECT 203.305 3017.285 203.955 3017.455 ;
        RECT 203.305 3016.615 203.475 3017.285 ;
        RECT 204.125 3017.115 204.295 3017.315 ;
        RECT 203.645 3017.025 204.295 3017.115 ;
        RECT 203.645 3016.855 204.125 3017.025 ;
        RECT 203.645 3016.785 204.295 3016.855 ;
        RECT 203.305 3016.445 203.950 3016.615 ;
        RECT 204.125 3016.565 204.295 3016.785 ;
        RECT 203.305 3016.210 203.475 3016.445 ;
        RECT 204.125 3016.275 204.295 3016.395 ;
        RECT 198.855 3015.985 199.335 3016.105 ;
        RECT 198.685 3015.645 198.855 3015.935 ;
        RECT 198.685 3015.185 199.335 3015.475 ;
        RECT 198.855 3015.145 199.335 3015.185 ;
        RECT 198.685 3014.725 198.855 3015.015 ;
        RECT 198.855 3014.555 199.335 3014.635 ;
        RECT 198.685 3014.305 199.335 3014.555 ;
        RECT 198.685 3014.265 198.855 3014.305 ;
        RECT 198.685 3013.805 198.855 3014.095 ;
        RECT 198.855 3013.635 199.335 3013.795 ;
        RECT 199.845 3013.705 200.015 3016.155 ;
        RECT 200.605 3016.105 202.375 3016.195 ;
        RECT 200.605 3015.985 201.405 3016.105 ;
        RECT 201.575 3016.025 202.375 3016.105 ;
        RECT 202.595 3016.035 203.475 3016.210 ;
        RECT 203.645 3016.105 204.295 3016.275 ;
        RECT 201.405 3015.645 201.575 3015.935 ;
      LAYER li1 ;
        RECT 201.745 3015.605 202.765 3015.775 ;
      LAYER li1 ;
        RECT 200.605 3015.435 201.575 3015.475 ;
        RECT 200.605 3015.185 202.375 3015.435 ;
        RECT 200.605 3015.145 201.405 3015.185 ;
        RECT 201.575 3015.105 202.375 3015.185 ;
        RECT 201.405 3014.725 201.575 3015.015 ;
      LAYER li1 ;
        RECT 202.595 3014.935 202.765 3015.605 ;
        RECT 201.745 3014.765 202.765 3014.935 ;
      LAYER li1 ;
        RECT 200.605 3014.555 201.405 3014.635 ;
        RECT 201.575 3014.555 202.375 3014.595 ;
        RECT 200.605 3014.305 202.375 3014.555 ;
        RECT 201.405 3014.265 202.375 3014.305 ;
      LAYER li1 ;
        RECT 202.595 3014.095 202.765 3014.765 ;
      LAYER li1 ;
        RECT 201.405 3013.805 201.575 3014.095 ;
      LAYER li1 ;
        RECT 201.745 3013.925 202.765 3014.095 ;
      LAYER li1 ;
        RECT 198.685 3013.465 199.335 3013.635 ;
        RECT 199.505 3013.530 200.385 3013.705 ;
        RECT 200.605 3013.635 201.405 3013.715 ;
        RECT 201.575 3013.635 202.375 3013.755 ;
        RECT 200.605 3013.545 202.375 3013.635 ;
        RECT 198.685 3013.345 198.855 3013.465 ;
        RECT 199.505 3013.295 199.675 3013.530 ;
        RECT 200.215 3013.375 200.385 3013.530 ;
        RECT 201.405 3013.425 202.375 3013.545 ;
        RECT 198.685 3012.955 198.855 3013.175 ;
        RECT 199.030 3013.125 199.675 3013.295 ;
        RECT 198.685 3012.885 199.335 3012.955 ;
        RECT 198.855 3012.715 199.335 3012.885 ;
        RECT 198.685 3012.625 199.335 3012.715 ;
        RECT 198.685 3012.425 198.855 3012.625 ;
        RECT 199.505 3012.455 199.675 3013.125 ;
        RECT 199.025 3012.285 199.675 3012.455 ;
        RECT 198.685 3012.025 198.855 3012.255 ;
      LAYER li1 ;
        RECT 199.845 3012.250 200.045 3013.350 ;
      LAYER li1 ;
        RECT 200.215 3013.045 201.235 3013.375 ;
        RECT 201.405 3013.345 201.575 3013.425 ;
      LAYER li1 ;
        RECT 202.595 3013.340 202.765 3013.925 ;
      LAYER li1 ;
        RECT 202.965 3013.585 203.135 3016.035 ;
        RECT 203.645 3015.945 204.125 3016.105 ;
      LAYER li1 ;
        RECT 203.305 3015.605 203.955 3015.775 ;
      LAYER li1 ;
        RECT 204.125 3015.645 204.295 3015.935 ;
      LAYER li1 ;
        RECT 203.305 3014.935 203.475 3015.605 ;
      LAYER li1 ;
        RECT 204.125 3015.435 204.295 3015.475 ;
        RECT 203.645 3015.185 204.295 3015.435 ;
        RECT 203.645 3015.105 204.125 3015.185 ;
      LAYER li1 ;
        RECT 203.305 3014.765 203.955 3014.935 ;
        RECT 203.305 3014.095 203.475 3014.765 ;
      LAYER li1 ;
        RECT 204.125 3014.725 204.295 3015.015 ;
        RECT 203.645 3014.555 204.125 3014.595 ;
        RECT 203.645 3014.265 204.295 3014.555 ;
      LAYER li1 ;
        RECT 203.305 3013.925 203.955 3014.095 ;
        RECT 203.305 3013.340 203.475 3013.925 ;
      LAYER li1 ;
        RECT 204.125 3013.805 204.295 3014.095 ;
        RECT 203.645 3013.635 204.125 3013.755 ;
        RECT 203.645 3013.425 204.295 3013.635 ;
        RECT 204.125 3013.345 204.295 3013.425 ;
      LAYER li1 ;
        RECT 202.595 3013.255 203.475 3013.340 ;
      LAYER li1 ;
        RECT 200.215 3012.535 200.385 3013.045 ;
        RECT 201.405 3012.915 201.575 3013.175 ;
      LAYER li1 ;
        RECT 201.745 3013.085 203.955 3013.255 ;
      LAYER li1 ;
        RECT 204.125 3012.915 204.295 3013.175 ;
        RECT 201.405 3012.885 202.725 3012.915 ;
        RECT 200.605 3012.715 201.405 3012.875 ;
        RECT 201.575 3012.715 202.725 3012.885 ;
        RECT 200.605 3012.705 202.725 3012.715 ;
        RECT 201.405 3012.585 202.725 3012.705 ;
        RECT 203.325 3012.885 204.295 3012.915 ;
        RECT 203.325 3012.715 204.125 3012.885 ;
        RECT 203.325 3012.585 204.295 3012.715 ;
        RECT 200.215 3012.205 201.235 3012.535 ;
        RECT 201.405 3012.425 201.575 3012.585 ;
        RECT 204.125 3012.425 204.295 3012.585 ;
        RECT 201.405 3012.025 201.575 3012.255 ;
        RECT 204.125 3012.025 204.295 3012.255 ;
        RECT 198.685 3011.965 199.580 3012.025 ;
        RECT 198.855 3011.795 199.580 3011.965 ;
        RECT 198.685 3011.735 199.580 3011.795 ;
        RECT 200.240 3011.965 202.740 3012.025 ;
        RECT 200.240 3011.795 201.405 3011.965 ;
        RECT 201.575 3011.795 202.740 3011.965 ;
        RECT 200.240 3011.735 202.740 3011.795 ;
        RECT 203.400 3011.965 204.295 3012.025 ;
        RECT 203.400 3011.795 204.125 3011.965 ;
        RECT 203.400 3011.735 204.295 3011.795 ;
        RECT 198.685 3011.505 198.855 3011.735 ;
        RECT 201.405 3011.505 201.575 3011.735 ;
        RECT 198.685 3011.175 198.855 3011.335 ;
        RECT 201.405 3011.175 201.575 3011.335 ;
        RECT 201.745 3011.225 202.765 3011.555 ;
        RECT 204.125 3011.505 204.295 3011.735 ;
        RECT 198.685 3011.045 199.655 3011.175 ;
        RECT 198.855 3010.875 199.655 3011.045 ;
        RECT 198.685 3010.845 199.655 3010.875 ;
        RECT 200.255 3011.055 201.575 3011.175 ;
        RECT 200.255 3011.045 202.375 3011.055 ;
        RECT 200.255 3010.875 201.405 3011.045 ;
        RECT 201.575 3010.885 202.375 3011.045 ;
        RECT 200.255 3010.845 201.575 3010.875 ;
        RECT 198.685 3010.585 198.855 3010.845 ;
        RECT 201.405 3010.585 201.575 3010.845 ;
        RECT 202.595 3010.715 202.765 3011.225 ;
        RECT 198.685 3010.335 198.855 3010.415 ;
        RECT 201.405 3010.335 201.575 3010.415 ;
        RECT 201.745 3010.385 202.765 3010.715 ;
        RECT 198.685 3010.125 199.335 3010.335 ;
        RECT 200.605 3010.215 201.575 3010.335 ;
        RECT 202.595 3010.230 202.765 3010.385 ;
        RECT 203.305 3011.305 203.955 3011.475 ;
        RECT 203.305 3010.635 203.475 3011.305 ;
        RECT 204.125 3011.135 204.295 3011.335 ;
        RECT 203.645 3011.045 204.295 3011.135 ;
        RECT 203.645 3010.875 204.125 3011.045 ;
        RECT 203.645 3010.805 204.295 3010.875 ;
        RECT 203.305 3010.465 203.950 3010.635 ;
        RECT 204.125 3010.585 204.295 3010.805 ;
        RECT 203.305 3010.230 203.475 3010.465 ;
        RECT 204.125 3010.295 204.295 3010.415 ;
        RECT 198.855 3010.005 199.335 3010.125 ;
        RECT 198.685 3009.665 198.855 3009.955 ;
        RECT 198.685 3009.205 199.335 3009.495 ;
        RECT 198.855 3009.165 199.335 3009.205 ;
        RECT 198.685 3008.745 198.855 3009.035 ;
        RECT 198.855 3008.575 199.335 3008.655 ;
        RECT 198.685 3008.325 199.335 3008.575 ;
        RECT 198.685 3008.285 198.855 3008.325 ;
        RECT 198.685 3007.825 198.855 3008.115 ;
        RECT 198.855 3007.655 199.335 3007.815 ;
        RECT 199.845 3007.725 200.015 3010.175 ;
        RECT 200.605 3010.125 202.375 3010.215 ;
        RECT 200.605 3010.005 201.405 3010.125 ;
        RECT 201.575 3010.045 202.375 3010.125 ;
        RECT 202.595 3010.055 203.475 3010.230 ;
        RECT 203.645 3010.125 204.295 3010.295 ;
        RECT 201.405 3009.665 201.575 3009.955 ;
      LAYER li1 ;
        RECT 201.745 3009.625 202.765 3009.795 ;
      LAYER li1 ;
        RECT 200.605 3009.455 201.575 3009.495 ;
        RECT 200.605 3009.205 202.375 3009.455 ;
        RECT 200.605 3009.165 201.405 3009.205 ;
        RECT 201.575 3009.125 202.375 3009.205 ;
        RECT 201.405 3008.745 201.575 3009.035 ;
      LAYER li1 ;
        RECT 202.595 3008.955 202.765 3009.625 ;
        RECT 201.745 3008.785 202.765 3008.955 ;
      LAYER li1 ;
        RECT 200.605 3008.575 201.405 3008.655 ;
        RECT 201.575 3008.575 202.375 3008.615 ;
        RECT 200.605 3008.325 202.375 3008.575 ;
        RECT 201.405 3008.285 202.375 3008.325 ;
      LAYER li1 ;
        RECT 202.595 3008.115 202.765 3008.785 ;
      LAYER li1 ;
        RECT 201.405 3007.825 201.575 3008.115 ;
      LAYER li1 ;
        RECT 201.745 3007.945 202.765 3008.115 ;
      LAYER li1 ;
        RECT 198.685 3007.485 199.335 3007.655 ;
        RECT 199.505 3007.550 200.385 3007.725 ;
        RECT 200.605 3007.655 201.405 3007.735 ;
        RECT 201.575 3007.655 202.375 3007.775 ;
        RECT 200.605 3007.565 202.375 3007.655 ;
        RECT 198.685 3007.365 198.855 3007.485 ;
        RECT 199.505 3007.315 199.675 3007.550 ;
        RECT 200.215 3007.395 200.385 3007.550 ;
        RECT 201.405 3007.445 202.375 3007.565 ;
        RECT 198.685 3006.975 198.855 3007.195 ;
        RECT 199.030 3007.145 199.675 3007.315 ;
        RECT 198.685 3006.905 199.335 3006.975 ;
        RECT 198.855 3006.735 199.335 3006.905 ;
        RECT 198.685 3006.645 199.335 3006.735 ;
        RECT 198.685 3006.445 198.855 3006.645 ;
        RECT 199.505 3006.475 199.675 3007.145 ;
        RECT 199.025 3006.305 199.675 3006.475 ;
        RECT 198.685 3006.045 198.855 3006.275 ;
      LAYER li1 ;
        RECT 199.845 3006.270 200.045 3007.370 ;
      LAYER li1 ;
        RECT 200.215 3007.065 201.235 3007.395 ;
        RECT 201.405 3007.365 201.575 3007.445 ;
      LAYER li1 ;
        RECT 202.595 3007.360 202.765 3007.945 ;
      LAYER li1 ;
        RECT 202.965 3007.605 203.135 3010.055 ;
        RECT 203.645 3009.965 204.125 3010.125 ;
      LAYER li1 ;
        RECT 203.305 3009.625 203.955 3009.795 ;
      LAYER li1 ;
        RECT 204.125 3009.665 204.295 3009.955 ;
      LAYER li1 ;
        RECT 203.305 3008.955 203.475 3009.625 ;
      LAYER li1 ;
        RECT 204.125 3009.455 204.295 3009.495 ;
        RECT 203.645 3009.205 204.295 3009.455 ;
        RECT 203.645 3009.125 204.125 3009.205 ;
      LAYER li1 ;
        RECT 203.305 3008.785 203.955 3008.955 ;
        RECT 203.305 3008.115 203.475 3008.785 ;
      LAYER li1 ;
        RECT 204.125 3008.745 204.295 3009.035 ;
        RECT 203.645 3008.575 204.125 3008.615 ;
        RECT 203.645 3008.285 204.295 3008.575 ;
      LAYER li1 ;
        RECT 203.305 3007.945 203.955 3008.115 ;
        RECT 203.305 3007.360 203.475 3007.945 ;
      LAYER li1 ;
        RECT 204.125 3007.825 204.295 3008.115 ;
        RECT 203.645 3007.655 204.125 3007.775 ;
        RECT 203.645 3007.445 204.295 3007.655 ;
        RECT 204.125 3007.365 204.295 3007.445 ;
      LAYER li1 ;
        RECT 202.595 3007.275 203.475 3007.360 ;
      LAYER li1 ;
        RECT 200.215 3006.555 200.385 3007.065 ;
        RECT 201.405 3006.935 201.575 3007.195 ;
      LAYER li1 ;
        RECT 201.745 3007.105 203.955 3007.275 ;
      LAYER li1 ;
        RECT 204.125 3006.935 204.295 3007.195 ;
        RECT 201.405 3006.905 202.725 3006.935 ;
        RECT 200.605 3006.735 201.405 3006.895 ;
        RECT 201.575 3006.735 202.725 3006.905 ;
        RECT 200.605 3006.725 202.725 3006.735 ;
        RECT 201.405 3006.605 202.725 3006.725 ;
        RECT 203.325 3006.905 204.295 3006.935 ;
        RECT 203.325 3006.735 204.125 3006.905 ;
        RECT 203.325 3006.605 204.295 3006.735 ;
        RECT 200.215 3006.225 201.235 3006.555 ;
        RECT 201.405 3006.445 201.575 3006.605 ;
        RECT 204.125 3006.445 204.295 3006.605 ;
        RECT 201.405 3006.045 201.575 3006.275 ;
        RECT 204.125 3006.045 204.295 3006.275 ;
        RECT 198.685 3005.985 199.580 3006.045 ;
        RECT 198.855 3005.815 199.580 3005.985 ;
        RECT 198.685 3005.755 199.580 3005.815 ;
        RECT 200.240 3005.985 202.740 3006.045 ;
        RECT 200.240 3005.815 201.405 3005.985 ;
        RECT 201.575 3005.815 202.740 3005.985 ;
        RECT 200.240 3005.755 202.740 3005.815 ;
        RECT 203.400 3005.985 204.295 3006.045 ;
        RECT 203.400 3005.815 204.125 3005.985 ;
        RECT 203.400 3005.755 204.295 3005.815 ;
        RECT 198.685 3005.525 198.855 3005.755 ;
        RECT 201.405 3005.525 201.575 3005.755 ;
        RECT 198.685 3005.195 198.855 3005.355 ;
        RECT 201.405 3005.195 201.575 3005.355 ;
        RECT 201.745 3005.245 202.765 3005.575 ;
        RECT 204.125 3005.525 204.295 3005.755 ;
        RECT 198.685 3005.065 199.655 3005.195 ;
        RECT 198.855 3004.895 199.655 3005.065 ;
        RECT 198.685 3004.865 199.655 3004.895 ;
        RECT 200.255 3005.075 201.575 3005.195 ;
        RECT 200.255 3005.065 202.375 3005.075 ;
        RECT 200.255 3004.895 201.405 3005.065 ;
        RECT 201.575 3004.905 202.375 3005.065 ;
        RECT 200.255 3004.865 201.575 3004.895 ;
        RECT 198.685 3004.605 198.855 3004.865 ;
        RECT 201.405 3004.605 201.575 3004.865 ;
        RECT 202.595 3004.735 202.765 3005.245 ;
        RECT 198.685 3004.355 198.855 3004.435 ;
        RECT 201.405 3004.355 201.575 3004.435 ;
        RECT 201.745 3004.405 202.765 3004.735 ;
        RECT 198.685 3004.145 199.335 3004.355 ;
        RECT 200.605 3004.235 201.575 3004.355 ;
        RECT 202.595 3004.250 202.765 3004.405 ;
        RECT 203.305 3005.325 203.955 3005.495 ;
        RECT 203.305 3004.655 203.475 3005.325 ;
        RECT 204.125 3005.155 204.295 3005.355 ;
        RECT 203.645 3005.065 204.295 3005.155 ;
        RECT 203.645 3004.895 204.125 3005.065 ;
        RECT 203.645 3004.825 204.295 3004.895 ;
        RECT 203.305 3004.485 203.950 3004.655 ;
        RECT 204.125 3004.605 204.295 3004.825 ;
        RECT 203.305 3004.250 203.475 3004.485 ;
        RECT 204.125 3004.315 204.295 3004.435 ;
        RECT 198.855 3004.025 199.335 3004.145 ;
        RECT 198.685 3003.685 198.855 3003.975 ;
        RECT 198.685 3003.225 199.335 3003.515 ;
        RECT 198.855 3003.185 199.335 3003.225 ;
        RECT 198.685 3002.765 198.855 3003.055 ;
        RECT 198.855 3002.595 199.335 3002.675 ;
        RECT 198.685 3002.345 199.335 3002.595 ;
        RECT 198.685 3002.305 198.855 3002.345 ;
        RECT 198.685 3001.845 198.855 3002.135 ;
        RECT 198.855 3001.675 199.335 3001.835 ;
        RECT 199.845 3001.745 200.015 3004.195 ;
        RECT 200.605 3004.145 202.375 3004.235 ;
        RECT 200.605 3004.025 201.405 3004.145 ;
        RECT 201.575 3004.065 202.375 3004.145 ;
        RECT 202.595 3004.075 203.475 3004.250 ;
        RECT 203.645 3004.145 204.295 3004.315 ;
        RECT 201.405 3003.685 201.575 3003.975 ;
      LAYER li1 ;
        RECT 201.745 3003.645 202.765 3003.815 ;
      LAYER li1 ;
        RECT 200.605 3003.475 201.575 3003.515 ;
        RECT 200.605 3003.225 202.375 3003.475 ;
        RECT 200.605 3003.185 201.405 3003.225 ;
        RECT 201.575 3003.145 202.375 3003.225 ;
        RECT 201.405 3002.765 201.575 3003.055 ;
      LAYER li1 ;
        RECT 202.595 3002.975 202.765 3003.645 ;
        RECT 201.745 3002.805 202.765 3002.975 ;
      LAYER li1 ;
        RECT 200.605 3002.595 201.405 3002.675 ;
        RECT 201.575 3002.595 202.375 3002.635 ;
        RECT 200.605 3002.345 202.375 3002.595 ;
        RECT 201.405 3002.305 202.375 3002.345 ;
      LAYER li1 ;
        RECT 202.595 3002.135 202.765 3002.805 ;
      LAYER li1 ;
        RECT 201.405 3001.845 201.575 3002.135 ;
      LAYER li1 ;
        RECT 201.745 3001.965 202.765 3002.135 ;
      LAYER li1 ;
        RECT 198.685 3001.505 199.335 3001.675 ;
        RECT 199.505 3001.570 200.385 3001.745 ;
        RECT 200.605 3001.675 201.405 3001.755 ;
        RECT 201.575 3001.675 202.375 3001.795 ;
        RECT 200.605 3001.585 202.375 3001.675 ;
        RECT 198.685 3001.385 198.855 3001.505 ;
        RECT 199.505 3001.335 199.675 3001.570 ;
        RECT 200.215 3001.415 200.385 3001.570 ;
        RECT 201.405 3001.465 202.375 3001.585 ;
        RECT 198.685 3000.995 198.855 3001.215 ;
        RECT 199.030 3001.165 199.675 3001.335 ;
        RECT 198.685 3000.925 199.335 3000.995 ;
        RECT 198.855 3000.755 199.335 3000.925 ;
        RECT 198.685 3000.665 199.335 3000.755 ;
        RECT 198.685 3000.465 198.855 3000.665 ;
        RECT 199.505 3000.495 199.675 3001.165 ;
        RECT 199.025 3000.325 199.675 3000.495 ;
        RECT 198.685 3000.065 198.855 3000.295 ;
      LAYER li1 ;
        RECT 199.845 3000.290 200.045 3001.390 ;
      LAYER li1 ;
        RECT 200.215 3001.085 201.235 3001.415 ;
        RECT 201.405 3001.385 201.575 3001.465 ;
      LAYER li1 ;
        RECT 202.595 3001.380 202.765 3001.965 ;
      LAYER li1 ;
        RECT 202.965 3001.625 203.135 3004.075 ;
        RECT 203.645 3003.985 204.125 3004.145 ;
      LAYER li1 ;
        RECT 203.305 3003.645 203.955 3003.815 ;
      LAYER li1 ;
        RECT 204.125 3003.685 204.295 3003.975 ;
      LAYER li1 ;
        RECT 203.305 3002.975 203.475 3003.645 ;
      LAYER li1 ;
        RECT 204.125 3003.475 204.295 3003.515 ;
        RECT 203.645 3003.225 204.295 3003.475 ;
        RECT 203.645 3003.145 204.125 3003.225 ;
      LAYER li1 ;
        RECT 203.305 3002.805 203.955 3002.975 ;
        RECT 203.305 3002.135 203.475 3002.805 ;
      LAYER li1 ;
        RECT 204.125 3002.765 204.295 3003.055 ;
        RECT 203.645 3002.595 204.125 3002.635 ;
        RECT 203.645 3002.305 204.295 3002.595 ;
      LAYER li1 ;
        RECT 203.305 3001.965 203.955 3002.135 ;
        RECT 203.305 3001.380 203.475 3001.965 ;
      LAYER li1 ;
        RECT 204.125 3001.845 204.295 3002.135 ;
        RECT 203.645 3001.675 204.125 3001.795 ;
        RECT 203.645 3001.465 204.295 3001.675 ;
        RECT 204.125 3001.385 204.295 3001.465 ;
      LAYER li1 ;
        RECT 202.595 3001.295 203.475 3001.380 ;
      LAYER li1 ;
        RECT 200.215 3000.575 200.385 3001.085 ;
        RECT 201.405 3000.955 201.575 3001.215 ;
      LAYER li1 ;
        RECT 201.745 3001.125 203.955 3001.295 ;
      LAYER li1 ;
        RECT 204.125 3000.955 204.295 3001.215 ;
        RECT 201.405 3000.925 202.725 3000.955 ;
        RECT 200.605 3000.755 201.405 3000.915 ;
        RECT 201.575 3000.755 202.725 3000.925 ;
        RECT 200.605 3000.745 202.725 3000.755 ;
        RECT 201.405 3000.625 202.725 3000.745 ;
        RECT 203.325 3000.925 204.295 3000.955 ;
        RECT 203.325 3000.755 204.125 3000.925 ;
        RECT 203.325 3000.625 204.295 3000.755 ;
        RECT 200.215 3000.245 201.235 3000.575 ;
        RECT 201.405 3000.465 201.575 3000.625 ;
        RECT 204.125 3000.465 204.295 3000.625 ;
        RECT 201.405 3000.065 201.575 3000.295 ;
        RECT 204.125 3000.065 204.295 3000.295 ;
        RECT 198.685 3000.005 199.580 3000.065 ;
        RECT 198.855 2999.835 199.580 3000.005 ;
        RECT 198.685 2999.775 199.580 2999.835 ;
        RECT 200.240 3000.005 202.740 3000.065 ;
        RECT 200.240 2999.835 201.405 3000.005 ;
        RECT 201.575 2999.835 202.740 3000.005 ;
        RECT 200.240 2999.775 202.740 2999.835 ;
        RECT 203.400 3000.005 204.295 3000.065 ;
        RECT 203.400 2999.835 204.125 3000.005 ;
        RECT 203.400 2999.775 204.295 2999.835 ;
        RECT 198.685 2999.545 198.855 2999.775 ;
        RECT 201.405 2999.545 201.575 2999.775 ;
        RECT 198.685 2999.215 198.855 2999.375 ;
        RECT 201.405 2999.215 201.575 2999.375 ;
        RECT 201.745 2999.265 202.765 2999.595 ;
        RECT 204.125 2999.545 204.295 2999.775 ;
        RECT 198.685 2999.085 199.655 2999.215 ;
        RECT 198.855 2998.915 199.655 2999.085 ;
        RECT 198.685 2998.885 199.655 2998.915 ;
        RECT 200.255 2999.095 201.575 2999.215 ;
        RECT 200.255 2999.085 202.375 2999.095 ;
        RECT 200.255 2998.915 201.405 2999.085 ;
        RECT 201.575 2998.925 202.375 2999.085 ;
        RECT 200.255 2998.885 201.575 2998.915 ;
        RECT 198.685 2998.625 198.855 2998.885 ;
        RECT 201.405 2998.625 201.575 2998.885 ;
        RECT 202.595 2998.755 202.765 2999.265 ;
        RECT 198.685 2998.375 198.855 2998.455 ;
        RECT 201.405 2998.375 201.575 2998.455 ;
        RECT 201.745 2998.425 202.765 2998.755 ;
        RECT 198.685 2998.165 199.335 2998.375 ;
        RECT 200.605 2998.255 201.575 2998.375 ;
        RECT 202.595 2998.270 202.765 2998.425 ;
        RECT 203.305 2999.345 203.955 2999.515 ;
        RECT 203.305 2998.675 203.475 2999.345 ;
        RECT 204.125 2999.175 204.295 2999.375 ;
        RECT 203.645 2999.085 204.295 2999.175 ;
        RECT 203.645 2998.915 204.125 2999.085 ;
        RECT 203.645 2998.845 204.295 2998.915 ;
        RECT 203.305 2998.505 203.950 2998.675 ;
        RECT 204.125 2998.625 204.295 2998.845 ;
        RECT 203.305 2998.270 203.475 2998.505 ;
        RECT 204.125 2998.335 204.295 2998.455 ;
        RECT 198.855 2998.045 199.335 2998.165 ;
        RECT 198.685 2997.705 198.855 2997.995 ;
        RECT 198.685 2997.245 199.335 2997.535 ;
        RECT 198.855 2997.205 199.335 2997.245 ;
        RECT 198.685 2996.785 198.855 2997.075 ;
        RECT 198.855 2996.615 199.335 2996.695 ;
        RECT 198.685 2996.365 199.335 2996.615 ;
        RECT 198.685 2996.325 198.855 2996.365 ;
        RECT 198.685 2995.865 198.855 2996.155 ;
        RECT 198.855 2995.695 199.335 2995.855 ;
        RECT 199.845 2995.765 200.015 2998.215 ;
        RECT 200.605 2998.165 202.375 2998.255 ;
        RECT 200.605 2998.045 201.405 2998.165 ;
        RECT 201.575 2998.085 202.375 2998.165 ;
        RECT 202.595 2998.095 203.475 2998.270 ;
        RECT 203.645 2998.165 204.295 2998.335 ;
        RECT 201.405 2997.705 201.575 2997.995 ;
      LAYER li1 ;
        RECT 201.745 2997.665 202.765 2997.835 ;
      LAYER li1 ;
        RECT 200.605 2997.495 201.575 2997.535 ;
        RECT 200.605 2997.245 202.375 2997.495 ;
        RECT 200.605 2997.205 201.405 2997.245 ;
        RECT 201.575 2997.165 202.375 2997.245 ;
        RECT 201.405 2996.785 201.575 2997.075 ;
      LAYER li1 ;
        RECT 202.595 2996.995 202.765 2997.665 ;
        RECT 201.745 2996.825 202.765 2996.995 ;
      LAYER li1 ;
        RECT 200.605 2996.615 201.405 2996.695 ;
        RECT 201.575 2996.615 202.375 2996.655 ;
        RECT 200.605 2996.365 202.375 2996.615 ;
        RECT 201.405 2996.325 202.375 2996.365 ;
      LAYER li1 ;
        RECT 202.595 2996.155 202.765 2996.825 ;
      LAYER li1 ;
        RECT 201.405 2995.865 201.575 2996.155 ;
      LAYER li1 ;
        RECT 201.745 2995.985 202.765 2996.155 ;
      LAYER li1 ;
        RECT 198.685 2995.525 199.335 2995.695 ;
        RECT 199.505 2995.590 200.385 2995.765 ;
        RECT 200.605 2995.695 201.405 2995.775 ;
        RECT 201.575 2995.695 202.375 2995.815 ;
        RECT 200.605 2995.605 202.375 2995.695 ;
        RECT 198.685 2995.405 198.855 2995.525 ;
        RECT 199.505 2995.355 199.675 2995.590 ;
        RECT 200.215 2995.435 200.385 2995.590 ;
        RECT 201.405 2995.485 202.375 2995.605 ;
        RECT 198.685 2995.015 198.855 2995.235 ;
        RECT 199.030 2995.185 199.675 2995.355 ;
        RECT 198.685 2994.945 199.335 2995.015 ;
        RECT 198.855 2994.775 199.335 2994.945 ;
        RECT 198.685 2994.685 199.335 2994.775 ;
        RECT 198.685 2994.485 198.855 2994.685 ;
        RECT 199.505 2994.515 199.675 2995.185 ;
        RECT 199.025 2994.345 199.675 2994.515 ;
        RECT 198.685 2994.085 198.855 2994.315 ;
      LAYER li1 ;
        RECT 199.845 2994.310 200.045 2995.410 ;
      LAYER li1 ;
        RECT 200.215 2995.105 201.235 2995.435 ;
        RECT 201.405 2995.405 201.575 2995.485 ;
      LAYER li1 ;
        RECT 202.595 2995.400 202.765 2995.985 ;
      LAYER li1 ;
        RECT 202.965 2995.645 203.135 2998.095 ;
        RECT 203.645 2998.005 204.125 2998.165 ;
      LAYER li1 ;
        RECT 203.305 2997.665 203.955 2997.835 ;
      LAYER li1 ;
        RECT 204.125 2997.705 204.295 2997.995 ;
      LAYER li1 ;
        RECT 203.305 2996.995 203.475 2997.665 ;
      LAYER li1 ;
        RECT 204.125 2997.495 204.295 2997.535 ;
        RECT 203.645 2997.245 204.295 2997.495 ;
        RECT 203.645 2997.165 204.125 2997.245 ;
      LAYER li1 ;
        RECT 203.305 2996.825 203.955 2996.995 ;
        RECT 203.305 2996.155 203.475 2996.825 ;
      LAYER li1 ;
        RECT 204.125 2996.785 204.295 2997.075 ;
        RECT 203.645 2996.615 204.125 2996.655 ;
        RECT 203.645 2996.325 204.295 2996.615 ;
      LAYER li1 ;
        RECT 203.305 2995.985 203.955 2996.155 ;
        RECT 203.305 2995.400 203.475 2995.985 ;
      LAYER li1 ;
        RECT 204.125 2995.865 204.295 2996.155 ;
        RECT 203.645 2995.695 204.125 2995.815 ;
        RECT 203.645 2995.485 204.295 2995.695 ;
        RECT 204.125 2995.405 204.295 2995.485 ;
      LAYER li1 ;
        RECT 202.595 2995.315 203.475 2995.400 ;
      LAYER li1 ;
        RECT 200.215 2994.595 200.385 2995.105 ;
        RECT 201.405 2994.975 201.575 2995.235 ;
      LAYER li1 ;
        RECT 201.745 2995.145 203.955 2995.315 ;
      LAYER li1 ;
        RECT 204.125 2994.975 204.295 2995.235 ;
        RECT 201.405 2994.945 202.725 2994.975 ;
        RECT 200.605 2994.775 201.405 2994.935 ;
        RECT 201.575 2994.775 202.725 2994.945 ;
        RECT 200.605 2994.765 202.725 2994.775 ;
        RECT 201.405 2994.645 202.725 2994.765 ;
        RECT 203.325 2994.945 204.295 2994.975 ;
        RECT 203.325 2994.775 204.125 2994.945 ;
        RECT 203.325 2994.645 204.295 2994.775 ;
        RECT 200.215 2994.265 201.235 2994.595 ;
        RECT 201.405 2994.485 201.575 2994.645 ;
        RECT 204.125 2994.485 204.295 2994.645 ;
        RECT 201.405 2994.085 201.575 2994.315 ;
        RECT 204.125 2994.085 204.295 2994.315 ;
        RECT 198.685 2994.025 199.580 2994.085 ;
        RECT 198.855 2993.855 199.580 2994.025 ;
        RECT 198.685 2993.795 199.580 2993.855 ;
        RECT 200.240 2994.025 202.740 2994.085 ;
        RECT 200.240 2993.855 201.405 2994.025 ;
        RECT 201.575 2993.855 202.740 2994.025 ;
        RECT 200.240 2993.795 202.740 2993.855 ;
        RECT 203.400 2994.025 204.295 2994.085 ;
        RECT 203.400 2993.855 204.125 2994.025 ;
        RECT 203.400 2993.795 204.295 2993.855 ;
        RECT 198.685 2993.565 198.855 2993.795 ;
        RECT 201.405 2993.565 201.575 2993.795 ;
        RECT 198.685 2993.235 198.855 2993.395 ;
        RECT 201.405 2993.235 201.575 2993.395 ;
        RECT 201.745 2993.285 202.765 2993.615 ;
        RECT 204.125 2993.565 204.295 2993.795 ;
        RECT 198.685 2993.105 199.655 2993.235 ;
        RECT 198.855 2992.935 199.655 2993.105 ;
        RECT 198.685 2992.905 199.655 2992.935 ;
        RECT 200.255 2993.115 201.575 2993.235 ;
        RECT 200.255 2993.105 202.375 2993.115 ;
        RECT 200.255 2992.935 201.405 2993.105 ;
        RECT 201.575 2992.945 202.375 2993.105 ;
        RECT 200.255 2992.905 201.575 2992.935 ;
        RECT 198.685 2992.645 198.855 2992.905 ;
        RECT 201.405 2992.645 201.575 2992.905 ;
        RECT 202.595 2992.775 202.765 2993.285 ;
        RECT 198.685 2992.395 198.855 2992.475 ;
        RECT 201.405 2992.395 201.575 2992.475 ;
        RECT 201.745 2992.445 202.765 2992.775 ;
        RECT 198.685 2992.185 199.335 2992.395 ;
        RECT 200.605 2992.275 201.575 2992.395 ;
        RECT 202.595 2992.290 202.765 2992.445 ;
        RECT 203.305 2993.365 203.955 2993.535 ;
        RECT 203.305 2992.695 203.475 2993.365 ;
        RECT 204.125 2993.195 204.295 2993.395 ;
        RECT 203.645 2993.105 204.295 2993.195 ;
        RECT 203.645 2992.935 204.125 2993.105 ;
        RECT 203.645 2992.865 204.295 2992.935 ;
        RECT 203.305 2992.525 203.950 2992.695 ;
        RECT 204.125 2992.645 204.295 2992.865 ;
        RECT 203.305 2992.290 203.475 2992.525 ;
        RECT 204.125 2992.355 204.295 2992.475 ;
        RECT 198.855 2992.065 199.335 2992.185 ;
        RECT 198.685 2991.725 198.855 2992.015 ;
        RECT 198.685 2991.265 199.335 2991.555 ;
        RECT 198.855 2991.225 199.335 2991.265 ;
        RECT 198.685 2990.805 198.855 2991.095 ;
        RECT 198.855 2990.635 199.335 2990.715 ;
        RECT 198.685 2990.385 199.335 2990.635 ;
        RECT 198.685 2990.345 198.855 2990.385 ;
        RECT 198.685 2989.885 198.855 2990.175 ;
        RECT 198.855 2989.715 199.335 2989.875 ;
        RECT 199.845 2989.785 200.015 2992.235 ;
        RECT 200.605 2992.185 202.375 2992.275 ;
        RECT 200.605 2992.065 201.405 2992.185 ;
        RECT 201.575 2992.105 202.375 2992.185 ;
        RECT 202.595 2992.115 203.475 2992.290 ;
        RECT 203.645 2992.185 204.295 2992.355 ;
        RECT 201.405 2991.725 201.575 2992.015 ;
      LAYER li1 ;
        RECT 201.745 2991.685 202.765 2991.855 ;
      LAYER li1 ;
        RECT 200.605 2991.515 201.575 2991.555 ;
        RECT 200.605 2991.265 202.375 2991.515 ;
        RECT 200.605 2991.225 201.405 2991.265 ;
        RECT 201.575 2991.185 202.375 2991.265 ;
        RECT 201.405 2990.805 201.575 2991.095 ;
      LAYER li1 ;
        RECT 202.595 2991.015 202.765 2991.685 ;
        RECT 201.745 2990.845 202.765 2991.015 ;
      LAYER li1 ;
        RECT 200.605 2990.635 201.405 2990.715 ;
        RECT 201.575 2990.635 202.375 2990.675 ;
        RECT 200.605 2990.385 202.375 2990.635 ;
        RECT 201.405 2990.345 202.375 2990.385 ;
      LAYER li1 ;
        RECT 202.595 2990.175 202.765 2990.845 ;
      LAYER li1 ;
        RECT 201.405 2989.885 201.575 2990.175 ;
      LAYER li1 ;
        RECT 201.745 2990.005 202.765 2990.175 ;
      LAYER li1 ;
        RECT 198.685 2989.545 199.335 2989.715 ;
        RECT 199.505 2989.610 200.385 2989.785 ;
        RECT 200.605 2989.715 201.405 2989.795 ;
        RECT 201.575 2989.715 202.375 2989.835 ;
        RECT 200.605 2989.625 202.375 2989.715 ;
        RECT 198.685 2989.425 198.855 2989.545 ;
        RECT 199.505 2989.375 199.675 2989.610 ;
        RECT 200.215 2989.455 200.385 2989.610 ;
        RECT 201.405 2989.505 202.375 2989.625 ;
        RECT 198.685 2989.035 198.855 2989.255 ;
        RECT 199.030 2989.205 199.675 2989.375 ;
        RECT 198.685 2988.965 199.335 2989.035 ;
        RECT 198.855 2988.795 199.335 2988.965 ;
        RECT 198.685 2988.705 199.335 2988.795 ;
        RECT 198.685 2988.505 198.855 2988.705 ;
        RECT 199.505 2988.535 199.675 2989.205 ;
        RECT 199.025 2988.365 199.675 2988.535 ;
        RECT 198.685 2988.105 198.855 2988.335 ;
      LAYER li1 ;
        RECT 199.845 2988.330 200.045 2989.430 ;
      LAYER li1 ;
        RECT 200.215 2989.125 201.235 2989.455 ;
        RECT 201.405 2989.425 201.575 2989.505 ;
      LAYER li1 ;
        RECT 202.595 2989.420 202.765 2990.005 ;
      LAYER li1 ;
        RECT 202.965 2989.665 203.135 2992.115 ;
        RECT 203.645 2992.025 204.125 2992.185 ;
      LAYER li1 ;
        RECT 203.305 2991.685 203.955 2991.855 ;
      LAYER li1 ;
        RECT 204.125 2991.725 204.295 2992.015 ;
      LAYER li1 ;
        RECT 203.305 2991.015 203.475 2991.685 ;
      LAYER li1 ;
        RECT 204.125 2991.515 204.295 2991.555 ;
        RECT 203.645 2991.265 204.295 2991.515 ;
        RECT 203.645 2991.185 204.125 2991.265 ;
      LAYER li1 ;
        RECT 203.305 2990.845 203.955 2991.015 ;
        RECT 203.305 2990.175 203.475 2990.845 ;
      LAYER li1 ;
        RECT 204.125 2990.805 204.295 2991.095 ;
        RECT 203.645 2990.635 204.125 2990.675 ;
        RECT 203.645 2990.345 204.295 2990.635 ;
      LAYER li1 ;
        RECT 203.305 2990.005 203.955 2990.175 ;
        RECT 203.305 2989.420 203.475 2990.005 ;
      LAYER li1 ;
        RECT 204.125 2989.885 204.295 2990.175 ;
        RECT 203.645 2989.715 204.125 2989.835 ;
        RECT 203.645 2989.505 204.295 2989.715 ;
        RECT 204.125 2989.425 204.295 2989.505 ;
      LAYER li1 ;
        RECT 202.595 2989.335 203.475 2989.420 ;
      LAYER li1 ;
        RECT 200.215 2988.615 200.385 2989.125 ;
        RECT 201.405 2988.995 201.575 2989.255 ;
      LAYER li1 ;
        RECT 201.745 2989.165 203.955 2989.335 ;
      LAYER li1 ;
        RECT 204.125 2988.995 204.295 2989.255 ;
        RECT 201.405 2988.965 202.725 2988.995 ;
        RECT 200.605 2988.795 201.405 2988.955 ;
        RECT 201.575 2988.795 202.725 2988.965 ;
        RECT 200.605 2988.785 202.725 2988.795 ;
        RECT 201.405 2988.665 202.725 2988.785 ;
        RECT 203.325 2988.965 204.295 2988.995 ;
        RECT 203.325 2988.795 204.125 2988.965 ;
        RECT 203.325 2988.665 204.295 2988.795 ;
        RECT 200.215 2988.285 201.235 2988.615 ;
        RECT 201.405 2988.505 201.575 2988.665 ;
        RECT 204.125 2988.505 204.295 2988.665 ;
        RECT 201.405 2988.105 201.575 2988.335 ;
        RECT 204.125 2988.105 204.295 2988.335 ;
        RECT 198.685 2988.045 199.580 2988.105 ;
        RECT 198.855 2987.875 199.580 2988.045 ;
        RECT 198.685 2987.815 199.580 2987.875 ;
        RECT 200.240 2988.045 202.740 2988.105 ;
        RECT 200.240 2987.875 201.405 2988.045 ;
        RECT 201.575 2987.875 202.740 2988.045 ;
        RECT 200.240 2987.815 202.740 2987.875 ;
        RECT 203.400 2988.045 204.295 2988.105 ;
        RECT 203.400 2987.875 204.125 2988.045 ;
        RECT 203.400 2987.815 204.295 2987.875 ;
        RECT 198.685 2987.730 198.855 2987.815 ;
        RECT 201.405 2987.730 201.575 2987.815 ;
        RECT 204.125 2987.730 204.295 2987.815 ;
        RECT 3383.500 2268.195 3383.670 2268.280 ;
        RECT 3386.220 2268.195 3386.390 2268.280 ;
        RECT 3388.940 2268.195 3389.110 2268.280 ;
        RECT 3383.500 2268.135 3384.395 2268.195 ;
        RECT 3383.670 2267.965 3384.395 2268.135 ;
        RECT 3383.500 2267.905 3384.395 2267.965 ;
        RECT 3383.500 2267.675 3383.670 2267.905 ;
        RECT 3383.500 2267.305 3383.670 2267.505 ;
        RECT 3383.840 2267.475 3384.490 2267.645 ;
        RECT 3383.500 2267.215 3384.150 2267.305 ;
        RECT 3383.670 2267.045 3384.150 2267.215 ;
        RECT 3383.500 2266.975 3384.150 2267.045 ;
        RECT 3383.500 2266.755 3383.670 2266.975 ;
        RECT 3384.320 2266.805 3384.490 2267.475 ;
        RECT 3383.845 2266.635 3384.490 2266.805 ;
        RECT 3383.500 2266.465 3383.670 2266.585 ;
        RECT 3383.500 2266.295 3384.150 2266.465 ;
        RECT 3383.670 2266.135 3384.150 2266.295 ;
        RECT 3384.320 2266.400 3384.490 2266.635 ;
      LAYER li1 ;
        RECT 3384.660 2266.580 3384.860 2268.170 ;
      LAYER li1 ;
        RECT 3385.055 2268.135 3387.555 2268.195 ;
        RECT 3385.055 2267.965 3386.220 2268.135 ;
        RECT 3386.390 2267.965 3387.555 2268.135 ;
        RECT 3385.055 2267.905 3387.555 2267.965 ;
        RECT 3388.215 2268.135 3389.110 2268.195 ;
        RECT 3388.215 2267.965 3388.940 2268.135 ;
        RECT 3388.215 2267.905 3389.110 2267.965 ;
        RECT 3385.030 2267.395 3386.050 2267.725 ;
        RECT 3386.220 2267.675 3386.390 2267.905 ;
        RECT 3388.940 2267.675 3389.110 2267.905 ;
        RECT 3385.030 2266.885 3385.200 2267.395 ;
        RECT 3386.220 2267.345 3386.390 2267.505 ;
        RECT 3388.940 2267.345 3389.110 2267.505 ;
        RECT 3386.220 2267.225 3387.540 2267.345 ;
        RECT 3385.420 2267.215 3387.540 2267.225 ;
        RECT 3385.420 2267.055 3386.220 2267.215 ;
        RECT 3386.390 2267.045 3387.540 2267.215 ;
        RECT 3386.220 2267.015 3387.540 2267.045 ;
        RECT 3388.140 2267.215 3389.110 2267.345 ;
        RECT 3388.140 2267.045 3388.940 2267.215 ;
        RECT 3388.140 2267.015 3389.110 2267.045 ;
        RECT 3385.030 2266.555 3386.050 2266.885 ;
        RECT 3386.220 2266.755 3386.390 2267.015 ;
      LAYER li1 ;
        RECT 3386.560 2266.675 3388.770 2266.845 ;
      LAYER li1 ;
        RECT 3388.940 2266.755 3389.110 2267.015 ;
      LAYER li1 ;
        RECT 3387.410 2266.590 3388.290 2266.675 ;
      LAYER li1 ;
        RECT 3385.030 2266.400 3385.200 2266.555 ;
        RECT 3384.320 2266.225 3385.200 2266.400 ;
        RECT 3386.220 2266.505 3386.390 2266.585 ;
        RECT 3386.220 2266.385 3387.190 2266.505 ;
        RECT 3385.420 2266.295 3387.190 2266.385 ;
        RECT 3383.500 2265.835 3383.670 2266.125 ;
        RECT 3383.500 2265.625 3383.670 2265.665 ;
        RECT 3383.500 2265.375 3384.150 2265.625 ;
        RECT 3383.670 2265.295 3384.150 2265.375 ;
        RECT 3383.500 2264.915 3383.670 2265.205 ;
        RECT 3383.670 2264.745 3384.150 2264.785 ;
        RECT 3383.500 2264.455 3384.150 2264.745 ;
        RECT 3383.500 2263.995 3383.670 2264.285 ;
        RECT 3383.670 2263.825 3384.150 2263.945 ;
        RECT 3383.500 2263.615 3384.150 2263.825 ;
        RECT 3384.660 2263.775 3384.830 2266.225 ;
        RECT 3385.420 2266.215 3386.220 2266.295 ;
        RECT 3386.390 2266.175 3387.190 2266.295 ;
        RECT 3386.220 2265.835 3386.390 2266.125 ;
      LAYER li1 ;
        RECT 3387.410 2266.005 3387.580 2266.590 ;
        RECT 3386.560 2265.835 3387.580 2266.005 ;
      LAYER li1 ;
        RECT 3386.220 2265.625 3387.190 2265.665 ;
        RECT 3385.420 2265.375 3387.190 2265.625 ;
        RECT 3385.420 2265.295 3386.220 2265.375 ;
        RECT 3386.390 2265.335 3387.190 2265.375 ;
        RECT 3386.220 2264.915 3386.390 2265.205 ;
      LAYER li1 ;
        RECT 3387.410 2265.165 3387.580 2265.835 ;
        RECT 3386.560 2264.995 3387.580 2265.165 ;
      LAYER li1 ;
        RECT 3385.420 2264.745 3386.220 2264.785 ;
        RECT 3386.390 2264.745 3387.190 2264.825 ;
        RECT 3385.420 2264.495 3387.190 2264.745 ;
        RECT 3385.420 2264.455 3386.390 2264.495 ;
      LAYER li1 ;
        RECT 3387.410 2264.325 3387.580 2264.995 ;
      LAYER li1 ;
        RECT 3386.220 2263.995 3386.390 2264.285 ;
      LAYER li1 ;
        RECT 3386.560 2264.155 3387.580 2264.325 ;
      LAYER li1 ;
        RECT 3385.420 2263.825 3386.220 2263.945 ;
        RECT 3386.390 2263.825 3387.190 2263.905 ;
        RECT 3387.780 2263.895 3387.950 2266.345 ;
      LAYER li1 ;
        RECT 3388.120 2266.005 3388.290 2266.590 ;
      LAYER li1 ;
        RECT 3388.940 2266.505 3389.110 2266.585 ;
        RECT 3388.460 2266.295 3389.110 2266.505 ;
        RECT 3388.460 2266.175 3388.940 2266.295 ;
      LAYER li1 ;
        RECT 3388.120 2265.835 3388.770 2266.005 ;
      LAYER li1 ;
        RECT 3388.940 2265.835 3389.110 2266.125 ;
      LAYER li1 ;
        RECT 3388.120 2265.165 3388.290 2265.835 ;
      LAYER li1 ;
        RECT 3388.460 2265.375 3389.110 2265.665 ;
        RECT 3388.460 2265.335 3388.940 2265.375 ;
      LAYER li1 ;
        RECT 3388.120 2264.995 3388.770 2265.165 ;
        RECT 3388.120 2264.325 3388.290 2264.995 ;
      LAYER li1 ;
        RECT 3388.940 2264.915 3389.110 2265.205 ;
        RECT 3388.460 2264.745 3388.940 2264.825 ;
        RECT 3388.460 2264.495 3389.110 2264.745 ;
        RECT 3388.940 2264.455 3389.110 2264.495 ;
      LAYER li1 ;
        RECT 3388.120 2264.155 3388.770 2264.325 ;
      LAYER li1 ;
        RECT 3388.940 2263.995 3389.110 2264.285 ;
        RECT 3385.420 2263.735 3387.190 2263.825 ;
        RECT 3385.420 2263.615 3386.390 2263.735 ;
        RECT 3383.500 2263.535 3383.670 2263.615 ;
        RECT 3386.220 2263.535 3386.390 2263.615 ;
        RECT 3387.410 2263.720 3388.290 2263.895 ;
        RECT 3387.410 2263.565 3387.580 2263.720 ;
        RECT 3383.500 2263.105 3383.670 2263.365 ;
        RECT 3386.220 2263.105 3386.390 2263.365 ;
        RECT 3386.560 2263.235 3387.580 2263.565 ;
        RECT 3383.500 2263.075 3384.470 2263.105 ;
        RECT 3383.670 2262.905 3384.470 2263.075 ;
        RECT 3383.500 2262.775 3384.470 2262.905 ;
        RECT 3385.070 2263.075 3386.390 2263.105 ;
        RECT 3385.070 2262.905 3386.220 2263.075 ;
        RECT 3386.390 2262.905 3387.190 2263.065 ;
        RECT 3385.070 2262.895 3387.190 2262.905 ;
        RECT 3385.070 2262.775 3386.390 2262.895 ;
        RECT 3383.500 2262.615 3383.670 2262.775 ;
        RECT 3386.220 2262.615 3386.390 2262.775 ;
        RECT 3387.410 2262.725 3387.580 2263.235 ;
        RECT 3383.500 2262.215 3383.670 2262.445 ;
        RECT 3386.220 2262.215 3386.390 2262.445 ;
        RECT 3386.560 2262.395 3387.580 2262.725 ;
        RECT 3388.120 2263.485 3388.290 2263.720 ;
        RECT 3388.460 2263.825 3388.940 2263.985 ;
        RECT 3388.460 2263.655 3389.110 2263.825 ;
        RECT 3388.940 2263.535 3389.110 2263.655 ;
        RECT 3388.120 2263.315 3388.765 2263.485 ;
        RECT 3388.120 2262.645 3388.290 2263.315 ;
        RECT 3388.940 2263.145 3389.110 2263.365 ;
        RECT 3388.460 2263.075 3389.110 2263.145 ;
        RECT 3388.460 2262.905 3388.940 2263.075 ;
        RECT 3388.460 2262.815 3389.110 2262.905 ;
        RECT 3388.120 2262.475 3388.770 2262.645 ;
        RECT 3388.940 2262.615 3389.110 2262.815 ;
        RECT 3388.940 2262.215 3389.110 2262.445 ;
        RECT 3383.500 2262.155 3384.395 2262.215 ;
        RECT 3383.670 2261.985 3384.395 2262.155 ;
        RECT 3383.500 2261.925 3384.395 2261.985 ;
        RECT 3383.500 2261.695 3383.670 2261.925 ;
        RECT 3383.500 2261.325 3383.670 2261.525 ;
        RECT 3383.840 2261.495 3384.490 2261.665 ;
        RECT 3383.500 2261.235 3384.150 2261.325 ;
        RECT 3383.670 2261.065 3384.150 2261.235 ;
        RECT 3383.500 2260.995 3384.150 2261.065 ;
        RECT 3383.500 2260.775 3383.670 2260.995 ;
        RECT 3384.320 2260.825 3384.490 2261.495 ;
        RECT 3383.845 2260.655 3384.490 2260.825 ;
        RECT 3383.500 2260.485 3383.670 2260.605 ;
        RECT 3383.500 2260.315 3384.150 2260.485 ;
        RECT 3383.670 2260.155 3384.150 2260.315 ;
        RECT 3384.320 2260.420 3384.490 2260.655 ;
      LAYER li1 ;
        RECT 3384.660 2260.600 3384.860 2262.190 ;
      LAYER li1 ;
        RECT 3385.055 2262.155 3387.555 2262.215 ;
        RECT 3385.055 2261.985 3386.220 2262.155 ;
        RECT 3386.390 2261.985 3387.555 2262.155 ;
        RECT 3385.055 2261.925 3387.555 2261.985 ;
        RECT 3388.215 2262.155 3389.110 2262.215 ;
        RECT 3388.215 2261.985 3388.940 2262.155 ;
        RECT 3388.215 2261.925 3389.110 2261.985 ;
        RECT 3385.030 2261.415 3386.050 2261.745 ;
        RECT 3386.220 2261.695 3386.390 2261.925 ;
        RECT 3388.940 2261.695 3389.110 2261.925 ;
        RECT 3385.030 2260.905 3385.200 2261.415 ;
        RECT 3386.220 2261.365 3386.390 2261.525 ;
        RECT 3388.940 2261.365 3389.110 2261.525 ;
        RECT 3386.220 2261.245 3387.540 2261.365 ;
        RECT 3385.420 2261.235 3387.540 2261.245 ;
        RECT 3385.420 2261.075 3386.220 2261.235 ;
        RECT 3386.390 2261.065 3387.540 2261.235 ;
        RECT 3386.220 2261.035 3387.540 2261.065 ;
        RECT 3388.140 2261.235 3389.110 2261.365 ;
        RECT 3388.140 2261.065 3388.940 2261.235 ;
        RECT 3388.140 2261.035 3389.110 2261.065 ;
        RECT 3385.030 2260.575 3386.050 2260.905 ;
        RECT 3386.220 2260.775 3386.390 2261.035 ;
      LAYER li1 ;
        RECT 3386.560 2260.695 3388.770 2260.865 ;
      LAYER li1 ;
        RECT 3388.940 2260.775 3389.110 2261.035 ;
      LAYER li1 ;
        RECT 3387.410 2260.610 3388.290 2260.695 ;
      LAYER li1 ;
        RECT 3385.030 2260.420 3385.200 2260.575 ;
        RECT 3384.320 2260.245 3385.200 2260.420 ;
        RECT 3386.220 2260.525 3386.390 2260.605 ;
        RECT 3386.220 2260.405 3387.190 2260.525 ;
        RECT 3385.420 2260.315 3387.190 2260.405 ;
        RECT 3383.500 2259.855 3383.670 2260.145 ;
        RECT 3383.500 2259.645 3383.670 2259.685 ;
        RECT 3383.500 2259.395 3384.150 2259.645 ;
        RECT 3383.670 2259.315 3384.150 2259.395 ;
        RECT 3383.500 2258.935 3383.670 2259.225 ;
        RECT 3383.670 2258.765 3384.150 2258.805 ;
        RECT 3383.500 2258.475 3384.150 2258.765 ;
        RECT 3383.500 2258.015 3383.670 2258.305 ;
        RECT 3383.670 2257.845 3384.150 2257.965 ;
        RECT 3383.500 2257.635 3384.150 2257.845 ;
        RECT 3384.660 2257.795 3384.830 2260.245 ;
        RECT 3385.420 2260.235 3386.220 2260.315 ;
        RECT 3386.390 2260.195 3387.190 2260.315 ;
        RECT 3386.220 2259.855 3386.390 2260.145 ;
      LAYER li1 ;
        RECT 3387.410 2260.025 3387.580 2260.610 ;
        RECT 3386.560 2259.855 3387.580 2260.025 ;
      LAYER li1 ;
        RECT 3386.220 2259.645 3387.190 2259.685 ;
        RECT 3385.420 2259.395 3387.190 2259.645 ;
        RECT 3385.420 2259.315 3386.220 2259.395 ;
        RECT 3386.390 2259.355 3387.190 2259.395 ;
        RECT 3386.220 2258.935 3386.390 2259.225 ;
      LAYER li1 ;
        RECT 3387.410 2259.185 3387.580 2259.855 ;
        RECT 3386.560 2259.015 3387.580 2259.185 ;
      LAYER li1 ;
        RECT 3385.420 2258.765 3386.220 2258.805 ;
        RECT 3386.390 2258.765 3387.190 2258.845 ;
        RECT 3385.420 2258.515 3387.190 2258.765 ;
        RECT 3385.420 2258.475 3386.390 2258.515 ;
      LAYER li1 ;
        RECT 3387.410 2258.345 3387.580 2259.015 ;
      LAYER li1 ;
        RECT 3386.220 2258.015 3386.390 2258.305 ;
      LAYER li1 ;
        RECT 3386.560 2258.175 3387.580 2258.345 ;
      LAYER li1 ;
        RECT 3385.420 2257.845 3386.220 2257.965 ;
        RECT 3386.390 2257.845 3387.190 2257.925 ;
        RECT 3387.780 2257.915 3387.950 2260.365 ;
      LAYER li1 ;
        RECT 3388.120 2260.025 3388.290 2260.610 ;
      LAYER li1 ;
        RECT 3388.940 2260.525 3389.110 2260.605 ;
        RECT 3388.460 2260.315 3389.110 2260.525 ;
        RECT 3388.460 2260.195 3388.940 2260.315 ;
      LAYER li1 ;
        RECT 3388.120 2259.855 3388.770 2260.025 ;
      LAYER li1 ;
        RECT 3388.940 2259.855 3389.110 2260.145 ;
      LAYER li1 ;
        RECT 3388.120 2259.185 3388.290 2259.855 ;
      LAYER li1 ;
        RECT 3388.460 2259.395 3389.110 2259.685 ;
        RECT 3388.460 2259.355 3388.940 2259.395 ;
      LAYER li1 ;
        RECT 3388.120 2259.015 3388.770 2259.185 ;
        RECT 3388.120 2258.345 3388.290 2259.015 ;
      LAYER li1 ;
        RECT 3388.940 2258.935 3389.110 2259.225 ;
        RECT 3388.460 2258.765 3388.940 2258.845 ;
        RECT 3388.460 2258.515 3389.110 2258.765 ;
        RECT 3388.940 2258.475 3389.110 2258.515 ;
      LAYER li1 ;
        RECT 3388.120 2258.175 3388.770 2258.345 ;
      LAYER li1 ;
        RECT 3388.940 2258.015 3389.110 2258.305 ;
        RECT 3385.420 2257.755 3387.190 2257.845 ;
        RECT 3385.420 2257.635 3386.390 2257.755 ;
        RECT 3383.500 2257.555 3383.670 2257.635 ;
        RECT 3386.220 2257.555 3386.390 2257.635 ;
        RECT 3387.410 2257.740 3388.290 2257.915 ;
        RECT 3387.410 2257.585 3387.580 2257.740 ;
        RECT 3383.500 2257.125 3383.670 2257.385 ;
        RECT 3386.220 2257.125 3386.390 2257.385 ;
        RECT 3386.560 2257.255 3387.580 2257.585 ;
        RECT 3383.500 2257.095 3384.470 2257.125 ;
        RECT 3383.670 2256.925 3384.470 2257.095 ;
        RECT 3383.500 2256.795 3384.470 2256.925 ;
        RECT 3385.070 2257.095 3386.390 2257.125 ;
        RECT 3385.070 2256.925 3386.220 2257.095 ;
        RECT 3386.390 2256.925 3387.190 2257.085 ;
        RECT 3385.070 2256.915 3387.190 2256.925 ;
        RECT 3385.070 2256.795 3386.390 2256.915 ;
        RECT 3383.500 2256.635 3383.670 2256.795 ;
        RECT 3386.220 2256.635 3386.390 2256.795 ;
        RECT 3387.410 2256.745 3387.580 2257.255 ;
        RECT 3383.500 2256.235 3383.670 2256.465 ;
        RECT 3386.220 2256.235 3386.390 2256.465 ;
        RECT 3386.560 2256.415 3387.580 2256.745 ;
        RECT 3388.120 2257.505 3388.290 2257.740 ;
        RECT 3388.460 2257.845 3388.940 2258.005 ;
        RECT 3388.460 2257.675 3389.110 2257.845 ;
        RECT 3388.940 2257.555 3389.110 2257.675 ;
        RECT 3388.120 2257.335 3388.765 2257.505 ;
        RECT 3388.120 2256.665 3388.290 2257.335 ;
        RECT 3388.940 2257.165 3389.110 2257.385 ;
        RECT 3388.460 2257.095 3389.110 2257.165 ;
        RECT 3388.460 2256.925 3388.940 2257.095 ;
        RECT 3388.460 2256.835 3389.110 2256.925 ;
        RECT 3388.120 2256.495 3388.770 2256.665 ;
        RECT 3388.940 2256.635 3389.110 2256.835 ;
        RECT 3388.940 2256.235 3389.110 2256.465 ;
        RECT 3383.500 2256.175 3384.395 2256.235 ;
        RECT 3383.670 2256.005 3384.395 2256.175 ;
        RECT 3383.500 2255.945 3384.395 2256.005 ;
        RECT 3383.500 2255.715 3383.670 2255.945 ;
        RECT 3383.500 2255.345 3383.670 2255.545 ;
        RECT 3383.840 2255.515 3384.490 2255.685 ;
        RECT 3383.500 2255.255 3384.150 2255.345 ;
        RECT 3383.670 2255.085 3384.150 2255.255 ;
        RECT 3383.500 2255.015 3384.150 2255.085 ;
        RECT 3383.500 2254.795 3383.670 2255.015 ;
        RECT 3384.320 2254.845 3384.490 2255.515 ;
        RECT 3383.845 2254.675 3384.490 2254.845 ;
        RECT 3383.500 2254.505 3383.670 2254.625 ;
        RECT 3383.500 2254.335 3384.150 2254.505 ;
        RECT 3383.670 2254.175 3384.150 2254.335 ;
        RECT 3384.320 2254.440 3384.490 2254.675 ;
      LAYER li1 ;
        RECT 3384.660 2254.620 3384.860 2256.210 ;
      LAYER li1 ;
        RECT 3385.055 2256.175 3387.555 2256.235 ;
        RECT 3385.055 2256.005 3386.220 2256.175 ;
        RECT 3386.390 2256.005 3387.555 2256.175 ;
        RECT 3385.055 2255.945 3387.555 2256.005 ;
        RECT 3388.215 2256.175 3389.110 2256.235 ;
        RECT 3388.215 2256.005 3388.940 2256.175 ;
        RECT 3388.215 2255.945 3389.110 2256.005 ;
        RECT 3385.030 2255.435 3386.050 2255.765 ;
        RECT 3386.220 2255.715 3386.390 2255.945 ;
        RECT 3388.940 2255.715 3389.110 2255.945 ;
        RECT 3385.030 2254.925 3385.200 2255.435 ;
        RECT 3386.220 2255.385 3386.390 2255.545 ;
        RECT 3388.940 2255.385 3389.110 2255.545 ;
        RECT 3386.220 2255.265 3387.540 2255.385 ;
        RECT 3385.420 2255.255 3387.540 2255.265 ;
        RECT 3385.420 2255.095 3386.220 2255.255 ;
        RECT 3386.390 2255.085 3387.540 2255.255 ;
        RECT 3386.220 2255.055 3387.540 2255.085 ;
        RECT 3388.140 2255.255 3389.110 2255.385 ;
        RECT 3388.140 2255.085 3388.940 2255.255 ;
        RECT 3388.140 2255.055 3389.110 2255.085 ;
        RECT 3385.030 2254.595 3386.050 2254.925 ;
        RECT 3386.220 2254.795 3386.390 2255.055 ;
      LAYER li1 ;
        RECT 3386.560 2254.715 3388.770 2254.885 ;
      LAYER li1 ;
        RECT 3388.940 2254.795 3389.110 2255.055 ;
      LAYER li1 ;
        RECT 3387.410 2254.630 3388.290 2254.715 ;
      LAYER li1 ;
        RECT 3385.030 2254.440 3385.200 2254.595 ;
        RECT 3384.320 2254.265 3385.200 2254.440 ;
        RECT 3386.220 2254.545 3386.390 2254.625 ;
        RECT 3386.220 2254.425 3387.190 2254.545 ;
        RECT 3385.420 2254.335 3387.190 2254.425 ;
        RECT 3383.500 2253.875 3383.670 2254.165 ;
        RECT 3383.500 2253.665 3383.670 2253.705 ;
        RECT 3383.500 2253.415 3384.150 2253.665 ;
        RECT 3383.670 2253.335 3384.150 2253.415 ;
        RECT 3383.500 2252.955 3383.670 2253.245 ;
        RECT 3383.670 2252.785 3384.150 2252.825 ;
        RECT 3383.500 2252.495 3384.150 2252.785 ;
        RECT 3383.500 2252.035 3383.670 2252.325 ;
        RECT 3383.670 2251.865 3384.150 2251.985 ;
        RECT 3383.500 2251.655 3384.150 2251.865 ;
        RECT 3384.660 2251.815 3384.830 2254.265 ;
        RECT 3385.420 2254.255 3386.220 2254.335 ;
        RECT 3386.390 2254.215 3387.190 2254.335 ;
        RECT 3386.220 2253.875 3386.390 2254.165 ;
      LAYER li1 ;
        RECT 3387.410 2254.045 3387.580 2254.630 ;
        RECT 3386.560 2253.875 3387.580 2254.045 ;
      LAYER li1 ;
        RECT 3386.220 2253.665 3387.190 2253.705 ;
        RECT 3385.420 2253.415 3387.190 2253.665 ;
        RECT 3385.420 2253.335 3386.220 2253.415 ;
        RECT 3386.390 2253.375 3387.190 2253.415 ;
        RECT 3386.220 2252.955 3386.390 2253.245 ;
      LAYER li1 ;
        RECT 3387.410 2253.205 3387.580 2253.875 ;
        RECT 3386.560 2253.035 3387.580 2253.205 ;
      LAYER li1 ;
        RECT 3385.420 2252.785 3386.220 2252.825 ;
        RECT 3386.390 2252.785 3387.190 2252.865 ;
        RECT 3385.420 2252.535 3387.190 2252.785 ;
        RECT 3385.420 2252.495 3386.390 2252.535 ;
      LAYER li1 ;
        RECT 3387.410 2252.365 3387.580 2253.035 ;
      LAYER li1 ;
        RECT 3386.220 2252.035 3386.390 2252.325 ;
      LAYER li1 ;
        RECT 3386.560 2252.195 3387.580 2252.365 ;
      LAYER li1 ;
        RECT 3385.420 2251.865 3386.220 2251.985 ;
        RECT 3386.390 2251.865 3387.190 2251.945 ;
        RECT 3387.780 2251.935 3387.950 2254.385 ;
      LAYER li1 ;
        RECT 3388.120 2254.045 3388.290 2254.630 ;
      LAYER li1 ;
        RECT 3388.940 2254.545 3389.110 2254.625 ;
        RECT 3388.460 2254.335 3389.110 2254.545 ;
        RECT 3388.460 2254.215 3388.940 2254.335 ;
      LAYER li1 ;
        RECT 3388.120 2253.875 3388.770 2254.045 ;
      LAYER li1 ;
        RECT 3388.940 2253.875 3389.110 2254.165 ;
      LAYER li1 ;
        RECT 3388.120 2253.205 3388.290 2253.875 ;
      LAYER li1 ;
        RECT 3388.460 2253.415 3389.110 2253.705 ;
        RECT 3388.460 2253.375 3388.940 2253.415 ;
      LAYER li1 ;
        RECT 3388.120 2253.035 3388.770 2253.205 ;
        RECT 3388.120 2252.365 3388.290 2253.035 ;
      LAYER li1 ;
        RECT 3388.940 2252.955 3389.110 2253.245 ;
        RECT 3388.460 2252.785 3388.940 2252.865 ;
        RECT 3388.460 2252.535 3389.110 2252.785 ;
        RECT 3388.940 2252.495 3389.110 2252.535 ;
      LAYER li1 ;
        RECT 3388.120 2252.195 3388.770 2252.365 ;
      LAYER li1 ;
        RECT 3388.940 2252.035 3389.110 2252.325 ;
        RECT 3385.420 2251.775 3387.190 2251.865 ;
        RECT 3385.420 2251.655 3386.390 2251.775 ;
        RECT 3383.500 2251.575 3383.670 2251.655 ;
        RECT 3386.220 2251.575 3386.390 2251.655 ;
        RECT 3387.410 2251.760 3388.290 2251.935 ;
        RECT 3387.410 2251.605 3387.580 2251.760 ;
        RECT 3383.500 2251.145 3383.670 2251.405 ;
        RECT 3386.220 2251.145 3386.390 2251.405 ;
        RECT 3386.560 2251.275 3387.580 2251.605 ;
        RECT 3383.500 2251.115 3384.470 2251.145 ;
        RECT 3383.670 2250.945 3384.470 2251.115 ;
        RECT 3383.500 2250.815 3384.470 2250.945 ;
        RECT 3385.070 2251.115 3386.390 2251.145 ;
        RECT 3385.070 2250.945 3386.220 2251.115 ;
        RECT 3386.390 2250.945 3387.190 2251.105 ;
        RECT 3385.070 2250.935 3387.190 2250.945 ;
        RECT 3385.070 2250.815 3386.390 2250.935 ;
        RECT 3383.500 2250.655 3383.670 2250.815 ;
        RECT 3386.220 2250.655 3386.390 2250.815 ;
        RECT 3387.410 2250.765 3387.580 2251.275 ;
        RECT 3383.500 2250.255 3383.670 2250.485 ;
        RECT 3386.220 2250.255 3386.390 2250.485 ;
        RECT 3386.560 2250.435 3387.580 2250.765 ;
        RECT 3388.120 2251.525 3388.290 2251.760 ;
        RECT 3388.460 2251.865 3388.940 2252.025 ;
        RECT 3388.460 2251.695 3389.110 2251.865 ;
        RECT 3388.940 2251.575 3389.110 2251.695 ;
        RECT 3388.120 2251.355 3388.765 2251.525 ;
        RECT 3388.120 2250.685 3388.290 2251.355 ;
        RECT 3388.940 2251.185 3389.110 2251.405 ;
        RECT 3388.460 2251.115 3389.110 2251.185 ;
        RECT 3388.460 2250.945 3388.940 2251.115 ;
        RECT 3388.460 2250.855 3389.110 2250.945 ;
        RECT 3388.120 2250.515 3388.770 2250.685 ;
        RECT 3388.940 2250.655 3389.110 2250.855 ;
        RECT 3388.940 2250.255 3389.110 2250.485 ;
        RECT 3383.500 2250.195 3384.395 2250.255 ;
        RECT 3383.670 2250.025 3384.395 2250.195 ;
        RECT 3383.500 2249.965 3384.395 2250.025 ;
        RECT 3383.500 2249.735 3383.670 2249.965 ;
        RECT 3383.500 2249.365 3383.670 2249.565 ;
        RECT 3383.840 2249.535 3384.490 2249.705 ;
        RECT 3383.500 2249.275 3384.150 2249.365 ;
        RECT 3383.670 2249.105 3384.150 2249.275 ;
        RECT 3383.500 2249.035 3384.150 2249.105 ;
        RECT 3383.500 2248.815 3383.670 2249.035 ;
        RECT 3384.320 2248.865 3384.490 2249.535 ;
        RECT 3383.845 2248.695 3384.490 2248.865 ;
        RECT 3383.500 2248.525 3383.670 2248.645 ;
        RECT 3383.500 2248.355 3384.150 2248.525 ;
        RECT 3383.670 2248.195 3384.150 2248.355 ;
        RECT 3384.320 2248.460 3384.490 2248.695 ;
      LAYER li1 ;
        RECT 3384.660 2248.640 3384.860 2250.230 ;
      LAYER li1 ;
        RECT 3385.055 2250.195 3387.555 2250.255 ;
        RECT 3385.055 2250.025 3386.220 2250.195 ;
        RECT 3386.390 2250.025 3387.555 2250.195 ;
        RECT 3385.055 2249.965 3387.555 2250.025 ;
        RECT 3388.215 2250.195 3389.110 2250.255 ;
        RECT 3388.215 2250.025 3388.940 2250.195 ;
        RECT 3388.215 2249.965 3389.110 2250.025 ;
        RECT 3385.030 2249.455 3386.050 2249.785 ;
        RECT 3386.220 2249.735 3386.390 2249.965 ;
        RECT 3388.940 2249.735 3389.110 2249.965 ;
        RECT 3385.030 2248.945 3385.200 2249.455 ;
        RECT 3386.220 2249.405 3386.390 2249.565 ;
        RECT 3388.940 2249.405 3389.110 2249.565 ;
        RECT 3386.220 2249.285 3387.540 2249.405 ;
        RECT 3385.420 2249.275 3387.540 2249.285 ;
        RECT 3385.420 2249.115 3386.220 2249.275 ;
        RECT 3386.390 2249.105 3387.540 2249.275 ;
        RECT 3386.220 2249.075 3387.540 2249.105 ;
        RECT 3388.140 2249.275 3389.110 2249.405 ;
        RECT 3388.140 2249.105 3388.940 2249.275 ;
        RECT 3388.140 2249.075 3389.110 2249.105 ;
        RECT 3385.030 2248.615 3386.050 2248.945 ;
        RECT 3386.220 2248.815 3386.390 2249.075 ;
      LAYER li1 ;
        RECT 3386.560 2248.735 3388.770 2248.905 ;
      LAYER li1 ;
        RECT 3388.940 2248.815 3389.110 2249.075 ;
      LAYER li1 ;
        RECT 3387.410 2248.650 3388.290 2248.735 ;
      LAYER li1 ;
        RECT 3385.030 2248.460 3385.200 2248.615 ;
        RECT 3384.320 2248.285 3385.200 2248.460 ;
        RECT 3386.220 2248.565 3386.390 2248.645 ;
        RECT 3386.220 2248.445 3387.190 2248.565 ;
        RECT 3385.420 2248.355 3387.190 2248.445 ;
        RECT 3383.500 2247.895 3383.670 2248.185 ;
        RECT 3383.500 2247.685 3383.670 2247.725 ;
        RECT 3383.500 2247.435 3384.150 2247.685 ;
        RECT 3383.670 2247.355 3384.150 2247.435 ;
        RECT 3383.500 2246.975 3383.670 2247.265 ;
        RECT 3383.670 2246.805 3384.150 2246.845 ;
        RECT 3383.500 2246.515 3384.150 2246.805 ;
        RECT 3383.500 2246.055 3383.670 2246.345 ;
        RECT 3383.670 2245.885 3384.150 2246.005 ;
        RECT 3383.500 2245.675 3384.150 2245.885 ;
        RECT 3384.660 2245.835 3384.830 2248.285 ;
        RECT 3385.420 2248.275 3386.220 2248.355 ;
        RECT 3386.390 2248.235 3387.190 2248.355 ;
        RECT 3386.220 2247.895 3386.390 2248.185 ;
      LAYER li1 ;
        RECT 3387.410 2248.065 3387.580 2248.650 ;
        RECT 3386.560 2247.895 3387.580 2248.065 ;
      LAYER li1 ;
        RECT 3386.220 2247.685 3387.190 2247.725 ;
        RECT 3385.420 2247.435 3387.190 2247.685 ;
        RECT 3385.420 2247.355 3386.220 2247.435 ;
        RECT 3386.390 2247.395 3387.190 2247.435 ;
        RECT 3386.220 2246.975 3386.390 2247.265 ;
      LAYER li1 ;
        RECT 3387.410 2247.225 3387.580 2247.895 ;
        RECT 3386.560 2247.055 3387.580 2247.225 ;
      LAYER li1 ;
        RECT 3385.420 2246.805 3386.220 2246.845 ;
        RECT 3386.390 2246.805 3387.190 2246.885 ;
        RECT 3385.420 2246.555 3387.190 2246.805 ;
        RECT 3385.420 2246.515 3386.390 2246.555 ;
      LAYER li1 ;
        RECT 3387.410 2246.385 3387.580 2247.055 ;
      LAYER li1 ;
        RECT 3386.220 2246.055 3386.390 2246.345 ;
      LAYER li1 ;
        RECT 3386.560 2246.215 3387.580 2246.385 ;
      LAYER li1 ;
        RECT 3385.420 2245.885 3386.220 2246.005 ;
        RECT 3386.390 2245.885 3387.190 2245.965 ;
        RECT 3387.780 2245.955 3387.950 2248.405 ;
      LAYER li1 ;
        RECT 3388.120 2248.065 3388.290 2248.650 ;
      LAYER li1 ;
        RECT 3388.940 2248.565 3389.110 2248.645 ;
        RECT 3388.460 2248.355 3389.110 2248.565 ;
        RECT 3388.460 2248.235 3388.940 2248.355 ;
      LAYER li1 ;
        RECT 3388.120 2247.895 3388.770 2248.065 ;
      LAYER li1 ;
        RECT 3388.940 2247.895 3389.110 2248.185 ;
      LAYER li1 ;
        RECT 3388.120 2247.225 3388.290 2247.895 ;
      LAYER li1 ;
        RECT 3388.460 2247.435 3389.110 2247.725 ;
        RECT 3388.460 2247.395 3388.940 2247.435 ;
      LAYER li1 ;
        RECT 3388.120 2247.055 3388.770 2247.225 ;
        RECT 3388.120 2246.385 3388.290 2247.055 ;
      LAYER li1 ;
        RECT 3388.940 2246.975 3389.110 2247.265 ;
        RECT 3388.460 2246.805 3388.940 2246.885 ;
        RECT 3388.460 2246.555 3389.110 2246.805 ;
        RECT 3388.940 2246.515 3389.110 2246.555 ;
      LAYER li1 ;
        RECT 3388.120 2246.215 3388.770 2246.385 ;
      LAYER li1 ;
        RECT 3388.940 2246.055 3389.110 2246.345 ;
        RECT 3385.420 2245.795 3387.190 2245.885 ;
        RECT 3385.420 2245.675 3386.390 2245.795 ;
        RECT 3383.500 2245.595 3383.670 2245.675 ;
        RECT 3386.220 2245.595 3386.390 2245.675 ;
        RECT 3387.410 2245.780 3388.290 2245.955 ;
        RECT 3387.410 2245.625 3387.580 2245.780 ;
        RECT 3383.500 2245.165 3383.670 2245.425 ;
        RECT 3386.220 2245.165 3386.390 2245.425 ;
        RECT 3386.560 2245.295 3387.580 2245.625 ;
        RECT 3383.500 2245.135 3384.470 2245.165 ;
        RECT 3383.670 2244.965 3384.470 2245.135 ;
        RECT 3383.500 2244.835 3384.470 2244.965 ;
        RECT 3385.070 2245.135 3386.390 2245.165 ;
        RECT 3385.070 2244.965 3386.220 2245.135 ;
        RECT 3386.390 2244.965 3387.190 2245.125 ;
        RECT 3385.070 2244.955 3387.190 2244.965 ;
        RECT 3385.070 2244.835 3386.390 2244.955 ;
        RECT 3383.500 2244.675 3383.670 2244.835 ;
        RECT 3386.220 2244.675 3386.390 2244.835 ;
        RECT 3387.410 2244.785 3387.580 2245.295 ;
        RECT 3383.500 2244.275 3383.670 2244.505 ;
        RECT 3386.220 2244.275 3386.390 2244.505 ;
        RECT 3386.560 2244.455 3387.580 2244.785 ;
        RECT 3388.120 2245.545 3388.290 2245.780 ;
        RECT 3388.460 2245.885 3388.940 2246.045 ;
        RECT 3388.460 2245.715 3389.110 2245.885 ;
        RECT 3388.940 2245.595 3389.110 2245.715 ;
        RECT 3388.120 2245.375 3388.765 2245.545 ;
        RECT 3388.120 2244.705 3388.290 2245.375 ;
        RECT 3388.940 2245.205 3389.110 2245.425 ;
        RECT 3388.460 2245.135 3389.110 2245.205 ;
        RECT 3388.460 2244.965 3388.940 2245.135 ;
        RECT 3388.460 2244.875 3389.110 2244.965 ;
        RECT 3388.120 2244.535 3388.770 2244.705 ;
        RECT 3388.940 2244.675 3389.110 2244.875 ;
        RECT 3388.940 2244.275 3389.110 2244.505 ;
        RECT 3383.500 2244.215 3384.395 2244.275 ;
        RECT 3383.670 2244.045 3384.395 2244.215 ;
        RECT 3383.500 2243.985 3384.395 2244.045 ;
        RECT 3383.500 2243.755 3383.670 2243.985 ;
        RECT 3383.500 2243.385 3383.670 2243.585 ;
        RECT 3383.840 2243.555 3384.490 2243.725 ;
        RECT 3383.500 2243.295 3384.150 2243.385 ;
        RECT 3383.670 2243.125 3384.150 2243.295 ;
        RECT 3383.500 2243.055 3384.150 2243.125 ;
        RECT 3383.500 2242.835 3383.670 2243.055 ;
        RECT 3384.320 2242.885 3384.490 2243.555 ;
        RECT 3383.845 2242.715 3384.490 2242.885 ;
        RECT 3383.500 2242.545 3383.670 2242.665 ;
        RECT 3383.500 2242.375 3384.150 2242.545 ;
        RECT 3383.670 2242.215 3384.150 2242.375 ;
        RECT 3384.320 2242.480 3384.490 2242.715 ;
      LAYER li1 ;
        RECT 3384.660 2242.660 3384.860 2244.250 ;
      LAYER li1 ;
        RECT 3385.055 2244.215 3387.555 2244.275 ;
        RECT 3385.055 2244.045 3386.220 2244.215 ;
        RECT 3386.390 2244.045 3387.555 2244.215 ;
        RECT 3385.055 2243.985 3387.555 2244.045 ;
        RECT 3388.215 2244.215 3389.110 2244.275 ;
        RECT 3388.215 2244.045 3388.940 2244.215 ;
        RECT 3388.215 2243.985 3389.110 2244.045 ;
        RECT 3385.030 2243.475 3386.050 2243.805 ;
        RECT 3386.220 2243.755 3386.390 2243.985 ;
        RECT 3388.940 2243.755 3389.110 2243.985 ;
        RECT 3385.030 2242.965 3385.200 2243.475 ;
        RECT 3386.220 2243.425 3386.390 2243.585 ;
        RECT 3388.940 2243.425 3389.110 2243.585 ;
        RECT 3386.220 2243.305 3387.540 2243.425 ;
        RECT 3385.420 2243.295 3387.540 2243.305 ;
        RECT 3385.420 2243.135 3386.220 2243.295 ;
        RECT 3386.390 2243.125 3387.540 2243.295 ;
        RECT 3386.220 2243.095 3387.540 2243.125 ;
        RECT 3388.140 2243.295 3389.110 2243.425 ;
        RECT 3388.140 2243.125 3388.940 2243.295 ;
        RECT 3388.140 2243.095 3389.110 2243.125 ;
        RECT 3385.030 2242.635 3386.050 2242.965 ;
        RECT 3386.220 2242.835 3386.390 2243.095 ;
      LAYER li1 ;
        RECT 3386.560 2242.755 3388.770 2242.925 ;
      LAYER li1 ;
        RECT 3388.940 2242.835 3389.110 2243.095 ;
      LAYER li1 ;
        RECT 3387.410 2242.670 3388.290 2242.755 ;
      LAYER li1 ;
        RECT 3385.030 2242.480 3385.200 2242.635 ;
        RECT 3384.320 2242.305 3385.200 2242.480 ;
        RECT 3386.220 2242.585 3386.390 2242.665 ;
        RECT 3386.220 2242.465 3387.190 2242.585 ;
        RECT 3385.420 2242.375 3387.190 2242.465 ;
        RECT 3383.500 2241.915 3383.670 2242.205 ;
        RECT 3383.500 2241.705 3383.670 2241.745 ;
        RECT 3383.500 2241.455 3384.150 2241.705 ;
        RECT 3383.670 2241.375 3384.150 2241.455 ;
        RECT 3383.500 2240.995 3383.670 2241.285 ;
        RECT 3383.670 2240.825 3384.150 2240.865 ;
        RECT 3383.500 2240.535 3384.150 2240.825 ;
        RECT 3383.500 2240.075 3383.670 2240.365 ;
        RECT 3383.670 2239.905 3384.150 2240.025 ;
        RECT 3383.500 2239.695 3384.150 2239.905 ;
        RECT 3384.660 2239.855 3384.830 2242.305 ;
        RECT 3385.420 2242.295 3386.220 2242.375 ;
        RECT 3386.390 2242.255 3387.190 2242.375 ;
        RECT 3386.220 2241.915 3386.390 2242.205 ;
      LAYER li1 ;
        RECT 3387.410 2242.085 3387.580 2242.670 ;
        RECT 3386.560 2241.915 3387.580 2242.085 ;
      LAYER li1 ;
        RECT 3386.220 2241.705 3387.190 2241.745 ;
        RECT 3385.420 2241.455 3387.190 2241.705 ;
        RECT 3385.420 2241.375 3386.220 2241.455 ;
        RECT 3386.390 2241.415 3387.190 2241.455 ;
        RECT 3386.220 2240.995 3386.390 2241.285 ;
      LAYER li1 ;
        RECT 3387.410 2241.245 3387.580 2241.915 ;
        RECT 3386.560 2241.075 3387.580 2241.245 ;
      LAYER li1 ;
        RECT 3385.420 2240.825 3386.220 2240.865 ;
        RECT 3386.390 2240.825 3387.190 2240.905 ;
        RECT 3385.420 2240.575 3387.190 2240.825 ;
        RECT 3385.420 2240.535 3386.390 2240.575 ;
      LAYER li1 ;
        RECT 3387.410 2240.405 3387.580 2241.075 ;
      LAYER li1 ;
        RECT 3386.220 2240.075 3386.390 2240.365 ;
      LAYER li1 ;
        RECT 3386.560 2240.235 3387.580 2240.405 ;
      LAYER li1 ;
        RECT 3385.420 2239.905 3386.220 2240.025 ;
        RECT 3386.390 2239.905 3387.190 2239.985 ;
        RECT 3387.780 2239.975 3387.950 2242.425 ;
      LAYER li1 ;
        RECT 3388.120 2242.085 3388.290 2242.670 ;
      LAYER li1 ;
        RECT 3388.940 2242.585 3389.110 2242.665 ;
        RECT 3388.460 2242.375 3389.110 2242.585 ;
        RECT 3388.460 2242.255 3388.940 2242.375 ;
      LAYER li1 ;
        RECT 3388.120 2241.915 3388.770 2242.085 ;
      LAYER li1 ;
        RECT 3388.940 2241.915 3389.110 2242.205 ;
      LAYER li1 ;
        RECT 3388.120 2241.245 3388.290 2241.915 ;
      LAYER li1 ;
        RECT 3388.460 2241.455 3389.110 2241.745 ;
        RECT 3388.460 2241.415 3388.940 2241.455 ;
      LAYER li1 ;
        RECT 3388.120 2241.075 3388.770 2241.245 ;
        RECT 3388.120 2240.405 3388.290 2241.075 ;
      LAYER li1 ;
        RECT 3388.940 2240.995 3389.110 2241.285 ;
        RECT 3388.460 2240.825 3388.940 2240.905 ;
        RECT 3388.460 2240.575 3389.110 2240.825 ;
        RECT 3388.940 2240.535 3389.110 2240.575 ;
      LAYER li1 ;
        RECT 3388.120 2240.235 3388.770 2240.405 ;
      LAYER li1 ;
        RECT 3388.940 2240.075 3389.110 2240.365 ;
        RECT 3385.420 2239.815 3387.190 2239.905 ;
        RECT 3385.420 2239.695 3386.390 2239.815 ;
        RECT 3383.500 2239.615 3383.670 2239.695 ;
        RECT 3386.220 2239.615 3386.390 2239.695 ;
        RECT 3387.410 2239.800 3388.290 2239.975 ;
        RECT 3387.410 2239.645 3387.580 2239.800 ;
        RECT 3383.500 2239.185 3383.670 2239.445 ;
        RECT 3386.220 2239.185 3386.390 2239.445 ;
        RECT 3386.560 2239.315 3387.580 2239.645 ;
        RECT 3383.500 2239.155 3384.470 2239.185 ;
        RECT 3383.670 2238.985 3384.470 2239.155 ;
        RECT 3383.500 2238.855 3384.470 2238.985 ;
        RECT 3385.070 2239.155 3386.390 2239.185 ;
        RECT 3385.070 2238.985 3386.220 2239.155 ;
        RECT 3386.390 2238.985 3387.190 2239.145 ;
        RECT 3385.070 2238.975 3387.190 2238.985 ;
        RECT 3385.070 2238.855 3386.390 2238.975 ;
        RECT 3383.500 2238.695 3383.670 2238.855 ;
        RECT 3386.220 2238.695 3386.390 2238.855 ;
        RECT 3387.410 2238.805 3387.580 2239.315 ;
        RECT 3383.500 2238.295 3383.670 2238.525 ;
        RECT 3386.220 2238.295 3386.390 2238.525 ;
        RECT 3386.560 2238.475 3387.580 2238.805 ;
        RECT 3388.120 2239.565 3388.290 2239.800 ;
        RECT 3388.460 2239.905 3388.940 2240.065 ;
        RECT 3388.460 2239.735 3389.110 2239.905 ;
        RECT 3388.940 2239.615 3389.110 2239.735 ;
        RECT 3388.120 2239.395 3388.765 2239.565 ;
        RECT 3388.120 2238.725 3388.290 2239.395 ;
        RECT 3388.940 2239.225 3389.110 2239.445 ;
        RECT 3388.460 2239.155 3389.110 2239.225 ;
        RECT 3388.460 2238.985 3388.940 2239.155 ;
        RECT 3388.460 2238.895 3389.110 2238.985 ;
        RECT 3388.120 2238.555 3388.770 2238.725 ;
        RECT 3388.940 2238.695 3389.110 2238.895 ;
        RECT 3388.940 2238.295 3389.110 2238.525 ;
        RECT 3383.500 2238.235 3384.395 2238.295 ;
        RECT 3383.670 2238.065 3384.395 2238.235 ;
        RECT 3383.500 2238.005 3384.395 2238.065 ;
        RECT 3383.500 2237.775 3383.670 2238.005 ;
        RECT 3383.500 2237.405 3383.670 2237.605 ;
        RECT 3383.840 2237.575 3384.490 2237.745 ;
        RECT 3383.500 2237.315 3384.150 2237.405 ;
        RECT 3383.670 2237.145 3384.150 2237.315 ;
        RECT 3383.500 2237.075 3384.150 2237.145 ;
        RECT 3383.500 2236.855 3383.670 2237.075 ;
        RECT 3384.320 2236.905 3384.490 2237.575 ;
        RECT 3383.845 2236.735 3384.490 2236.905 ;
        RECT 3383.500 2236.565 3383.670 2236.685 ;
        RECT 3383.500 2236.395 3384.150 2236.565 ;
        RECT 3383.670 2236.235 3384.150 2236.395 ;
        RECT 3384.320 2236.500 3384.490 2236.735 ;
      LAYER li1 ;
        RECT 3384.660 2236.680 3384.860 2238.270 ;
      LAYER li1 ;
        RECT 3385.055 2238.235 3387.555 2238.295 ;
        RECT 3385.055 2238.065 3386.220 2238.235 ;
        RECT 3386.390 2238.065 3387.555 2238.235 ;
        RECT 3385.055 2238.005 3387.555 2238.065 ;
        RECT 3388.215 2238.235 3389.110 2238.295 ;
        RECT 3388.215 2238.065 3388.940 2238.235 ;
        RECT 3388.215 2238.005 3389.110 2238.065 ;
        RECT 3385.030 2237.495 3386.050 2237.825 ;
        RECT 3386.220 2237.775 3386.390 2238.005 ;
        RECT 3388.940 2237.775 3389.110 2238.005 ;
        RECT 3385.030 2236.985 3385.200 2237.495 ;
        RECT 3386.220 2237.445 3386.390 2237.605 ;
        RECT 3388.940 2237.445 3389.110 2237.605 ;
        RECT 3386.220 2237.325 3387.540 2237.445 ;
        RECT 3385.420 2237.315 3387.540 2237.325 ;
        RECT 3385.420 2237.155 3386.220 2237.315 ;
        RECT 3386.390 2237.145 3387.540 2237.315 ;
        RECT 3386.220 2237.115 3387.540 2237.145 ;
        RECT 3388.140 2237.315 3389.110 2237.445 ;
        RECT 3388.140 2237.145 3388.940 2237.315 ;
        RECT 3388.140 2237.115 3389.110 2237.145 ;
        RECT 3385.030 2236.655 3386.050 2236.985 ;
        RECT 3386.220 2236.855 3386.390 2237.115 ;
      LAYER li1 ;
        RECT 3386.560 2236.775 3388.770 2236.945 ;
      LAYER li1 ;
        RECT 3388.940 2236.855 3389.110 2237.115 ;
      LAYER li1 ;
        RECT 3387.410 2236.690 3388.290 2236.775 ;
      LAYER li1 ;
        RECT 3385.030 2236.500 3385.200 2236.655 ;
        RECT 3384.320 2236.325 3385.200 2236.500 ;
        RECT 3386.220 2236.605 3386.390 2236.685 ;
        RECT 3386.220 2236.485 3387.190 2236.605 ;
        RECT 3385.420 2236.395 3387.190 2236.485 ;
        RECT 3383.500 2235.935 3383.670 2236.225 ;
        RECT 3383.500 2235.725 3383.670 2235.765 ;
        RECT 3383.500 2235.475 3384.150 2235.725 ;
        RECT 3383.670 2235.395 3384.150 2235.475 ;
        RECT 3383.500 2235.015 3383.670 2235.305 ;
        RECT 3383.670 2234.845 3384.150 2234.885 ;
        RECT 3383.500 2234.555 3384.150 2234.845 ;
        RECT 3383.500 2234.095 3383.670 2234.385 ;
        RECT 3383.670 2233.925 3384.150 2234.045 ;
        RECT 3383.500 2233.715 3384.150 2233.925 ;
        RECT 3384.660 2233.875 3384.830 2236.325 ;
        RECT 3385.420 2236.315 3386.220 2236.395 ;
        RECT 3386.390 2236.275 3387.190 2236.395 ;
        RECT 3386.220 2235.935 3386.390 2236.225 ;
      LAYER li1 ;
        RECT 3387.410 2236.105 3387.580 2236.690 ;
        RECT 3386.560 2235.935 3387.580 2236.105 ;
      LAYER li1 ;
        RECT 3386.220 2235.725 3387.190 2235.765 ;
        RECT 3385.420 2235.475 3387.190 2235.725 ;
        RECT 3385.420 2235.395 3386.220 2235.475 ;
        RECT 3386.390 2235.435 3387.190 2235.475 ;
        RECT 3386.220 2235.015 3386.390 2235.305 ;
      LAYER li1 ;
        RECT 3387.410 2235.265 3387.580 2235.935 ;
        RECT 3386.560 2235.095 3387.580 2235.265 ;
      LAYER li1 ;
        RECT 3385.420 2234.845 3386.220 2234.885 ;
        RECT 3386.390 2234.845 3387.190 2234.925 ;
        RECT 3385.420 2234.595 3387.190 2234.845 ;
        RECT 3385.420 2234.555 3386.390 2234.595 ;
      LAYER li1 ;
        RECT 3387.410 2234.425 3387.580 2235.095 ;
      LAYER li1 ;
        RECT 3386.220 2234.095 3386.390 2234.385 ;
      LAYER li1 ;
        RECT 3386.560 2234.255 3387.580 2234.425 ;
      LAYER li1 ;
        RECT 3385.420 2233.925 3386.220 2234.045 ;
        RECT 3386.390 2233.925 3387.190 2234.005 ;
        RECT 3387.780 2233.995 3387.950 2236.445 ;
      LAYER li1 ;
        RECT 3388.120 2236.105 3388.290 2236.690 ;
      LAYER li1 ;
        RECT 3388.940 2236.605 3389.110 2236.685 ;
        RECT 3388.460 2236.395 3389.110 2236.605 ;
        RECT 3388.460 2236.275 3388.940 2236.395 ;
      LAYER li1 ;
        RECT 3388.120 2235.935 3388.770 2236.105 ;
      LAYER li1 ;
        RECT 3388.940 2235.935 3389.110 2236.225 ;
      LAYER li1 ;
        RECT 3388.120 2235.265 3388.290 2235.935 ;
      LAYER li1 ;
        RECT 3388.460 2235.475 3389.110 2235.765 ;
        RECT 3388.460 2235.435 3388.940 2235.475 ;
      LAYER li1 ;
        RECT 3388.120 2235.095 3388.770 2235.265 ;
        RECT 3388.120 2234.425 3388.290 2235.095 ;
      LAYER li1 ;
        RECT 3388.940 2235.015 3389.110 2235.305 ;
        RECT 3388.460 2234.845 3388.940 2234.925 ;
        RECT 3388.460 2234.595 3389.110 2234.845 ;
        RECT 3388.940 2234.555 3389.110 2234.595 ;
      LAYER li1 ;
        RECT 3388.120 2234.255 3388.770 2234.425 ;
      LAYER li1 ;
        RECT 3388.940 2234.095 3389.110 2234.385 ;
        RECT 3385.420 2233.835 3387.190 2233.925 ;
        RECT 3385.420 2233.715 3386.390 2233.835 ;
        RECT 3383.500 2233.635 3383.670 2233.715 ;
        RECT 3386.220 2233.635 3386.390 2233.715 ;
        RECT 3387.410 2233.820 3388.290 2233.995 ;
        RECT 3387.410 2233.665 3387.580 2233.820 ;
        RECT 3383.500 2233.205 3383.670 2233.465 ;
        RECT 3386.220 2233.205 3386.390 2233.465 ;
        RECT 3386.560 2233.335 3387.580 2233.665 ;
        RECT 3383.500 2233.175 3384.470 2233.205 ;
        RECT 3383.670 2233.005 3384.470 2233.175 ;
        RECT 3383.500 2232.875 3384.470 2233.005 ;
        RECT 3385.070 2233.175 3386.390 2233.205 ;
        RECT 3385.070 2233.005 3386.220 2233.175 ;
        RECT 3386.390 2233.005 3387.190 2233.165 ;
        RECT 3385.070 2232.995 3387.190 2233.005 ;
        RECT 3385.070 2232.875 3386.390 2232.995 ;
        RECT 3383.500 2232.715 3383.670 2232.875 ;
        RECT 3386.220 2232.715 3386.390 2232.875 ;
        RECT 3387.410 2232.825 3387.580 2233.335 ;
        RECT 3383.500 2232.315 3383.670 2232.545 ;
        RECT 3386.220 2232.315 3386.390 2232.545 ;
        RECT 3386.560 2232.495 3387.580 2232.825 ;
        RECT 3388.120 2233.585 3388.290 2233.820 ;
        RECT 3388.460 2233.925 3388.940 2234.085 ;
        RECT 3388.460 2233.755 3389.110 2233.925 ;
        RECT 3388.940 2233.635 3389.110 2233.755 ;
        RECT 3388.120 2233.415 3388.765 2233.585 ;
        RECT 3388.120 2232.745 3388.290 2233.415 ;
        RECT 3388.940 2233.245 3389.110 2233.465 ;
        RECT 3388.460 2233.175 3389.110 2233.245 ;
        RECT 3388.460 2233.005 3388.940 2233.175 ;
        RECT 3388.460 2232.915 3389.110 2233.005 ;
        RECT 3388.120 2232.575 3388.770 2232.745 ;
        RECT 3388.940 2232.715 3389.110 2232.915 ;
        RECT 3388.940 2232.315 3389.110 2232.545 ;
        RECT 3383.500 2232.255 3384.395 2232.315 ;
        RECT 3383.670 2232.085 3384.395 2232.255 ;
        RECT 3383.500 2232.025 3384.395 2232.085 ;
        RECT 3385.055 2232.255 3387.555 2232.315 ;
        RECT 3385.055 2232.085 3386.220 2232.255 ;
        RECT 3386.390 2232.085 3387.555 2232.255 ;
        RECT 3385.055 2232.025 3387.555 2232.085 ;
        RECT 3388.215 2232.255 3389.110 2232.315 ;
        RECT 3388.215 2232.085 3388.940 2232.255 ;
        RECT 3388.215 2232.025 3389.110 2232.085 ;
        RECT 3383.500 2231.795 3383.670 2232.025 ;
        RECT 3383.500 2231.425 3383.670 2231.625 ;
        RECT 3383.840 2231.595 3384.490 2231.765 ;
        RECT 3383.500 2231.335 3384.150 2231.425 ;
        RECT 3383.670 2231.165 3384.150 2231.335 ;
        RECT 3383.500 2231.095 3384.150 2231.165 ;
        RECT 3383.500 2230.875 3383.670 2231.095 ;
        RECT 3384.320 2230.925 3384.490 2231.595 ;
        RECT 3383.845 2230.755 3384.490 2230.925 ;
        RECT 3383.500 2230.585 3383.670 2230.705 ;
        RECT 3383.500 2230.415 3384.150 2230.585 ;
        RECT 3383.670 2230.255 3384.150 2230.415 ;
        RECT 3384.320 2230.520 3384.490 2230.755 ;
        RECT 3385.030 2231.515 3386.050 2231.845 ;
        RECT 3386.220 2231.795 3386.390 2232.025 ;
        RECT 3388.940 2231.795 3389.110 2232.025 ;
        RECT 3385.030 2231.005 3385.200 2231.515 ;
        RECT 3386.220 2231.465 3386.390 2231.625 ;
        RECT 3388.940 2231.465 3389.110 2231.625 ;
        RECT 3386.220 2231.345 3387.540 2231.465 ;
        RECT 3385.420 2231.335 3387.540 2231.345 ;
        RECT 3385.420 2231.175 3386.220 2231.335 ;
        RECT 3386.390 2231.165 3387.540 2231.335 ;
        RECT 3386.220 2231.135 3387.540 2231.165 ;
        RECT 3388.140 2231.335 3389.110 2231.465 ;
        RECT 3388.140 2231.165 3388.940 2231.335 ;
        RECT 3388.140 2231.135 3389.110 2231.165 ;
        RECT 3385.030 2230.675 3386.050 2231.005 ;
        RECT 3386.220 2230.875 3386.390 2231.135 ;
        RECT 3388.940 2230.875 3389.110 2231.135 ;
        RECT 3385.030 2230.520 3385.200 2230.675 ;
        RECT 3384.320 2230.345 3385.200 2230.520 ;
        RECT 3386.220 2230.625 3386.390 2230.705 ;
        RECT 3388.940 2230.625 3389.110 2230.705 ;
        RECT 3386.220 2230.505 3387.190 2230.625 ;
        RECT 3385.420 2230.415 3387.190 2230.505 ;
        RECT 3383.500 2229.955 3383.670 2230.245 ;
        RECT 3383.500 2229.745 3383.670 2229.785 ;
        RECT 3383.500 2229.495 3384.150 2229.745 ;
        RECT 3383.670 2229.415 3384.150 2229.495 ;
        RECT 3383.500 2229.035 3383.670 2229.325 ;
        RECT 3383.670 2228.865 3384.150 2228.905 ;
        RECT 3383.500 2228.575 3384.150 2228.865 ;
        RECT 3383.500 2228.115 3383.670 2228.405 ;
        RECT 3383.670 2227.945 3384.150 2228.065 ;
        RECT 3383.500 2227.735 3384.150 2227.945 ;
        RECT 3384.660 2227.895 3384.830 2230.345 ;
        RECT 3385.420 2230.335 3386.220 2230.415 ;
        RECT 3386.390 2230.295 3387.190 2230.415 ;
        RECT 3386.220 2229.955 3386.390 2230.245 ;
        RECT 3386.220 2229.745 3387.190 2229.785 ;
        RECT 3385.420 2229.495 3387.190 2229.745 ;
        RECT 3385.420 2229.415 3386.220 2229.495 ;
        RECT 3386.390 2229.455 3387.190 2229.495 ;
        RECT 3386.220 2229.035 3386.390 2229.325 ;
        RECT 3385.420 2228.865 3386.220 2228.905 ;
        RECT 3386.390 2228.865 3387.190 2228.945 ;
        RECT 3385.420 2228.615 3387.190 2228.865 ;
        RECT 3385.420 2228.575 3386.390 2228.615 ;
        RECT 3386.220 2228.115 3386.390 2228.405 ;
        RECT 3385.420 2227.945 3386.220 2228.065 ;
        RECT 3386.390 2227.945 3387.190 2228.025 ;
        RECT 3387.780 2228.015 3387.950 2230.465 ;
        RECT 3388.460 2230.415 3389.110 2230.625 ;
        RECT 3388.460 2230.295 3388.940 2230.415 ;
        RECT 3388.940 2229.955 3389.110 2230.245 ;
        RECT 3388.460 2229.495 3389.110 2229.785 ;
        RECT 3388.460 2229.455 3388.940 2229.495 ;
        RECT 3388.940 2229.035 3389.110 2229.325 ;
        RECT 3388.460 2228.865 3388.940 2228.945 ;
        RECT 3388.460 2228.615 3389.110 2228.865 ;
        RECT 3388.940 2228.575 3389.110 2228.615 ;
        RECT 3388.940 2228.115 3389.110 2228.405 ;
        RECT 3385.420 2227.855 3387.190 2227.945 ;
        RECT 3385.420 2227.735 3386.390 2227.855 ;
        RECT 3383.500 2227.655 3383.670 2227.735 ;
        RECT 3386.220 2227.655 3386.390 2227.735 ;
        RECT 3387.410 2227.840 3388.290 2228.015 ;
        RECT 3387.410 2227.685 3387.580 2227.840 ;
        RECT 3383.500 2227.225 3383.670 2227.485 ;
        RECT 3386.220 2227.225 3386.390 2227.485 ;
        RECT 3386.560 2227.355 3387.580 2227.685 ;
        RECT 3383.500 2227.195 3384.470 2227.225 ;
        RECT 3383.670 2227.025 3384.470 2227.195 ;
        RECT 3383.500 2226.895 3384.470 2227.025 ;
        RECT 3385.070 2227.195 3386.390 2227.225 ;
        RECT 3385.070 2227.025 3386.220 2227.195 ;
        RECT 3386.390 2227.025 3387.190 2227.185 ;
        RECT 3385.070 2227.015 3387.190 2227.025 ;
        RECT 3385.070 2226.895 3386.390 2227.015 ;
        RECT 3383.500 2226.735 3383.670 2226.895 ;
        RECT 3386.220 2226.735 3386.390 2226.895 ;
        RECT 3387.410 2226.845 3387.580 2227.355 ;
        RECT 3383.500 2226.335 3383.670 2226.565 ;
        RECT 3386.220 2226.335 3386.390 2226.565 ;
        RECT 3386.560 2226.515 3387.580 2226.845 ;
        RECT 3388.120 2227.605 3388.290 2227.840 ;
        RECT 3388.460 2227.945 3388.940 2228.105 ;
        RECT 3388.460 2227.775 3389.110 2227.945 ;
        RECT 3388.940 2227.655 3389.110 2227.775 ;
        RECT 3388.120 2227.435 3388.765 2227.605 ;
        RECT 3388.120 2226.765 3388.290 2227.435 ;
        RECT 3388.940 2227.265 3389.110 2227.485 ;
        RECT 3388.460 2227.195 3389.110 2227.265 ;
        RECT 3388.460 2227.025 3388.940 2227.195 ;
        RECT 3388.460 2226.935 3389.110 2227.025 ;
        RECT 3388.120 2226.595 3388.770 2226.765 ;
        RECT 3388.940 2226.735 3389.110 2226.935 ;
        RECT 3388.940 2226.335 3389.110 2226.565 ;
        RECT 3383.500 2226.275 3384.395 2226.335 ;
        RECT 3383.670 2226.105 3384.395 2226.275 ;
        RECT 3383.500 2226.045 3384.395 2226.105 ;
        RECT 3385.055 2226.275 3387.555 2226.335 ;
        RECT 3385.055 2226.105 3386.220 2226.275 ;
        RECT 3386.390 2226.105 3387.555 2226.275 ;
        RECT 3385.055 2226.045 3387.555 2226.105 ;
        RECT 3388.215 2226.275 3389.110 2226.335 ;
        RECT 3388.215 2226.105 3388.940 2226.275 ;
        RECT 3388.215 2226.045 3389.110 2226.105 ;
        RECT 3383.500 2225.815 3383.670 2226.045 ;
        RECT 3383.500 2225.445 3383.670 2225.645 ;
        RECT 3383.840 2225.615 3384.490 2225.785 ;
        RECT 3383.500 2225.355 3384.150 2225.445 ;
        RECT 3383.670 2225.185 3384.150 2225.355 ;
        RECT 3383.500 2225.115 3384.150 2225.185 ;
        RECT 3383.500 2224.895 3383.670 2225.115 ;
        RECT 3384.320 2224.945 3384.490 2225.615 ;
        RECT 3383.845 2224.775 3384.490 2224.945 ;
        RECT 3383.500 2224.605 3383.670 2224.725 ;
        RECT 3383.500 2224.435 3384.150 2224.605 ;
        RECT 3383.670 2224.275 3384.150 2224.435 ;
        RECT 3384.320 2224.540 3384.490 2224.775 ;
        RECT 3385.030 2225.535 3386.050 2225.865 ;
        RECT 3386.220 2225.815 3386.390 2226.045 ;
        RECT 3388.940 2225.815 3389.110 2226.045 ;
        RECT 3385.030 2225.025 3385.200 2225.535 ;
        RECT 3386.220 2225.485 3386.390 2225.645 ;
        RECT 3388.940 2225.485 3389.110 2225.645 ;
        RECT 3386.220 2225.365 3387.540 2225.485 ;
        RECT 3385.420 2225.355 3387.540 2225.365 ;
        RECT 3385.420 2225.195 3386.220 2225.355 ;
        RECT 3386.390 2225.185 3387.540 2225.355 ;
        RECT 3386.220 2225.155 3387.540 2225.185 ;
        RECT 3388.140 2225.355 3389.110 2225.485 ;
        RECT 3388.140 2225.185 3388.940 2225.355 ;
        RECT 3388.140 2225.155 3389.110 2225.185 ;
        RECT 3385.030 2224.695 3386.050 2225.025 ;
        RECT 3386.220 2224.895 3386.390 2225.155 ;
        RECT 3388.940 2224.895 3389.110 2225.155 ;
        RECT 3385.030 2224.540 3385.200 2224.695 ;
        RECT 3384.320 2224.365 3385.200 2224.540 ;
        RECT 3386.220 2224.645 3386.390 2224.725 ;
        RECT 3388.940 2224.645 3389.110 2224.725 ;
        RECT 3386.220 2224.525 3387.190 2224.645 ;
        RECT 3385.420 2224.435 3387.190 2224.525 ;
        RECT 3383.500 2223.975 3383.670 2224.265 ;
        RECT 3383.500 2223.765 3383.670 2223.805 ;
        RECT 3383.500 2223.515 3384.150 2223.765 ;
        RECT 3383.670 2223.435 3384.150 2223.515 ;
        RECT 3383.500 2223.055 3383.670 2223.345 ;
        RECT 3383.670 2222.885 3384.150 2222.925 ;
        RECT 3383.500 2222.595 3384.150 2222.885 ;
        RECT 3383.500 2222.135 3383.670 2222.425 ;
        RECT 3383.670 2221.965 3384.150 2222.085 ;
        RECT 3383.500 2221.755 3384.150 2221.965 ;
        RECT 3384.660 2221.915 3384.830 2224.365 ;
        RECT 3385.420 2224.355 3386.220 2224.435 ;
        RECT 3386.390 2224.315 3387.190 2224.435 ;
        RECT 3386.220 2223.975 3386.390 2224.265 ;
        RECT 3386.220 2223.765 3387.190 2223.805 ;
        RECT 3385.420 2223.515 3387.190 2223.765 ;
        RECT 3385.420 2223.435 3386.220 2223.515 ;
        RECT 3386.390 2223.475 3387.190 2223.515 ;
        RECT 3386.220 2223.055 3386.390 2223.345 ;
        RECT 3385.420 2222.885 3386.220 2222.925 ;
        RECT 3386.390 2222.885 3387.190 2222.965 ;
        RECT 3385.420 2222.635 3387.190 2222.885 ;
        RECT 3385.420 2222.595 3386.390 2222.635 ;
        RECT 3386.220 2222.135 3386.390 2222.425 ;
        RECT 3385.420 2221.965 3386.220 2222.085 ;
        RECT 3386.390 2221.965 3387.190 2222.045 ;
        RECT 3387.780 2222.035 3387.950 2224.485 ;
        RECT 3388.460 2224.435 3389.110 2224.645 ;
        RECT 3388.460 2224.315 3388.940 2224.435 ;
        RECT 3388.940 2223.975 3389.110 2224.265 ;
        RECT 3388.460 2223.515 3389.110 2223.805 ;
        RECT 3388.460 2223.475 3388.940 2223.515 ;
        RECT 3388.940 2223.055 3389.110 2223.345 ;
        RECT 3388.460 2222.885 3388.940 2222.965 ;
        RECT 3388.460 2222.635 3389.110 2222.885 ;
        RECT 3388.940 2222.595 3389.110 2222.635 ;
        RECT 3388.940 2222.135 3389.110 2222.425 ;
        RECT 3385.420 2221.875 3387.190 2221.965 ;
        RECT 3385.420 2221.755 3386.390 2221.875 ;
        RECT 3383.500 2221.675 3383.670 2221.755 ;
        RECT 3386.220 2221.675 3386.390 2221.755 ;
        RECT 3387.410 2221.860 3388.290 2222.035 ;
        RECT 3387.410 2221.705 3387.580 2221.860 ;
        RECT 3383.500 2221.245 3383.670 2221.505 ;
        RECT 3386.220 2221.245 3386.390 2221.505 ;
        RECT 3386.560 2221.375 3387.580 2221.705 ;
        RECT 3383.500 2221.215 3384.470 2221.245 ;
        RECT 3383.670 2221.045 3384.470 2221.215 ;
        RECT 3383.500 2220.915 3384.470 2221.045 ;
        RECT 3385.070 2221.215 3386.390 2221.245 ;
        RECT 3385.070 2221.045 3386.220 2221.215 ;
        RECT 3386.390 2221.045 3387.190 2221.205 ;
        RECT 3385.070 2221.035 3387.190 2221.045 ;
        RECT 3385.070 2220.915 3386.390 2221.035 ;
        RECT 3383.500 2220.755 3383.670 2220.915 ;
        RECT 3386.220 2220.755 3386.390 2220.915 ;
        RECT 3387.410 2220.865 3387.580 2221.375 ;
        RECT 3383.500 2220.355 3383.670 2220.585 ;
        RECT 3386.220 2220.355 3386.390 2220.585 ;
        RECT 3386.560 2220.535 3387.580 2220.865 ;
        RECT 3388.120 2221.625 3388.290 2221.860 ;
        RECT 3388.460 2221.965 3388.940 2222.125 ;
        RECT 3388.460 2221.795 3389.110 2221.965 ;
        RECT 3388.940 2221.675 3389.110 2221.795 ;
        RECT 3388.120 2221.455 3388.765 2221.625 ;
        RECT 3388.120 2220.785 3388.290 2221.455 ;
        RECT 3388.940 2221.285 3389.110 2221.505 ;
        RECT 3388.460 2221.215 3389.110 2221.285 ;
        RECT 3388.460 2221.045 3388.940 2221.215 ;
        RECT 3388.460 2220.955 3389.110 2221.045 ;
        RECT 3388.120 2220.615 3388.770 2220.785 ;
        RECT 3388.940 2220.755 3389.110 2220.955 ;
        RECT 3388.940 2220.355 3389.110 2220.585 ;
        RECT 3383.500 2220.295 3384.395 2220.355 ;
        RECT 3383.670 2220.125 3384.395 2220.295 ;
        RECT 3383.500 2220.065 3384.395 2220.125 ;
        RECT 3385.055 2220.295 3387.555 2220.355 ;
        RECT 3385.055 2220.125 3386.220 2220.295 ;
        RECT 3386.390 2220.125 3387.555 2220.295 ;
        RECT 3385.055 2220.065 3387.555 2220.125 ;
        RECT 3388.215 2220.295 3389.110 2220.355 ;
        RECT 3388.215 2220.125 3388.940 2220.295 ;
        RECT 3388.215 2220.065 3389.110 2220.125 ;
        RECT 3383.500 2219.835 3383.670 2220.065 ;
        RECT 3383.500 2219.465 3383.670 2219.665 ;
        RECT 3383.840 2219.635 3384.490 2219.805 ;
        RECT 3383.500 2219.375 3384.150 2219.465 ;
        RECT 3383.670 2219.205 3384.150 2219.375 ;
        RECT 3383.500 2219.135 3384.150 2219.205 ;
        RECT 3383.500 2218.915 3383.670 2219.135 ;
        RECT 3384.320 2218.965 3384.490 2219.635 ;
        RECT 3383.845 2218.795 3384.490 2218.965 ;
        RECT 3383.500 2218.625 3383.670 2218.745 ;
        RECT 3383.500 2218.455 3384.150 2218.625 ;
        RECT 3383.670 2218.295 3384.150 2218.455 ;
        RECT 3384.320 2218.560 3384.490 2218.795 ;
        RECT 3385.030 2219.555 3386.050 2219.885 ;
        RECT 3386.220 2219.835 3386.390 2220.065 ;
        RECT 3388.940 2219.835 3389.110 2220.065 ;
        RECT 3385.030 2219.045 3385.200 2219.555 ;
        RECT 3386.220 2219.505 3386.390 2219.665 ;
        RECT 3388.940 2219.505 3389.110 2219.665 ;
        RECT 3386.220 2219.385 3387.540 2219.505 ;
        RECT 3385.420 2219.375 3387.540 2219.385 ;
        RECT 3385.420 2219.215 3386.220 2219.375 ;
        RECT 3386.390 2219.205 3387.540 2219.375 ;
        RECT 3386.220 2219.175 3387.540 2219.205 ;
        RECT 3388.140 2219.375 3389.110 2219.505 ;
        RECT 3388.140 2219.205 3388.940 2219.375 ;
        RECT 3388.140 2219.175 3389.110 2219.205 ;
        RECT 3385.030 2218.715 3386.050 2219.045 ;
        RECT 3386.220 2218.915 3386.390 2219.175 ;
        RECT 3388.940 2218.915 3389.110 2219.175 ;
        RECT 3385.030 2218.560 3385.200 2218.715 ;
        RECT 3384.320 2218.385 3385.200 2218.560 ;
        RECT 3386.220 2218.665 3386.390 2218.745 ;
        RECT 3388.940 2218.665 3389.110 2218.745 ;
        RECT 3386.220 2218.545 3387.190 2218.665 ;
        RECT 3385.420 2218.455 3387.190 2218.545 ;
        RECT 3383.500 2217.995 3383.670 2218.285 ;
        RECT 3383.500 2217.785 3383.670 2217.825 ;
        RECT 3383.500 2217.535 3384.150 2217.785 ;
        RECT 3383.670 2217.455 3384.150 2217.535 ;
        RECT 3383.500 2217.075 3383.670 2217.365 ;
        RECT 3383.670 2216.905 3384.150 2216.945 ;
        RECT 3383.500 2216.615 3384.150 2216.905 ;
        RECT 3383.500 2216.155 3383.670 2216.445 ;
        RECT 3383.670 2215.985 3384.150 2216.105 ;
        RECT 3383.500 2215.775 3384.150 2215.985 ;
        RECT 3384.660 2215.935 3384.830 2218.385 ;
        RECT 3385.420 2218.375 3386.220 2218.455 ;
        RECT 3386.390 2218.335 3387.190 2218.455 ;
        RECT 3386.220 2217.995 3386.390 2218.285 ;
        RECT 3386.220 2217.785 3387.190 2217.825 ;
        RECT 3385.420 2217.535 3387.190 2217.785 ;
        RECT 3385.420 2217.455 3386.220 2217.535 ;
        RECT 3386.390 2217.495 3387.190 2217.535 ;
        RECT 3386.220 2217.075 3386.390 2217.365 ;
        RECT 3385.420 2216.905 3386.220 2216.945 ;
        RECT 3386.390 2216.905 3387.190 2216.985 ;
        RECT 3385.420 2216.655 3387.190 2216.905 ;
        RECT 3385.420 2216.615 3386.390 2216.655 ;
        RECT 3386.220 2216.155 3386.390 2216.445 ;
        RECT 3385.420 2215.985 3386.220 2216.105 ;
        RECT 3386.390 2215.985 3387.190 2216.065 ;
        RECT 3387.780 2216.055 3387.950 2218.505 ;
        RECT 3388.460 2218.455 3389.110 2218.665 ;
        RECT 3388.460 2218.335 3388.940 2218.455 ;
        RECT 3388.940 2217.995 3389.110 2218.285 ;
        RECT 3388.460 2217.535 3389.110 2217.825 ;
        RECT 3388.460 2217.495 3388.940 2217.535 ;
        RECT 3388.940 2217.075 3389.110 2217.365 ;
        RECT 3388.460 2216.905 3388.940 2216.985 ;
        RECT 3388.460 2216.655 3389.110 2216.905 ;
        RECT 3388.940 2216.615 3389.110 2216.655 ;
        RECT 3388.940 2216.155 3389.110 2216.445 ;
        RECT 3385.420 2215.895 3387.190 2215.985 ;
        RECT 3385.420 2215.775 3386.390 2215.895 ;
        RECT 3383.500 2215.695 3383.670 2215.775 ;
        RECT 3386.220 2215.695 3386.390 2215.775 ;
        RECT 3387.410 2215.880 3388.290 2216.055 ;
        RECT 3387.410 2215.725 3387.580 2215.880 ;
        RECT 3383.500 2215.265 3383.670 2215.525 ;
        RECT 3386.220 2215.265 3386.390 2215.525 ;
        RECT 3386.560 2215.395 3387.580 2215.725 ;
        RECT 3383.500 2215.235 3384.470 2215.265 ;
        RECT 3383.670 2215.065 3384.470 2215.235 ;
        RECT 3383.500 2214.935 3384.470 2215.065 ;
        RECT 3385.070 2215.235 3386.390 2215.265 ;
        RECT 3385.070 2215.065 3386.220 2215.235 ;
        RECT 3386.390 2215.065 3387.190 2215.225 ;
        RECT 3385.070 2215.055 3387.190 2215.065 ;
        RECT 3385.070 2214.935 3386.390 2215.055 ;
        RECT 3383.500 2214.775 3383.670 2214.935 ;
        RECT 3386.220 2214.775 3386.390 2214.935 ;
        RECT 3387.410 2214.885 3387.580 2215.395 ;
        RECT 3383.500 2214.375 3383.670 2214.605 ;
        RECT 3386.220 2214.375 3386.390 2214.605 ;
        RECT 3386.560 2214.555 3387.580 2214.885 ;
        RECT 3388.120 2215.645 3388.290 2215.880 ;
        RECT 3388.460 2215.985 3388.940 2216.145 ;
        RECT 3388.460 2215.815 3389.110 2215.985 ;
        RECT 3388.940 2215.695 3389.110 2215.815 ;
        RECT 3388.120 2215.475 3388.765 2215.645 ;
        RECT 3388.120 2214.805 3388.290 2215.475 ;
        RECT 3388.940 2215.305 3389.110 2215.525 ;
        RECT 3388.460 2215.235 3389.110 2215.305 ;
        RECT 3388.460 2215.065 3388.940 2215.235 ;
        RECT 3388.460 2214.975 3389.110 2215.065 ;
        RECT 3388.120 2214.635 3388.770 2214.805 ;
        RECT 3388.940 2214.775 3389.110 2214.975 ;
        RECT 3388.940 2214.375 3389.110 2214.605 ;
        RECT 3383.500 2214.315 3384.395 2214.375 ;
        RECT 3383.670 2214.145 3384.395 2214.315 ;
        RECT 3383.500 2214.085 3384.395 2214.145 ;
        RECT 3385.055 2214.315 3387.555 2214.375 ;
        RECT 3385.055 2214.145 3386.220 2214.315 ;
        RECT 3386.390 2214.145 3387.555 2214.315 ;
        RECT 3385.055 2214.085 3387.555 2214.145 ;
        RECT 3388.215 2214.315 3389.110 2214.375 ;
        RECT 3388.215 2214.145 3388.940 2214.315 ;
        RECT 3388.215 2214.085 3389.110 2214.145 ;
        RECT 3383.500 2213.855 3383.670 2214.085 ;
        RECT 3383.500 2213.485 3383.670 2213.685 ;
        RECT 3383.840 2213.655 3384.490 2213.825 ;
        RECT 3383.500 2213.395 3384.150 2213.485 ;
        RECT 3383.670 2213.225 3384.150 2213.395 ;
        RECT 3383.500 2213.155 3384.150 2213.225 ;
        RECT 3383.500 2212.935 3383.670 2213.155 ;
        RECT 3384.320 2212.985 3384.490 2213.655 ;
        RECT 3383.845 2212.815 3384.490 2212.985 ;
        RECT 3383.500 2212.645 3383.670 2212.765 ;
        RECT 3383.500 2212.475 3384.150 2212.645 ;
        RECT 3383.670 2212.315 3384.150 2212.475 ;
        RECT 3384.320 2212.580 3384.490 2212.815 ;
        RECT 3385.030 2213.575 3386.050 2213.905 ;
        RECT 3386.220 2213.855 3386.390 2214.085 ;
        RECT 3388.940 2213.855 3389.110 2214.085 ;
        RECT 3385.030 2213.065 3385.200 2213.575 ;
        RECT 3386.220 2213.525 3386.390 2213.685 ;
        RECT 3388.940 2213.525 3389.110 2213.685 ;
        RECT 3386.220 2213.405 3387.540 2213.525 ;
        RECT 3385.420 2213.395 3387.540 2213.405 ;
        RECT 3385.420 2213.235 3386.220 2213.395 ;
        RECT 3386.390 2213.225 3387.540 2213.395 ;
        RECT 3386.220 2213.195 3387.540 2213.225 ;
        RECT 3388.140 2213.395 3389.110 2213.525 ;
        RECT 3388.140 2213.225 3388.940 2213.395 ;
        RECT 3388.140 2213.195 3389.110 2213.225 ;
        RECT 3385.030 2212.735 3386.050 2213.065 ;
        RECT 3386.220 2212.935 3386.390 2213.195 ;
        RECT 3388.940 2212.935 3389.110 2213.195 ;
        RECT 3385.030 2212.580 3385.200 2212.735 ;
        RECT 3384.320 2212.405 3385.200 2212.580 ;
        RECT 3386.220 2212.685 3386.390 2212.765 ;
        RECT 3388.940 2212.685 3389.110 2212.765 ;
        RECT 3386.220 2212.565 3387.190 2212.685 ;
        RECT 3385.420 2212.475 3387.190 2212.565 ;
        RECT 3383.500 2212.015 3383.670 2212.305 ;
        RECT 3383.500 2211.805 3383.670 2211.845 ;
        RECT 3383.500 2211.555 3384.150 2211.805 ;
        RECT 3383.670 2211.475 3384.150 2211.555 ;
        RECT 3383.500 2211.095 3383.670 2211.385 ;
        RECT 3383.670 2210.925 3384.150 2210.965 ;
        RECT 3383.500 2210.635 3384.150 2210.925 ;
        RECT 3383.500 2210.175 3383.670 2210.465 ;
        RECT 3383.670 2210.005 3384.150 2210.125 ;
        RECT 3383.500 2209.795 3384.150 2210.005 ;
        RECT 3384.660 2209.955 3384.830 2212.405 ;
        RECT 3385.420 2212.395 3386.220 2212.475 ;
        RECT 3386.390 2212.355 3387.190 2212.475 ;
        RECT 3386.220 2212.015 3386.390 2212.305 ;
        RECT 3386.220 2211.805 3387.190 2211.845 ;
        RECT 3385.420 2211.555 3387.190 2211.805 ;
        RECT 3385.420 2211.475 3386.220 2211.555 ;
        RECT 3386.390 2211.515 3387.190 2211.555 ;
        RECT 3386.220 2211.095 3386.390 2211.385 ;
        RECT 3385.420 2210.925 3386.220 2210.965 ;
        RECT 3386.390 2210.925 3387.190 2211.005 ;
        RECT 3385.420 2210.675 3387.190 2210.925 ;
        RECT 3385.420 2210.635 3386.390 2210.675 ;
        RECT 3386.220 2210.175 3386.390 2210.465 ;
        RECT 3385.420 2210.005 3386.220 2210.125 ;
        RECT 3386.390 2210.005 3387.190 2210.085 ;
        RECT 3387.780 2210.075 3387.950 2212.525 ;
        RECT 3388.460 2212.475 3389.110 2212.685 ;
        RECT 3388.460 2212.355 3388.940 2212.475 ;
        RECT 3388.940 2212.015 3389.110 2212.305 ;
        RECT 3388.460 2211.555 3389.110 2211.845 ;
        RECT 3388.460 2211.515 3388.940 2211.555 ;
        RECT 3388.940 2211.095 3389.110 2211.385 ;
        RECT 3388.460 2210.925 3388.940 2211.005 ;
        RECT 3388.460 2210.675 3389.110 2210.925 ;
        RECT 3388.940 2210.635 3389.110 2210.675 ;
        RECT 3388.940 2210.175 3389.110 2210.465 ;
        RECT 3385.420 2209.915 3387.190 2210.005 ;
        RECT 3385.420 2209.795 3386.390 2209.915 ;
        RECT 3383.500 2209.715 3383.670 2209.795 ;
        RECT 3386.220 2209.715 3386.390 2209.795 ;
        RECT 3387.410 2209.900 3388.290 2210.075 ;
        RECT 3387.410 2209.745 3387.580 2209.900 ;
        RECT 3383.500 2209.285 3383.670 2209.545 ;
        RECT 3386.220 2209.285 3386.390 2209.545 ;
        RECT 3386.560 2209.415 3387.580 2209.745 ;
        RECT 3383.500 2209.255 3384.470 2209.285 ;
        RECT 3383.670 2209.085 3384.470 2209.255 ;
        RECT 3383.500 2208.955 3384.470 2209.085 ;
        RECT 3385.070 2209.255 3386.390 2209.285 ;
        RECT 3385.070 2209.085 3386.220 2209.255 ;
        RECT 3386.390 2209.085 3387.190 2209.245 ;
        RECT 3385.070 2209.075 3387.190 2209.085 ;
        RECT 3385.070 2208.955 3386.390 2209.075 ;
        RECT 3383.500 2208.795 3383.670 2208.955 ;
        RECT 3386.220 2208.795 3386.390 2208.955 ;
        RECT 3387.410 2208.905 3387.580 2209.415 ;
        RECT 3383.500 2208.395 3383.670 2208.625 ;
        RECT 3386.220 2208.395 3386.390 2208.625 ;
        RECT 3386.560 2208.575 3387.580 2208.905 ;
        RECT 3388.120 2209.665 3388.290 2209.900 ;
        RECT 3388.460 2210.005 3388.940 2210.165 ;
        RECT 3388.460 2209.835 3389.110 2210.005 ;
        RECT 3388.940 2209.715 3389.110 2209.835 ;
        RECT 3388.120 2209.495 3388.765 2209.665 ;
        RECT 3388.120 2208.825 3388.290 2209.495 ;
        RECT 3388.940 2209.325 3389.110 2209.545 ;
        RECT 3388.460 2209.255 3389.110 2209.325 ;
        RECT 3388.460 2209.085 3388.940 2209.255 ;
        RECT 3388.460 2208.995 3389.110 2209.085 ;
        RECT 3388.120 2208.655 3388.770 2208.825 ;
        RECT 3388.940 2208.795 3389.110 2208.995 ;
        RECT 3388.940 2208.395 3389.110 2208.625 ;
        RECT 3383.500 2208.335 3384.395 2208.395 ;
        RECT 3383.670 2208.165 3384.395 2208.335 ;
        RECT 3383.500 2208.105 3384.395 2208.165 ;
        RECT 3385.055 2208.335 3387.555 2208.395 ;
        RECT 3385.055 2208.165 3386.220 2208.335 ;
        RECT 3386.390 2208.165 3387.555 2208.335 ;
        RECT 3385.055 2208.105 3387.555 2208.165 ;
        RECT 3388.215 2208.335 3389.110 2208.395 ;
        RECT 3388.215 2208.165 3388.940 2208.335 ;
        RECT 3388.215 2208.105 3389.110 2208.165 ;
        RECT 3383.500 2207.875 3383.670 2208.105 ;
        RECT 3383.500 2207.505 3383.670 2207.705 ;
        RECT 3383.840 2207.675 3384.490 2207.845 ;
        RECT 3383.500 2207.415 3384.150 2207.505 ;
        RECT 3383.670 2207.245 3384.150 2207.415 ;
        RECT 3383.500 2207.175 3384.150 2207.245 ;
        RECT 3383.500 2206.955 3383.670 2207.175 ;
        RECT 3384.320 2207.005 3384.490 2207.675 ;
        RECT 3383.845 2206.835 3384.490 2207.005 ;
        RECT 3383.500 2206.665 3383.670 2206.785 ;
        RECT 3383.500 2206.495 3384.150 2206.665 ;
        RECT 3383.670 2206.335 3384.150 2206.495 ;
        RECT 3384.320 2206.600 3384.490 2206.835 ;
        RECT 3385.030 2207.595 3386.050 2207.925 ;
        RECT 3386.220 2207.875 3386.390 2208.105 ;
        RECT 3388.940 2207.875 3389.110 2208.105 ;
        RECT 3385.030 2207.085 3385.200 2207.595 ;
        RECT 3386.220 2207.545 3386.390 2207.705 ;
        RECT 3388.940 2207.545 3389.110 2207.705 ;
        RECT 3386.220 2207.425 3387.540 2207.545 ;
        RECT 3385.420 2207.415 3387.540 2207.425 ;
        RECT 3385.420 2207.255 3386.220 2207.415 ;
        RECT 3386.390 2207.245 3387.540 2207.415 ;
        RECT 3386.220 2207.215 3387.540 2207.245 ;
        RECT 3388.140 2207.415 3389.110 2207.545 ;
        RECT 3388.140 2207.245 3388.940 2207.415 ;
        RECT 3388.140 2207.215 3389.110 2207.245 ;
        RECT 3385.030 2206.755 3386.050 2207.085 ;
        RECT 3386.220 2206.955 3386.390 2207.215 ;
        RECT 3388.940 2206.955 3389.110 2207.215 ;
        RECT 3385.030 2206.600 3385.200 2206.755 ;
        RECT 3384.320 2206.425 3385.200 2206.600 ;
        RECT 3386.220 2206.705 3386.390 2206.785 ;
        RECT 3388.940 2206.705 3389.110 2206.785 ;
        RECT 3386.220 2206.585 3387.190 2206.705 ;
        RECT 3385.420 2206.495 3387.190 2206.585 ;
        RECT 3383.500 2206.035 3383.670 2206.325 ;
        RECT 3383.500 2205.825 3383.670 2205.865 ;
        RECT 3383.500 2205.575 3384.150 2205.825 ;
        RECT 3383.670 2205.495 3384.150 2205.575 ;
        RECT 3383.500 2205.115 3383.670 2205.405 ;
        RECT 3383.670 2204.945 3384.150 2204.985 ;
        RECT 3383.500 2204.655 3384.150 2204.945 ;
        RECT 3383.500 2204.195 3383.670 2204.485 ;
        RECT 3383.670 2204.025 3384.150 2204.145 ;
        RECT 3383.500 2203.815 3384.150 2204.025 ;
        RECT 3384.660 2203.975 3384.830 2206.425 ;
        RECT 3385.420 2206.415 3386.220 2206.495 ;
        RECT 3386.390 2206.375 3387.190 2206.495 ;
        RECT 3386.220 2206.035 3386.390 2206.325 ;
        RECT 3386.220 2205.825 3387.190 2205.865 ;
        RECT 3385.420 2205.575 3387.190 2205.825 ;
        RECT 3385.420 2205.495 3386.220 2205.575 ;
        RECT 3386.390 2205.535 3387.190 2205.575 ;
        RECT 3386.220 2205.115 3386.390 2205.405 ;
        RECT 3385.420 2204.945 3386.220 2204.985 ;
        RECT 3386.390 2204.945 3387.190 2205.025 ;
        RECT 3385.420 2204.695 3387.190 2204.945 ;
        RECT 3385.420 2204.655 3386.390 2204.695 ;
        RECT 3386.220 2204.195 3386.390 2204.485 ;
        RECT 3385.420 2204.025 3386.220 2204.145 ;
        RECT 3386.390 2204.025 3387.190 2204.105 ;
        RECT 3387.780 2204.095 3387.950 2206.545 ;
        RECT 3388.460 2206.495 3389.110 2206.705 ;
        RECT 3388.460 2206.375 3388.940 2206.495 ;
        RECT 3388.940 2206.035 3389.110 2206.325 ;
        RECT 3388.460 2205.575 3389.110 2205.865 ;
        RECT 3388.460 2205.535 3388.940 2205.575 ;
        RECT 3388.940 2205.115 3389.110 2205.405 ;
        RECT 3388.460 2204.945 3388.940 2205.025 ;
        RECT 3388.460 2204.695 3389.110 2204.945 ;
        RECT 3388.940 2204.655 3389.110 2204.695 ;
        RECT 3388.940 2204.195 3389.110 2204.485 ;
        RECT 3385.420 2203.935 3387.190 2204.025 ;
        RECT 3385.420 2203.815 3386.390 2203.935 ;
        RECT 3383.500 2203.735 3383.670 2203.815 ;
        RECT 3386.220 2203.735 3386.390 2203.815 ;
        RECT 3387.410 2203.920 3388.290 2204.095 ;
        RECT 3387.410 2203.765 3387.580 2203.920 ;
        RECT 3383.500 2203.305 3383.670 2203.565 ;
        RECT 3386.220 2203.305 3386.390 2203.565 ;
        RECT 3386.560 2203.435 3387.580 2203.765 ;
        RECT 3383.500 2203.275 3384.470 2203.305 ;
        RECT 3383.670 2203.105 3384.470 2203.275 ;
        RECT 3383.500 2202.975 3384.470 2203.105 ;
        RECT 3385.070 2203.275 3386.390 2203.305 ;
        RECT 3385.070 2203.105 3386.220 2203.275 ;
        RECT 3386.390 2203.105 3387.190 2203.265 ;
        RECT 3385.070 2203.095 3387.190 2203.105 ;
        RECT 3385.070 2202.975 3386.390 2203.095 ;
        RECT 3383.500 2202.815 3383.670 2202.975 ;
        RECT 3386.220 2202.815 3386.390 2202.975 ;
        RECT 3387.410 2202.925 3387.580 2203.435 ;
        RECT 3383.500 2202.415 3383.670 2202.645 ;
        RECT 3386.220 2202.415 3386.390 2202.645 ;
        RECT 3386.560 2202.595 3387.580 2202.925 ;
        RECT 3388.120 2203.685 3388.290 2203.920 ;
        RECT 3388.460 2204.025 3388.940 2204.185 ;
        RECT 3388.460 2203.855 3389.110 2204.025 ;
        RECT 3388.940 2203.735 3389.110 2203.855 ;
        RECT 3388.120 2203.515 3388.765 2203.685 ;
        RECT 3388.120 2202.845 3388.290 2203.515 ;
        RECT 3388.940 2203.345 3389.110 2203.565 ;
        RECT 3388.460 2203.275 3389.110 2203.345 ;
        RECT 3388.460 2203.105 3388.940 2203.275 ;
        RECT 3388.460 2203.015 3389.110 2203.105 ;
        RECT 3388.120 2202.675 3388.770 2202.845 ;
        RECT 3388.940 2202.815 3389.110 2203.015 ;
        RECT 3388.940 2202.415 3389.110 2202.645 ;
        RECT 3383.500 2202.355 3384.395 2202.415 ;
        RECT 3383.670 2202.185 3384.395 2202.355 ;
        RECT 3383.500 2202.125 3384.395 2202.185 ;
        RECT 3385.055 2202.355 3387.555 2202.415 ;
        RECT 3385.055 2202.185 3386.220 2202.355 ;
        RECT 3386.390 2202.185 3387.555 2202.355 ;
        RECT 3385.055 2202.125 3387.555 2202.185 ;
        RECT 3388.215 2202.355 3389.110 2202.415 ;
        RECT 3388.215 2202.185 3388.940 2202.355 ;
        RECT 3388.215 2202.125 3389.110 2202.185 ;
        RECT 3383.500 2201.895 3383.670 2202.125 ;
        RECT 3383.500 2201.525 3383.670 2201.725 ;
        RECT 3383.840 2201.695 3384.490 2201.865 ;
        RECT 3383.500 2201.435 3384.150 2201.525 ;
        RECT 3383.670 2201.265 3384.150 2201.435 ;
        RECT 3383.500 2201.195 3384.150 2201.265 ;
        RECT 3383.500 2200.975 3383.670 2201.195 ;
        RECT 3384.320 2201.025 3384.490 2201.695 ;
        RECT 3383.845 2200.855 3384.490 2201.025 ;
        RECT 3383.500 2200.685 3383.670 2200.805 ;
        RECT 3383.500 2200.515 3384.150 2200.685 ;
        RECT 3383.670 2200.355 3384.150 2200.515 ;
        RECT 3384.320 2200.620 3384.490 2200.855 ;
        RECT 3385.030 2201.615 3386.050 2201.945 ;
        RECT 3386.220 2201.895 3386.390 2202.125 ;
        RECT 3388.940 2201.895 3389.110 2202.125 ;
        RECT 3385.030 2201.105 3385.200 2201.615 ;
        RECT 3386.220 2201.565 3386.390 2201.725 ;
        RECT 3388.940 2201.565 3389.110 2201.725 ;
        RECT 3386.220 2201.445 3387.540 2201.565 ;
        RECT 3385.420 2201.435 3387.540 2201.445 ;
        RECT 3385.420 2201.275 3386.220 2201.435 ;
        RECT 3386.390 2201.265 3387.540 2201.435 ;
        RECT 3386.220 2201.235 3387.540 2201.265 ;
        RECT 3388.140 2201.435 3389.110 2201.565 ;
        RECT 3388.140 2201.265 3388.940 2201.435 ;
        RECT 3388.140 2201.235 3389.110 2201.265 ;
        RECT 3385.030 2200.775 3386.050 2201.105 ;
        RECT 3386.220 2200.975 3386.390 2201.235 ;
        RECT 3388.940 2200.975 3389.110 2201.235 ;
        RECT 3385.030 2200.620 3385.200 2200.775 ;
        RECT 3384.320 2200.445 3385.200 2200.620 ;
        RECT 3386.220 2200.725 3386.390 2200.805 ;
        RECT 3388.940 2200.725 3389.110 2200.805 ;
        RECT 3386.220 2200.605 3387.190 2200.725 ;
        RECT 3385.420 2200.515 3387.190 2200.605 ;
        RECT 3383.500 2200.055 3383.670 2200.345 ;
        RECT 3383.500 2199.845 3383.670 2199.885 ;
        RECT 3383.500 2199.595 3384.150 2199.845 ;
        RECT 3383.670 2199.515 3384.150 2199.595 ;
        RECT 3383.500 2199.135 3383.670 2199.425 ;
        RECT 3383.670 2198.965 3384.150 2199.005 ;
        RECT 3383.500 2198.675 3384.150 2198.965 ;
        RECT 3383.500 2198.215 3383.670 2198.505 ;
        RECT 3383.670 2198.045 3384.150 2198.165 ;
        RECT 3383.500 2197.835 3384.150 2198.045 ;
        RECT 3384.660 2197.995 3384.830 2200.445 ;
        RECT 3385.420 2200.435 3386.220 2200.515 ;
        RECT 3386.390 2200.395 3387.190 2200.515 ;
        RECT 3386.220 2200.055 3386.390 2200.345 ;
        RECT 3386.220 2199.845 3387.190 2199.885 ;
        RECT 3385.420 2199.595 3387.190 2199.845 ;
        RECT 3385.420 2199.515 3386.220 2199.595 ;
        RECT 3386.390 2199.555 3387.190 2199.595 ;
        RECT 3386.220 2199.135 3386.390 2199.425 ;
        RECT 3385.420 2198.965 3386.220 2199.005 ;
        RECT 3386.390 2198.965 3387.190 2199.045 ;
        RECT 3385.420 2198.715 3387.190 2198.965 ;
        RECT 3385.420 2198.675 3386.390 2198.715 ;
        RECT 3386.220 2198.215 3386.390 2198.505 ;
        RECT 3385.420 2198.045 3386.220 2198.165 ;
        RECT 3386.390 2198.045 3387.190 2198.125 ;
        RECT 3387.780 2198.115 3387.950 2200.565 ;
        RECT 3388.460 2200.515 3389.110 2200.725 ;
        RECT 3388.460 2200.395 3388.940 2200.515 ;
        RECT 3388.940 2200.055 3389.110 2200.345 ;
        RECT 3388.460 2199.595 3389.110 2199.885 ;
        RECT 3388.460 2199.555 3388.940 2199.595 ;
        RECT 3388.940 2199.135 3389.110 2199.425 ;
        RECT 3388.460 2198.965 3388.940 2199.045 ;
        RECT 3388.460 2198.715 3389.110 2198.965 ;
        RECT 3388.940 2198.675 3389.110 2198.715 ;
        RECT 3388.940 2198.215 3389.110 2198.505 ;
        RECT 3385.420 2197.955 3387.190 2198.045 ;
        RECT 3385.420 2197.835 3386.390 2197.955 ;
        RECT 3383.500 2197.755 3383.670 2197.835 ;
        RECT 3386.220 2197.755 3386.390 2197.835 ;
        RECT 3387.410 2197.940 3388.290 2198.115 ;
        RECT 3387.410 2197.785 3387.580 2197.940 ;
        RECT 3383.500 2197.325 3383.670 2197.585 ;
        RECT 3386.220 2197.325 3386.390 2197.585 ;
        RECT 3386.560 2197.455 3387.580 2197.785 ;
        RECT 3383.500 2197.295 3384.470 2197.325 ;
        RECT 3383.670 2197.125 3384.470 2197.295 ;
        RECT 3383.500 2196.995 3384.470 2197.125 ;
        RECT 3385.070 2197.295 3386.390 2197.325 ;
        RECT 3385.070 2197.125 3386.220 2197.295 ;
        RECT 3386.390 2197.125 3387.190 2197.285 ;
        RECT 3385.070 2197.115 3387.190 2197.125 ;
        RECT 3385.070 2196.995 3386.390 2197.115 ;
        RECT 3383.500 2196.835 3383.670 2196.995 ;
        RECT 3386.220 2196.835 3386.390 2196.995 ;
        RECT 3387.410 2196.945 3387.580 2197.455 ;
        RECT 3383.500 2196.435 3383.670 2196.665 ;
        RECT 3386.220 2196.435 3386.390 2196.665 ;
        RECT 3386.560 2196.615 3387.580 2196.945 ;
        RECT 3388.120 2197.705 3388.290 2197.940 ;
        RECT 3388.460 2198.045 3388.940 2198.205 ;
        RECT 3388.460 2197.875 3389.110 2198.045 ;
        RECT 3388.940 2197.755 3389.110 2197.875 ;
        RECT 3388.120 2197.535 3388.765 2197.705 ;
        RECT 3388.120 2196.865 3388.290 2197.535 ;
        RECT 3388.940 2197.365 3389.110 2197.585 ;
        RECT 3388.460 2197.295 3389.110 2197.365 ;
        RECT 3388.460 2197.125 3388.940 2197.295 ;
        RECT 3388.460 2197.035 3389.110 2197.125 ;
        RECT 3388.120 2196.695 3388.770 2196.865 ;
        RECT 3388.940 2196.835 3389.110 2197.035 ;
        RECT 3388.940 2196.435 3389.110 2196.665 ;
        RECT 3383.500 2196.375 3384.395 2196.435 ;
        RECT 3383.670 2196.205 3384.395 2196.375 ;
        RECT 3383.500 2196.145 3384.395 2196.205 ;
        RECT 3385.055 2196.375 3387.555 2196.435 ;
        RECT 3385.055 2196.205 3386.220 2196.375 ;
        RECT 3386.390 2196.205 3387.555 2196.375 ;
        RECT 3385.055 2196.145 3387.555 2196.205 ;
        RECT 3388.215 2196.375 3389.110 2196.435 ;
        RECT 3388.215 2196.205 3388.940 2196.375 ;
        RECT 3388.215 2196.145 3389.110 2196.205 ;
        RECT 3383.500 2196.060 3383.670 2196.145 ;
        RECT 3386.220 2196.060 3386.390 2196.145 ;
        RECT 3388.940 2196.060 3389.110 2196.145 ;
        RECT 198.795 1762.980 198.965 1763.065 ;
        RECT 201.515 1762.980 201.685 1763.065 ;
        RECT 204.235 1762.980 204.405 1763.065 ;
        RECT 198.795 1762.920 199.690 1762.980 ;
        RECT 198.965 1762.750 199.690 1762.920 ;
        RECT 198.795 1762.690 199.690 1762.750 ;
        RECT 200.350 1762.920 202.850 1762.980 ;
        RECT 200.350 1762.750 201.515 1762.920 ;
        RECT 201.685 1762.750 202.850 1762.920 ;
        RECT 200.350 1762.690 202.850 1762.750 ;
        RECT 198.795 1762.460 198.965 1762.690 ;
        RECT 201.515 1762.460 201.685 1762.690 ;
        RECT 198.795 1762.130 198.965 1762.290 ;
        RECT 201.515 1762.130 201.685 1762.290 ;
        RECT 201.855 1762.180 202.875 1762.510 ;
        RECT 198.795 1762.000 199.765 1762.130 ;
        RECT 198.965 1761.830 199.765 1762.000 ;
        RECT 198.795 1761.800 199.765 1761.830 ;
        RECT 200.365 1762.010 201.685 1762.130 ;
        RECT 200.365 1762.000 202.485 1762.010 ;
        RECT 200.365 1761.830 201.515 1762.000 ;
        RECT 201.685 1761.840 202.485 1762.000 ;
        RECT 200.365 1761.800 201.685 1761.830 ;
        RECT 198.795 1761.540 198.965 1761.800 ;
      LAYER li1 ;
        RECT 199.135 1761.460 201.345 1761.630 ;
      LAYER li1 ;
        RECT 201.515 1761.540 201.685 1761.800 ;
        RECT 202.705 1761.670 202.875 1762.180 ;
      LAYER li1 ;
        RECT 199.615 1761.375 200.495 1761.460 ;
      LAYER li1 ;
        RECT 198.795 1761.290 198.965 1761.370 ;
        RECT 198.795 1761.080 199.445 1761.290 ;
        RECT 198.965 1760.960 199.445 1761.080 ;
        RECT 198.795 1760.620 198.965 1760.910 ;
      LAYER li1 ;
        RECT 199.615 1760.790 199.785 1761.375 ;
        RECT 199.135 1760.620 199.785 1760.790 ;
      LAYER li1 ;
        RECT 198.795 1760.160 199.445 1760.450 ;
        RECT 198.965 1760.120 199.445 1760.160 ;
        RECT 198.795 1759.700 198.965 1759.990 ;
      LAYER li1 ;
        RECT 199.615 1759.950 199.785 1760.620 ;
        RECT 199.135 1759.780 199.785 1759.950 ;
      LAYER li1 ;
        RECT 198.965 1759.530 199.445 1759.610 ;
        RECT 198.795 1759.280 199.445 1759.530 ;
        RECT 198.795 1759.240 198.965 1759.280 ;
      LAYER li1 ;
        RECT 199.615 1759.110 199.785 1759.780 ;
      LAYER li1 ;
        RECT 198.795 1758.780 198.965 1759.070 ;
      LAYER li1 ;
        RECT 199.135 1758.940 199.785 1759.110 ;
      LAYER li1 ;
        RECT 198.965 1758.610 199.445 1758.770 ;
        RECT 199.955 1758.680 200.125 1761.130 ;
      LAYER li1 ;
        RECT 200.325 1760.790 200.495 1761.375 ;
      LAYER li1 ;
        RECT 201.515 1761.290 201.685 1761.370 ;
        RECT 201.855 1761.340 202.875 1761.670 ;
      LAYER li1 ;
        RECT 203.045 1761.365 203.245 1762.955 ;
      LAYER li1 ;
        RECT 203.510 1762.920 204.405 1762.980 ;
        RECT 203.510 1762.750 204.235 1762.920 ;
        RECT 203.510 1762.690 204.405 1762.750 ;
        RECT 204.235 1762.460 204.405 1762.690 ;
        RECT 203.415 1762.260 204.065 1762.430 ;
        RECT 203.415 1761.590 203.585 1762.260 ;
        RECT 204.235 1762.090 204.405 1762.290 ;
        RECT 203.755 1762.000 204.405 1762.090 ;
        RECT 203.755 1761.830 204.235 1762.000 ;
        RECT 203.755 1761.760 204.405 1761.830 ;
        RECT 203.415 1761.420 204.060 1761.590 ;
        RECT 204.235 1761.540 204.405 1761.760 ;
        RECT 200.715 1761.170 201.685 1761.290 ;
        RECT 202.705 1761.185 202.875 1761.340 ;
        RECT 203.415 1761.185 203.585 1761.420 ;
        RECT 204.235 1761.250 204.405 1761.370 ;
        RECT 200.715 1761.080 202.485 1761.170 ;
        RECT 200.715 1760.960 201.515 1761.080 ;
        RECT 201.685 1761.000 202.485 1761.080 ;
        RECT 202.705 1761.010 203.585 1761.185 ;
        RECT 203.755 1761.080 204.405 1761.250 ;
      LAYER li1 ;
        RECT 200.325 1760.620 201.345 1760.790 ;
      LAYER li1 ;
        RECT 201.515 1760.620 201.685 1760.910 ;
      LAYER li1 ;
        RECT 200.325 1759.950 200.495 1760.620 ;
        RECT 201.855 1760.580 202.875 1760.750 ;
      LAYER li1 ;
        RECT 200.715 1760.410 201.685 1760.450 ;
        RECT 200.715 1760.160 202.485 1760.410 ;
        RECT 200.715 1760.120 201.515 1760.160 ;
        RECT 201.685 1760.080 202.485 1760.160 ;
      LAYER li1 ;
        RECT 200.325 1759.780 201.345 1759.950 ;
        RECT 200.325 1759.110 200.495 1759.780 ;
      LAYER li1 ;
        RECT 201.515 1759.700 201.685 1759.990 ;
      LAYER li1 ;
        RECT 202.705 1759.910 202.875 1760.580 ;
        RECT 201.855 1759.740 202.875 1759.910 ;
      LAYER li1 ;
        RECT 200.715 1759.530 201.515 1759.610 ;
        RECT 201.685 1759.530 202.485 1759.570 ;
        RECT 200.715 1759.280 202.485 1759.530 ;
        RECT 201.515 1759.240 202.485 1759.280 ;
      LAYER li1 ;
        RECT 200.325 1758.940 201.345 1759.110 ;
        RECT 202.705 1759.070 202.875 1759.740 ;
      LAYER li1 ;
        RECT 201.515 1758.780 201.685 1759.070 ;
      LAYER li1 ;
        RECT 201.855 1758.900 202.875 1759.070 ;
      LAYER li1 ;
        RECT 198.795 1758.440 199.445 1758.610 ;
        RECT 199.615 1758.505 200.495 1758.680 ;
        RECT 200.715 1758.610 201.515 1758.690 ;
        RECT 201.685 1758.610 202.485 1758.730 ;
        RECT 200.715 1758.520 202.485 1758.610 ;
        RECT 198.795 1758.320 198.965 1758.440 ;
        RECT 199.615 1758.270 199.785 1758.505 ;
        RECT 200.325 1758.350 200.495 1758.505 ;
        RECT 201.515 1758.400 202.485 1758.520 ;
        RECT 198.795 1757.930 198.965 1758.150 ;
        RECT 199.140 1758.100 199.785 1758.270 ;
        RECT 198.795 1757.860 199.445 1757.930 ;
        RECT 198.965 1757.690 199.445 1757.860 ;
        RECT 198.795 1757.600 199.445 1757.690 ;
        RECT 198.795 1757.400 198.965 1757.600 ;
        RECT 199.615 1757.430 199.785 1758.100 ;
        RECT 199.135 1757.260 199.785 1757.430 ;
        RECT 198.795 1757.000 198.965 1757.230 ;
      LAYER li1 ;
        RECT 199.955 1757.225 200.155 1758.325 ;
      LAYER li1 ;
        RECT 200.325 1758.020 201.345 1758.350 ;
        RECT 201.515 1758.320 201.685 1758.400 ;
      LAYER li1 ;
        RECT 202.705 1758.315 202.875 1758.900 ;
      LAYER li1 ;
        RECT 203.075 1758.560 203.245 1761.010 ;
        RECT 203.755 1760.920 204.235 1761.080 ;
      LAYER li1 ;
        RECT 203.415 1760.580 204.065 1760.750 ;
      LAYER li1 ;
        RECT 204.235 1760.620 204.405 1760.910 ;
      LAYER li1 ;
        RECT 203.415 1759.910 203.585 1760.580 ;
      LAYER li1 ;
        RECT 204.235 1760.410 204.405 1760.450 ;
        RECT 203.755 1760.160 204.405 1760.410 ;
        RECT 203.755 1760.080 204.235 1760.160 ;
      LAYER li1 ;
        RECT 203.415 1759.740 204.065 1759.910 ;
        RECT 203.415 1759.070 203.585 1759.740 ;
      LAYER li1 ;
        RECT 204.235 1759.700 204.405 1759.990 ;
        RECT 203.755 1759.530 204.235 1759.570 ;
        RECT 203.755 1759.240 204.405 1759.530 ;
      LAYER li1 ;
        RECT 203.415 1758.900 204.065 1759.070 ;
        RECT 203.415 1758.315 203.585 1758.900 ;
      LAYER li1 ;
        RECT 204.235 1758.780 204.405 1759.070 ;
        RECT 203.755 1758.610 204.235 1758.730 ;
        RECT 203.755 1758.400 204.405 1758.610 ;
        RECT 204.235 1758.320 204.405 1758.400 ;
      LAYER li1 ;
        RECT 202.705 1758.230 203.585 1758.315 ;
      LAYER li1 ;
        RECT 200.325 1757.510 200.495 1758.020 ;
        RECT 201.515 1757.890 201.685 1758.150 ;
      LAYER li1 ;
        RECT 201.855 1758.060 204.065 1758.230 ;
      LAYER li1 ;
        RECT 204.235 1757.890 204.405 1758.150 ;
        RECT 201.515 1757.860 202.835 1757.890 ;
        RECT 200.715 1757.690 201.515 1757.850 ;
        RECT 201.685 1757.690 202.835 1757.860 ;
        RECT 200.715 1757.680 202.835 1757.690 ;
        RECT 201.515 1757.560 202.835 1757.680 ;
        RECT 203.435 1757.860 204.405 1757.890 ;
        RECT 203.435 1757.690 204.235 1757.860 ;
        RECT 203.435 1757.560 204.405 1757.690 ;
        RECT 200.325 1757.180 201.345 1757.510 ;
        RECT 201.515 1757.400 201.685 1757.560 ;
        RECT 204.235 1757.400 204.405 1757.560 ;
        RECT 201.515 1757.000 201.685 1757.230 ;
        RECT 204.235 1757.000 204.405 1757.230 ;
        RECT 198.795 1756.940 199.690 1757.000 ;
        RECT 198.965 1756.770 199.690 1756.940 ;
        RECT 198.795 1756.710 199.690 1756.770 ;
        RECT 200.350 1756.940 202.850 1757.000 ;
        RECT 200.350 1756.770 201.515 1756.940 ;
        RECT 201.685 1756.770 202.850 1756.940 ;
        RECT 200.350 1756.710 202.850 1756.770 ;
        RECT 198.795 1756.480 198.965 1756.710 ;
        RECT 201.515 1756.480 201.685 1756.710 ;
        RECT 198.795 1756.150 198.965 1756.310 ;
        RECT 201.515 1756.150 201.685 1756.310 ;
        RECT 201.855 1756.200 202.875 1756.530 ;
        RECT 198.795 1756.020 199.765 1756.150 ;
        RECT 198.965 1755.850 199.765 1756.020 ;
        RECT 198.795 1755.820 199.765 1755.850 ;
        RECT 200.365 1756.030 201.685 1756.150 ;
        RECT 200.365 1756.020 202.485 1756.030 ;
        RECT 200.365 1755.850 201.515 1756.020 ;
        RECT 201.685 1755.860 202.485 1756.020 ;
        RECT 200.365 1755.820 201.685 1755.850 ;
        RECT 198.795 1755.560 198.965 1755.820 ;
      LAYER li1 ;
        RECT 199.135 1755.480 201.345 1755.650 ;
      LAYER li1 ;
        RECT 201.515 1755.560 201.685 1755.820 ;
        RECT 202.705 1755.690 202.875 1756.200 ;
      LAYER li1 ;
        RECT 199.615 1755.395 200.495 1755.480 ;
      LAYER li1 ;
        RECT 198.795 1755.310 198.965 1755.390 ;
        RECT 198.795 1755.100 199.445 1755.310 ;
        RECT 198.965 1754.980 199.445 1755.100 ;
        RECT 198.795 1754.640 198.965 1754.930 ;
      LAYER li1 ;
        RECT 199.615 1754.810 199.785 1755.395 ;
        RECT 199.135 1754.640 199.785 1754.810 ;
      LAYER li1 ;
        RECT 198.795 1754.180 199.445 1754.470 ;
        RECT 198.965 1754.140 199.445 1754.180 ;
        RECT 198.795 1753.720 198.965 1754.010 ;
      LAYER li1 ;
        RECT 199.615 1753.970 199.785 1754.640 ;
        RECT 199.135 1753.800 199.785 1753.970 ;
      LAYER li1 ;
        RECT 198.965 1753.550 199.445 1753.630 ;
        RECT 198.795 1753.300 199.445 1753.550 ;
        RECT 198.795 1753.260 198.965 1753.300 ;
      LAYER li1 ;
        RECT 199.615 1753.130 199.785 1753.800 ;
      LAYER li1 ;
        RECT 198.795 1752.800 198.965 1753.090 ;
      LAYER li1 ;
        RECT 199.135 1752.960 199.785 1753.130 ;
      LAYER li1 ;
        RECT 198.965 1752.630 199.445 1752.790 ;
        RECT 199.955 1752.700 200.125 1755.150 ;
      LAYER li1 ;
        RECT 200.325 1754.810 200.495 1755.395 ;
      LAYER li1 ;
        RECT 201.515 1755.310 201.685 1755.390 ;
        RECT 201.855 1755.360 202.875 1755.690 ;
      LAYER li1 ;
        RECT 203.045 1755.385 203.245 1756.975 ;
      LAYER li1 ;
        RECT 203.510 1756.940 204.405 1757.000 ;
        RECT 203.510 1756.770 204.235 1756.940 ;
        RECT 203.510 1756.710 204.405 1756.770 ;
        RECT 204.235 1756.480 204.405 1756.710 ;
        RECT 203.415 1756.280 204.065 1756.450 ;
        RECT 203.415 1755.610 203.585 1756.280 ;
        RECT 204.235 1756.110 204.405 1756.310 ;
        RECT 203.755 1756.020 204.405 1756.110 ;
        RECT 203.755 1755.850 204.235 1756.020 ;
        RECT 203.755 1755.780 204.405 1755.850 ;
        RECT 203.415 1755.440 204.060 1755.610 ;
        RECT 204.235 1755.560 204.405 1755.780 ;
        RECT 200.715 1755.190 201.685 1755.310 ;
        RECT 202.705 1755.205 202.875 1755.360 ;
        RECT 203.415 1755.205 203.585 1755.440 ;
        RECT 204.235 1755.270 204.405 1755.390 ;
        RECT 200.715 1755.100 202.485 1755.190 ;
        RECT 200.715 1754.980 201.515 1755.100 ;
        RECT 201.685 1755.020 202.485 1755.100 ;
        RECT 202.705 1755.030 203.585 1755.205 ;
        RECT 203.755 1755.100 204.405 1755.270 ;
      LAYER li1 ;
        RECT 200.325 1754.640 201.345 1754.810 ;
      LAYER li1 ;
        RECT 201.515 1754.640 201.685 1754.930 ;
      LAYER li1 ;
        RECT 200.325 1753.970 200.495 1754.640 ;
        RECT 201.855 1754.600 202.875 1754.770 ;
      LAYER li1 ;
        RECT 200.715 1754.430 201.685 1754.470 ;
        RECT 200.715 1754.180 202.485 1754.430 ;
        RECT 200.715 1754.140 201.515 1754.180 ;
        RECT 201.685 1754.100 202.485 1754.180 ;
      LAYER li1 ;
        RECT 200.325 1753.800 201.345 1753.970 ;
        RECT 200.325 1753.130 200.495 1753.800 ;
      LAYER li1 ;
        RECT 201.515 1753.720 201.685 1754.010 ;
      LAYER li1 ;
        RECT 202.705 1753.930 202.875 1754.600 ;
        RECT 201.855 1753.760 202.875 1753.930 ;
      LAYER li1 ;
        RECT 200.715 1753.550 201.515 1753.630 ;
        RECT 201.685 1753.550 202.485 1753.590 ;
        RECT 200.715 1753.300 202.485 1753.550 ;
        RECT 201.515 1753.260 202.485 1753.300 ;
      LAYER li1 ;
        RECT 200.325 1752.960 201.345 1753.130 ;
        RECT 202.705 1753.090 202.875 1753.760 ;
      LAYER li1 ;
        RECT 201.515 1752.800 201.685 1753.090 ;
      LAYER li1 ;
        RECT 201.855 1752.920 202.875 1753.090 ;
      LAYER li1 ;
        RECT 198.795 1752.460 199.445 1752.630 ;
        RECT 199.615 1752.525 200.495 1752.700 ;
        RECT 200.715 1752.630 201.515 1752.710 ;
        RECT 201.685 1752.630 202.485 1752.750 ;
        RECT 200.715 1752.540 202.485 1752.630 ;
        RECT 198.795 1752.340 198.965 1752.460 ;
        RECT 199.615 1752.290 199.785 1752.525 ;
        RECT 200.325 1752.370 200.495 1752.525 ;
        RECT 201.515 1752.420 202.485 1752.540 ;
        RECT 198.795 1751.950 198.965 1752.170 ;
        RECT 199.140 1752.120 199.785 1752.290 ;
        RECT 198.795 1751.880 199.445 1751.950 ;
        RECT 198.965 1751.710 199.445 1751.880 ;
        RECT 198.795 1751.620 199.445 1751.710 ;
        RECT 198.795 1751.420 198.965 1751.620 ;
        RECT 199.615 1751.450 199.785 1752.120 ;
        RECT 199.135 1751.280 199.785 1751.450 ;
        RECT 198.795 1751.020 198.965 1751.250 ;
      LAYER li1 ;
        RECT 199.955 1751.245 200.155 1752.345 ;
      LAYER li1 ;
        RECT 200.325 1752.040 201.345 1752.370 ;
        RECT 201.515 1752.340 201.685 1752.420 ;
      LAYER li1 ;
        RECT 202.705 1752.335 202.875 1752.920 ;
      LAYER li1 ;
        RECT 203.075 1752.580 203.245 1755.030 ;
        RECT 203.755 1754.940 204.235 1755.100 ;
      LAYER li1 ;
        RECT 203.415 1754.600 204.065 1754.770 ;
      LAYER li1 ;
        RECT 204.235 1754.640 204.405 1754.930 ;
      LAYER li1 ;
        RECT 203.415 1753.930 203.585 1754.600 ;
      LAYER li1 ;
        RECT 204.235 1754.430 204.405 1754.470 ;
        RECT 203.755 1754.180 204.405 1754.430 ;
        RECT 203.755 1754.100 204.235 1754.180 ;
      LAYER li1 ;
        RECT 203.415 1753.760 204.065 1753.930 ;
        RECT 203.415 1753.090 203.585 1753.760 ;
      LAYER li1 ;
        RECT 204.235 1753.720 204.405 1754.010 ;
        RECT 203.755 1753.550 204.235 1753.590 ;
        RECT 203.755 1753.260 204.405 1753.550 ;
      LAYER li1 ;
        RECT 203.415 1752.920 204.065 1753.090 ;
        RECT 203.415 1752.335 203.585 1752.920 ;
      LAYER li1 ;
        RECT 204.235 1752.800 204.405 1753.090 ;
        RECT 203.755 1752.630 204.235 1752.750 ;
        RECT 203.755 1752.420 204.405 1752.630 ;
        RECT 204.235 1752.340 204.405 1752.420 ;
      LAYER li1 ;
        RECT 202.705 1752.250 203.585 1752.335 ;
      LAYER li1 ;
        RECT 200.325 1751.530 200.495 1752.040 ;
        RECT 201.515 1751.910 201.685 1752.170 ;
      LAYER li1 ;
        RECT 201.855 1752.080 204.065 1752.250 ;
      LAYER li1 ;
        RECT 204.235 1751.910 204.405 1752.170 ;
        RECT 201.515 1751.880 202.835 1751.910 ;
        RECT 200.715 1751.710 201.515 1751.870 ;
        RECT 201.685 1751.710 202.835 1751.880 ;
        RECT 200.715 1751.700 202.835 1751.710 ;
        RECT 201.515 1751.580 202.835 1751.700 ;
        RECT 203.435 1751.880 204.405 1751.910 ;
        RECT 203.435 1751.710 204.235 1751.880 ;
        RECT 203.435 1751.580 204.405 1751.710 ;
        RECT 200.325 1751.200 201.345 1751.530 ;
        RECT 201.515 1751.420 201.685 1751.580 ;
        RECT 204.235 1751.420 204.405 1751.580 ;
        RECT 201.515 1751.020 201.685 1751.250 ;
        RECT 204.235 1751.020 204.405 1751.250 ;
        RECT 198.795 1750.960 199.690 1751.020 ;
        RECT 198.965 1750.790 199.690 1750.960 ;
        RECT 198.795 1750.730 199.690 1750.790 ;
        RECT 200.350 1750.960 202.850 1751.020 ;
        RECT 200.350 1750.790 201.515 1750.960 ;
        RECT 201.685 1750.790 202.850 1750.960 ;
        RECT 200.350 1750.730 202.850 1750.790 ;
        RECT 198.795 1750.500 198.965 1750.730 ;
        RECT 201.515 1750.500 201.685 1750.730 ;
        RECT 198.795 1750.170 198.965 1750.330 ;
        RECT 201.515 1750.170 201.685 1750.330 ;
        RECT 201.855 1750.220 202.875 1750.550 ;
        RECT 198.795 1750.040 199.765 1750.170 ;
        RECT 198.965 1749.870 199.765 1750.040 ;
        RECT 198.795 1749.840 199.765 1749.870 ;
        RECT 200.365 1750.050 201.685 1750.170 ;
        RECT 200.365 1750.040 202.485 1750.050 ;
        RECT 200.365 1749.870 201.515 1750.040 ;
        RECT 201.685 1749.880 202.485 1750.040 ;
        RECT 200.365 1749.840 201.685 1749.870 ;
        RECT 198.795 1749.580 198.965 1749.840 ;
      LAYER li1 ;
        RECT 199.135 1749.500 201.345 1749.670 ;
      LAYER li1 ;
        RECT 201.515 1749.580 201.685 1749.840 ;
        RECT 202.705 1749.710 202.875 1750.220 ;
      LAYER li1 ;
        RECT 199.615 1749.415 200.495 1749.500 ;
      LAYER li1 ;
        RECT 198.795 1749.330 198.965 1749.410 ;
        RECT 198.795 1749.120 199.445 1749.330 ;
        RECT 198.965 1749.000 199.445 1749.120 ;
        RECT 198.795 1748.660 198.965 1748.950 ;
      LAYER li1 ;
        RECT 199.615 1748.830 199.785 1749.415 ;
        RECT 199.135 1748.660 199.785 1748.830 ;
      LAYER li1 ;
        RECT 198.795 1748.200 199.445 1748.490 ;
        RECT 198.965 1748.160 199.445 1748.200 ;
        RECT 198.795 1747.740 198.965 1748.030 ;
      LAYER li1 ;
        RECT 199.615 1747.990 199.785 1748.660 ;
        RECT 199.135 1747.820 199.785 1747.990 ;
      LAYER li1 ;
        RECT 198.965 1747.570 199.445 1747.650 ;
        RECT 198.795 1747.320 199.445 1747.570 ;
        RECT 198.795 1747.280 198.965 1747.320 ;
      LAYER li1 ;
        RECT 199.615 1747.150 199.785 1747.820 ;
      LAYER li1 ;
        RECT 198.795 1746.820 198.965 1747.110 ;
      LAYER li1 ;
        RECT 199.135 1746.980 199.785 1747.150 ;
      LAYER li1 ;
        RECT 198.965 1746.650 199.445 1746.810 ;
        RECT 199.955 1746.720 200.125 1749.170 ;
      LAYER li1 ;
        RECT 200.325 1748.830 200.495 1749.415 ;
      LAYER li1 ;
        RECT 201.515 1749.330 201.685 1749.410 ;
        RECT 201.855 1749.380 202.875 1749.710 ;
      LAYER li1 ;
        RECT 203.045 1749.405 203.245 1750.995 ;
      LAYER li1 ;
        RECT 203.510 1750.960 204.405 1751.020 ;
        RECT 203.510 1750.790 204.235 1750.960 ;
        RECT 203.510 1750.730 204.405 1750.790 ;
        RECT 204.235 1750.500 204.405 1750.730 ;
        RECT 203.415 1750.300 204.065 1750.470 ;
        RECT 203.415 1749.630 203.585 1750.300 ;
        RECT 204.235 1750.130 204.405 1750.330 ;
        RECT 203.755 1750.040 204.405 1750.130 ;
        RECT 203.755 1749.870 204.235 1750.040 ;
        RECT 203.755 1749.800 204.405 1749.870 ;
        RECT 203.415 1749.460 204.060 1749.630 ;
        RECT 204.235 1749.580 204.405 1749.800 ;
        RECT 200.715 1749.210 201.685 1749.330 ;
        RECT 202.705 1749.225 202.875 1749.380 ;
        RECT 203.415 1749.225 203.585 1749.460 ;
        RECT 204.235 1749.290 204.405 1749.410 ;
        RECT 200.715 1749.120 202.485 1749.210 ;
        RECT 200.715 1749.000 201.515 1749.120 ;
        RECT 201.685 1749.040 202.485 1749.120 ;
        RECT 202.705 1749.050 203.585 1749.225 ;
        RECT 203.755 1749.120 204.405 1749.290 ;
      LAYER li1 ;
        RECT 200.325 1748.660 201.345 1748.830 ;
      LAYER li1 ;
        RECT 201.515 1748.660 201.685 1748.950 ;
      LAYER li1 ;
        RECT 200.325 1747.990 200.495 1748.660 ;
        RECT 201.855 1748.620 202.875 1748.790 ;
      LAYER li1 ;
        RECT 200.715 1748.450 201.685 1748.490 ;
        RECT 200.715 1748.200 202.485 1748.450 ;
        RECT 200.715 1748.160 201.515 1748.200 ;
        RECT 201.685 1748.120 202.485 1748.200 ;
      LAYER li1 ;
        RECT 200.325 1747.820 201.345 1747.990 ;
        RECT 200.325 1747.150 200.495 1747.820 ;
      LAYER li1 ;
        RECT 201.515 1747.740 201.685 1748.030 ;
      LAYER li1 ;
        RECT 202.705 1747.950 202.875 1748.620 ;
        RECT 201.855 1747.780 202.875 1747.950 ;
      LAYER li1 ;
        RECT 200.715 1747.570 201.515 1747.650 ;
        RECT 201.685 1747.570 202.485 1747.610 ;
        RECT 200.715 1747.320 202.485 1747.570 ;
        RECT 201.515 1747.280 202.485 1747.320 ;
      LAYER li1 ;
        RECT 200.325 1746.980 201.345 1747.150 ;
        RECT 202.705 1747.110 202.875 1747.780 ;
      LAYER li1 ;
        RECT 201.515 1746.820 201.685 1747.110 ;
      LAYER li1 ;
        RECT 201.855 1746.940 202.875 1747.110 ;
      LAYER li1 ;
        RECT 198.795 1746.480 199.445 1746.650 ;
        RECT 199.615 1746.545 200.495 1746.720 ;
        RECT 200.715 1746.650 201.515 1746.730 ;
        RECT 201.685 1746.650 202.485 1746.770 ;
        RECT 200.715 1746.560 202.485 1746.650 ;
        RECT 198.795 1746.360 198.965 1746.480 ;
        RECT 199.615 1746.310 199.785 1746.545 ;
        RECT 200.325 1746.390 200.495 1746.545 ;
        RECT 201.515 1746.440 202.485 1746.560 ;
        RECT 198.795 1745.970 198.965 1746.190 ;
        RECT 199.140 1746.140 199.785 1746.310 ;
        RECT 198.795 1745.900 199.445 1745.970 ;
        RECT 198.965 1745.730 199.445 1745.900 ;
        RECT 198.795 1745.640 199.445 1745.730 ;
        RECT 198.795 1745.440 198.965 1745.640 ;
        RECT 199.615 1745.470 199.785 1746.140 ;
        RECT 199.135 1745.300 199.785 1745.470 ;
        RECT 198.795 1745.040 198.965 1745.270 ;
      LAYER li1 ;
        RECT 199.955 1745.265 200.155 1746.365 ;
      LAYER li1 ;
        RECT 200.325 1746.060 201.345 1746.390 ;
        RECT 201.515 1746.360 201.685 1746.440 ;
      LAYER li1 ;
        RECT 202.705 1746.355 202.875 1746.940 ;
      LAYER li1 ;
        RECT 203.075 1746.600 203.245 1749.050 ;
        RECT 203.755 1748.960 204.235 1749.120 ;
      LAYER li1 ;
        RECT 203.415 1748.620 204.065 1748.790 ;
      LAYER li1 ;
        RECT 204.235 1748.660 204.405 1748.950 ;
      LAYER li1 ;
        RECT 203.415 1747.950 203.585 1748.620 ;
      LAYER li1 ;
        RECT 204.235 1748.450 204.405 1748.490 ;
        RECT 203.755 1748.200 204.405 1748.450 ;
        RECT 203.755 1748.120 204.235 1748.200 ;
      LAYER li1 ;
        RECT 203.415 1747.780 204.065 1747.950 ;
        RECT 203.415 1747.110 203.585 1747.780 ;
      LAYER li1 ;
        RECT 204.235 1747.740 204.405 1748.030 ;
        RECT 203.755 1747.570 204.235 1747.610 ;
        RECT 203.755 1747.280 204.405 1747.570 ;
      LAYER li1 ;
        RECT 203.415 1746.940 204.065 1747.110 ;
        RECT 203.415 1746.355 203.585 1746.940 ;
      LAYER li1 ;
        RECT 204.235 1746.820 204.405 1747.110 ;
        RECT 203.755 1746.650 204.235 1746.770 ;
        RECT 203.755 1746.440 204.405 1746.650 ;
        RECT 204.235 1746.360 204.405 1746.440 ;
      LAYER li1 ;
        RECT 202.705 1746.270 203.585 1746.355 ;
      LAYER li1 ;
        RECT 200.325 1745.550 200.495 1746.060 ;
        RECT 201.515 1745.930 201.685 1746.190 ;
      LAYER li1 ;
        RECT 201.855 1746.100 204.065 1746.270 ;
      LAYER li1 ;
        RECT 204.235 1745.930 204.405 1746.190 ;
        RECT 201.515 1745.900 202.835 1745.930 ;
        RECT 200.715 1745.730 201.515 1745.890 ;
        RECT 201.685 1745.730 202.835 1745.900 ;
        RECT 200.715 1745.720 202.835 1745.730 ;
        RECT 201.515 1745.600 202.835 1745.720 ;
        RECT 203.435 1745.900 204.405 1745.930 ;
        RECT 203.435 1745.730 204.235 1745.900 ;
        RECT 203.435 1745.600 204.405 1745.730 ;
        RECT 200.325 1745.220 201.345 1745.550 ;
        RECT 201.515 1745.440 201.685 1745.600 ;
        RECT 204.235 1745.440 204.405 1745.600 ;
        RECT 201.515 1745.040 201.685 1745.270 ;
        RECT 204.235 1745.040 204.405 1745.270 ;
        RECT 198.795 1744.980 199.690 1745.040 ;
        RECT 198.965 1744.810 199.690 1744.980 ;
        RECT 198.795 1744.750 199.690 1744.810 ;
        RECT 200.350 1744.980 202.850 1745.040 ;
        RECT 200.350 1744.810 201.515 1744.980 ;
        RECT 201.685 1744.810 202.850 1744.980 ;
        RECT 200.350 1744.750 202.850 1744.810 ;
        RECT 198.795 1744.520 198.965 1744.750 ;
        RECT 201.515 1744.520 201.685 1744.750 ;
        RECT 198.795 1744.190 198.965 1744.350 ;
        RECT 201.515 1744.190 201.685 1744.350 ;
        RECT 201.855 1744.240 202.875 1744.570 ;
        RECT 198.795 1744.060 199.765 1744.190 ;
        RECT 198.965 1743.890 199.765 1744.060 ;
        RECT 198.795 1743.860 199.765 1743.890 ;
        RECT 200.365 1744.070 201.685 1744.190 ;
        RECT 200.365 1744.060 202.485 1744.070 ;
        RECT 200.365 1743.890 201.515 1744.060 ;
        RECT 201.685 1743.900 202.485 1744.060 ;
        RECT 200.365 1743.860 201.685 1743.890 ;
        RECT 198.795 1743.600 198.965 1743.860 ;
      LAYER li1 ;
        RECT 199.135 1743.520 201.345 1743.690 ;
      LAYER li1 ;
        RECT 201.515 1743.600 201.685 1743.860 ;
        RECT 202.705 1743.730 202.875 1744.240 ;
      LAYER li1 ;
        RECT 199.615 1743.435 200.495 1743.520 ;
      LAYER li1 ;
        RECT 198.795 1743.350 198.965 1743.430 ;
        RECT 198.795 1743.140 199.445 1743.350 ;
        RECT 198.965 1743.020 199.445 1743.140 ;
        RECT 198.795 1742.680 198.965 1742.970 ;
      LAYER li1 ;
        RECT 199.615 1742.850 199.785 1743.435 ;
        RECT 199.135 1742.680 199.785 1742.850 ;
      LAYER li1 ;
        RECT 198.795 1742.220 199.445 1742.510 ;
        RECT 198.965 1742.180 199.445 1742.220 ;
        RECT 198.795 1741.760 198.965 1742.050 ;
      LAYER li1 ;
        RECT 199.615 1742.010 199.785 1742.680 ;
        RECT 199.135 1741.840 199.785 1742.010 ;
      LAYER li1 ;
        RECT 198.965 1741.590 199.445 1741.670 ;
        RECT 198.795 1741.340 199.445 1741.590 ;
        RECT 198.795 1741.300 198.965 1741.340 ;
      LAYER li1 ;
        RECT 199.615 1741.170 199.785 1741.840 ;
      LAYER li1 ;
        RECT 198.795 1740.840 198.965 1741.130 ;
      LAYER li1 ;
        RECT 199.135 1741.000 199.785 1741.170 ;
      LAYER li1 ;
        RECT 198.965 1740.670 199.445 1740.830 ;
        RECT 199.955 1740.740 200.125 1743.190 ;
      LAYER li1 ;
        RECT 200.325 1742.850 200.495 1743.435 ;
      LAYER li1 ;
        RECT 201.515 1743.350 201.685 1743.430 ;
        RECT 201.855 1743.400 202.875 1743.730 ;
      LAYER li1 ;
        RECT 203.045 1743.425 203.245 1745.015 ;
      LAYER li1 ;
        RECT 203.510 1744.980 204.405 1745.040 ;
        RECT 203.510 1744.810 204.235 1744.980 ;
        RECT 203.510 1744.750 204.405 1744.810 ;
        RECT 204.235 1744.520 204.405 1744.750 ;
        RECT 203.415 1744.320 204.065 1744.490 ;
        RECT 203.415 1743.650 203.585 1744.320 ;
        RECT 204.235 1744.150 204.405 1744.350 ;
        RECT 203.755 1744.060 204.405 1744.150 ;
        RECT 203.755 1743.890 204.235 1744.060 ;
        RECT 203.755 1743.820 204.405 1743.890 ;
        RECT 203.415 1743.480 204.060 1743.650 ;
        RECT 204.235 1743.600 204.405 1743.820 ;
        RECT 200.715 1743.230 201.685 1743.350 ;
        RECT 202.705 1743.245 202.875 1743.400 ;
        RECT 203.415 1743.245 203.585 1743.480 ;
        RECT 204.235 1743.310 204.405 1743.430 ;
        RECT 200.715 1743.140 202.485 1743.230 ;
        RECT 200.715 1743.020 201.515 1743.140 ;
        RECT 201.685 1743.060 202.485 1743.140 ;
        RECT 202.705 1743.070 203.585 1743.245 ;
        RECT 203.755 1743.140 204.405 1743.310 ;
      LAYER li1 ;
        RECT 200.325 1742.680 201.345 1742.850 ;
      LAYER li1 ;
        RECT 201.515 1742.680 201.685 1742.970 ;
      LAYER li1 ;
        RECT 200.325 1742.010 200.495 1742.680 ;
        RECT 201.855 1742.640 202.875 1742.810 ;
      LAYER li1 ;
        RECT 200.715 1742.470 201.685 1742.510 ;
        RECT 200.715 1742.220 202.485 1742.470 ;
        RECT 200.715 1742.180 201.515 1742.220 ;
        RECT 201.685 1742.140 202.485 1742.220 ;
      LAYER li1 ;
        RECT 200.325 1741.840 201.345 1742.010 ;
        RECT 200.325 1741.170 200.495 1741.840 ;
      LAYER li1 ;
        RECT 201.515 1741.760 201.685 1742.050 ;
      LAYER li1 ;
        RECT 202.705 1741.970 202.875 1742.640 ;
        RECT 201.855 1741.800 202.875 1741.970 ;
      LAYER li1 ;
        RECT 200.715 1741.590 201.515 1741.670 ;
        RECT 201.685 1741.590 202.485 1741.630 ;
        RECT 200.715 1741.340 202.485 1741.590 ;
        RECT 201.515 1741.300 202.485 1741.340 ;
      LAYER li1 ;
        RECT 200.325 1741.000 201.345 1741.170 ;
        RECT 202.705 1741.130 202.875 1741.800 ;
      LAYER li1 ;
        RECT 201.515 1740.840 201.685 1741.130 ;
      LAYER li1 ;
        RECT 201.855 1740.960 202.875 1741.130 ;
      LAYER li1 ;
        RECT 198.795 1740.500 199.445 1740.670 ;
        RECT 199.615 1740.565 200.495 1740.740 ;
        RECT 200.715 1740.670 201.515 1740.750 ;
        RECT 201.685 1740.670 202.485 1740.790 ;
        RECT 200.715 1740.580 202.485 1740.670 ;
        RECT 198.795 1740.380 198.965 1740.500 ;
        RECT 199.615 1740.330 199.785 1740.565 ;
        RECT 200.325 1740.410 200.495 1740.565 ;
        RECT 201.515 1740.460 202.485 1740.580 ;
        RECT 198.795 1739.990 198.965 1740.210 ;
        RECT 199.140 1740.160 199.785 1740.330 ;
        RECT 198.795 1739.920 199.445 1739.990 ;
        RECT 198.965 1739.750 199.445 1739.920 ;
        RECT 198.795 1739.660 199.445 1739.750 ;
        RECT 198.795 1739.460 198.965 1739.660 ;
        RECT 199.615 1739.490 199.785 1740.160 ;
        RECT 199.135 1739.320 199.785 1739.490 ;
        RECT 198.795 1739.060 198.965 1739.290 ;
      LAYER li1 ;
        RECT 199.955 1739.285 200.155 1740.385 ;
      LAYER li1 ;
        RECT 200.325 1740.080 201.345 1740.410 ;
        RECT 201.515 1740.380 201.685 1740.460 ;
      LAYER li1 ;
        RECT 202.705 1740.375 202.875 1740.960 ;
      LAYER li1 ;
        RECT 203.075 1740.620 203.245 1743.070 ;
        RECT 203.755 1742.980 204.235 1743.140 ;
      LAYER li1 ;
        RECT 203.415 1742.640 204.065 1742.810 ;
      LAYER li1 ;
        RECT 204.235 1742.680 204.405 1742.970 ;
      LAYER li1 ;
        RECT 203.415 1741.970 203.585 1742.640 ;
      LAYER li1 ;
        RECT 204.235 1742.470 204.405 1742.510 ;
        RECT 203.755 1742.220 204.405 1742.470 ;
        RECT 203.755 1742.140 204.235 1742.220 ;
      LAYER li1 ;
        RECT 203.415 1741.800 204.065 1741.970 ;
        RECT 203.415 1741.130 203.585 1741.800 ;
      LAYER li1 ;
        RECT 204.235 1741.760 204.405 1742.050 ;
        RECT 203.755 1741.590 204.235 1741.630 ;
        RECT 203.755 1741.300 204.405 1741.590 ;
      LAYER li1 ;
        RECT 203.415 1740.960 204.065 1741.130 ;
        RECT 203.415 1740.375 203.585 1740.960 ;
      LAYER li1 ;
        RECT 204.235 1740.840 204.405 1741.130 ;
        RECT 203.755 1740.670 204.235 1740.790 ;
        RECT 203.755 1740.460 204.405 1740.670 ;
        RECT 204.235 1740.380 204.405 1740.460 ;
      LAYER li1 ;
        RECT 202.705 1740.290 203.585 1740.375 ;
      LAYER li1 ;
        RECT 200.325 1739.570 200.495 1740.080 ;
        RECT 201.515 1739.950 201.685 1740.210 ;
      LAYER li1 ;
        RECT 201.855 1740.120 204.065 1740.290 ;
      LAYER li1 ;
        RECT 204.235 1739.950 204.405 1740.210 ;
        RECT 201.515 1739.920 202.835 1739.950 ;
        RECT 200.715 1739.750 201.515 1739.910 ;
        RECT 201.685 1739.750 202.835 1739.920 ;
        RECT 200.715 1739.740 202.835 1739.750 ;
        RECT 201.515 1739.620 202.835 1739.740 ;
        RECT 203.435 1739.920 204.405 1739.950 ;
        RECT 203.435 1739.750 204.235 1739.920 ;
        RECT 203.435 1739.620 204.405 1739.750 ;
        RECT 200.325 1739.240 201.345 1739.570 ;
        RECT 201.515 1739.460 201.685 1739.620 ;
        RECT 204.235 1739.460 204.405 1739.620 ;
        RECT 201.515 1739.060 201.685 1739.290 ;
        RECT 204.235 1739.060 204.405 1739.290 ;
        RECT 198.795 1739.000 199.690 1739.060 ;
        RECT 198.965 1738.830 199.690 1739.000 ;
        RECT 198.795 1738.770 199.690 1738.830 ;
        RECT 200.350 1739.000 202.850 1739.060 ;
        RECT 200.350 1738.830 201.515 1739.000 ;
        RECT 201.685 1738.830 202.850 1739.000 ;
        RECT 200.350 1738.770 202.850 1738.830 ;
        RECT 198.795 1738.540 198.965 1738.770 ;
        RECT 201.515 1738.540 201.685 1738.770 ;
        RECT 198.795 1738.210 198.965 1738.370 ;
        RECT 201.515 1738.210 201.685 1738.370 ;
        RECT 201.855 1738.260 202.875 1738.590 ;
        RECT 198.795 1738.080 199.765 1738.210 ;
        RECT 198.965 1737.910 199.765 1738.080 ;
        RECT 198.795 1737.880 199.765 1737.910 ;
        RECT 200.365 1738.090 201.685 1738.210 ;
        RECT 200.365 1738.080 202.485 1738.090 ;
        RECT 200.365 1737.910 201.515 1738.080 ;
        RECT 201.685 1737.920 202.485 1738.080 ;
        RECT 200.365 1737.880 201.685 1737.910 ;
        RECT 198.795 1737.620 198.965 1737.880 ;
      LAYER li1 ;
        RECT 199.135 1737.540 201.345 1737.710 ;
      LAYER li1 ;
        RECT 201.515 1737.620 201.685 1737.880 ;
        RECT 202.705 1737.750 202.875 1738.260 ;
      LAYER li1 ;
        RECT 199.615 1737.455 200.495 1737.540 ;
      LAYER li1 ;
        RECT 198.795 1737.370 198.965 1737.450 ;
        RECT 198.795 1737.160 199.445 1737.370 ;
        RECT 198.965 1737.040 199.445 1737.160 ;
        RECT 198.795 1736.700 198.965 1736.990 ;
      LAYER li1 ;
        RECT 199.615 1736.870 199.785 1737.455 ;
        RECT 199.135 1736.700 199.785 1736.870 ;
      LAYER li1 ;
        RECT 198.795 1736.240 199.445 1736.530 ;
        RECT 198.965 1736.200 199.445 1736.240 ;
        RECT 198.795 1735.780 198.965 1736.070 ;
      LAYER li1 ;
        RECT 199.615 1736.030 199.785 1736.700 ;
        RECT 199.135 1735.860 199.785 1736.030 ;
      LAYER li1 ;
        RECT 198.965 1735.610 199.445 1735.690 ;
        RECT 198.795 1735.360 199.445 1735.610 ;
        RECT 198.795 1735.320 198.965 1735.360 ;
      LAYER li1 ;
        RECT 199.615 1735.190 199.785 1735.860 ;
      LAYER li1 ;
        RECT 198.795 1734.860 198.965 1735.150 ;
      LAYER li1 ;
        RECT 199.135 1735.020 199.785 1735.190 ;
      LAYER li1 ;
        RECT 198.965 1734.690 199.445 1734.850 ;
        RECT 199.955 1734.760 200.125 1737.210 ;
      LAYER li1 ;
        RECT 200.325 1736.870 200.495 1737.455 ;
      LAYER li1 ;
        RECT 201.515 1737.370 201.685 1737.450 ;
        RECT 201.855 1737.420 202.875 1737.750 ;
      LAYER li1 ;
        RECT 203.045 1737.445 203.245 1739.035 ;
      LAYER li1 ;
        RECT 203.510 1739.000 204.405 1739.060 ;
        RECT 203.510 1738.830 204.235 1739.000 ;
        RECT 203.510 1738.770 204.405 1738.830 ;
        RECT 204.235 1738.540 204.405 1738.770 ;
        RECT 203.415 1738.340 204.065 1738.510 ;
        RECT 203.415 1737.670 203.585 1738.340 ;
        RECT 204.235 1738.170 204.405 1738.370 ;
        RECT 203.755 1738.080 204.405 1738.170 ;
        RECT 203.755 1737.910 204.235 1738.080 ;
        RECT 203.755 1737.840 204.405 1737.910 ;
        RECT 203.415 1737.500 204.060 1737.670 ;
        RECT 204.235 1737.620 204.405 1737.840 ;
        RECT 200.715 1737.250 201.685 1737.370 ;
        RECT 202.705 1737.265 202.875 1737.420 ;
        RECT 203.415 1737.265 203.585 1737.500 ;
        RECT 204.235 1737.330 204.405 1737.450 ;
        RECT 200.715 1737.160 202.485 1737.250 ;
        RECT 200.715 1737.040 201.515 1737.160 ;
        RECT 201.685 1737.080 202.485 1737.160 ;
        RECT 202.705 1737.090 203.585 1737.265 ;
        RECT 203.755 1737.160 204.405 1737.330 ;
      LAYER li1 ;
        RECT 200.325 1736.700 201.345 1736.870 ;
      LAYER li1 ;
        RECT 201.515 1736.700 201.685 1736.990 ;
      LAYER li1 ;
        RECT 200.325 1736.030 200.495 1736.700 ;
        RECT 201.855 1736.660 202.875 1736.830 ;
      LAYER li1 ;
        RECT 200.715 1736.490 201.685 1736.530 ;
        RECT 200.715 1736.240 202.485 1736.490 ;
        RECT 200.715 1736.200 201.515 1736.240 ;
        RECT 201.685 1736.160 202.485 1736.240 ;
      LAYER li1 ;
        RECT 200.325 1735.860 201.345 1736.030 ;
        RECT 200.325 1735.190 200.495 1735.860 ;
      LAYER li1 ;
        RECT 201.515 1735.780 201.685 1736.070 ;
      LAYER li1 ;
        RECT 202.705 1735.990 202.875 1736.660 ;
        RECT 201.855 1735.820 202.875 1735.990 ;
      LAYER li1 ;
        RECT 200.715 1735.610 201.515 1735.690 ;
        RECT 201.685 1735.610 202.485 1735.650 ;
        RECT 200.715 1735.360 202.485 1735.610 ;
        RECT 201.515 1735.320 202.485 1735.360 ;
      LAYER li1 ;
        RECT 200.325 1735.020 201.345 1735.190 ;
        RECT 202.705 1735.150 202.875 1735.820 ;
      LAYER li1 ;
        RECT 201.515 1734.860 201.685 1735.150 ;
      LAYER li1 ;
        RECT 201.855 1734.980 202.875 1735.150 ;
      LAYER li1 ;
        RECT 198.795 1734.520 199.445 1734.690 ;
        RECT 199.615 1734.585 200.495 1734.760 ;
        RECT 200.715 1734.690 201.515 1734.770 ;
        RECT 201.685 1734.690 202.485 1734.810 ;
        RECT 200.715 1734.600 202.485 1734.690 ;
        RECT 198.795 1734.400 198.965 1734.520 ;
        RECT 199.615 1734.350 199.785 1734.585 ;
        RECT 200.325 1734.430 200.495 1734.585 ;
        RECT 201.515 1734.480 202.485 1734.600 ;
        RECT 198.795 1734.010 198.965 1734.230 ;
        RECT 199.140 1734.180 199.785 1734.350 ;
        RECT 198.795 1733.940 199.445 1734.010 ;
        RECT 198.965 1733.770 199.445 1733.940 ;
        RECT 198.795 1733.680 199.445 1733.770 ;
        RECT 198.795 1733.480 198.965 1733.680 ;
        RECT 199.615 1733.510 199.785 1734.180 ;
        RECT 199.135 1733.340 199.785 1733.510 ;
        RECT 198.795 1733.080 198.965 1733.310 ;
      LAYER li1 ;
        RECT 199.955 1733.305 200.155 1734.405 ;
      LAYER li1 ;
        RECT 200.325 1734.100 201.345 1734.430 ;
        RECT 201.515 1734.400 201.685 1734.480 ;
      LAYER li1 ;
        RECT 202.705 1734.395 202.875 1734.980 ;
      LAYER li1 ;
        RECT 203.075 1734.640 203.245 1737.090 ;
        RECT 203.755 1737.000 204.235 1737.160 ;
      LAYER li1 ;
        RECT 203.415 1736.660 204.065 1736.830 ;
      LAYER li1 ;
        RECT 204.235 1736.700 204.405 1736.990 ;
      LAYER li1 ;
        RECT 203.415 1735.990 203.585 1736.660 ;
      LAYER li1 ;
        RECT 204.235 1736.490 204.405 1736.530 ;
        RECT 203.755 1736.240 204.405 1736.490 ;
        RECT 203.755 1736.160 204.235 1736.240 ;
      LAYER li1 ;
        RECT 203.415 1735.820 204.065 1735.990 ;
        RECT 203.415 1735.150 203.585 1735.820 ;
      LAYER li1 ;
        RECT 204.235 1735.780 204.405 1736.070 ;
        RECT 203.755 1735.610 204.235 1735.650 ;
        RECT 203.755 1735.320 204.405 1735.610 ;
      LAYER li1 ;
        RECT 203.415 1734.980 204.065 1735.150 ;
        RECT 203.415 1734.395 203.585 1734.980 ;
      LAYER li1 ;
        RECT 204.235 1734.860 204.405 1735.150 ;
        RECT 203.755 1734.690 204.235 1734.810 ;
        RECT 203.755 1734.480 204.405 1734.690 ;
        RECT 204.235 1734.400 204.405 1734.480 ;
      LAYER li1 ;
        RECT 202.705 1734.310 203.585 1734.395 ;
      LAYER li1 ;
        RECT 200.325 1733.590 200.495 1734.100 ;
        RECT 201.515 1733.970 201.685 1734.230 ;
      LAYER li1 ;
        RECT 201.855 1734.140 204.065 1734.310 ;
      LAYER li1 ;
        RECT 204.235 1733.970 204.405 1734.230 ;
        RECT 201.515 1733.940 202.835 1733.970 ;
        RECT 200.715 1733.770 201.515 1733.930 ;
        RECT 201.685 1733.770 202.835 1733.940 ;
        RECT 200.715 1733.760 202.835 1733.770 ;
        RECT 201.515 1733.640 202.835 1733.760 ;
        RECT 203.435 1733.940 204.405 1733.970 ;
        RECT 203.435 1733.770 204.235 1733.940 ;
        RECT 203.435 1733.640 204.405 1733.770 ;
        RECT 200.325 1733.260 201.345 1733.590 ;
        RECT 201.515 1733.480 201.685 1733.640 ;
        RECT 204.235 1733.480 204.405 1733.640 ;
        RECT 201.515 1733.080 201.685 1733.310 ;
        RECT 204.235 1733.080 204.405 1733.310 ;
        RECT 198.795 1733.020 199.690 1733.080 ;
        RECT 198.965 1732.850 199.690 1733.020 ;
        RECT 198.795 1732.790 199.690 1732.850 ;
        RECT 200.350 1733.020 202.850 1733.080 ;
        RECT 200.350 1732.850 201.515 1733.020 ;
        RECT 201.685 1732.850 202.850 1733.020 ;
        RECT 200.350 1732.790 202.850 1732.850 ;
        RECT 198.795 1732.560 198.965 1732.790 ;
        RECT 201.515 1732.560 201.685 1732.790 ;
        RECT 198.795 1732.230 198.965 1732.390 ;
        RECT 201.515 1732.230 201.685 1732.390 ;
        RECT 201.855 1732.280 202.875 1732.610 ;
        RECT 198.795 1732.100 199.765 1732.230 ;
        RECT 198.965 1731.930 199.765 1732.100 ;
        RECT 198.795 1731.900 199.765 1731.930 ;
        RECT 200.365 1732.110 201.685 1732.230 ;
        RECT 200.365 1732.100 202.485 1732.110 ;
        RECT 200.365 1731.930 201.515 1732.100 ;
        RECT 201.685 1731.940 202.485 1732.100 ;
        RECT 200.365 1731.900 201.685 1731.930 ;
        RECT 198.795 1731.640 198.965 1731.900 ;
      LAYER li1 ;
        RECT 199.135 1731.560 201.345 1731.730 ;
      LAYER li1 ;
        RECT 201.515 1731.640 201.685 1731.900 ;
        RECT 202.705 1731.770 202.875 1732.280 ;
      LAYER li1 ;
        RECT 199.615 1731.475 200.495 1731.560 ;
      LAYER li1 ;
        RECT 198.795 1731.390 198.965 1731.470 ;
        RECT 198.795 1731.180 199.445 1731.390 ;
        RECT 198.965 1731.060 199.445 1731.180 ;
        RECT 198.795 1730.720 198.965 1731.010 ;
      LAYER li1 ;
        RECT 199.615 1730.890 199.785 1731.475 ;
        RECT 199.135 1730.720 199.785 1730.890 ;
      LAYER li1 ;
        RECT 198.795 1730.260 199.445 1730.550 ;
        RECT 198.965 1730.220 199.445 1730.260 ;
        RECT 198.795 1729.800 198.965 1730.090 ;
      LAYER li1 ;
        RECT 199.615 1730.050 199.785 1730.720 ;
        RECT 199.135 1729.880 199.785 1730.050 ;
      LAYER li1 ;
        RECT 198.965 1729.630 199.445 1729.710 ;
        RECT 198.795 1729.380 199.445 1729.630 ;
        RECT 198.795 1729.340 198.965 1729.380 ;
      LAYER li1 ;
        RECT 199.615 1729.210 199.785 1729.880 ;
      LAYER li1 ;
        RECT 198.795 1728.880 198.965 1729.170 ;
      LAYER li1 ;
        RECT 199.135 1729.040 199.785 1729.210 ;
      LAYER li1 ;
        RECT 198.965 1728.710 199.445 1728.870 ;
        RECT 199.955 1728.780 200.125 1731.230 ;
      LAYER li1 ;
        RECT 200.325 1730.890 200.495 1731.475 ;
      LAYER li1 ;
        RECT 201.515 1731.390 201.685 1731.470 ;
        RECT 201.855 1731.440 202.875 1731.770 ;
      LAYER li1 ;
        RECT 203.045 1731.465 203.245 1733.055 ;
      LAYER li1 ;
        RECT 203.510 1733.020 204.405 1733.080 ;
        RECT 203.510 1732.850 204.235 1733.020 ;
        RECT 203.510 1732.790 204.405 1732.850 ;
        RECT 204.235 1732.560 204.405 1732.790 ;
        RECT 203.415 1732.360 204.065 1732.530 ;
        RECT 203.415 1731.690 203.585 1732.360 ;
        RECT 204.235 1732.190 204.405 1732.390 ;
        RECT 203.755 1732.100 204.405 1732.190 ;
        RECT 203.755 1731.930 204.235 1732.100 ;
        RECT 203.755 1731.860 204.405 1731.930 ;
        RECT 203.415 1731.520 204.060 1731.690 ;
        RECT 204.235 1731.640 204.405 1731.860 ;
        RECT 200.715 1731.270 201.685 1731.390 ;
        RECT 202.705 1731.285 202.875 1731.440 ;
        RECT 203.415 1731.285 203.585 1731.520 ;
        RECT 204.235 1731.350 204.405 1731.470 ;
        RECT 200.715 1731.180 202.485 1731.270 ;
        RECT 200.715 1731.060 201.515 1731.180 ;
        RECT 201.685 1731.100 202.485 1731.180 ;
        RECT 202.705 1731.110 203.585 1731.285 ;
        RECT 203.755 1731.180 204.405 1731.350 ;
      LAYER li1 ;
        RECT 200.325 1730.720 201.345 1730.890 ;
      LAYER li1 ;
        RECT 201.515 1730.720 201.685 1731.010 ;
      LAYER li1 ;
        RECT 200.325 1730.050 200.495 1730.720 ;
        RECT 201.855 1730.680 202.875 1730.850 ;
      LAYER li1 ;
        RECT 200.715 1730.510 201.685 1730.550 ;
        RECT 200.715 1730.260 202.485 1730.510 ;
        RECT 200.715 1730.220 201.515 1730.260 ;
        RECT 201.685 1730.180 202.485 1730.260 ;
      LAYER li1 ;
        RECT 200.325 1729.880 201.345 1730.050 ;
        RECT 200.325 1729.210 200.495 1729.880 ;
      LAYER li1 ;
        RECT 201.515 1729.800 201.685 1730.090 ;
      LAYER li1 ;
        RECT 202.705 1730.010 202.875 1730.680 ;
        RECT 201.855 1729.840 202.875 1730.010 ;
      LAYER li1 ;
        RECT 200.715 1729.630 201.515 1729.710 ;
        RECT 201.685 1729.630 202.485 1729.670 ;
        RECT 200.715 1729.380 202.485 1729.630 ;
        RECT 201.515 1729.340 202.485 1729.380 ;
      LAYER li1 ;
        RECT 200.325 1729.040 201.345 1729.210 ;
        RECT 202.705 1729.170 202.875 1729.840 ;
      LAYER li1 ;
        RECT 201.515 1728.880 201.685 1729.170 ;
      LAYER li1 ;
        RECT 201.855 1729.000 202.875 1729.170 ;
      LAYER li1 ;
        RECT 198.795 1728.540 199.445 1728.710 ;
        RECT 199.615 1728.605 200.495 1728.780 ;
        RECT 200.715 1728.710 201.515 1728.790 ;
        RECT 201.685 1728.710 202.485 1728.830 ;
        RECT 200.715 1728.620 202.485 1728.710 ;
        RECT 198.795 1728.420 198.965 1728.540 ;
        RECT 199.615 1728.370 199.785 1728.605 ;
        RECT 200.325 1728.450 200.495 1728.605 ;
        RECT 201.515 1728.500 202.485 1728.620 ;
        RECT 198.795 1728.030 198.965 1728.250 ;
        RECT 199.140 1728.200 199.785 1728.370 ;
        RECT 198.795 1727.960 199.445 1728.030 ;
        RECT 198.965 1727.790 199.445 1727.960 ;
        RECT 198.795 1727.700 199.445 1727.790 ;
        RECT 198.795 1727.500 198.965 1727.700 ;
        RECT 199.615 1727.530 199.785 1728.200 ;
        RECT 199.135 1727.360 199.785 1727.530 ;
        RECT 198.795 1727.100 198.965 1727.330 ;
      LAYER li1 ;
        RECT 199.955 1727.325 200.155 1728.425 ;
      LAYER li1 ;
        RECT 200.325 1728.120 201.345 1728.450 ;
        RECT 201.515 1728.420 201.685 1728.500 ;
      LAYER li1 ;
        RECT 202.705 1728.415 202.875 1729.000 ;
      LAYER li1 ;
        RECT 203.075 1728.660 203.245 1731.110 ;
        RECT 203.755 1731.020 204.235 1731.180 ;
      LAYER li1 ;
        RECT 203.415 1730.680 204.065 1730.850 ;
      LAYER li1 ;
        RECT 204.235 1730.720 204.405 1731.010 ;
      LAYER li1 ;
        RECT 203.415 1730.010 203.585 1730.680 ;
      LAYER li1 ;
        RECT 204.235 1730.510 204.405 1730.550 ;
        RECT 203.755 1730.260 204.405 1730.510 ;
        RECT 203.755 1730.180 204.235 1730.260 ;
      LAYER li1 ;
        RECT 203.415 1729.840 204.065 1730.010 ;
        RECT 203.415 1729.170 203.585 1729.840 ;
      LAYER li1 ;
        RECT 204.235 1729.800 204.405 1730.090 ;
        RECT 203.755 1729.630 204.235 1729.670 ;
        RECT 203.755 1729.340 204.405 1729.630 ;
      LAYER li1 ;
        RECT 203.415 1729.000 204.065 1729.170 ;
        RECT 203.415 1728.415 203.585 1729.000 ;
      LAYER li1 ;
        RECT 204.235 1728.880 204.405 1729.170 ;
        RECT 203.755 1728.710 204.235 1728.830 ;
        RECT 203.755 1728.500 204.405 1728.710 ;
        RECT 204.235 1728.420 204.405 1728.500 ;
      LAYER li1 ;
        RECT 202.705 1728.330 203.585 1728.415 ;
      LAYER li1 ;
        RECT 200.325 1727.610 200.495 1728.120 ;
        RECT 201.515 1727.990 201.685 1728.250 ;
      LAYER li1 ;
        RECT 201.855 1728.160 204.065 1728.330 ;
      LAYER li1 ;
        RECT 204.235 1727.990 204.405 1728.250 ;
        RECT 201.515 1727.960 202.835 1727.990 ;
        RECT 200.715 1727.790 201.515 1727.950 ;
        RECT 201.685 1727.790 202.835 1727.960 ;
        RECT 200.715 1727.780 202.835 1727.790 ;
        RECT 201.515 1727.660 202.835 1727.780 ;
        RECT 203.435 1727.960 204.405 1727.990 ;
        RECT 203.435 1727.790 204.235 1727.960 ;
        RECT 203.435 1727.660 204.405 1727.790 ;
        RECT 200.325 1727.280 201.345 1727.610 ;
        RECT 201.515 1727.500 201.685 1727.660 ;
        RECT 204.235 1727.500 204.405 1727.660 ;
        RECT 201.515 1727.100 201.685 1727.330 ;
        RECT 204.235 1727.100 204.405 1727.330 ;
        RECT 198.795 1727.040 199.690 1727.100 ;
        RECT 198.965 1726.870 199.690 1727.040 ;
        RECT 198.795 1726.810 199.690 1726.870 ;
        RECT 200.350 1727.040 202.850 1727.100 ;
        RECT 200.350 1726.870 201.515 1727.040 ;
        RECT 201.685 1726.870 202.850 1727.040 ;
        RECT 200.350 1726.810 202.850 1726.870 ;
        RECT 198.795 1726.580 198.965 1726.810 ;
        RECT 201.515 1726.580 201.685 1726.810 ;
        RECT 198.795 1726.250 198.965 1726.410 ;
        RECT 201.515 1726.250 201.685 1726.410 ;
        RECT 201.855 1726.300 202.875 1726.630 ;
        RECT 198.795 1726.120 199.765 1726.250 ;
        RECT 198.965 1725.950 199.765 1726.120 ;
        RECT 198.795 1725.920 199.765 1725.950 ;
        RECT 200.365 1726.130 201.685 1726.250 ;
        RECT 200.365 1726.120 202.485 1726.130 ;
        RECT 200.365 1725.950 201.515 1726.120 ;
        RECT 201.685 1725.960 202.485 1726.120 ;
        RECT 200.365 1725.920 201.685 1725.950 ;
        RECT 198.795 1725.660 198.965 1725.920 ;
      LAYER li1 ;
        RECT 199.135 1725.580 201.345 1725.750 ;
      LAYER li1 ;
        RECT 201.515 1725.660 201.685 1725.920 ;
        RECT 202.705 1725.790 202.875 1726.300 ;
      LAYER li1 ;
        RECT 199.615 1725.495 200.495 1725.580 ;
      LAYER li1 ;
        RECT 198.795 1725.410 198.965 1725.490 ;
        RECT 198.795 1725.200 199.445 1725.410 ;
        RECT 198.965 1725.080 199.445 1725.200 ;
        RECT 198.795 1724.740 198.965 1725.030 ;
      LAYER li1 ;
        RECT 199.615 1724.910 199.785 1725.495 ;
        RECT 199.135 1724.740 199.785 1724.910 ;
      LAYER li1 ;
        RECT 198.795 1724.280 199.445 1724.570 ;
        RECT 198.965 1724.240 199.445 1724.280 ;
        RECT 198.795 1723.820 198.965 1724.110 ;
      LAYER li1 ;
        RECT 199.615 1724.070 199.785 1724.740 ;
        RECT 199.135 1723.900 199.785 1724.070 ;
      LAYER li1 ;
        RECT 198.965 1723.650 199.445 1723.730 ;
        RECT 198.795 1723.400 199.445 1723.650 ;
        RECT 198.795 1723.360 198.965 1723.400 ;
      LAYER li1 ;
        RECT 199.615 1723.230 199.785 1723.900 ;
      LAYER li1 ;
        RECT 198.795 1722.900 198.965 1723.190 ;
      LAYER li1 ;
        RECT 199.135 1723.060 199.785 1723.230 ;
      LAYER li1 ;
        RECT 198.965 1722.730 199.445 1722.890 ;
        RECT 199.955 1722.800 200.125 1725.250 ;
      LAYER li1 ;
        RECT 200.325 1724.910 200.495 1725.495 ;
      LAYER li1 ;
        RECT 201.515 1725.410 201.685 1725.490 ;
        RECT 201.855 1725.460 202.875 1725.790 ;
      LAYER li1 ;
        RECT 203.045 1725.485 203.245 1727.075 ;
      LAYER li1 ;
        RECT 203.510 1727.040 204.405 1727.100 ;
        RECT 203.510 1726.870 204.235 1727.040 ;
        RECT 203.510 1726.810 204.405 1726.870 ;
        RECT 204.235 1726.580 204.405 1726.810 ;
        RECT 203.415 1726.380 204.065 1726.550 ;
        RECT 203.415 1725.710 203.585 1726.380 ;
        RECT 204.235 1726.210 204.405 1726.410 ;
        RECT 203.755 1726.120 204.405 1726.210 ;
        RECT 203.755 1725.950 204.235 1726.120 ;
        RECT 203.755 1725.880 204.405 1725.950 ;
        RECT 203.415 1725.540 204.060 1725.710 ;
        RECT 204.235 1725.660 204.405 1725.880 ;
        RECT 200.715 1725.290 201.685 1725.410 ;
        RECT 202.705 1725.305 202.875 1725.460 ;
        RECT 203.415 1725.305 203.585 1725.540 ;
        RECT 204.235 1725.370 204.405 1725.490 ;
        RECT 200.715 1725.200 202.485 1725.290 ;
        RECT 200.715 1725.080 201.515 1725.200 ;
        RECT 201.685 1725.120 202.485 1725.200 ;
        RECT 202.705 1725.130 203.585 1725.305 ;
        RECT 203.755 1725.200 204.405 1725.370 ;
      LAYER li1 ;
        RECT 200.325 1724.740 201.345 1724.910 ;
      LAYER li1 ;
        RECT 201.515 1724.740 201.685 1725.030 ;
      LAYER li1 ;
        RECT 200.325 1724.070 200.495 1724.740 ;
        RECT 201.855 1724.700 202.875 1724.870 ;
      LAYER li1 ;
        RECT 200.715 1724.530 201.685 1724.570 ;
        RECT 200.715 1724.280 202.485 1724.530 ;
        RECT 200.715 1724.240 201.515 1724.280 ;
        RECT 201.685 1724.200 202.485 1724.280 ;
      LAYER li1 ;
        RECT 200.325 1723.900 201.345 1724.070 ;
        RECT 200.325 1723.230 200.495 1723.900 ;
      LAYER li1 ;
        RECT 201.515 1723.820 201.685 1724.110 ;
      LAYER li1 ;
        RECT 202.705 1724.030 202.875 1724.700 ;
        RECT 201.855 1723.860 202.875 1724.030 ;
      LAYER li1 ;
        RECT 200.715 1723.650 201.515 1723.730 ;
        RECT 201.685 1723.650 202.485 1723.690 ;
        RECT 200.715 1723.400 202.485 1723.650 ;
        RECT 201.515 1723.360 202.485 1723.400 ;
      LAYER li1 ;
        RECT 200.325 1723.060 201.345 1723.230 ;
        RECT 202.705 1723.190 202.875 1723.860 ;
      LAYER li1 ;
        RECT 201.515 1722.900 201.685 1723.190 ;
      LAYER li1 ;
        RECT 201.855 1723.020 202.875 1723.190 ;
      LAYER li1 ;
        RECT 198.795 1722.560 199.445 1722.730 ;
        RECT 199.615 1722.625 200.495 1722.800 ;
        RECT 200.715 1722.730 201.515 1722.810 ;
        RECT 201.685 1722.730 202.485 1722.850 ;
        RECT 200.715 1722.640 202.485 1722.730 ;
        RECT 198.795 1722.440 198.965 1722.560 ;
        RECT 199.615 1722.390 199.785 1722.625 ;
        RECT 200.325 1722.470 200.495 1722.625 ;
        RECT 201.515 1722.520 202.485 1722.640 ;
        RECT 198.795 1722.050 198.965 1722.270 ;
        RECT 199.140 1722.220 199.785 1722.390 ;
        RECT 198.795 1721.980 199.445 1722.050 ;
        RECT 198.965 1721.810 199.445 1721.980 ;
        RECT 198.795 1721.720 199.445 1721.810 ;
        RECT 198.795 1721.520 198.965 1721.720 ;
        RECT 199.615 1721.550 199.785 1722.220 ;
        RECT 199.135 1721.380 199.785 1721.550 ;
        RECT 198.795 1721.120 198.965 1721.350 ;
      LAYER li1 ;
        RECT 199.955 1721.345 200.155 1722.445 ;
      LAYER li1 ;
        RECT 200.325 1722.140 201.345 1722.470 ;
        RECT 201.515 1722.440 201.685 1722.520 ;
      LAYER li1 ;
        RECT 202.705 1722.435 202.875 1723.020 ;
      LAYER li1 ;
        RECT 203.075 1722.680 203.245 1725.130 ;
        RECT 203.755 1725.040 204.235 1725.200 ;
      LAYER li1 ;
        RECT 203.415 1724.700 204.065 1724.870 ;
      LAYER li1 ;
        RECT 204.235 1724.740 204.405 1725.030 ;
      LAYER li1 ;
        RECT 203.415 1724.030 203.585 1724.700 ;
      LAYER li1 ;
        RECT 204.235 1724.530 204.405 1724.570 ;
        RECT 203.755 1724.280 204.405 1724.530 ;
        RECT 203.755 1724.200 204.235 1724.280 ;
      LAYER li1 ;
        RECT 203.415 1723.860 204.065 1724.030 ;
        RECT 203.415 1723.190 203.585 1723.860 ;
      LAYER li1 ;
        RECT 204.235 1723.820 204.405 1724.110 ;
        RECT 203.755 1723.650 204.235 1723.690 ;
        RECT 203.755 1723.360 204.405 1723.650 ;
      LAYER li1 ;
        RECT 203.415 1723.020 204.065 1723.190 ;
        RECT 203.415 1722.435 203.585 1723.020 ;
      LAYER li1 ;
        RECT 204.235 1722.900 204.405 1723.190 ;
        RECT 203.755 1722.730 204.235 1722.850 ;
        RECT 203.755 1722.520 204.405 1722.730 ;
        RECT 204.235 1722.440 204.405 1722.520 ;
      LAYER li1 ;
        RECT 202.705 1722.350 203.585 1722.435 ;
      LAYER li1 ;
        RECT 200.325 1721.630 200.495 1722.140 ;
        RECT 201.515 1722.010 201.685 1722.270 ;
      LAYER li1 ;
        RECT 201.855 1722.180 204.065 1722.350 ;
      LAYER li1 ;
        RECT 204.235 1722.010 204.405 1722.270 ;
        RECT 201.515 1721.980 202.835 1722.010 ;
        RECT 200.715 1721.810 201.515 1721.970 ;
        RECT 201.685 1721.810 202.835 1721.980 ;
        RECT 200.715 1721.800 202.835 1721.810 ;
        RECT 201.515 1721.680 202.835 1721.800 ;
        RECT 203.435 1721.980 204.405 1722.010 ;
        RECT 203.435 1721.810 204.235 1721.980 ;
        RECT 203.435 1721.680 204.405 1721.810 ;
        RECT 200.325 1721.300 201.345 1721.630 ;
        RECT 201.515 1721.520 201.685 1721.680 ;
        RECT 204.235 1721.520 204.405 1721.680 ;
        RECT 201.515 1721.120 201.685 1721.350 ;
        RECT 204.235 1721.120 204.405 1721.350 ;
        RECT 198.795 1721.060 199.690 1721.120 ;
        RECT 198.965 1720.890 199.690 1721.060 ;
        RECT 198.795 1720.830 199.690 1720.890 ;
        RECT 200.350 1721.060 202.850 1721.120 ;
        RECT 200.350 1720.890 201.515 1721.060 ;
        RECT 201.685 1720.890 202.850 1721.060 ;
        RECT 200.350 1720.830 202.850 1720.890 ;
        RECT 198.795 1720.600 198.965 1720.830 ;
        RECT 201.515 1720.600 201.685 1720.830 ;
        RECT 198.795 1720.270 198.965 1720.430 ;
        RECT 201.515 1720.270 201.685 1720.430 ;
        RECT 201.855 1720.320 202.875 1720.650 ;
        RECT 198.795 1720.140 199.765 1720.270 ;
        RECT 198.965 1719.970 199.765 1720.140 ;
        RECT 198.795 1719.940 199.765 1719.970 ;
        RECT 200.365 1720.150 201.685 1720.270 ;
        RECT 200.365 1720.140 202.485 1720.150 ;
        RECT 200.365 1719.970 201.515 1720.140 ;
        RECT 201.685 1719.980 202.485 1720.140 ;
        RECT 200.365 1719.940 201.685 1719.970 ;
        RECT 198.795 1719.680 198.965 1719.940 ;
      LAYER li1 ;
        RECT 199.135 1719.600 201.345 1719.770 ;
      LAYER li1 ;
        RECT 201.515 1719.680 201.685 1719.940 ;
        RECT 202.705 1719.810 202.875 1720.320 ;
      LAYER li1 ;
        RECT 199.615 1719.515 200.495 1719.600 ;
      LAYER li1 ;
        RECT 198.795 1719.430 198.965 1719.510 ;
        RECT 198.795 1719.220 199.445 1719.430 ;
        RECT 198.965 1719.100 199.445 1719.220 ;
        RECT 198.795 1718.760 198.965 1719.050 ;
      LAYER li1 ;
        RECT 199.615 1718.930 199.785 1719.515 ;
        RECT 199.135 1718.760 199.785 1718.930 ;
      LAYER li1 ;
        RECT 198.795 1718.300 199.445 1718.590 ;
        RECT 198.965 1718.260 199.445 1718.300 ;
        RECT 198.795 1717.840 198.965 1718.130 ;
      LAYER li1 ;
        RECT 199.615 1718.090 199.785 1718.760 ;
        RECT 199.135 1717.920 199.785 1718.090 ;
      LAYER li1 ;
        RECT 198.965 1717.670 199.445 1717.750 ;
        RECT 198.795 1717.420 199.445 1717.670 ;
        RECT 198.795 1717.380 198.965 1717.420 ;
      LAYER li1 ;
        RECT 199.615 1717.250 199.785 1717.920 ;
      LAYER li1 ;
        RECT 198.795 1716.920 198.965 1717.210 ;
      LAYER li1 ;
        RECT 199.135 1717.080 199.785 1717.250 ;
      LAYER li1 ;
        RECT 198.965 1716.750 199.445 1716.910 ;
        RECT 199.955 1716.820 200.125 1719.270 ;
      LAYER li1 ;
        RECT 200.325 1718.930 200.495 1719.515 ;
      LAYER li1 ;
        RECT 201.515 1719.430 201.685 1719.510 ;
        RECT 201.855 1719.480 202.875 1719.810 ;
      LAYER li1 ;
        RECT 203.045 1719.505 203.245 1721.095 ;
      LAYER li1 ;
        RECT 203.510 1721.060 204.405 1721.120 ;
        RECT 203.510 1720.890 204.235 1721.060 ;
        RECT 203.510 1720.830 204.405 1720.890 ;
        RECT 204.235 1720.600 204.405 1720.830 ;
        RECT 203.415 1720.400 204.065 1720.570 ;
        RECT 203.415 1719.730 203.585 1720.400 ;
        RECT 204.235 1720.230 204.405 1720.430 ;
        RECT 203.755 1720.140 204.405 1720.230 ;
        RECT 203.755 1719.970 204.235 1720.140 ;
        RECT 203.755 1719.900 204.405 1719.970 ;
        RECT 203.415 1719.560 204.060 1719.730 ;
        RECT 204.235 1719.680 204.405 1719.900 ;
        RECT 200.715 1719.310 201.685 1719.430 ;
        RECT 202.705 1719.325 202.875 1719.480 ;
        RECT 203.415 1719.325 203.585 1719.560 ;
        RECT 204.235 1719.390 204.405 1719.510 ;
        RECT 200.715 1719.220 202.485 1719.310 ;
        RECT 200.715 1719.100 201.515 1719.220 ;
        RECT 201.685 1719.140 202.485 1719.220 ;
        RECT 202.705 1719.150 203.585 1719.325 ;
        RECT 203.755 1719.220 204.405 1719.390 ;
      LAYER li1 ;
        RECT 200.325 1718.760 201.345 1718.930 ;
      LAYER li1 ;
        RECT 201.515 1718.760 201.685 1719.050 ;
      LAYER li1 ;
        RECT 200.325 1718.090 200.495 1718.760 ;
        RECT 201.855 1718.720 202.875 1718.890 ;
      LAYER li1 ;
        RECT 200.715 1718.550 201.685 1718.590 ;
        RECT 200.715 1718.300 202.485 1718.550 ;
        RECT 200.715 1718.260 201.515 1718.300 ;
        RECT 201.685 1718.220 202.485 1718.300 ;
      LAYER li1 ;
        RECT 200.325 1717.920 201.345 1718.090 ;
        RECT 200.325 1717.250 200.495 1717.920 ;
      LAYER li1 ;
        RECT 201.515 1717.840 201.685 1718.130 ;
      LAYER li1 ;
        RECT 202.705 1718.050 202.875 1718.720 ;
        RECT 201.855 1717.880 202.875 1718.050 ;
      LAYER li1 ;
        RECT 200.715 1717.670 201.515 1717.750 ;
        RECT 201.685 1717.670 202.485 1717.710 ;
        RECT 200.715 1717.420 202.485 1717.670 ;
        RECT 201.515 1717.380 202.485 1717.420 ;
      LAYER li1 ;
        RECT 200.325 1717.080 201.345 1717.250 ;
        RECT 202.705 1717.210 202.875 1717.880 ;
      LAYER li1 ;
        RECT 201.515 1716.920 201.685 1717.210 ;
      LAYER li1 ;
        RECT 201.855 1717.040 202.875 1717.210 ;
      LAYER li1 ;
        RECT 198.795 1716.580 199.445 1716.750 ;
        RECT 199.615 1716.645 200.495 1716.820 ;
        RECT 200.715 1716.750 201.515 1716.830 ;
        RECT 201.685 1716.750 202.485 1716.870 ;
        RECT 200.715 1716.660 202.485 1716.750 ;
        RECT 198.795 1716.460 198.965 1716.580 ;
        RECT 199.615 1716.410 199.785 1716.645 ;
        RECT 200.325 1716.490 200.495 1716.645 ;
        RECT 201.515 1716.540 202.485 1716.660 ;
        RECT 198.795 1716.070 198.965 1716.290 ;
        RECT 199.140 1716.240 199.785 1716.410 ;
        RECT 198.795 1716.000 199.445 1716.070 ;
        RECT 198.965 1715.830 199.445 1716.000 ;
        RECT 198.795 1715.740 199.445 1715.830 ;
        RECT 198.795 1715.540 198.965 1715.740 ;
        RECT 199.615 1715.570 199.785 1716.240 ;
        RECT 199.135 1715.400 199.785 1715.570 ;
        RECT 198.795 1715.140 198.965 1715.370 ;
      LAYER li1 ;
        RECT 199.955 1715.365 200.155 1716.465 ;
      LAYER li1 ;
        RECT 200.325 1716.160 201.345 1716.490 ;
        RECT 201.515 1716.460 201.685 1716.540 ;
      LAYER li1 ;
        RECT 202.705 1716.455 202.875 1717.040 ;
      LAYER li1 ;
        RECT 203.075 1716.700 203.245 1719.150 ;
        RECT 203.755 1719.060 204.235 1719.220 ;
      LAYER li1 ;
        RECT 203.415 1718.720 204.065 1718.890 ;
      LAYER li1 ;
        RECT 204.235 1718.760 204.405 1719.050 ;
      LAYER li1 ;
        RECT 203.415 1718.050 203.585 1718.720 ;
      LAYER li1 ;
        RECT 204.235 1718.550 204.405 1718.590 ;
        RECT 203.755 1718.300 204.405 1718.550 ;
        RECT 203.755 1718.220 204.235 1718.300 ;
      LAYER li1 ;
        RECT 203.415 1717.880 204.065 1718.050 ;
        RECT 203.415 1717.210 203.585 1717.880 ;
      LAYER li1 ;
        RECT 204.235 1717.840 204.405 1718.130 ;
        RECT 203.755 1717.670 204.235 1717.710 ;
        RECT 203.755 1717.380 204.405 1717.670 ;
      LAYER li1 ;
        RECT 203.415 1717.040 204.065 1717.210 ;
        RECT 203.415 1716.455 203.585 1717.040 ;
      LAYER li1 ;
        RECT 204.235 1716.920 204.405 1717.210 ;
        RECT 203.755 1716.750 204.235 1716.870 ;
        RECT 203.755 1716.540 204.405 1716.750 ;
        RECT 204.235 1716.460 204.405 1716.540 ;
      LAYER li1 ;
        RECT 202.705 1716.370 203.585 1716.455 ;
      LAYER li1 ;
        RECT 200.325 1715.650 200.495 1716.160 ;
        RECT 201.515 1716.030 201.685 1716.290 ;
      LAYER li1 ;
        RECT 201.855 1716.200 204.065 1716.370 ;
      LAYER li1 ;
        RECT 204.235 1716.030 204.405 1716.290 ;
        RECT 201.515 1716.000 202.835 1716.030 ;
        RECT 200.715 1715.830 201.515 1715.990 ;
        RECT 201.685 1715.830 202.835 1716.000 ;
        RECT 200.715 1715.820 202.835 1715.830 ;
        RECT 201.515 1715.700 202.835 1715.820 ;
        RECT 203.435 1716.000 204.405 1716.030 ;
        RECT 203.435 1715.830 204.235 1716.000 ;
        RECT 203.435 1715.700 204.405 1715.830 ;
        RECT 200.325 1715.320 201.345 1715.650 ;
        RECT 201.515 1715.540 201.685 1715.700 ;
        RECT 204.235 1715.540 204.405 1715.700 ;
        RECT 201.515 1715.140 201.685 1715.370 ;
        RECT 204.235 1715.140 204.405 1715.370 ;
        RECT 198.795 1715.080 199.690 1715.140 ;
        RECT 198.965 1714.910 199.690 1715.080 ;
        RECT 198.795 1714.850 199.690 1714.910 ;
        RECT 200.350 1715.080 202.850 1715.140 ;
        RECT 200.350 1714.910 201.515 1715.080 ;
        RECT 201.685 1714.910 202.850 1715.080 ;
        RECT 200.350 1714.850 202.850 1714.910 ;
        RECT 198.795 1714.620 198.965 1714.850 ;
        RECT 201.515 1714.620 201.685 1714.850 ;
        RECT 198.795 1714.290 198.965 1714.450 ;
        RECT 201.515 1714.290 201.685 1714.450 ;
        RECT 201.855 1714.340 202.875 1714.670 ;
        RECT 198.795 1714.160 199.765 1714.290 ;
        RECT 198.965 1713.990 199.765 1714.160 ;
        RECT 198.795 1713.960 199.765 1713.990 ;
        RECT 200.365 1714.170 201.685 1714.290 ;
        RECT 200.365 1714.160 202.485 1714.170 ;
        RECT 200.365 1713.990 201.515 1714.160 ;
        RECT 201.685 1714.000 202.485 1714.160 ;
        RECT 200.365 1713.960 201.685 1713.990 ;
        RECT 198.795 1713.700 198.965 1713.960 ;
      LAYER li1 ;
        RECT 199.135 1713.620 201.345 1713.790 ;
      LAYER li1 ;
        RECT 201.515 1713.700 201.685 1713.960 ;
        RECT 202.705 1713.830 202.875 1714.340 ;
      LAYER li1 ;
        RECT 199.615 1713.535 200.495 1713.620 ;
      LAYER li1 ;
        RECT 198.795 1713.450 198.965 1713.530 ;
        RECT 198.795 1713.240 199.445 1713.450 ;
        RECT 198.965 1713.120 199.445 1713.240 ;
        RECT 198.795 1712.780 198.965 1713.070 ;
      LAYER li1 ;
        RECT 199.615 1712.950 199.785 1713.535 ;
        RECT 199.135 1712.780 199.785 1712.950 ;
      LAYER li1 ;
        RECT 198.795 1712.320 199.445 1712.610 ;
        RECT 198.965 1712.280 199.445 1712.320 ;
        RECT 198.795 1711.860 198.965 1712.150 ;
      LAYER li1 ;
        RECT 199.615 1712.110 199.785 1712.780 ;
        RECT 199.135 1711.940 199.785 1712.110 ;
      LAYER li1 ;
        RECT 198.965 1711.690 199.445 1711.770 ;
        RECT 198.795 1711.440 199.445 1711.690 ;
        RECT 198.795 1711.400 198.965 1711.440 ;
      LAYER li1 ;
        RECT 199.615 1711.270 199.785 1711.940 ;
      LAYER li1 ;
        RECT 198.795 1710.940 198.965 1711.230 ;
      LAYER li1 ;
        RECT 199.135 1711.100 199.785 1711.270 ;
      LAYER li1 ;
        RECT 198.965 1710.770 199.445 1710.930 ;
        RECT 199.955 1710.840 200.125 1713.290 ;
      LAYER li1 ;
        RECT 200.325 1712.950 200.495 1713.535 ;
      LAYER li1 ;
        RECT 201.515 1713.450 201.685 1713.530 ;
        RECT 201.855 1713.500 202.875 1713.830 ;
      LAYER li1 ;
        RECT 203.045 1713.525 203.245 1715.115 ;
      LAYER li1 ;
        RECT 203.510 1715.080 204.405 1715.140 ;
        RECT 203.510 1714.910 204.235 1715.080 ;
        RECT 203.510 1714.850 204.405 1714.910 ;
        RECT 204.235 1714.620 204.405 1714.850 ;
        RECT 203.415 1714.420 204.065 1714.590 ;
        RECT 203.415 1713.750 203.585 1714.420 ;
        RECT 204.235 1714.250 204.405 1714.450 ;
        RECT 203.755 1714.160 204.405 1714.250 ;
        RECT 203.755 1713.990 204.235 1714.160 ;
        RECT 203.755 1713.920 204.405 1713.990 ;
        RECT 203.415 1713.580 204.060 1713.750 ;
        RECT 204.235 1713.700 204.405 1713.920 ;
        RECT 200.715 1713.330 201.685 1713.450 ;
        RECT 202.705 1713.345 202.875 1713.500 ;
        RECT 203.415 1713.345 203.585 1713.580 ;
        RECT 204.235 1713.410 204.405 1713.530 ;
        RECT 200.715 1713.240 202.485 1713.330 ;
        RECT 200.715 1713.120 201.515 1713.240 ;
        RECT 201.685 1713.160 202.485 1713.240 ;
        RECT 202.705 1713.170 203.585 1713.345 ;
        RECT 203.755 1713.240 204.405 1713.410 ;
      LAYER li1 ;
        RECT 200.325 1712.780 201.345 1712.950 ;
      LAYER li1 ;
        RECT 201.515 1712.780 201.685 1713.070 ;
      LAYER li1 ;
        RECT 200.325 1712.110 200.495 1712.780 ;
        RECT 201.855 1712.740 202.875 1712.910 ;
      LAYER li1 ;
        RECT 200.715 1712.570 201.685 1712.610 ;
        RECT 200.715 1712.320 202.485 1712.570 ;
        RECT 200.715 1712.280 201.515 1712.320 ;
        RECT 201.685 1712.240 202.485 1712.320 ;
      LAYER li1 ;
        RECT 200.325 1711.940 201.345 1712.110 ;
        RECT 200.325 1711.270 200.495 1711.940 ;
      LAYER li1 ;
        RECT 201.515 1711.860 201.685 1712.150 ;
      LAYER li1 ;
        RECT 202.705 1712.070 202.875 1712.740 ;
        RECT 201.855 1711.900 202.875 1712.070 ;
      LAYER li1 ;
        RECT 200.715 1711.690 201.515 1711.770 ;
        RECT 201.685 1711.690 202.485 1711.730 ;
        RECT 200.715 1711.440 202.485 1711.690 ;
        RECT 201.515 1711.400 202.485 1711.440 ;
      LAYER li1 ;
        RECT 200.325 1711.100 201.345 1711.270 ;
        RECT 202.705 1711.230 202.875 1711.900 ;
      LAYER li1 ;
        RECT 201.515 1710.940 201.685 1711.230 ;
      LAYER li1 ;
        RECT 201.855 1711.060 202.875 1711.230 ;
      LAYER li1 ;
        RECT 198.795 1710.600 199.445 1710.770 ;
        RECT 199.615 1710.665 200.495 1710.840 ;
        RECT 200.715 1710.770 201.515 1710.850 ;
        RECT 201.685 1710.770 202.485 1710.890 ;
        RECT 200.715 1710.680 202.485 1710.770 ;
        RECT 198.795 1710.480 198.965 1710.600 ;
        RECT 199.615 1710.430 199.785 1710.665 ;
        RECT 200.325 1710.510 200.495 1710.665 ;
        RECT 201.515 1710.560 202.485 1710.680 ;
        RECT 198.795 1710.090 198.965 1710.310 ;
        RECT 199.140 1710.260 199.785 1710.430 ;
        RECT 198.795 1710.020 199.445 1710.090 ;
        RECT 198.965 1709.850 199.445 1710.020 ;
        RECT 198.795 1709.760 199.445 1709.850 ;
        RECT 198.795 1709.560 198.965 1709.760 ;
        RECT 199.615 1709.590 199.785 1710.260 ;
        RECT 199.135 1709.420 199.785 1709.590 ;
        RECT 198.795 1709.160 198.965 1709.390 ;
      LAYER li1 ;
        RECT 199.955 1709.385 200.155 1710.485 ;
      LAYER li1 ;
        RECT 200.325 1710.180 201.345 1710.510 ;
        RECT 201.515 1710.480 201.685 1710.560 ;
      LAYER li1 ;
        RECT 202.705 1710.475 202.875 1711.060 ;
      LAYER li1 ;
        RECT 203.075 1710.720 203.245 1713.170 ;
        RECT 203.755 1713.080 204.235 1713.240 ;
      LAYER li1 ;
        RECT 203.415 1712.740 204.065 1712.910 ;
      LAYER li1 ;
        RECT 204.235 1712.780 204.405 1713.070 ;
      LAYER li1 ;
        RECT 203.415 1712.070 203.585 1712.740 ;
      LAYER li1 ;
        RECT 204.235 1712.570 204.405 1712.610 ;
        RECT 203.755 1712.320 204.405 1712.570 ;
        RECT 203.755 1712.240 204.235 1712.320 ;
      LAYER li1 ;
        RECT 203.415 1711.900 204.065 1712.070 ;
        RECT 203.415 1711.230 203.585 1711.900 ;
      LAYER li1 ;
        RECT 204.235 1711.860 204.405 1712.150 ;
        RECT 203.755 1711.690 204.235 1711.730 ;
        RECT 203.755 1711.400 204.405 1711.690 ;
      LAYER li1 ;
        RECT 203.415 1711.060 204.065 1711.230 ;
        RECT 203.415 1710.475 203.585 1711.060 ;
      LAYER li1 ;
        RECT 204.235 1710.940 204.405 1711.230 ;
        RECT 203.755 1710.770 204.235 1710.890 ;
        RECT 203.755 1710.560 204.405 1710.770 ;
        RECT 204.235 1710.480 204.405 1710.560 ;
      LAYER li1 ;
        RECT 202.705 1710.390 203.585 1710.475 ;
      LAYER li1 ;
        RECT 200.325 1709.670 200.495 1710.180 ;
        RECT 201.515 1710.050 201.685 1710.310 ;
      LAYER li1 ;
        RECT 201.855 1710.220 204.065 1710.390 ;
      LAYER li1 ;
        RECT 204.235 1710.050 204.405 1710.310 ;
        RECT 201.515 1710.020 202.835 1710.050 ;
        RECT 200.715 1709.850 201.515 1710.010 ;
        RECT 201.685 1709.850 202.835 1710.020 ;
        RECT 200.715 1709.840 202.835 1709.850 ;
        RECT 201.515 1709.720 202.835 1709.840 ;
        RECT 203.435 1710.020 204.405 1710.050 ;
        RECT 203.435 1709.850 204.235 1710.020 ;
        RECT 203.435 1709.720 204.405 1709.850 ;
        RECT 200.325 1709.340 201.345 1709.670 ;
        RECT 201.515 1709.560 201.685 1709.720 ;
        RECT 204.235 1709.560 204.405 1709.720 ;
        RECT 201.515 1709.160 201.685 1709.390 ;
        RECT 204.235 1709.160 204.405 1709.390 ;
        RECT 198.795 1709.100 199.690 1709.160 ;
        RECT 198.965 1708.930 199.690 1709.100 ;
        RECT 198.795 1708.870 199.690 1708.930 ;
        RECT 200.350 1709.100 202.850 1709.160 ;
        RECT 200.350 1708.930 201.515 1709.100 ;
        RECT 201.685 1708.930 202.850 1709.100 ;
        RECT 200.350 1708.870 202.850 1708.930 ;
        RECT 198.795 1708.640 198.965 1708.870 ;
        RECT 201.515 1708.640 201.685 1708.870 ;
        RECT 198.795 1708.310 198.965 1708.470 ;
        RECT 201.515 1708.310 201.685 1708.470 ;
        RECT 201.855 1708.360 202.875 1708.690 ;
        RECT 198.795 1708.180 199.765 1708.310 ;
        RECT 198.965 1708.010 199.765 1708.180 ;
        RECT 198.795 1707.980 199.765 1708.010 ;
        RECT 200.365 1708.190 201.685 1708.310 ;
        RECT 200.365 1708.180 202.485 1708.190 ;
        RECT 200.365 1708.010 201.515 1708.180 ;
        RECT 201.685 1708.020 202.485 1708.180 ;
        RECT 200.365 1707.980 201.685 1708.010 ;
        RECT 198.795 1707.720 198.965 1707.980 ;
      LAYER li1 ;
        RECT 199.135 1707.640 201.345 1707.810 ;
      LAYER li1 ;
        RECT 201.515 1707.720 201.685 1707.980 ;
        RECT 202.705 1707.850 202.875 1708.360 ;
      LAYER li1 ;
        RECT 199.615 1707.555 200.495 1707.640 ;
      LAYER li1 ;
        RECT 198.795 1707.470 198.965 1707.550 ;
        RECT 198.795 1707.260 199.445 1707.470 ;
        RECT 198.965 1707.140 199.445 1707.260 ;
        RECT 198.795 1706.800 198.965 1707.090 ;
      LAYER li1 ;
        RECT 199.615 1706.970 199.785 1707.555 ;
        RECT 199.135 1706.800 199.785 1706.970 ;
      LAYER li1 ;
        RECT 198.795 1706.340 199.445 1706.630 ;
        RECT 198.965 1706.300 199.445 1706.340 ;
        RECT 198.795 1705.880 198.965 1706.170 ;
      LAYER li1 ;
        RECT 199.615 1706.130 199.785 1706.800 ;
        RECT 199.135 1705.960 199.785 1706.130 ;
      LAYER li1 ;
        RECT 198.965 1705.710 199.445 1705.790 ;
        RECT 198.795 1705.460 199.445 1705.710 ;
        RECT 198.795 1705.420 198.965 1705.460 ;
      LAYER li1 ;
        RECT 199.615 1705.290 199.785 1705.960 ;
      LAYER li1 ;
        RECT 198.795 1704.960 198.965 1705.250 ;
      LAYER li1 ;
        RECT 199.135 1705.120 199.785 1705.290 ;
      LAYER li1 ;
        RECT 198.965 1704.790 199.445 1704.950 ;
        RECT 199.955 1704.860 200.125 1707.310 ;
      LAYER li1 ;
        RECT 200.325 1706.970 200.495 1707.555 ;
      LAYER li1 ;
        RECT 201.515 1707.470 201.685 1707.550 ;
        RECT 201.855 1707.520 202.875 1707.850 ;
      LAYER li1 ;
        RECT 203.045 1707.545 203.245 1709.135 ;
      LAYER li1 ;
        RECT 203.510 1709.100 204.405 1709.160 ;
        RECT 203.510 1708.930 204.235 1709.100 ;
        RECT 203.510 1708.870 204.405 1708.930 ;
        RECT 204.235 1708.640 204.405 1708.870 ;
        RECT 203.415 1708.440 204.065 1708.610 ;
        RECT 203.415 1707.770 203.585 1708.440 ;
        RECT 204.235 1708.270 204.405 1708.470 ;
        RECT 203.755 1708.180 204.405 1708.270 ;
        RECT 203.755 1708.010 204.235 1708.180 ;
        RECT 203.755 1707.940 204.405 1708.010 ;
        RECT 203.415 1707.600 204.060 1707.770 ;
        RECT 204.235 1707.720 204.405 1707.940 ;
        RECT 200.715 1707.350 201.685 1707.470 ;
        RECT 202.705 1707.365 202.875 1707.520 ;
        RECT 203.415 1707.365 203.585 1707.600 ;
        RECT 204.235 1707.430 204.405 1707.550 ;
        RECT 200.715 1707.260 202.485 1707.350 ;
        RECT 200.715 1707.140 201.515 1707.260 ;
        RECT 201.685 1707.180 202.485 1707.260 ;
        RECT 202.705 1707.190 203.585 1707.365 ;
        RECT 203.755 1707.260 204.405 1707.430 ;
      LAYER li1 ;
        RECT 200.325 1706.800 201.345 1706.970 ;
      LAYER li1 ;
        RECT 201.515 1706.800 201.685 1707.090 ;
      LAYER li1 ;
        RECT 200.325 1706.130 200.495 1706.800 ;
        RECT 201.855 1706.760 202.875 1706.930 ;
      LAYER li1 ;
        RECT 200.715 1706.590 201.685 1706.630 ;
        RECT 200.715 1706.340 202.485 1706.590 ;
        RECT 200.715 1706.300 201.515 1706.340 ;
        RECT 201.685 1706.260 202.485 1706.340 ;
      LAYER li1 ;
        RECT 200.325 1705.960 201.345 1706.130 ;
        RECT 200.325 1705.290 200.495 1705.960 ;
      LAYER li1 ;
        RECT 201.515 1705.880 201.685 1706.170 ;
      LAYER li1 ;
        RECT 202.705 1706.090 202.875 1706.760 ;
        RECT 201.855 1705.920 202.875 1706.090 ;
      LAYER li1 ;
        RECT 200.715 1705.710 201.515 1705.790 ;
        RECT 201.685 1705.710 202.485 1705.750 ;
        RECT 200.715 1705.460 202.485 1705.710 ;
        RECT 201.515 1705.420 202.485 1705.460 ;
      LAYER li1 ;
        RECT 200.325 1705.120 201.345 1705.290 ;
        RECT 202.705 1705.250 202.875 1705.920 ;
      LAYER li1 ;
        RECT 201.515 1704.960 201.685 1705.250 ;
      LAYER li1 ;
        RECT 201.855 1705.080 202.875 1705.250 ;
      LAYER li1 ;
        RECT 198.795 1704.620 199.445 1704.790 ;
        RECT 199.615 1704.685 200.495 1704.860 ;
        RECT 200.715 1704.790 201.515 1704.870 ;
        RECT 201.685 1704.790 202.485 1704.910 ;
        RECT 200.715 1704.700 202.485 1704.790 ;
        RECT 198.795 1704.500 198.965 1704.620 ;
        RECT 199.615 1704.450 199.785 1704.685 ;
        RECT 200.325 1704.530 200.495 1704.685 ;
        RECT 201.515 1704.580 202.485 1704.700 ;
        RECT 198.795 1704.110 198.965 1704.330 ;
        RECT 199.140 1704.280 199.785 1704.450 ;
        RECT 198.795 1704.040 199.445 1704.110 ;
        RECT 198.965 1703.870 199.445 1704.040 ;
        RECT 198.795 1703.780 199.445 1703.870 ;
        RECT 198.795 1703.580 198.965 1703.780 ;
        RECT 199.615 1703.610 199.785 1704.280 ;
        RECT 199.135 1703.440 199.785 1703.610 ;
        RECT 198.795 1703.180 198.965 1703.410 ;
      LAYER li1 ;
        RECT 199.955 1703.405 200.155 1704.505 ;
      LAYER li1 ;
        RECT 200.325 1704.200 201.345 1704.530 ;
        RECT 201.515 1704.500 201.685 1704.580 ;
      LAYER li1 ;
        RECT 202.705 1704.495 202.875 1705.080 ;
      LAYER li1 ;
        RECT 203.075 1704.740 203.245 1707.190 ;
        RECT 203.755 1707.100 204.235 1707.260 ;
      LAYER li1 ;
        RECT 203.415 1706.760 204.065 1706.930 ;
      LAYER li1 ;
        RECT 204.235 1706.800 204.405 1707.090 ;
      LAYER li1 ;
        RECT 203.415 1706.090 203.585 1706.760 ;
      LAYER li1 ;
        RECT 204.235 1706.590 204.405 1706.630 ;
        RECT 203.755 1706.340 204.405 1706.590 ;
        RECT 203.755 1706.260 204.235 1706.340 ;
      LAYER li1 ;
        RECT 203.415 1705.920 204.065 1706.090 ;
        RECT 203.415 1705.250 203.585 1705.920 ;
      LAYER li1 ;
        RECT 204.235 1705.880 204.405 1706.170 ;
        RECT 203.755 1705.710 204.235 1705.750 ;
        RECT 203.755 1705.420 204.405 1705.710 ;
      LAYER li1 ;
        RECT 203.415 1705.080 204.065 1705.250 ;
        RECT 203.415 1704.495 203.585 1705.080 ;
      LAYER li1 ;
        RECT 204.235 1704.960 204.405 1705.250 ;
        RECT 203.755 1704.790 204.235 1704.910 ;
        RECT 203.755 1704.580 204.405 1704.790 ;
        RECT 204.235 1704.500 204.405 1704.580 ;
      LAYER li1 ;
        RECT 202.705 1704.410 203.585 1704.495 ;
      LAYER li1 ;
        RECT 200.325 1703.690 200.495 1704.200 ;
        RECT 201.515 1704.070 201.685 1704.330 ;
      LAYER li1 ;
        RECT 201.855 1704.240 204.065 1704.410 ;
      LAYER li1 ;
        RECT 204.235 1704.070 204.405 1704.330 ;
        RECT 201.515 1704.040 202.835 1704.070 ;
        RECT 200.715 1703.870 201.515 1704.030 ;
        RECT 201.685 1703.870 202.835 1704.040 ;
        RECT 200.715 1703.860 202.835 1703.870 ;
        RECT 201.515 1703.740 202.835 1703.860 ;
        RECT 203.435 1704.040 204.405 1704.070 ;
        RECT 203.435 1703.870 204.235 1704.040 ;
        RECT 203.435 1703.740 204.405 1703.870 ;
        RECT 200.325 1703.360 201.345 1703.690 ;
        RECT 201.515 1703.580 201.685 1703.740 ;
        RECT 204.235 1703.580 204.405 1703.740 ;
        RECT 201.515 1703.180 201.685 1703.410 ;
        RECT 204.235 1703.180 204.405 1703.410 ;
        RECT 198.795 1703.120 199.690 1703.180 ;
        RECT 198.965 1702.950 199.690 1703.120 ;
        RECT 198.795 1702.890 199.690 1702.950 ;
        RECT 200.350 1703.120 202.850 1703.180 ;
        RECT 200.350 1702.950 201.515 1703.120 ;
        RECT 201.685 1702.950 202.850 1703.120 ;
        RECT 200.350 1702.890 202.850 1702.950 ;
        RECT 198.795 1702.660 198.965 1702.890 ;
        RECT 201.515 1702.660 201.685 1702.890 ;
        RECT 198.795 1702.330 198.965 1702.490 ;
        RECT 201.515 1702.330 201.685 1702.490 ;
        RECT 201.855 1702.380 202.875 1702.710 ;
        RECT 198.795 1702.200 199.765 1702.330 ;
        RECT 198.965 1702.030 199.765 1702.200 ;
        RECT 198.795 1702.000 199.765 1702.030 ;
        RECT 200.365 1702.210 201.685 1702.330 ;
        RECT 200.365 1702.200 202.485 1702.210 ;
        RECT 200.365 1702.030 201.515 1702.200 ;
        RECT 201.685 1702.040 202.485 1702.200 ;
        RECT 200.365 1702.000 201.685 1702.030 ;
        RECT 198.795 1701.740 198.965 1702.000 ;
      LAYER li1 ;
        RECT 199.135 1701.660 201.345 1701.830 ;
      LAYER li1 ;
        RECT 201.515 1701.740 201.685 1702.000 ;
        RECT 202.705 1701.870 202.875 1702.380 ;
      LAYER li1 ;
        RECT 199.615 1701.575 200.495 1701.660 ;
      LAYER li1 ;
        RECT 198.795 1701.490 198.965 1701.570 ;
        RECT 198.795 1701.280 199.445 1701.490 ;
        RECT 198.965 1701.160 199.445 1701.280 ;
        RECT 198.795 1700.820 198.965 1701.110 ;
      LAYER li1 ;
        RECT 199.615 1700.990 199.785 1701.575 ;
        RECT 199.135 1700.820 199.785 1700.990 ;
      LAYER li1 ;
        RECT 198.795 1700.360 199.445 1700.650 ;
        RECT 198.965 1700.320 199.445 1700.360 ;
        RECT 198.795 1699.900 198.965 1700.190 ;
      LAYER li1 ;
        RECT 199.615 1700.150 199.785 1700.820 ;
        RECT 199.135 1699.980 199.785 1700.150 ;
      LAYER li1 ;
        RECT 198.965 1699.730 199.445 1699.810 ;
        RECT 198.795 1699.480 199.445 1699.730 ;
        RECT 198.795 1699.440 198.965 1699.480 ;
      LAYER li1 ;
        RECT 199.615 1699.310 199.785 1699.980 ;
      LAYER li1 ;
        RECT 198.795 1698.980 198.965 1699.270 ;
      LAYER li1 ;
        RECT 199.135 1699.140 199.785 1699.310 ;
      LAYER li1 ;
        RECT 198.965 1698.810 199.445 1698.970 ;
        RECT 199.955 1698.880 200.125 1701.330 ;
      LAYER li1 ;
        RECT 200.325 1700.990 200.495 1701.575 ;
      LAYER li1 ;
        RECT 201.515 1701.490 201.685 1701.570 ;
        RECT 201.855 1701.540 202.875 1701.870 ;
      LAYER li1 ;
        RECT 203.045 1701.565 203.245 1703.155 ;
      LAYER li1 ;
        RECT 203.510 1703.120 204.405 1703.180 ;
        RECT 203.510 1702.950 204.235 1703.120 ;
        RECT 203.510 1702.890 204.405 1702.950 ;
        RECT 204.235 1702.660 204.405 1702.890 ;
        RECT 203.415 1702.460 204.065 1702.630 ;
        RECT 203.415 1701.790 203.585 1702.460 ;
        RECT 204.235 1702.290 204.405 1702.490 ;
        RECT 203.755 1702.200 204.405 1702.290 ;
        RECT 203.755 1702.030 204.235 1702.200 ;
        RECT 203.755 1701.960 204.405 1702.030 ;
        RECT 203.415 1701.620 204.060 1701.790 ;
        RECT 204.235 1701.740 204.405 1701.960 ;
        RECT 200.715 1701.370 201.685 1701.490 ;
        RECT 202.705 1701.385 202.875 1701.540 ;
        RECT 203.415 1701.385 203.585 1701.620 ;
        RECT 204.235 1701.450 204.405 1701.570 ;
        RECT 200.715 1701.280 202.485 1701.370 ;
        RECT 200.715 1701.160 201.515 1701.280 ;
        RECT 201.685 1701.200 202.485 1701.280 ;
        RECT 202.705 1701.210 203.585 1701.385 ;
        RECT 203.755 1701.280 204.405 1701.450 ;
      LAYER li1 ;
        RECT 200.325 1700.820 201.345 1700.990 ;
      LAYER li1 ;
        RECT 201.515 1700.820 201.685 1701.110 ;
      LAYER li1 ;
        RECT 200.325 1700.150 200.495 1700.820 ;
        RECT 201.855 1700.780 202.875 1700.950 ;
      LAYER li1 ;
        RECT 200.715 1700.610 201.685 1700.650 ;
        RECT 200.715 1700.360 202.485 1700.610 ;
        RECT 200.715 1700.320 201.515 1700.360 ;
        RECT 201.685 1700.280 202.485 1700.360 ;
      LAYER li1 ;
        RECT 200.325 1699.980 201.345 1700.150 ;
        RECT 200.325 1699.310 200.495 1699.980 ;
      LAYER li1 ;
        RECT 201.515 1699.900 201.685 1700.190 ;
      LAYER li1 ;
        RECT 202.705 1700.110 202.875 1700.780 ;
        RECT 201.855 1699.940 202.875 1700.110 ;
      LAYER li1 ;
        RECT 200.715 1699.730 201.515 1699.810 ;
        RECT 201.685 1699.730 202.485 1699.770 ;
        RECT 200.715 1699.480 202.485 1699.730 ;
        RECT 201.515 1699.440 202.485 1699.480 ;
      LAYER li1 ;
        RECT 200.325 1699.140 201.345 1699.310 ;
        RECT 202.705 1699.270 202.875 1699.940 ;
      LAYER li1 ;
        RECT 201.515 1698.980 201.685 1699.270 ;
      LAYER li1 ;
        RECT 201.855 1699.100 202.875 1699.270 ;
      LAYER li1 ;
        RECT 198.795 1698.640 199.445 1698.810 ;
        RECT 199.615 1698.705 200.495 1698.880 ;
        RECT 200.715 1698.810 201.515 1698.890 ;
        RECT 201.685 1698.810 202.485 1698.930 ;
        RECT 200.715 1698.720 202.485 1698.810 ;
        RECT 198.795 1698.520 198.965 1698.640 ;
        RECT 199.615 1698.470 199.785 1698.705 ;
        RECT 200.325 1698.550 200.495 1698.705 ;
        RECT 201.515 1698.600 202.485 1698.720 ;
        RECT 198.795 1698.130 198.965 1698.350 ;
        RECT 199.140 1698.300 199.785 1698.470 ;
        RECT 198.795 1698.060 199.445 1698.130 ;
        RECT 198.965 1697.890 199.445 1698.060 ;
        RECT 198.795 1697.800 199.445 1697.890 ;
        RECT 198.795 1697.600 198.965 1697.800 ;
        RECT 199.615 1697.630 199.785 1698.300 ;
        RECT 199.135 1697.460 199.785 1697.630 ;
        RECT 198.795 1697.200 198.965 1697.430 ;
      LAYER li1 ;
        RECT 199.955 1697.425 200.155 1698.525 ;
      LAYER li1 ;
        RECT 200.325 1698.220 201.345 1698.550 ;
        RECT 201.515 1698.520 201.685 1698.600 ;
      LAYER li1 ;
        RECT 202.705 1698.515 202.875 1699.100 ;
      LAYER li1 ;
        RECT 203.075 1698.760 203.245 1701.210 ;
        RECT 203.755 1701.120 204.235 1701.280 ;
      LAYER li1 ;
        RECT 203.415 1700.780 204.065 1700.950 ;
      LAYER li1 ;
        RECT 204.235 1700.820 204.405 1701.110 ;
      LAYER li1 ;
        RECT 203.415 1700.110 203.585 1700.780 ;
      LAYER li1 ;
        RECT 204.235 1700.610 204.405 1700.650 ;
        RECT 203.755 1700.360 204.405 1700.610 ;
        RECT 203.755 1700.280 204.235 1700.360 ;
      LAYER li1 ;
        RECT 203.415 1699.940 204.065 1700.110 ;
        RECT 203.415 1699.270 203.585 1699.940 ;
      LAYER li1 ;
        RECT 204.235 1699.900 204.405 1700.190 ;
        RECT 203.755 1699.730 204.235 1699.770 ;
        RECT 203.755 1699.440 204.405 1699.730 ;
      LAYER li1 ;
        RECT 203.415 1699.100 204.065 1699.270 ;
        RECT 203.415 1698.515 203.585 1699.100 ;
      LAYER li1 ;
        RECT 204.235 1698.980 204.405 1699.270 ;
        RECT 203.755 1698.810 204.235 1698.930 ;
        RECT 203.755 1698.600 204.405 1698.810 ;
        RECT 204.235 1698.520 204.405 1698.600 ;
      LAYER li1 ;
        RECT 202.705 1698.430 203.585 1698.515 ;
      LAYER li1 ;
        RECT 200.325 1697.710 200.495 1698.220 ;
        RECT 201.515 1698.090 201.685 1698.350 ;
      LAYER li1 ;
        RECT 201.855 1698.260 204.065 1698.430 ;
      LAYER li1 ;
        RECT 204.235 1698.090 204.405 1698.350 ;
        RECT 201.515 1698.060 202.835 1698.090 ;
        RECT 200.715 1697.890 201.515 1698.050 ;
        RECT 201.685 1697.890 202.835 1698.060 ;
        RECT 200.715 1697.880 202.835 1697.890 ;
        RECT 201.515 1697.760 202.835 1697.880 ;
        RECT 203.435 1698.060 204.405 1698.090 ;
        RECT 203.435 1697.890 204.235 1698.060 ;
        RECT 203.435 1697.760 204.405 1697.890 ;
        RECT 200.325 1697.380 201.345 1697.710 ;
        RECT 201.515 1697.600 201.685 1697.760 ;
        RECT 204.235 1697.600 204.405 1697.760 ;
        RECT 201.515 1697.200 201.685 1697.430 ;
        RECT 204.235 1697.200 204.405 1697.430 ;
        RECT 198.795 1697.140 199.690 1697.200 ;
        RECT 198.965 1696.970 199.690 1697.140 ;
        RECT 198.795 1696.910 199.690 1696.970 ;
        RECT 200.350 1697.140 202.850 1697.200 ;
        RECT 200.350 1696.970 201.515 1697.140 ;
        RECT 201.685 1696.970 202.850 1697.140 ;
        RECT 200.350 1696.910 202.850 1696.970 ;
        RECT 203.510 1697.140 204.405 1697.200 ;
        RECT 203.510 1696.970 204.235 1697.140 ;
        RECT 203.510 1696.910 204.405 1696.970 ;
        RECT 198.795 1696.680 198.965 1696.910 ;
        RECT 201.515 1696.680 201.685 1696.910 ;
        RECT 198.795 1696.350 198.965 1696.510 ;
        RECT 201.515 1696.350 201.685 1696.510 ;
        RECT 201.855 1696.400 202.875 1696.730 ;
        RECT 204.235 1696.680 204.405 1696.910 ;
        RECT 198.795 1696.220 199.765 1696.350 ;
        RECT 198.965 1696.050 199.765 1696.220 ;
        RECT 198.795 1696.020 199.765 1696.050 ;
        RECT 200.365 1696.230 201.685 1696.350 ;
        RECT 200.365 1696.220 202.485 1696.230 ;
        RECT 200.365 1696.050 201.515 1696.220 ;
        RECT 201.685 1696.060 202.485 1696.220 ;
        RECT 200.365 1696.020 201.685 1696.050 ;
        RECT 198.795 1695.760 198.965 1696.020 ;
        RECT 201.515 1695.760 201.685 1696.020 ;
        RECT 202.705 1695.890 202.875 1696.400 ;
        RECT 198.795 1695.510 198.965 1695.590 ;
        RECT 201.515 1695.510 201.685 1695.590 ;
        RECT 201.855 1695.560 202.875 1695.890 ;
        RECT 198.795 1695.300 199.445 1695.510 ;
        RECT 200.715 1695.390 201.685 1695.510 ;
        RECT 202.705 1695.405 202.875 1695.560 ;
        RECT 203.415 1696.480 204.065 1696.650 ;
        RECT 203.415 1695.810 203.585 1696.480 ;
        RECT 204.235 1696.310 204.405 1696.510 ;
        RECT 203.755 1696.220 204.405 1696.310 ;
        RECT 203.755 1696.050 204.235 1696.220 ;
        RECT 203.755 1695.980 204.405 1696.050 ;
        RECT 203.415 1695.640 204.060 1695.810 ;
        RECT 204.235 1695.760 204.405 1695.980 ;
        RECT 203.415 1695.405 203.585 1695.640 ;
        RECT 204.235 1695.470 204.405 1695.590 ;
        RECT 198.965 1695.180 199.445 1695.300 ;
        RECT 198.795 1694.840 198.965 1695.130 ;
        RECT 198.795 1694.380 199.445 1694.670 ;
        RECT 198.965 1694.340 199.445 1694.380 ;
        RECT 198.795 1693.920 198.965 1694.210 ;
        RECT 198.965 1693.750 199.445 1693.830 ;
        RECT 198.795 1693.500 199.445 1693.750 ;
        RECT 198.795 1693.460 198.965 1693.500 ;
        RECT 198.795 1693.000 198.965 1693.290 ;
        RECT 198.965 1692.830 199.445 1692.990 ;
        RECT 199.955 1692.900 200.125 1695.350 ;
        RECT 200.715 1695.300 202.485 1695.390 ;
        RECT 200.715 1695.180 201.515 1695.300 ;
        RECT 201.685 1695.220 202.485 1695.300 ;
        RECT 202.705 1695.230 203.585 1695.405 ;
        RECT 203.755 1695.300 204.405 1695.470 ;
        RECT 201.515 1694.840 201.685 1695.130 ;
      LAYER li1 ;
        RECT 201.855 1694.800 202.875 1694.970 ;
      LAYER li1 ;
        RECT 200.715 1694.630 201.685 1694.670 ;
        RECT 200.715 1694.380 202.485 1694.630 ;
        RECT 200.715 1694.340 201.515 1694.380 ;
        RECT 201.685 1694.300 202.485 1694.380 ;
        RECT 201.515 1693.920 201.685 1694.210 ;
      LAYER li1 ;
        RECT 202.705 1694.130 202.875 1694.800 ;
        RECT 201.855 1693.960 202.875 1694.130 ;
      LAYER li1 ;
        RECT 200.715 1693.750 201.515 1693.830 ;
        RECT 201.685 1693.750 202.485 1693.790 ;
        RECT 200.715 1693.500 202.485 1693.750 ;
        RECT 201.515 1693.460 202.485 1693.500 ;
      LAYER li1 ;
        RECT 202.705 1693.290 202.875 1693.960 ;
      LAYER li1 ;
        RECT 201.515 1693.000 201.685 1693.290 ;
      LAYER li1 ;
        RECT 201.855 1693.120 202.875 1693.290 ;
      LAYER li1 ;
        RECT 198.795 1692.660 199.445 1692.830 ;
        RECT 199.615 1692.725 200.495 1692.900 ;
        RECT 200.715 1692.830 201.515 1692.910 ;
        RECT 201.685 1692.830 202.485 1692.950 ;
        RECT 200.715 1692.740 202.485 1692.830 ;
        RECT 198.795 1692.540 198.965 1692.660 ;
        RECT 199.615 1692.490 199.785 1692.725 ;
        RECT 200.325 1692.570 200.495 1692.725 ;
        RECT 201.515 1692.620 202.485 1692.740 ;
        RECT 198.795 1692.150 198.965 1692.370 ;
        RECT 199.140 1692.320 199.785 1692.490 ;
        RECT 198.795 1692.080 199.445 1692.150 ;
        RECT 198.965 1691.910 199.445 1692.080 ;
        RECT 198.795 1691.820 199.445 1691.910 ;
        RECT 198.795 1691.620 198.965 1691.820 ;
        RECT 199.615 1691.650 199.785 1692.320 ;
        RECT 199.135 1691.480 199.785 1691.650 ;
        RECT 198.795 1691.220 198.965 1691.450 ;
      LAYER li1 ;
        RECT 199.955 1691.445 200.155 1692.545 ;
      LAYER li1 ;
        RECT 200.325 1692.240 201.345 1692.570 ;
        RECT 201.515 1692.540 201.685 1692.620 ;
      LAYER li1 ;
        RECT 202.705 1692.535 202.875 1693.120 ;
      LAYER li1 ;
        RECT 203.075 1692.780 203.245 1695.230 ;
        RECT 203.755 1695.140 204.235 1695.300 ;
      LAYER li1 ;
        RECT 203.415 1694.800 204.065 1694.970 ;
      LAYER li1 ;
        RECT 204.235 1694.840 204.405 1695.130 ;
      LAYER li1 ;
        RECT 203.415 1694.130 203.585 1694.800 ;
      LAYER li1 ;
        RECT 204.235 1694.630 204.405 1694.670 ;
        RECT 203.755 1694.380 204.405 1694.630 ;
        RECT 203.755 1694.300 204.235 1694.380 ;
      LAYER li1 ;
        RECT 203.415 1693.960 204.065 1694.130 ;
        RECT 203.415 1693.290 203.585 1693.960 ;
      LAYER li1 ;
        RECT 204.235 1693.920 204.405 1694.210 ;
        RECT 203.755 1693.750 204.235 1693.790 ;
        RECT 203.755 1693.460 204.405 1693.750 ;
      LAYER li1 ;
        RECT 203.415 1693.120 204.065 1693.290 ;
        RECT 203.415 1692.535 203.585 1693.120 ;
      LAYER li1 ;
        RECT 204.235 1693.000 204.405 1693.290 ;
        RECT 203.755 1692.830 204.235 1692.950 ;
        RECT 203.755 1692.620 204.405 1692.830 ;
        RECT 204.235 1692.540 204.405 1692.620 ;
      LAYER li1 ;
        RECT 202.705 1692.450 203.585 1692.535 ;
      LAYER li1 ;
        RECT 200.325 1691.730 200.495 1692.240 ;
        RECT 201.515 1692.110 201.685 1692.370 ;
      LAYER li1 ;
        RECT 201.855 1692.280 204.065 1692.450 ;
      LAYER li1 ;
        RECT 204.235 1692.110 204.405 1692.370 ;
        RECT 201.515 1692.080 202.835 1692.110 ;
        RECT 200.715 1691.910 201.515 1692.070 ;
        RECT 201.685 1691.910 202.835 1692.080 ;
        RECT 200.715 1691.900 202.835 1691.910 ;
        RECT 201.515 1691.780 202.835 1691.900 ;
        RECT 203.435 1692.080 204.405 1692.110 ;
        RECT 203.435 1691.910 204.235 1692.080 ;
        RECT 203.435 1691.780 204.405 1691.910 ;
        RECT 200.325 1691.400 201.345 1691.730 ;
        RECT 201.515 1691.620 201.685 1691.780 ;
        RECT 204.235 1691.620 204.405 1691.780 ;
        RECT 201.515 1691.220 201.685 1691.450 ;
        RECT 204.235 1691.220 204.405 1691.450 ;
        RECT 198.795 1691.160 199.690 1691.220 ;
        RECT 198.965 1690.990 199.690 1691.160 ;
        RECT 198.795 1690.930 199.690 1690.990 ;
        RECT 200.350 1691.160 202.850 1691.220 ;
        RECT 200.350 1690.990 201.515 1691.160 ;
        RECT 201.685 1690.990 202.850 1691.160 ;
        RECT 200.350 1690.930 202.850 1690.990 ;
        RECT 203.510 1691.160 204.405 1691.220 ;
        RECT 203.510 1690.990 204.235 1691.160 ;
        RECT 203.510 1690.930 204.405 1690.990 ;
        RECT 198.795 1690.700 198.965 1690.930 ;
        RECT 201.515 1690.700 201.685 1690.930 ;
        RECT 198.795 1690.370 198.965 1690.530 ;
        RECT 201.515 1690.370 201.685 1690.530 ;
        RECT 201.855 1690.420 202.875 1690.750 ;
        RECT 204.235 1690.700 204.405 1690.930 ;
        RECT 198.795 1690.240 199.765 1690.370 ;
        RECT 198.965 1690.070 199.765 1690.240 ;
        RECT 198.795 1690.040 199.765 1690.070 ;
        RECT 200.365 1690.250 201.685 1690.370 ;
        RECT 200.365 1690.240 202.485 1690.250 ;
        RECT 200.365 1690.070 201.515 1690.240 ;
        RECT 201.685 1690.080 202.485 1690.240 ;
        RECT 200.365 1690.040 201.685 1690.070 ;
        RECT 198.795 1689.780 198.965 1690.040 ;
        RECT 201.515 1689.780 201.685 1690.040 ;
        RECT 202.705 1689.910 202.875 1690.420 ;
        RECT 198.795 1689.530 198.965 1689.610 ;
        RECT 201.515 1689.530 201.685 1689.610 ;
        RECT 201.855 1689.580 202.875 1689.910 ;
        RECT 198.795 1689.320 199.445 1689.530 ;
        RECT 200.715 1689.410 201.685 1689.530 ;
        RECT 202.705 1689.425 202.875 1689.580 ;
        RECT 203.415 1690.500 204.065 1690.670 ;
        RECT 203.415 1689.830 203.585 1690.500 ;
        RECT 204.235 1690.330 204.405 1690.530 ;
        RECT 203.755 1690.240 204.405 1690.330 ;
        RECT 203.755 1690.070 204.235 1690.240 ;
        RECT 203.755 1690.000 204.405 1690.070 ;
        RECT 203.415 1689.660 204.060 1689.830 ;
        RECT 204.235 1689.780 204.405 1690.000 ;
        RECT 203.415 1689.425 203.585 1689.660 ;
        RECT 204.235 1689.490 204.405 1689.610 ;
        RECT 198.965 1689.200 199.445 1689.320 ;
        RECT 198.795 1688.860 198.965 1689.150 ;
        RECT 198.795 1688.400 199.445 1688.690 ;
        RECT 198.965 1688.360 199.445 1688.400 ;
        RECT 198.795 1687.940 198.965 1688.230 ;
        RECT 198.965 1687.770 199.445 1687.850 ;
        RECT 198.795 1687.520 199.445 1687.770 ;
        RECT 198.795 1687.480 198.965 1687.520 ;
        RECT 198.795 1687.020 198.965 1687.310 ;
        RECT 198.965 1686.850 199.445 1687.010 ;
        RECT 199.955 1686.920 200.125 1689.370 ;
        RECT 200.715 1689.320 202.485 1689.410 ;
        RECT 200.715 1689.200 201.515 1689.320 ;
        RECT 201.685 1689.240 202.485 1689.320 ;
        RECT 202.705 1689.250 203.585 1689.425 ;
        RECT 203.755 1689.320 204.405 1689.490 ;
        RECT 201.515 1688.860 201.685 1689.150 ;
      LAYER li1 ;
        RECT 201.855 1688.820 202.875 1688.990 ;
      LAYER li1 ;
        RECT 200.715 1688.650 201.685 1688.690 ;
        RECT 200.715 1688.400 202.485 1688.650 ;
        RECT 200.715 1688.360 201.515 1688.400 ;
        RECT 201.685 1688.320 202.485 1688.400 ;
        RECT 201.515 1687.940 201.685 1688.230 ;
      LAYER li1 ;
        RECT 202.705 1688.150 202.875 1688.820 ;
        RECT 201.855 1687.980 202.875 1688.150 ;
      LAYER li1 ;
        RECT 200.715 1687.770 201.515 1687.850 ;
        RECT 201.685 1687.770 202.485 1687.810 ;
        RECT 200.715 1687.520 202.485 1687.770 ;
        RECT 201.515 1687.480 202.485 1687.520 ;
      LAYER li1 ;
        RECT 202.705 1687.310 202.875 1687.980 ;
      LAYER li1 ;
        RECT 201.515 1687.020 201.685 1687.310 ;
      LAYER li1 ;
        RECT 201.855 1687.140 202.875 1687.310 ;
      LAYER li1 ;
        RECT 198.795 1686.680 199.445 1686.850 ;
        RECT 199.615 1686.745 200.495 1686.920 ;
        RECT 200.715 1686.850 201.515 1686.930 ;
        RECT 201.685 1686.850 202.485 1686.970 ;
        RECT 200.715 1686.760 202.485 1686.850 ;
        RECT 198.795 1686.560 198.965 1686.680 ;
        RECT 199.615 1686.510 199.785 1686.745 ;
        RECT 200.325 1686.590 200.495 1686.745 ;
        RECT 201.515 1686.640 202.485 1686.760 ;
        RECT 198.795 1686.170 198.965 1686.390 ;
        RECT 199.140 1686.340 199.785 1686.510 ;
        RECT 198.795 1686.100 199.445 1686.170 ;
        RECT 198.965 1685.930 199.445 1686.100 ;
        RECT 198.795 1685.840 199.445 1685.930 ;
        RECT 198.795 1685.640 198.965 1685.840 ;
        RECT 199.615 1685.670 199.785 1686.340 ;
        RECT 199.135 1685.500 199.785 1685.670 ;
        RECT 198.795 1685.240 198.965 1685.470 ;
      LAYER li1 ;
        RECT 199.955 1685.465 200.155 1686.565 ;
      LAYER li1 ;
        RECT 200.325 1686.260 201.345 1686.590 ;
        RECT 201.515 1686.560 201.685 1686.640 ;
      LAYER li1 ;
        RECT 202.705 1686.555 202.875 1687.140 ;
      LAYER li1 ;
        RECT 203.075 1686.800 203.245 1689.250 ;
        RECT 203.755 1689.160 204.235 1689.320 ;
      LAYER li1 ;
        RECT 203.415 1688.820 204.065 1688.990 ;
      LAYER li1 ;
        RECT 204.235 1688.860 204.405 1689.150 ;
      LAYER li1 ;
        RECT 203.415 1688.150 203.585 1688.820 ;
      LAYER li1 ;
        RECT 204.235 1688.650 204.405 1688.690 ;
        RECT 203.755 1688.400 204.405 1688.650 ;
        RECT 203.755 1688.320 204.235 1688.400 ;
      LAYER li1 ;
        RECT 203.415 1687.980 204.065 1688.150 ;
        RECT 203.415 1687.310 203.585 1687.980 ;
      LAYER li1 ;
        RECT 204.235 1687.940 204.405 1688.230 ;
        RECT 203.755 1687.770 204.235 1687.810 ;
        RECT 203.755 1687.480 204.405 1687.770 ;
      LAYER li1 ;
        RECT 203.415 1687.140 204.065 1687.310 ;
        RECT 203.415 1686.555 203.585 1687.140 ;
      LAYER li1 ;
        RECT 204.235 1687.020 204.405 1687.310 ;
        RECT 203.755 1686.850 204.235 1686.970 ;
        RECT 203.755 1686.640 204.405 1686.850 ;
        RECT 204.235 1686.560 204.405 1686.640 ;
      LAYER li1 ;
        RECT 202.705 1686.470 203.585 1686.555 ;
      LAYER li1 ;
        RECT 200.325 1685.750 200.495 1686.260 ;
        RECT 201.515 1686.130 201.685 1686.390 ;
      LAYER li1 ;
        RECT 201.855 1686.300 204.065 1686.470 ;
      LAYER li1 ;
        RECT 204.235 1686.130 204.405 1686.390 ;
        RECT 201.515 1686.100 202.835 1686.130 ;
        RECT 200.715 1685.930 201.515 1686.090 ;
        RECT 201.685 1685.930 202.835 1686.100 ;
        RECT 200.715 1685.920 202.835 1685.930 ;
        RECT 201.515 1685.800 202.835 1685.920 ;
        RECT 203.435 1686.100 204.405 1686.130 ;
        RECT 203.435 1685.930 204.235 1686.100 ;
        RECT 203.435 1685.800 204.405 1685.930 ;
        RECT 200.325 1685.420 201.345 1685.750 ;
        RECT 201.515 1685.640 201.685 1685.800 ;
        RECT 204.235 1685.640 204.405 1685.800 ;
        RECT 201.515 1685.240 201.685 1685.470 ;
        RECT 204.235 1685.240 204.405 1685.470 ;
        RECT 198.795 1685.180 199.690 1685.240 ;
        RECT 198.965 1685.010 199.690 1685.180 ;
        RECT 198.795 1684.950 199.690 1685.010 ;
        RECT 200.350 1685.180 202.850 1685.240 ;
        RECT 200.350 1685.010 201.515 1685.180 ;
        RECT 201.685 1685.010 202.850 1685.180 ;
        RECT 200.350 1684.950 202.850 1685.010 ;
        RECT 203.510 1685.180 204.405 1685.240 ;
        RECT 203.510 1685.010 204.235 1685.180 ;
        RECT 203.510 1684.950 204.405 1685.010 ;
        RECT 198.795 1684.720 198.965 1684.950 ;
        RECT 201.515 1684.720 201.685 1684.950 ;
        RECT 198.795 1684.390 198.965 1684.550 ;
        RECT 201.515 1684.390 201.685 1684.550 ;
        RECT 201.855 1684.440 202.875 1684.770 ;
        RECT 204.235 1684.720 204.405 1684.950 ;
        RECT 198.795 1684.260 199.765 1684.390 ;
        RECT 198.965 1684.090 199.765 1684.260 ;
        RECT 198.795 1684.060 199.765 1684.090 ;
        RECT 200.365 1684.270 201.685 1684.390 ;
        RECT 200.365 1684.260 202.485 1684.270 ;
        RECT 200.365 1684.090 201.515 1684.260 ;
        RECT 201.685 1684.100 202.485 1684.260 ;
        RECT 200.365 1684.060 201.685 1684.090 ;
        RECT 198.795 1683.800 198.965 1684.060 ;
        RECT 201.515 1683.800 201.685 1684.060 ;
        RECT 202.705 1683.930 202.875 1684.440 ;
        RECT 198.795 1683.550 198.965 1683.630 ;
        RECT 201.515 1683.550 201.685 1683.630 ;
        RECT 201.855 1683.600 202.875 1683.930 ;
        RECT 198.795 1683.340 199.445 1683.550 ;
        RECT 200.715 1683.430 201.685 1683.550 ;
        RECT 202.705 1683.445 202.875 1683.600 ;
        RECT 203.415 1684.520 204.065 1684.690 ;
        RECT 203.415 1683.850 203.585 1684.520 ;
        RECT 204.235 1684.350 204.405 1684.550 ;
        RECT 203.755 1684.260 204.405 1684.350 ;
        RECT 203.755 1684.090 204.235 1684.260 ;
        RECT 203.755 1684.020 204.405 1684.090 ;
        RECT 203.415 1683.680 204.060 1683.850 ;
        RECT 204.235 1683.800 204.405 1684.020 ;
        RECT 203.415 1683.445 203.585 1683.680 ;
        RECT 204.235 1683.510 204.405 1683.630 ;
        RECT 198.965 1683.220 199.445 1683.340 ;
        RECT 198.795 1682.880 198.965 1683.170 ;
        RECT 198.795 1682.420 199.445 1682.710 ;
        RECT 198.965 1682.380 199.445 1682.420 ;
        RECT 198.795 1681.960 198.965 1682.250 ;
        RECT 198.965 1681.790 199.445 1681.870 ;
        RECT 198.795 1681.540 199.445 1681.790 ;
        RECT 198.795 1681.500 198.965 1681.540 ;
        RECT 198.795 1681.040 198.965 1681.330 ;
        RECT 198.965 1680.870 199.445 1681.030 ;
        RECT 199.955 1680.940 200.125 1683.390 ;
        RECT 200.715 1683.340 202.485 1683.430 ;
        RECT 200.715 1683.220 201.515 1683.340 ;
        RECT 201.685 1683.260 202.485 1683.340 ;
        RECT 202.705 1683.270 203.585 1683.445 ;
        RECT 203.755 1683.340 204.405 1683.510 ;
        RECT 201.515 1682.880 201.685 1683.170 ;
      LAYER li1 ;
        RECT 201.855 1682.840 202.875 1683.010 ;
      LAYER li1 ;
        RECT 200.715 1682.670 201.685 1682.710 ;
        RECT 200.715 1682.420 202.485 1682.670 ;
        RECT 200.715 1682.380 201.515 1682.420 ;
        RECT 201.685 1682.340 202.485 1682.420 ;
        RECT 201.515 1681.960 201.685 1682.250 ;
      LAYER li1 ;
        RECT 202.705 1682.170 202.875 1682.840 ;
        RECT 201.855 1682.000 202.875 1682.170 ;
      LAYER li1 ;
        RECT 200.715 1681.790 201.515 1681.870 ;
        RECT 201.685 1681.790 202.485 1681.830 ;
        RECT 200.715 1681.540 202.485 1681.790 ;
        RECT 201.515 1681.500 202.485 1681.540 ;
      LAYER li1 ;
        RECT 202.705 1681.330 202.875 1682.000 ;
      LAYER li1 ;
        RECT 201.515 1681.040 201.685 1681.330 ;
      LAYER li1 ;
        RECT 201.855 1681.160 202.875 1681.330 ;
      LAYER li1 ;
        RECT 198.795 1680.700 199.445 1680.870 ;
        RECT 199.615 1680.765 200.495 1680.940 ;
        RECT 200.715 1680.870 201.515 1680.950 ;
        RECT 201.685 1680.870 202.485 1680.990 ;
        RECT 200.715 1680.780 202.485 1680.870 ;
        RECT 198.795 1680.580 198.965 1680.700 ;
        RECT 199.615 1680.530 199.785 1680.765 ;
        RECT 200.325 1680.610 200.495 1680.765 ;
        RECT 201.515 1680.660 202.485 1680.780 ;
        RECT 198.795 1680.190 198.965 1680.410 ;
        RECT 199.140 1680.360 199.785 1680.530 ;
        RECT 198.795 1680.120 199.445 1680.190 ;
        RECT 198.965 1679.950 199.445 1680.120 ;
        RECT 198.795 1679.860 199.445 1679.950 ;
        RECT 198.795 1679.660 198.965 1679.860 ;
        RECT 199.615 1679.690 199.785 1680.360 ;
        RECT 199.135 1679.520 199.785 1679.690 ;
        RECT 198.795 1679.260 198.965 1679.490 ;
      LAYER li1 ;
        RECT 199.955 1679.485 200.155 1680.585 ;
      LAYER li1 ;
        RECT 200.325 1680.280 201.345 1680.610 ;
        RECT 201.515 1680.580 201.685 1680.660 ;
      LAYER li1 ;
        RECT 202.705 1680.575 202.875 1681.160 ;
      LAYER li1 ;
        RECT 203.075 1680.820 203.245 1683.270 ;
        RECT 203.755 1683.180 204.235 1683.340 ;
      LAYER li1 ;
        RECT 203.415 1682.840 204.065 1683.010 ;
      LAYER li1 ;
        RECT 204.235 1682.880 204.405 1683.170 ;
      LAYER li1 ;
        RECT 203.415 1682.170 203.585 1682.840 ;
      LAYER li1 ;
        RECT 204.235 1682.670 204.405 1682.710 ;
        RECT 203.755 1682.420 204.405 1682.670 ;
        RECT 203.755 1682.340 204.235 1682.420 ;
      LAYER li1 ;
        RECT 203.415 1682.000 204.065 1682.170 ;
        RECT 203.415 1681.330 203.585 1682.000 ;
      LAYER li1 ;
        RECT 204.235 1681.960 204.405 1682.250 ;
        RECT 203.755 1681.790 204.235 1681.830 ;
        RECT 203.755 1681.500 204.405 1681.790 ;
      LAYER li1 ;
        RECT 203.415 1681.160 204.065 1681.330 ;
        RECT 203.415 1680.575 203.585 1681.160 ;
      LAYER li1 ;
        RECT 204.235 1681.040 204.405 1681.330 ;
        RECT 203.755 1680.870 204.235 1680.990 ;
        RECT 203.755 1680.660 204.405 1680.870 ;
        RECT 204.235 1680.580 204.405 1680.660 ;
      LAYER li1 ;
        RECT 202.705 1680.490 203.585 1680.575 ;
      LAYER li1 ;
        RECT 200.325 1679.770 200.495 1680.280 ;
        RECT 201.515 1680.150 201.685 1680.410 ;
      LAYER li1 ;
        RECT 201.855 1680.320 204.065 1680.490 ;
      LAYER li1 ;
        RECT 204.235 1680.150 204.405 1680.410 ;
        RECT 201.515 1680.120 202.835 1680.150 ;
        RECT 200.715 1679.950 201.515 1680.110 ;
        RECT 201.685 1679.950 202.835 1680.120 ;
        RECT 200.715 1679.940 202.835 1679.950 ;
        RECT 201.515 1679.820 202.835 1679.940 ;
        RECT 203.435 1680.120 204.405 1680.150 ;
        RECT 203.435 1679.950 204.235 1680.120 ;
        RECT 203.435 1679.820 204.405 1679.950 ;
        RECT 200.325 1679.440 201.345 1679.770 ;
        RECT 201.515 1679.660 201.685 1679.820 ;
        RECT 204.235 1679.660 204.405 1679.820 ;
        RECT 201.515 1679.260 201.685 1679.490 ;
        RECT 204.235 1679.260 204.405 1679.490 ;
        RECT 198.795 1679.200 199.690 1679.260 ;
        RECT 198.965 1679.030 199.690 1679.200 ;
        RECT 198.795 1678.970 199.690 1679.030 ;
        RECT 200.350 1679.200 202.850 1679.260 ;
        RECT 200.350 1679.030 201.515 1679.200 ;
        RECT 201.685 1679.030 202.850 1679.200 ;
        RECT 200.350 1678.970 202.850 1679.030 ;
        RECT 203.510 1679.200 204.405 1679.260 ;
        RECT 203.510 1679.030 204.235 1679.200 ;
        RECT 203.510 1678.970 204.405 1679.030 ;
        RECT 198.795 1678.740 198.965 1678.970 ;
        RECT 201.515 1678.740 201.685 1678.970 ;
        RECT 198.795 1678.410 198.965 1678.570 ;
        RECT 201.515 1678.410 201.685 1678.570 ;
        RECT 201.855 1678.460 202.875 1678.790 ;
        RECT 204.235 1678.740 204.405 1678.970 ;
        RECT 198.795 1678.280 199.765 1678.410 ;
        RECT 198.965 1678.110 199.765 1678.280 ;
        RECT 198.795 1678.080 199.765 1678.110 ;
        RECT 200.365 1678.290 201.685 1678.410 ;
        RECT 200.365 1678.280 202.485 1678.290 ;
        RECT 200.365 1678.110 201.515 1678.280 ;
        RECT 201.685 1678.120 202.485 1678.280 ;
        RECT 200.365 1678.080 201.685 1678.110 ;
        RECT 198.795 1677.820 198.965 1678.080 ;
        RECT 201.515 1677.820 201.685 1678.080 ;
        RECT 202.705 1677.950 202.875 1678.460 ;
        RECT 198.795 1677.570 198.965 1677.650 ;
        RECT 201.515 1677.570 201.685 1677.650 ;
        RECT 201.855 1677.620 202.875 1677.950 ;
        RECT 198.795 1677.360 199.445 1677.570 ;
        RECT 200.715 1677.450 201.685 1677.570 ;
        RECT 202.705 1677.465 202.875 1677.620 ;
        RECT 203.415 1678.540 204.065 1678.710 ;
        RECT 203.415 1677.870 203.585 1678.540 ;
        RECT 204.235 1678.370 204.405 1678.570 ;
        RECT 203.755 1678.280 204.405 1678.370 ;
        RECT 203.755 1678.110 204.235 1678.280 ;
        RECT 203.755 1678.040 204.405 1678.110 ;
        RECT 203.415 1677.700 204.060 1677.870 ;
        RECT 204.235 1677.820 204.405 1678.040 ;
        RECT 203.415 1677.465 203.585 1677.700 ;
        RECT 204.235 1677.530 204.405 1677.650 ;
        RECT 198.965 1677.240 199.445 1677.360 ;
        RECT 198.795 1676.900 198.965 1677.190 ;
        RECT 198.795 1676.440 199.445 1676.730 ;
        RECT 198.965 1676.400 199.445 1676.440 ;
        RECT 198.795 1675.980 198.965 1676.270 ;
        RECT 198.965 1675.810 199.445 1675.890 ;
        RECT 198.795 1675.560 199.445 1675.810 ;
        RECT 198.795 1675.520 198.965 1675.560 ;
        RECT 198.795 1675.060 198.965 1675.350 ;
        RECT 198.965 1674.890 199.445 1675.050 ;
        RECT 199.955 1674.960 200.125 1677.410 ;
        RECT 200.715 1677.360 202.485 1677.450 ;
        RECT 200.715 1677.240 201.515 1677.360 ;
        RECT 201.685 1677.280 202.485 1677.360 ;
        RECT 202.705 1677.290 203.585 1677.465 ;
        RECT 203.755 1677.360 204.405 1677.530 ;
        RECT 201.515 1676.900 201.685 1677.190 ;
      LAYER li1 ;
        RECT 201.855 1676.860 202.875 1677.030 ;
      LAYER li1 ;
        RECT 200.715 1676.690 201.685 1676.730 ;
        RECT 200.715 1676.440 202.485 1676.690 ;
        RECT 200.715 1676.400 201.515 1676.440 ;
        RECT 201.685 1676.360 202.485 1676.440 ;
        RECT 201.515 1675.980 201.685 1676.270 ;
      LAYER li1 ;
        RECT 202.705 1676.190 202.875 1676.860 ;
        RECT 201.855 1676.020 202.875 1676.190 ;
      LAYER li1 ;
        RECT 200.715 1675.810 201.515 1675.890 ;
        RECT 201.685 1675.810 202.485 1675.850 ;
        RECT 200.715 1675.560 202.485 1675.810 ;
        RECT 201.515 1675.520 202.485 1675.560 ;
      LAYER li1 ;
        RECT 202.705 1675.350 202.875 1676.020 ;
      LAYER li1 ;
        RECT 201.515 1675.060 201.685 1675.350 ;
      LAYER li1 ;
        RECT 201.855 1675.180 202.875 1675.350 ;
      LAYER li1 ;
        RECT 198.795 1674.720 199.445 1674.890 ;
        RECT 199.615 1674.785 200.495 1674.960 ;
        RECT 200.715 1674.890 201.515 1674.970 ;
        RECT 201.685 1674.890 202.485 1675.010 ;
        RECT 200.715 1674.800 202.485 1674.890 ;
        RECT 198.795 1674.600 198.965 1674.720 ;
        RECT 199.615 1674.550 199.785 1674.785 ;
        RECT 200.325 1674.630 200.495 1674.785 ;
        RECT 201.515 1674.680 202.485 1674.800 ;
        RECT 198.795 1674.210 198.965 1674.430 ;
        RECT 199.140 1674.380 199.785 1674.550 ;
        RECT 198.795 1674.140 199.445 1674.210 ;
        RECT 198.965 1673.970 199.445 1674.140 ;
        RECT 198.795 1673.880 199.445 1673.970 ;
        RECT 198.795 1673.680 198.965 1673.880 ;
        RECT 199.615 1673.710 199.785 1674.380 ;
        RECT 199.135 1673.540 199.785 1673.710 ;
        RECT 198.795 1673.280 198.965 1673.510 ;
      LAYER li1 ;
        RECT 199.955 1673.505 200.155 1674.605 ;
      LAYER li1 ;
        RECT 200.325 1674.300 201.345 1674.630 ;
        RECT 201.515 1674.600 201.685 1674.680 ;
      LAYER li1 ;
        RECT 202.705 1674.595 202.875 1675.180 ;
      LAYER li1 ;
        RECT 203.075 1674.840 203.245 1677.290 ;
        RECT 203.755 1677.200 204.235 1677.360 ;
      LAYER li1 ;
        RECT 203.415 1676.860 204.065 1677.030 ;
      LAYER li1 ;
        RECT 204.235 1676.900 204.405 1677.190 ;
      LAYER li1 ;
        RECT 203.415 1676.190 203.585 1676.860 ;
      LAYER li1 ;
        RECT 204.235 1676.690 204.405 1676.730 ;
        RECT 203.755 1676.440 204.405 1676.690 ;
        RECT 203.755 1676.360 204.235 1676.440 ;
      LAYER li1 ;
        RECT 203.415 1676.020 204.065 1676.190 ;
        RECT 203.415 1675.350 203.585 1676.020 ;
      LAYER li1 ;
        RECT 204.235 1675.980 204.405 1676.270 ;
        RECT 203.755 1675.810 204.235 1675.850 ;
        RECT 203.755 1675.520 204.405 1675.810 ;
      LAYER li1 ;
        RECT 203.415 1675.180 204.065 1675.350 ;
        RECT 203.415 1674.595 203.585 1675.180 ;
      LAYER li1 ;
        RECT 204.235 1675.060 204.405 1675.350 ;
        RECT 203.755 1674.890 204.235 1675.010 ;
        RECT 203.755 1674.680 204.405 1674.890 ;
        RECT 204.235 1674.600 204.405 1674.680 ;
      LAYER li1 ;
        RECT 202.705 1674.510 203.585 1674.595 ;
      LAYER li1 ;
        RECT 200.325 1673.790 200.495 1674.300 ;
        RECT 201.515 1674.170 201.685 1674.430 ;
      LAYER li1 ;
        RECT 201.855 1674.340 204.065 1674.510 ;
      LAYER li1 ;
        RECT 204.235 1674.170 204.405 1674.430 ;
        RECT 201.515 1674.140 202.835 1674.170 ;
        RECT 200.715 1673.970 201.515 1674.130 ;
        RECT 201.685 1673.970 202.835 1674.140 ;
        RECT 200.715 1673.960 202.835 1673.970 ;
        RECT 201.515 1673.840 202.835 1673.960 ;
        RECT 203.435 1674.140 204.405 1674.170 ;
        RECT 203.435 1673.970 204.235 1674.140 ;
        RECT 203.435 1673.840 204.405 1673.970 ;
        RECT 200.325 1673.460 201.345 1673.790 ;
        RECT 201.515 1673.680 201.685 1673.840 ;
        RECT 204.235 1673.680 204.405 1673.840 ;
        RECT 201.515 1673.280 201.685 1673.510 ;
        RECT 204.235 1673.280 204.405 1673.510 ;
        RECT 198.795 1673.220 199.690 1673.280 ;
        RECT 198.965 1673.050 199.690 1673.220 ;
        RECT 198.795 1672.990 199.690 1673.050 ;
        RECT 200.350 1673.220 202.850 1673.280 ;
        RECT 200.350 1673.050 201.515 1673.220 ;
        RECT 201.685 1673.050 202.850 1673.220 ;
        RECT 200.350 1672.990 202.850 1673.050 ;
        RECT 203.510 1673.220 204.405 1673.280 ;
        RECT 203.510 1673.050 204.235 1673.220 ;
        RECT 203.510 1672.990 204.405 1673.050 ;
        RECT 198.795 1672.905 198.965 1672.990 ;
        RECT 201.515 1672.905 201.685 1672.990 ;
        RECT 204.235 1672.905 204.405 1672.990 ;
        RECT 669.000 1117.040 669.145 1117.210 ;
        RECT 669.315 1117.040 669.605 1117.210 ;
        RECT 669.775 1117.040 670.065 1117.210 ;
        RECT 670.235 1117.040 670.525 1117.210 ;
        RECT 670.695 1117.040 670.985 1117.210 ;
        RECT 671.155 1117.040 671.445 1117.210 ;
        RECT 671.615 1117.040 671.905 1117.210 ;
        RECT 672.075 1117.040 672.365 1117.210 ;
        RECT 672.535 1117.040 672.825 1117.210 ;
        RECT 672.995 1117.040 673.285 1117.210 ;
        RECT 673.455 1117.040 673.745 1117.210 ;
        RECT 673.915 1117.040 674.205 1117.210 ;
        RECT 674.375 1117.040 674.665 1117.210 ;
        RECT 674.835 1117.040 675.125 1117.210 ;
        RECT 675.295 1117.040 675.585 1117.210 ;
        RECT 675.755 1117.040 676.045 1117.210 ;
        RECT 676.215 1117.040 676.505 1117.210 ;
        RECT 676.675 1117.040 676.965 1117.210 ;
        RECT 677.135 1117.040 677.425 1117.210 ;
        RECT 677.595 1117.040 677.885 1117.210 ;
        RECT 678.055 1117.040 678.345 1117.210 ;
        RECT 678.515 1117.040 678.805 1117.210 ;
        RECT 678.975 1117.040 679.265 1117.210 ;
        RECT 679.435 1117.040 679.725 1117.210 ;
        RECT 679.895 1117.040 680.185 1117.210 ;
        RECT 680.355 1117.040 680.645 1117.210 ;
        RECT 680.815 1117.040 681.105 1117.210 ;
        RECT 681.275 1117.040 681.565 1117.210 ;
        RECT 681.735 1117.040 682.025 1117.210 ;
        RECT 682.195 1117.040 682.485 1117.210 ;
        RECT 682.655 1117.040 682.945 1117.210 ;
        RECT 683.115 1117.040 683.405 1117.210 ;
        RECT 683.575 1117.040 683.865 1117.210 ;
        RECT 684.035 1117.040 684.325 1117.210 ;
        RECT 684.495 1117.040 684.785 1117.210 ;
        RECT 684.955 1117.040 685.245 1117.210 ;
        RECT 685.415 1117.040 685.705 1117.210 ;
        RECT 685.875 1117.040 686.165 1117.210 ;
        RECT 686.335 1117.040 686.625 1117.210 ;
        RECT 686.795 1117.040 687.085 1117.210 ;
        RECT 687.255 1117.040 687.545 1117.210 ;
        RECT 687.715 1117.040 688.005 1117.210 ;
        RECT 688.175 1117.040 688.465 1117.210 ;
        RECT 688.635 1117.040 688.925 1117.210 ;
        RECT 689.095 1117.040 689.385 1117.210 ;
        RECT 689.555 1117.040 689.845 1117.210 ;
        RECT 690.015 1117.040 690.305 1117.210 ;
        RECT 690.475 1117.040 690.765 1117.210 ;
        RECT 690.935 1117.040 691.225 1117.210 ;
        RECT 691.395 1117.040 691.685 1117.210 ;
        RECT 691.855 1117.040 692.145 1117.210 ;
        RECT 692.315 1117.040 692.605 1117.210 ;
        RECT 692.775 1117.040 693.065 1117.210 ;
        RECT 693.235 1117.040 693.525 1117.210 ;
        RECT 693.695 1117.040 693.985 1117.210 ;
        RECT 694.155 1117.040 694.445 1117.210 ;
        RECT 694.615 1117.040 694.905 1117.210 ;
        RECT 695.075 1117.040 695.365 1117.210 ;
        RECT 695.535 1117.040 695.825 1117.210 ;
        RECT 695.995 1117.040 696.285 1117.210 ;
        RECT 696.455 1117.040 696.745 1117.210 ;
        RECT 696.915 1117.040 697.205 1117.210 ;
        RECT 697.375 1117.040 697.665 1117.210 ;
        RECT 697.835 1117.040 698.125 1117.210 ;
        RECT 698.295 1117.040 698.585 1117.210 ;
        RECT 698.755 1117.040 699.045 1117.210 ;
        RECT 699.215 1117.040 699.505 1117.210 ;
        RECT 699.675 1117.040 699.965 1117.210 ;
        RECT 700.135 1117.040 700.425 1117.210 ;
        RECT 700.595 1117.040 700.885 1117.210 ;
        RECT 701.055 1117.040 701.345 1117.210 ;
        RECT 701.515 1117.040 701.805 1117.210 ;
        RECT 701.975 1117.040 702.265 1117.210 ;
        RECT 702.435 1117.040 702.725 1117.210 ;
        RECT 702.895 1117.040 703.185 1117.210 ;
        RECT 703.355 1117.040 703.645 1117.210 ;
        RECT 703.815 1117.040 704.105 1117.210 ;
        RECT 704.275 1117.040 704.565 1117.210 ;
        RECT 704.735 1117.040 705.025 1117.210 ;
        RECT 705.195 1117.040 705.485 1117.210 ;
        RECT 705.655 1117.040 705.945 1117.210 ;
        RECT 706.115 1117.040 706.405 1117.210 ;
        RECT 706.575 1117.040 706.865 1117.210 ;
        RECT 707.035 1117.040 707.325 1117.210 ;
        RECT 707.495 1117.040 707.785 1117.210 ;
        RECT 707.955 1117.040 708.245 1117.210 ;
        RECT 708.415 1117.040 708.705 1117.210 ;
        RECT 708.875 1117.040 709.165 1117.210 ;
        RECT 709.335 1117.040 709.625 1117.210 ;
        RECT 709.795 1117.040 710.085 1117.210 ;
        RECT 710.255 1117.040 710.545 1117.210 ;
        RECT 710.715 1117.040 711.005 1117.210 ;
        RECT 711.175 1117.040 711.465 1117.210 ;
        RECT 711.635 1117.040 711.925 1117.210 ;
        RECT 712.095 1117.040 712.385 1117.210 ;
        RECT 712.555 1117.040 712.845 1117.210 ;
        RECT 713.015 1117.040 713.305 1117.210 ;
        RECT 713.475 1117.040 713.765 1117.210 ;
        RECT 713.935 1117.040 714.225 1117.210 ;
        RECT 714.395 1117.040 714.685 1117.210 ;
        RECT 714.855 1117.040 715.145 1117.210 ;
        RECT 715.315 1117.040 715.605 1117.210 ;
        RECT 715.775 1117.040 716.065 1117.210 ;
        RECT 716.235 1117.040 716.525 1117.210 ;
        RECT 716.695 1117.040 716.985 1117.210 ;
        RECT 717.155 1117.040 717.445 1117.210 ;
        RECT 717.615 1117.040 717.905 1117.210 ;
        RECT 718.075 1117.040 718.365 1117.210 ;
        RECT 718.535 1117.040 718.825 1117.210 ;
        RECT 718.995 1117.040 719.285 1117.210 ;
        RECT 719.455 1117.040 719.745 1117.210 ;
        RECT 719.915 1117.040 720.205 1117.210 ;
        RECT 720.375 1117.040 720.665 1117.210 ;
        RECT 720.835 1117.040 721.125 1117.210 ;
        RECT 721.295 1117.040 721.585 1117.210 ;
        RECT 721.755 1117.040 722.045 1117.210 ;
        RECT 722.215 1117.040 722.505 1117.210 ;
        RECT 722.675 1117.040 722.965 1117.210 ;
        RECT 723.135 1117.040 723.425 1117.210 ;
        RECT 723.595 1117.040 723.885 1117.210 ;
        RECT 724.055 1117.040 724.345 1117.210 ;
        RECT 724.515 1117.040 724.805 1117.210 ;
        RECT 724.975 1117.040 725.265 1117.210 ;
        RECT 725.435 1117.040 725.725 1117.210 ;
        RECT 725.895 1117.040 726.185 1117.210 ;
        RECT 726.355 1117.040 726.645 1117.210 ;
        RECT 726.815 1117.040 727.105 1117.210 ;
        RECT 727.275 1117.040 727.565 1117.210 ;
        RECT 727.735 1117.040 728.025 1117.210 ;
        RECT 728.195 1117.040 728.485 1117.210 ;
        RECT 728.655 1117.040 728.945 1117.210 ;
        RECT 729.115 1117.040 729.405 1117.210 ;
        RECT 729.575 1117.040 729.865 1117.210 ;
        RECT 730.035 1117.040 730.325 1117.210 ;
        RECT 730.495 1117.040 730.785 1117.210 ;
        RECT 730.955 1117.040 731.245 1117.210 ;
        RECT 731.415 1117.040 731.705 1117.210 ;
        RECT 731.875 1117.040 732.165 1117.210 ;
        RECT 732.335 1117.040 732.625 1117.210 ;
        RECT 732.795 1117.040 733.085 1117.210 ;
        RECT 733.255 1117.040 733.545 1117.210 ;
        RECT 733.715 1117.040 734.005 1117.210 ;
        RECT 734.175 1117.040 734.465 1117.210 ;
        RECT 734.635 1117.040 734.925 1117.210 ;
        RECT 735.095 1117.040 735.385 1117.210 ;
        RECT 735.555 1117.040 735.845 1117.210 ;
        RECT 736.015 1117.040 736.305 1117.210 ;
        RECT 736.475 1117.040 736.765 1117.210 ;
        RECT 736.935 1117.040 737.225 1117.210 ;
        RECT 737.395 1117.040 737.685 1117.210 ;
        RECT 737.855 1117.040 738.145 1117.210 ;
        RECT 738.315 1117.040 738.605 1117.210 ;
        RECT 738.775 1117.040 739.065 1117.210 ;
        RECT 739.235 1117.040 739.525 1117.210 ;
        RECT 739.695 1117.040 739.985 1117.210 ;
        RECT 740.155 1117.040 740.445 1117.210 ;
        RECT 740.615 1117.040 740.905 1117.210 ;
        RECT 741.075 1117.040 741.365 1117.210 ;
        RECT 741.535 1117.040 741.825 1117.210 ;
        RECT 741.995 1117.040 742.285 1117.210 ;
        RECT 742.455 1117.040 742.745 1117.210 ;
        RECT 742.915 1117.040 743.205 1117.210 ;
        RECT 743.375 1117.040 743.665 1117.210 ;
        RECT 743.835 1117.040 744.125 1117.210 ;
        RECT 744.295 1117.040 744.585 1117.210 ;
        RECT 744.755 1117.040 745.045 1117.210 ;
        RECT 745.215 1117.040 745.505 1117.210 ;
        RECT 745.675 1117.040 745.965 1117.210 ;
        RECT 746.135 1117.040 746.425 1117.210 ;
        RECT 746.595 1117.040 746.885 1117.210 ;
        RECT 747.055 1117.040 747.345 1117.210 ;
        RECT 747.515 1117.040 747.805 1117.210 ;
        RECT 747.975 1117.040 748.265 1117.210 ;
        RECT 748.435 1117.040 748.725 1117.210 ;
        RECT 748.895 1117.040 749.185 1117.210 ;
        RECT 749.355 1117.040 749.645 1117.210 ;
        RECT 749.815 1117.040 750.105 1117.210 ;
        RECT 750.275 1117.040 750.565 1117.210 ;
        RECT 750.735 1117.040 751.025 1117.210 ;
        RECT 751.195 1117.040 751.485 1117.210 ;
        RECT 751.655 1117.040 751.945 1117.210 ;
        RECT 752.115 1117.040 752.405 1117.210 ;
        RECT 752.575 1117.040 752.865 1117.210 ;
        RECT 753.035 1117.040 753.325 1117.210 ;
        RECT 753.495 1117.040 753.785 1117.210 ;
        RECT 753.955 1117.040 754.245 1117.210 ;
        RECT 754.415 1117.040 754.705 1117.210 ;
        RECT 754.875 1117.040 755.165 1117.210 ;
        RECT 755.335 1117.040 755.625 1117.210 ;
        RECT 755.795 1117.040 756.085 1117.210 ;
        RECT 756.255 1117.040 756.545 1117.210 ;
        RECT 756.715 1117.040 757.005 1117.210 ;
        RECT 757.175 1117.040 757.465 1117.210 ;
        RECT 757.635 1117.040 757.925 1117.210 ;
        RECT 758.095 1117.040 758.385 1117.210 ;
        RECT 758.555 1117.040 758.845 1117.210 ;
        RECT 759.015 1117.040 759.305 1117.210 ;
        RECT 759.475 1117.040 759.765 1117.210 ;
        RECT 759.935 1117.040 760.225 1117.210 ;
        RECT 760.395 1117.040 760.685 1117.210 ;
        RECT 760.855 1117.040 761.145 1117.210 ;
        RECT 761.315 1117.040 761.605 1117.210 ;
        RECT 761.775 1117.040 762.065 1117.210 ;
        RECT 762.235 1117.040 762.525 1117.210 ;
        RECT 762.695 1117.040 762.985 1117.210 ;
        RECT 763.155 1117.040 763.445 1117.210 ;
        RECT 763.615 1117.040 763.905 1117.210 ;
        RECT 764.075 1117.040 764.365 1117.210 ;
        RECT 764.535 1117.040 764.825 1117.210 ;
        RECT 764.995 1117.040 765.285 1117.210 ;
        RECT 765.455 1117.040 765.745 1117.210 ;
        RECT 765.915 1117.040 766.205 1117.210 ;
        RECT 766.375 1117.040 766.665 1117.210 ;
        RECT 766.835 1117.040 767.125 1117.210 ;
        RECT 767.295 1117.040 767.585 1117.210 ;
        RECT 767.755 1117.040 768.045 1117.210 ;
        RECT 768.215 1117.040 768.505 1117.210 ;
        RECT 768.675 1117.040 768.965 1117.210 ;
        RECT 769.135 1117.040 769.425 1117.210 ;
        RECT 769.595 1117.040 769.885 1117.210 ;
        RECT 770.055 1117.040 770.345 1117.210 ;
        RECT 770.515 1117.040 770.805 1117.210 ;
        RECT 770.975 1117.040 771.265 1117.210 ;
        RECT 771.435 1117.040 771.725 1117.210 ;
        RECT 771.895 1117.040 772.185 1117.210 ;
        RECT 772.355 1117.040 772.645 1117.210 ;
        RECT 772.815 1117.040 773.105 1117.210 ;
        RECT 773.275 1117.040 773.565 1117.210 ;
        RECT 773.735 1117.040 774.025 1117.210 ;
        RECT 774.195 1117.040 774.485 1117.210 ;
        RECT 774.655 1117.040 774.945 1117.210 ;
        RECT 775.115 1117.040 775.405 1117.210 ;
        RECT 775.575 1117.040 775.865 1117.210 ;
        RECT 776.035 1117.040 776.325 1117.210 ;
        RECT 776.495 1117.040 776.785 1117.210 ;
        RECT 776.955 1117.040 777.245 1117.210 ;
        RECT 777.415 1117.040 777.705 1117.210 ;
        RECT 777.875 1117.040 778.165 1117.210 ;
        RECT 778.335 1117.040 778.625 1117.210 ;
        RECT 778.795 1117.040 779.085 1117.210 ;
        RECT 779.255 1117.040 779.545 1117.210 ;
        RECT 779.715 1117.040 780.005 1117.210 ;
        RECT 780.175 1117.040 780.465 1117.210 ;
        RECT 780.635 1117.040 780.925 1117.210 ;
        RECT 781.095 1117.040 781.385 1117.210 ;
        RECT 781.555 1117.040 781.845 1117.210 ;
        RECT 782.015 1117.040 782.305 1117.210 ;
        RECT 782.475 1117.040 782.765 1117.210 ;
        RECT 782.935 1117.040 783.225 1117.210 ;
        RECT 783.395 1117.040 783.685 1117.210 ;
        RECT 783.855 1117.040 784.145 1117.210 ;
        RECT 784.315 1117.040 784.605 1117.210 ;
        RECT 784.775 1117.040 785.065 1117.210 ;
        RECT 785.235 1117.040 785.525 1117.210 ;
        RECT 785.695 1117.040 785.985 1117.210 ;
        RECT 786.155 1117.040 786.445 1117.210 ;
        RECT 786.615 1117.040 786.905 1117.210 ;
        RECT 787.075 1117.040 787.365 1117.210 ;
        RECT 787.535 1117.040 787.825 1117.210 ;
        RECT 787.995 1117.040 788.285 1117.210 ;
        RECT 788.455 1117.040 788.745 1117.210 ;
        RECT 788.915 1117.040 789.205 1117.210 ;
        RECT 789.375 1117.040 789.665 1117.210 ;
        RECT 789.835 1117.040 790.125 1117.210 ;
        RECT 790.295 1117.040 790.585 1117.210 ;
        RECT 790.755 1117.040 791.045 1117.210 ;
        RECT 791.215 1117.040 791.505 1117.210 ;
        RECT 791.675 1117.040 791.965 1117.210 ;
        RECT 792.135 1117.040 792.425 1117.210 ;
        RECT 792.595 1117.040 792.885 1117.210 ;
        RECT 793.055 1117.040 793.345 1117.210 ;
        RECT 793.515 1117.040 793.805 1117.210 ;
        RECT 793.975 1117.040 794.265 1117.210 ;
        RECT 794.435 1117.040 794.725 1117.210 ;
        RECT 794.895 1117.040 795.040 1117.210 ;
        RECT 1969.000 1117.040 1969.145 1117.210 ;
        RECT 1969.315 1117.040 1969.605 1117.210 ;
        RECT 1969.775 1117.040 1970.065 1117.210 ;
        RECT 1970.235 1117.040 1970.525 1117.210 ;
        RECT 1970.695 1117.040 1970.985 1117.210 ;
        RECT 1971.155 1117.040 1971.445 1117.210 ;
        RECT 1971.615 1117.040 1971.905 1117.210 ;
        RECT 1972.075 1117.040 1972.365 1117.210 ;
        RECT 1972.535 1117.040 1972.825 1117.210 ;
        RECT 1972.995 1117.040 1973.285 1117.210 ;
        RECT 1973.455 1117.040 1973.745 1117.210 ;
        RECT 1973.915 1117.040 1974.205 1117.210 ;
        RECT 1974.375 1117.040 1974.665 1117.210 ;
        RECT 1974.835 1117.040 1975.125 1117.210 ;
        RECT 1975.295 1117.040 1975.585 1117.210 ;
        RECT 1975.755 1117.040 1976.045 1117.210 ;
        RECT 1976.215 1117.040 1976.505 1117.210 ;
        RECT 1976.675 1117.040 1976.965 1117.210 ;
        RECT 1977.135 1117.040 1977.425 1117.210 ;
        RECT 1977.595 1117.040 1977.885 1117.210 ;
        RECT 1978.055 1117.040 1978.345 1117.210 ;
        RECT 1978.515 1117.040 1978.805 1117.210 ;
        RECT 1978.975 1117.040 1979.265 1117.210 ;
        RECT 1979.435 1117.040 1979.725 1117.210 ;
        RECT 1979.895 1117.040 1980.185 1117.210 ;
        RECT 1980.355 1117.040 1980.645 1117.210 ;
        RECT 1980.815 1117.040 1981.105 1117.210 ;
        RECT 1981.275 1117.040 1981.565 1117.210 ;
        RECT 1981.735 1117.040 1982.025 1117.210 ;
        RECT 1982.195 1117.040 1982.485 1117.210 ;
        RECT 1982.655 1117.040 1982.945 1117.210 ;
        RECT 1983.115 1117.040 1983.405 1117.210 ;
        RECT 1983.575 1117.040 1983.865 1117.210 ;
        RECT 1984.035 1117.040 1984.325 1117.210 ;
        RECT 1984.495 1117.040 1984.785 1117.210 ;
        RECT 1984.955 1117.040 1985.245 1117.210 ;
        RECT 1985.415 1117.040 1985.705 1117.210 ;
        RECT 1985.875 1117.040 1986.165 1117.210 ;
        RECT 1986.335 1117.040 1986.625 1117.210 ;
        RECT 1986.795 1117.040 1987.085 1117.210 ;
        RECT 1987.255 1117.040 1987.545 1117.210 ;
        RECT 1987.715 1117.040 1988.005 1117.210 ;
        RECT 1988.175 1117.040 1988.465 1117.210 ;
        RECT 1988.635 1117.040 1988.925 1117.210 ;
        RECT 1989.095 1117.040 1989.385 1117.210 ;
        RECT 1989.555 1117.040 1989.845 1117.210 ;
        RECT 1990.015 1117.040 1990.305 1117.210 ;
        RECT 1990.475 1117.040 1990.765 1117.210 ;
        RECT 1990.935 1117.040 1991.225 1117.210 ;
        RECT 1991.395 1117.040 1991.685 1117.210 ;
        RECT 1991.855 1117.040 1992.145 1117.210 ;
        RECT 1992.315 1117.040 1992.605 1117.210 ;
        RECT 1992.775 1117.040 1993.065 1117.210 ;
        RECT 1993.235 1117.040 1993.525 1117.210 ;
        RECT 1993.695 1117.040 1993.985 1117.210 ;
        RECT 1994.155 1117.040 1994.445 1117.210 ;
        RECT 1994.615 1117.040 1994.905 1117.210 ;
        RECT 1995.075 1117.040 1995.365 1117.210 ;
        RECT 1995.535 1117.040 1995.825 1117.210 ;
        RECT 1995.995 1117.040 1996.285 1117.210 ;
        RECT 1996.455 1117.040 1996.745 1117.210 ;
        RECT 1996.915 1117.040 1997.205 1117.210 ;
        RECT 1997.375 1117.040 1997.665 1117.210 ;
        RECT 1997.835 1117.040 1998.125 1117.210 ;
        RECT 1998.295 1117.040 1998.585 1117.210 ;
        RECT 1998.755 1117.040 1999.045 1117.210 ;
        RECT 1999.215 1117.040 1999.505 1117.210 ;
        RECT 1999.675 1117.040 1999.965 1117.210 ;
        RECT 2000.135 1117.040 2000.425 1117.210 ;
        RECT 2000.595 1117.040 2000.885 1117.210 ;
        RECT 2001.055 1117.040 2001.345 1117.210 ;
        RECT 2001.515 1117.040 2001.805 1117.210 ;
        RECT 2001.975 1117.040 2002.265 1117.210 ;
        RECT 2002.435 1117.040 2002.725 1117.210 ;
        RECT 2002.895 1117.040 2003.185 1117.210 ;
        RECT 2003.355 1117.040 2003.645 1117.210 ;
        RECT 2003.815 1117.040 2004.105 1117.210 ;
        RECT 2004.275 1117.040 2004.565 1117.210 ;
        RECT 2004.735 1117.040 2005.025 1117.210 ;
        RECT 2005.195 1117.040 2005.485 1117.210 ;
        RECT 2005.655 1117.040 2005.945 1117.210 ;
        RECT 2006.115 1117.040 2006.405 1117.210 ;
        RECT 2006.575 1117.040 2006.865 1117.210 ;
        RECT 2007.035 1117.040 2007.325 1117.210 ;
        RECT 2007.495 1117.040 2007.785 1117.210 ;
        RECT 2007.955 1117.040 2008.245 1117.210 ;
        RECT 2008.415 1117.040 2008.705 1117.210 ;
        RECT 2008.875 1117.040 2009.165 1117.210 ;
        RECT 2009.335 1117.040 2009.625 1117.210 ;
        RECT 2009.795 1117.040 2010.085 1117.210 ;
        RECT 2010.255 1117.040 2010.545 1117.210 ;
        RECT 2010.715 1117.040 2011.005 1117.210 ;
        RECT 2011.175 1117.040 2011.465 1117.210 ;
        RECT 2011.635 1117.040 2011.925 1117.210 ;
        RECT 2012.095 1117.040 2012.385 1117.210 ;
        RECT 2012.555 1117.040 2012.845 1117.210 ;
        RECT 2013.015 1117.040 2013.305 1117.210 ;
        RECT 2013.475 1117.040 2013.765 1117.210 ;
        RECT 2013.935 1117.040 2014.225 1117.210 ;
        RECT 2014.395 1117.040 2014.685 1117.210 ;
        RECT 2014.855 1117.040 2015.145 1117.210 ;
        RECT 2015.315 1117.040 2015.605 1117.210 ;
        RECT 2015.775 1117.040 2016.065 1117.210 ;
        RECT 2016.235 1117.040 2016.525 1117.210 ;
        RECT 2016.695 1117.040 2016.985 1117.210 ;
        RECT 2017.155 1117.040 2017.445 1117.210 ;
        RECT 2017.615 1117.040 2017.905 1117.210 ;
        RECT 2018.075 1117.040 2018.365 1117.210 ;
        RECT 2018.535 1117.040 2018.825 1117.210 ;
        RECT 2018.995 1117.040 2019.285 1117.210 ;
        RECT 2019.455 1117.040 2019.745 1117.210 ;
        RECT 2019.915 1117.040 2020.205 1117.210 ;
        RECT 2020.375 1117.040 2020.665 1117.210 ;
        RECT 2020.835 1117.040 2021.125 1117.210 ;
        RECT 2021.295 1117.040 2021.585 1117.210 ;
        RECT 2021.755 1117.040 2022.045 1117.210 ;
        RECT 2022.215 1117.040 2022.505 1117.210 ;
        RECT 2022.675 1117.040 2022.965 1117.210 ;
        RECT 2023.135 1117.040 2023.425 1117.210 ;
        RECT 2023.595 1117.040 2023.885 1117.210 ;
        RECT 2024.055 1117.040 2024.345 1117.210 ;
        RECT 2024.515 1117.040 2024.805 1117.210 ;
        RECT 2024.975 1117.040 2025.265 1117.210 ;
        RECT 2025.435 1117.040 2025.725 1117.210 ;
        RECT 2025.895 1117.040 2026.185 1117.210 ;
        RECT 2026.355 1117.040 2026.645 1117.210 ;
        RECT 2026.815 1117.040 2027.105 1117.210 ;
        RECT 2027.275 1117.040 2027.565 1117.210 ;
        RECT 2027.735 1117.040 2028.025 1117.210 ;
        RECT 2028.195 1117.040 2028.485 1117.210 ;
        RECT 2028.655 1117.040 2028.945 1117.210 ;
        RECT 2029.115 1117.040 2029.405 1117.210 ;
        RECT 2029.575 1117.040 2029.865 1117.210 ;
        RECT 2030.035 1117.040 2030.325 1117.210 ;
        RECT 2030.495 1117.040 2030.785 1117.210 ;
        RECT 2030.955 1117.040 2031.245 1117.210 ;
        RECT 2031.415 1117.040 2031.705 1117.210 ;
        RECT 2031.875 1117.040 2032.165 1117.210 ;
        RECT 2032.335 1117.040 2032.625 1117.210 ;
        RECT 2032.795 1117.040 2033.085 1117.210 ;
        RECT 2033.255 1117.040 2033.545 1117.210 ;
        RECT 2033.715 1117.040 2034.005 1117.210 ;
        RECT 2034.175 1117.040 2034.465 1117.210 ;
        RECT 2034.635 1117.040 2034.925 1117.210 ;
        RECT 2035.095 1117.040 2035.385 1117.210 ;
        RECT 2035.555 1117.040 2035.845 1117.210 ;
        RECT 2036.015 1117.040 2036.305 1117.210 ;
        RECT 2036.475 1117.040 2036.765 1117.210 ;
        RECT 2036.935 1117.040 2037.225 1117.210 ;
        RECT 2037.395 1117.040 2037.685 1117.210 ;
        RECT 2037.855 1117.040 2038.145 1117.210 ;
        RECT 2038.315 1117.040 2038.605 1117.210 ;
        RECT 2038.775 1117.040 2039.065 1117.210 ;
        RECT 2039.235 1117.040 2039.525 1117.210 ;
        RECT 2039.695 1117.040 2039.985 1117.210 ;
        RECT 2040.155 1117.040 2040.445 1117.210 ;
        RECT 2040.615 1117.040 2040.905 1117.210 ;
        RECT 2041.075 1117.040 2041.365 1117.210 ;
        RECT 2041.535 1117.040 2041.825 1117.210 ;
        RECT 2041.995 1117.040 2042.285 1117.210 ;
        RECT 2042.455 1117.040 2042.745 1117.210 ;
        RECT 2042.915 1117.040 2043.205 1117.210 ;
        RECT 2043.375 1117.040 2043.665 1117.210 ;
        RECT 2043.835 1117.040 2044.125 1117.210 ;
        RECT 2044.295 1117.040 2044.585 1117.210 ;
        RECT 2044.755 1117.040 2045.045 1117.210 ;
        RECT 2045.215 1117.040 2045.505 1117.210 ;
        RECT 2045.675 1117.040 2045.965 1117.210 ;
        RECT 2046.135 1117.040 2046.425 1117.210 ;
        RECT 2046.595 1117.040 2046.885 1117.210 ;
        RECT 2047.055 1117.040 2047.345 1117.210 ;
        RECT 2047.515 1117.040 2047.805 1117.210 ;
        RECT 2047.975 1117.040 2048.265 1117.210 ;
        RECT 2048.435 1117.040 2048.725 1117.210 ;
        RECT 2048.895 1117.040 2049.185 1117.210 ;
        RECT 2049.355 1117.040 2049.645 1117.210 ;
        RECT 2049.815 1117.040 2050.105 1117.210 ;
        RECT 2050.275 1117.040 2050.565 1117.210 ;
        RECT 2050.735 1117.040 2051.025 1117.210 ;
        RECT 2051.195 1117.040 2051.485 1117.210 ;
        RECT 2051.655 1117.040 2051.945 1117.210 ;
        RECT 2052.115 1117.040 2052.405 1117.210 ;
        RECT 2052.575 1117.040 2052.865 1117.210 ;
        RECT 2053.035 1117.040 2053.325 1117.210 ;
        RECT 2053.495 1117.040 2053.785 1117.210 ;
        RECT 2053.955 1117.040 2054.245 1117.210 ;
        RECT 2054.415 1117.040 2054.705 1117.210 ;
        RECT 2054.875 1117.040 2055.165 1117.210 ;
        RECT 2055.335 1117.040 2055.625 1117.210 ;
        RECT 2055.795 1117.040 2056.085 1117.210 ;
        RECT 2056.255 1117.040 2056.545 1117.210 ;
        RECT 2056.715 1117.040 2057.005 1117.210 ;
        RECT 2057.175 1117.040 2057.465 1117.210 ;
        RECT 2057.635 1117.040 2057.925 1117.210 ;
        RECT 2058.095 1117.040 2058.385 1117.210 ;
        RECT 2058.555 1117.040 2058.845 1117.210 ;
        RECT 2059.015 1117.040 2059.305 1117.210 ;
        RECT 2059.475 1117.040 2059.765 1117.210 ;
        RECT 2059.935 1117.040 2060.225 1117.210 ;
        RECT 2060.395 1117.040 2060.685 1117.210 ;
        RECT 2060.855 1117.040 2061.145 1117.210 ;
        RECT 2061.315 1117.040 2061.605 1117.210 ;
        RECT 2061.775 1117.040 2062.065 1117.210 ;
        RECT 2062.235 1117.040 2062.525 1117.210 ;
        RECT 2062.695 1117.040 2062.985 1117.210 ;
        RECT 2063.155 1117.040 2063.445 1117.210 ;
        RECT 2063.615 1117.040 2063.905 1117.210 ;
        RECT 2064.075 1117.040 2064.365 1117.210 ;
        RECT 2064.535 1117.040 2064.825 1117.210 ;
        RECT 2064.995 1117.040 2065.285 1117.210 ;
        RECT 2065.455 1117.040 2065.745 1117.210 ;
        RECT 2065.915 1117.040 2066.205 1117.210 ;
        RECT 2066.375 1117.040 2066.665 1117.210 ;
        RECT 2066.835 1117.040 2067.125 1117.210 ;
        RECT 2067.295 1117.040 2067.585 1117.210 ;
        RECT 2067.755 1117.040 2068.045 1117.210 ;
        RECT 2068.215 1117.040 2068.505 1117.210 ;
        RECT 2068.675 1117.040 2068.965 1117.210 ;
        RECT 2069.135 1117.040 2069.425 1117.210 ;
        RECT 2069.595 1117.040 2069.885 1117.210 ;
        RECT 2070.055 1117.040 2070.345 1117.210 ;
        RECT 2070.515 1117.040 2070.805 1117.210 ;
        RECT 2070.975 1117.040 2071.265 1117.210 ;
        RECT 2071.435 1117.040 2071.725 1117.210 ;
        RECT 2071.895 1117.040 2072.185 1117.210 ;
        RECT 2072.355 1117.040 2072.645 1117.210 ;
        RECT 2072.815 1117.040 2073.105 1117.210 ;
        RECT 2073.275 1117.040 2073.565 1117.210 ;
        RECT 2073.735 1117.040 2074.025 1117.210 ;
        RECT 2074.195 1117.040 2074.485 1117.210 ;
        RECT 2074.655 1117.040 2074.945 1117.210 ;
        RECT 2075.115 1117.040 2075.405 1117.210 ;
        RECT 2075.575 1117.040 2075.865 1117.210 ;
        RECT 2076.035 1117.040 2076.325 1117.210 ;
        RECT 2076.495 1117.040 2076.785 1117.210 ;
        RECT 2076.955 1117.040 2077.245 1117.210 ;
        RECT 2077.415 1117.040 2077.705 1117.210 ;
        RECT 2077.875 1117.040 2078.165 1117.210 ;
        RECT 2078.335 1117.040 2078.625 1117.210 ;
        RECT 2078.795 1117.040 2079.085 1117.210 ;
        RECT 2079.255 1117.040 2079.545 1117.210 ;
        RECT 2079.715 1117.040 2080.005 1117.210 ;
        RECT 2080.175 1117.040 2080.465 1117.210 ;
        RECT 2080.635 1117.040 2080.925 1117.210 ;
        RECT 2081.095 1117.040 2081.385 1117.210 ;
        RECT 2081.555 1117.040 2081.845 1117.210 ;
        RECT 2082.015 1117.040 2082.305 1117.210 ;
        RECT 2082.475 1117.040 2082.765 1117.210 ;
        RECT 2082.935 1117.040 2083.225 1117.210 ;
        RECT 2083.395 1117.040 2083.685 1117.210 ;
        RECT 2083.855 1117.040 2084.145 1117.210 ;
        RECT 2084.315 1117.040 2084.605 1117.210 ;
        RECT 2084.775 1117.040 2085.065 1117.210 ;
        RECT 2085.235 1117.040 2085.525 1117.210 ;
        RECT 2085.695 1117.040 2085.985 1117.210 ;
        RECT 2086.155 1117.040 2086.445 1117.210 ;
        RECT 2086.615 1117.040 2086.905 1117.210 ;
        RECT 2087.075 1117.040 2087.365 1117.210 ;
        RECT 2087.535 1117.040 2087.825 1117.210 ;
        RECT 2087.995 1117.040 2088.285 1117.210 ;
        RECT 2088.455 1117.040 2088.745 1117.210 ;
        RECT 2088.915 1117.040 2089.205 1117.210 ;
        RECT 2089.375 1117.040 2089.665 1117.210 ;
        RECT 2089.835 1117.040 2090.125 1117.210 ;
        RECT 2090.295 1117.040 2090.585 1117.210 ;
        RECT 2090.755 1117.040 2091.045 1117.210 ;
        RECT 2091.215 1117.040 2091.505 1117.210 ;
        RECT 2091.675 1117.040 2091.965 1117.210 ;
        RECT 2092.135 1117.040 2092.425 1117.210 ;
        RECT 2092.595 1117.040 2092.885 1117.210 ;
        RECT 2093.055 1117.040 2093.345 1117.210 ;
        RECT 2093.515 1117.040 2093.805 1117.210 ;
        RECT 2093.975 1117.040 2094.265 1117.210 ;
        RECT 2094.435 1117.040 2094.725 1117.210 ;
        RECT 2094.895 1117.040 2095.040 1117.210 ;
        RECT 669.085 1116.315 669.375 1117.040 ;
        RECT 669.935 1116.240 670.265 1117.040 ;
      LAYER li1 ;
        RECT 670.435 1116.390 670.605 1116.870 ;
      LAYER li1 ;
        RECT 670.775 1116.560 671.105 1117.040 ;
      LAYER li1 ;
        RECT 671.275 1116.390 671.445 1116.870 ;
      LAYER li1 ;
        RECT 671.615 1116.560 671.945 1117.040 ;
      LAYER li1 ;
        RECT 672.115 1116.390 672.285 1116.870 ;
      LAYER li1 ;
        RECT 672.455 1116.560 672.785 1117.040 ;
      LAYER li1 ;
        RECT 672.955 1116.390 673.125 1116.870 ;
      LAYER li1 ;
        RECT 673.295 1116.560 673.625 1117.040 ;
        RECT 673.795 1116.390 673.965 1116.865 ;
        RECT 674.135 1116.560 674.465 1117.040 ;
        RECT 674.635 1116.390 674.805 1116.870 ;
      LAYER li1 ;
        RECT 670.435 1116.220 673.125 1116.390 ;
      LAYER li1 ;
        RECT 673.385 1116.220 674.805 1116.390 ;
        RECT 675.065 1116.315 675.355 1117.040 ;
        RECT 675.915 1116.240 676.245 1117.040 ;
      LAYER li1 ;
        RECT 676.415 1116.390 676.585 1116.870 ;
      LAYER li1 ;
        RECT 676.755 1116.560 677.085 1117.040 ;
      LAYER li1 ;
        RECT 677.255 1116.390 677.425 1116.870 ;
      LAYER li1 ;
        RECT 677.595 1116.560 677.925 1117.040 ;
      LAYER li1 ;
        RECT 678.095 1116.390 678.265 1116.870 ;
      LAYER li1 ;
        RECT 678.435 1116.560 678.765 1117.040 ;
      LAYER li1 ;
        RECT 678.935 1116.390 679.105 1116.870 ;
      LAYER li1 ;
        RECT 679.275 1116.560 679.605 1117.040 ;
        RECT 679.775 1116.390 679.945 1116.865 ;
        RECT 680.115 1116.560 680.445 1117.040 ;
        RECT 680.615 1116.390 680.785 1116.870 ;
      LAYER li1 ;
        RECT 676.415 1116.220 679.105 1116.390 ;
      LAYER li1 ;
        RECT 679.365 1116.220 680.785 1116.390 ;
        RECT 681.045 1116.315 681.335 1117.040 ;
        RECT 681.895 1116.240 682.225 1117.040 ;
      LAYER li1 ;
        RECT 682.395 1116.390 682.565 1116.870 ;
      LAYER li1 ;
        RECT 682.735 1116.560 683.065 1117.040 ;
      LAYER li1 ;
        RECT 683.235 1116.390 683.405 1116.870 ;
      LAYER li1 ;
        RECT 683.575 1116.560 683.905 1117.040 ;
      LAYER li1 ;
        RECT 684.075 1116.390 684.245 1116.870 ;
      LAYER li1 ;
        RECT 684.415 1116.560 684.745 1117.040 ;
      LAYER li1 ;
        RECT 684.915 1116.390 685.085 1116.870 ;
      LAYER li1 ;
        RECT 685.255 1116.560 685.585 1117.040 ;
        RECT 685.755 1116.390 685.925 1116.865 ;
        RECT 686.095 1116.560 686.425 1117.040 ;
        RECT 686.595 1116.390 686.765 1116.870 ;
      LAYER li1 ;
        RECT 682.395 1116.220 685.085 1116.390 ;
      LAYER li1 ;
        RECT 685.345 1116.220 686.765 1116.390 ;
        RECT 687.025 1116.315 687.315 1117.040 ;
        RECT 687.875 1116.240 688.205 1117.040 ;
      LAYER li1 ;
        RECT 688.375 1116.390 688.545 1116.870 ;
      LAYER li1 ;
        RECT 688.715 1116.560 689.045 1117.040 ;
      LAYER li1 ;
        RECT 689.215 1116.390 689.385 1116.870 ;
      LAYER li1 ;
        RECT 689.555 1116.560 689.885 1117.040 ;
      LAYER li1 ;
        RECT 690.055 1116.390 690.225 1116.870 ;
      LAYER li1 ;
        RECT 690.395 1116.560 690.725 1117.040 ;
      LAYER li1 ;
        RECT 690.895 1116.390 691.065 1116.870 ;
      LAYER li1 ;
        RECT 691.235 1116.560 691.565 1117.040 ;
        RECT 691.735 1116.390 691.905 1116.865 ;
        RECT 692.075 1116.560 692.405 1117.040 ;
        RECT 692.575 1116.390 692.745 1116.870 ;
      LAYER li1 ;
        RECT 688.375 1116.220 691.065 1116.390 ;
      LAYER li1 ;
        RECT 691.325 1116.220 692.745 1116.390 ;
        RECT 693.005 1116.315 693.295 1117.040 ;
        RECT 693.855 1116.240 694.185 1117.040 ;
      LAYER li1 ;
        RECT 694.355 1116.390 694.525 1116.870 ;
      LAYER li1 ;
        RECT 694.695 1116.560 695.025 1117.040 ;
      LAYER li1 ;
        RECT 695.195 1116.390 695.365 1116.870 ;
      LAYER li1 ;
        RECT 695.535 1116.560 695.865 1117.040 ;
      LAYER li1 ;
        RECT 696.035 1116.390 696.205 1116.870 ;
      LAYER li1 ;
        RECT 696.375 1116.560 696.705 1117.040 ;
      LAYER li1 ;
        RECT 696.875 1116.390 697.045 1116.870 ;
      LAYER li1 ;
        RECT 697.215 1116.560 697.545 1117.040 ;
        RECT 697.715 1116.390 697.885 1116.865 ;
        RECT 698.055 1116.560 698.385 1117.040 ;
        RECT 698.555 1116.390 698.725 1116.870 ;
      LAYER li1 ;
        RECT 694.355 1116.220 697.045 1116.390 ;
      LAYER li1 ;
        RECT 697.305 1116.220 698.725 1116.390 ;
        RECT 698.985 1116.315 699.275 1117.040 ;
        RECT 699.835 1116.240 700.165 1117.040 ;
      LAYER li1 ;
        RECT 700.335 1116.390 700.505 1116.870 ;
      LAYER li1 ;
        RECT 700.675 1116.560 701.005 1117.040 ;
      LAYER li1 ;
        RECT 701.175 1116.390 701.345 1116.870 ;
      LAYER li1 ;
        RECT 701.515 1116.560 701.845 1117.040 ;
      LAYER li1 ;
        RECT 702.015 1116.390 702.185 1116.870 ;
      LAYER li1 ;
        RECT 702.355 1116.560 702.685 1117.040 ;
      LAYER li1 ;
        RECT 702.855 1116.390 703.025 1116.870 ;
      LAYER li1 ;
        RECT 703.195 1116.560 703.525 1117.040 ;
        RECT 703.695 1116.390 703.865 1116.865 ;
        RECT 704.035 1116.560 704.365 1117.040 ;
        RECT 704.535 1116.390 704.705 1116.870 ;
      LAYER li1 ;
        RECT 700.335 1116.220 703.025 1116.390 ;
      LAYER li1 ;
        RECT 703.285 1116.220 704.705 1116.390 ;
        RECT 704.965 1116.315 705.255 1117.040 ;
        RECT 705.815 1116.240 706.145 1117.040 ;
      LAYER li1 ;
        RECT 706.315 1116.390 706.485 1116.870 ;
      LAYER li1 ;
        RECT 706.655 1116.560 706.985 1117.040 ;
      LAYER li1 ;
        RECT 707.155 1116.390 707.325 1116.870 ;
      LAYER li1 ;
        RECT 707.495 1116.560 707.825 1117.040 ;
      LAYER li1 ;
        RECT 707.995 1116.390 708.165 1116.870 ;
      LAYER li1 ;
        RECT 708.335 1116.560 708.665 1117.040 ;
      LAYER li1 ;
        RECT 708.835 1116.390 709.005 1116.870 ;
      LAYER li1 ;
        RECT 709.175 1116.560 709.505 1117.040 ;
        RECT 709.675 1116.390 709.845 1116.865 ;
        RECT 710.015 1116.560 710.345 1117.040 ;
        RECT 710.515 1116.390 710.685 1116.870 ;
      LAYER li1 ;
        RECT 706.315 1116.220 709.005 1116.390 ;
      LAYER li1 ;
        RECT 709.265 1116.220 710.685 1116.390 ;
        RECT 710.945 1116.315 711.235 1117.040 ;
        RECT 711.795 1116.240 712.125 1117.040 ;
      LAYER li1 ;
        RECT 712.295 1116.390 712.465 1116.870 ;
      LAYER li1 ;
        RECT 712.635 1116.560 712.965 1117.040 ;
      LAYER li1 ;
        RECT 713.135 1116.390 713.305 1116.870 ;
      LAYER li1 ;
        RECT 713.475 1116.560 713.805 1117.040 ;
      LAYER li1 ;
        RECT 713.975 1116.390 714.145 1116.870 ;
      LAYER li1 ;
        RECT 714.315 1116.560 714.645 1117.040 ;
      LAYER li1 ;
        RECT 714.815 1116.390 714.985 1116.870 ;
      LAYER li1 ;
        RECT 715.155 1116.560 715.485 1117.040 ;
        RECT 715.655 1116.390 715.825 1116.865 ;
        RECT 715.995 1116.560 716.325 1117.040 ;
        RECT 716.495 1116.390 716.665 1116.870 ;
      LAYER li1 ;
        RECT 712.295 1116.220 714.985 1116.390 ;
      LAYER li1 ;
        RECT 715.245 1116.220 716.665 1116.390 ;
        RECT 716.925 1116.315 717.215 1117.040 ;
        RECT 717.775 1116.240 718.105 1117.040 ;
      LAYER li1 ;
        RECT 718.275 1116.390 718.445 1116.870 ;
      LAYER li1 ;
        RECT 718.615 1116.560 718.945 1117.040 ;
      LAYER li1 ;
        RECT 719.115 1116.390 719.285 1116.870 ;
      LAYER li1 ;
        RECT 719.455 1116.560 719.785 1117.040 ;
      LAYER li1 ;
        RECT 719.955 1116.390 720.125 1116.870 ;
      LAYER li1 ;
        RECT 720.295 1116.560 720.625 1117.040 ;
      LAYER li1 ;
        RECT 720.795 1116.390 720.965 1116.870 ;
      LAYER li1 ;
        RECT 721.135 1116.560 721.465 1117.040 ;
        RECT 721.635 1116.390 721.805 1116.865 ;
        RECT 721.975 1116.560 722.305 1117.040 ;
        RECT 722.475 1116.390 722.645 1116.870 ;
      LAYER li1 ;
        RECT 718.275 1116.220 720.965 1116.390 ;
      LAYER li1 ;
        RECT 721.225 1116.220 722.645 1116.390 ;
        RECT 722.905 1116.315 723.195 1117.040 ;
        RECT 723.755 1116.240 724.085 1117.040 ;
      LAYER li1 ;
        RECT 724.255 1116.390 724.425 1116.870 ;
      LAYER li1 ;
        RECT 724.595 1116.560 724.925 1117.040 ;
      LAYER li1 ;
        RECT 725.095 1116.390 725.265 1116.870 ;
      LAYER li1 ;
        RECT 725.435 1116.560 725.765 1117.040 ;
      LAYER li1 ;
        RECT 725.935 1116.390 726.105 1116.870 ;
      LAYER li1 ;
        RECT 726.275 1116.560 726.605 1117.040 ;
      LAYER li1 ;
        RECT 726.775 1116.390 726.945 1116.870 ;
      LAYER li1 ;
        RECT 727.115 1116.560 727.445 1117.040 ;
        RECT 727.615 1116.390 727.785 1116.865 ;
        RECT 727.955 1116.560 728.285 1117.040 ;
        RECT 728.455 1116.390 728.625 1116.870 ;
      LAYER li1 ;
        RECT 724.255 1116.220 726.945 1116.390 ;
      LAYER li1 ;
        RECT 727.205 1116.220 728.625 1116.390 ;
        RECT 728.885 1116.315 729.175 1117.040 ;
        RECT 729.735 1116.240 730.065 1117.040 ;
      LAYER li1 ;
        RECT 730.235 1116.390 730.405 1116.870 ;
      LAYER li1 ;
        RECT 730.575 1116.560 730.905 1117.040 ;
      LAYER li1 ;
        RECT 731.075 1116.390 731.245 1116.870 ;
      LAYER li1 ;
        RECT 731.415 1116.560 731.745 1117.040 ;
      LAYER li1 ;
        RECT 731.915 1116.390 732.085 1116.870 ;
      LAYER li1 ;
        RECT 732.255 1116.560 732.585 1117.040 ;
      LAYER li1 ;
        RECT 732.755 1116.390 732.925 1116.870 ;
      LAYER li1 ;
        RECT 733.095 1116.560 733.425 1117.040 ;
        RECT 733.595 1116.390 733.765 1116.865 ;
        RECT 733.935 1116.560 734.265 1117.040 ;
        RECT 734.435 1116.390 734.605 1116.870 ;
      LAYER li1 ;
        RECT 730.235 1116.220 732.925 1116.390 ;
      LAYER li1 ;
        RECT 733.185 1116.220 734.605 1116.390 ;
        RECT 734.865 1116.315 735.155 1117.040 ;
        RECT 735.715 1116.240 736.045 1117.040 ;
      LAYER li1 ;
        RECT 736.215 1116.390 736.385 1116.870 ;
      LAYER li1 ;
        RECT 736.555 1116.560 736.885 1117.040 ;
      LAYER li1 ;
        RECT 737.055 1116.390 737.225 1116.870 ;
      LAYER li1 ;
        RECT 737.395 1116.560 737.725 1117.040 ;
      LAYER li1 ;
        RECT 737.895 1116.390 738.065 1116.870 ;
      LAYER li1 ;
        RECT 738.235 1116.560 738.565 1117.040 ;
      LAYER li1 ;
        RECT 738.735 1116.390 738.905 1116.870 ;
      LAYER li1 ;
        RECT 739.075 1116.560 739.405 1117.040 ;
        RECT 739.575 1116.390 739.745 1116.865 ;
        RECT 739.915 1116.560 740.245 1117.040 ;
        RECT 740.415 1116.390 740.585 1116.870 ;
      LAYER li1 ;
        RECT 736.215 1116.220 738.905 1116.390 ;
      LAYER li1 ;
        RECT 739.165 1116.220 740.585 1116.390 ;
        RECT 740.845 1116.315 741.135 1117.040 ;
        RECT 741.695 1116.240 742.025 1117.040 ;
      LAYER li1 ;
        RECT 742.195 1116.390 742.365 1116.870 ;
      LAYER li1 ;
        RECT 742.535 1116.560 742.865 1117.040 ;
      LAYER li1 ;
        RECT 743.035 1116.390 743.205 1116.870 ;
      LAYER li1 ;
        RECT 743.375 1116.560 743.705 1117.040 ;
      LAYER li1 ;
        RECT 743.875 1116.390 744.045 1116.870 ;
      LAYER li1 ;
        RECT 744.215 1116.560 744.545 1117.040 ;
      LAYER li1 ;
        RECT 744.715 1116.390 744.885 1116.870 ;
      LAYER li1 ;
        RECT 745.055 1116.560 745.385 1117.040 ;
        RECT 745.555 1116.390 745.725 1116.865 ;
        RECT 745.895 1116.560 746.225 1117.040 ;
        RECT 746.395 1116.390 746.565 1116.870 ;
      LAYER li1 ;
        RECT 742.195 1116.220 744.885 1116.390 ;
      LAYER li1 ;
        RECT 745.145 1116.220 746.565 1116.390 ;
        RECT 746.825 1116.315 747.115 1117.040 ;
        RECT 747.675 1116.240 748.005 1117.040 ;
      LAYER li1 ;
        RECT 748.175 1116.390 748.345 1116.870 ;
      LAYER li1 ;
        RECT 748.515 1116.560 748.845 1117.040 ;
      LAYER li1 ;
        RECT 749.015 1116.390 749.185 1116.870 ;
      LAYER li1 ;
        RECT 749.355 1116.560 749.685 1117.040 ;
      LAYER li1 ;
        RECT 749.855 1116.390 750.025 1116.870 ;
      LAYER li1 ;
        RECT 750.195 1116.560 750.525 1117.040 ;
      LAYER li1 ;
        RECT 750.695 1116.390 750.865 1116.870 ;
      LAYER li1 ;
        RECT 751.035 1116.560 751.365 1117.040 ;
        RECT 751.535 1116.390 751.705 1116.865 ;
        RECT 751.875 1116.560 752.205 1117.040 ;
        RECT 752.375 1116.390 752.545 1116.870 ;
      LAYER li1 ;
        RECT 748.175 1116.220 750.865 1116.390 ;
      LAYER li1 ;
        RECT 751.125 1116.220 752.545 1116.390 ;
        RECT 752.805 1116.315 753.095 1117.040 ;
        RECT 753.655 1116.240 753.985 1117.040 ;
      LAYER li1 ;
        RECT 754.155 1116.390 754.325 1116.870 ;
      LAYER li1 ;
        RECT 754.495 1116.560 754.825 1117.040 ;
      LAYER li1 ;
        RECT 754.995 1116.390 755.165 1116.870 ;
      LAYER li1 ;
        RECT 755.335 1116.560 755.665 1117.040 ;
      LAYER li1 ;
        RECT 755.835 1116.390 756.005 1116.870 ;
      LAYER li1 ;
        RECT 756.175 1116.560 756.505 1117.040 ;
      LAYER li1 ;
        RECT 756.675 1116.390 756.845 1116.870 ;
      LAYER li1 ;
        RECT 757.015 1116.560 757.345 1117.040 ;
        RECT 757.515 1116.390 757.685 1116.865 ;
        RECT 757.855 1116.560 758.185 1117.040 ;
        RECT 758.355 1116.390 758.525 1116.870 ;
      LAYER li1 ;
        RECT 754.155 1116.220 756.845 1116.390 ;
      LAYER li1 ;
        RECT 757.105 1116.220 758.525 1116.390 ;
        RECT 758.785 1116.315 759.075 1117.040 ;
        RECT 759.635 1116.240 759.965 1117.040 ;
        RECT 760.475 1116.560 760.805 1117.040 ;
        RECT 761.315 1116.560 761.645 1117.040 ;
        RECT 762.155 1116.560 762.485 1117.040 ;
        RECT 762.995 1116.560 763.325 1117.040 ;
        RECT 763.495 1116.390 763.665 1116.865 ;
        RECT 763.835 1116.560 764.165 1117.040 ;
        RECT 764.335 1116.390 764.505 1116.870 ;
        RECT 763.085 1116.220 764.505 1116.390 ;
        RECT 764.765 1116.315 765.055 1117.040 ;
        RECT 765.615 1116.240 765.945 1117.040 ;
        RECT 766.455 1116.560 766.785 1117.040 ;
        RECT 767.295 1116.560 767.625 1117.040 ;
        RECT 768.135 1116.560 768.465 1117.040 ;
        RECT 768.975 1116.560 769.305 1117.040 ;
        RECT 769.475 1116.390 769.645 1116.865 ;
        RECT 769.815 1116.560 770.145 1117.040 ;
        RECT 770.315 1116.390 770.485 1116.870 ;
        RECT 769.065 1116.220 770.485 1116.390 ;
        RECT 770.745 1116.315 771.035 1117.040 ;
        RECT 771.595 1116.240 771.925 1117.040 ;
        RECT 772.435 1116.560 772.765 1117.040 ;
        RECT 773.275 1116.560 773.605 1117.040 ;
        RECT 774.115 1116.560 774.445 1117.040 ;
        RECT 774.955 1116.560 775.285 1117.040 ;
        RECT 775.455 1116.390 775.625 1116.865 ;
        RECT 775.795 1116.560 776.125 1117.040 ;
        RECT 776.295 1116.390 776.465 1116.870 ;
        RECT 775.045 1116.220 776.465 1116.390 ;
        RECT 776.725 1116.315 777.015 1117.040 ;
        RECT 777.575 1116.240 777.905 1117.040 ;
        RECT 778.415 1116.560 778.745 1117.040 ;
        RECT 779.255 1116.560 779.585 1117.040 ;
        RECT 780.095 1116.560 780.425 1117.040 ;
        RECT 780.935 1116.560 781.265 1117.040 ;
        RECT 781.435 1116.390 781.605 1116.865 ;
        RECT 781.775 1116.560 782.105 1117.040 ;
        RECT 782.275 1116.390 782.445 1116.870 ;
        RECT 781.025 1116.220 782.445 1116.390 ;
        RECT 782.705 1116.315 782.995 1117.040 ;
        RECT 783.555 1116.240 783.885 1117.040 ;
        RECT 784.395 1116.560 784.725 1117.040 ;
        RECT 785.235 1116.560 785.565 1117.040 ;
        RECT 786.075 1116.560 786.405 1117.040 ;
        RECT 786.915 1116.560 787.245 1117.040 ;
        RECT 787.415 1116.390 787.585 1116.865 ;
        RECT 787.755 1116.560 788.085 1117.040 ;
        RECT 788.255 1116.390 788.425 1116.870 ;
        RECT 787.005 1116.220 788.425 1116.390 ;
        RECT 788.685 1116.315 788.975 1117.040 ;
        RECT 789.535 1116.240 789.865 1117.040 ;
        RECT 790.375 1116.560 790.705 1117.040 ;
        RECT 791.215 1116.560 791.545 1117.040 ;
        RECT 792.055 1116.560 792.385 1117.040 ;
        RECT 792.895 1116.560 793.225 1117.040 ;
        RECT 793.395 1116.390 793.565 1116.865 ;
        RECT 793.735 1116.560 794.065 1117.040 ;
        RECT 794.235 1116.390 794.405 1116.870 ;
        RECT 792.985 1116.220 794.405 1116.390 ;
        RECT 794.665 1116.315 794.955 1117.040 ;
        RECT 1969.085 1116.315 1969.375 1117.040 ;
        RECT 1969.935 1116.240 1970.265 1117.040 ;
      LAYER li1 ;
        RECT 1970.435 1116.390 1970.605 1116.870 ;
      LAYER li1 ;
        RECT 1970.775 1116.560 1971.105 1117.040 ;
      LAYER li1 ;
        RECT 1971.275 1116.390 1971.445 1116.870 ;
      LAYER li1 ;
        RECT 1971.615 1116.560 1971.945 1117.040 ;
      LAYER li1 ;
        RECT 1972.115 1116.390 1972.285 1116.870 ;
      LAYER li1 ;
        RECT 1972.455 1116.560 1972.785 1117.040 ;
      LAYER li1 ;
        RECT 1972.955 1116.390 1973.125 1116.870 ;
      LAYER li1 ;
        RECT 1973.295 1116.560 1973.625 1117.040 ;
        RECT 1973.795 1116.390 1973.965 1116.865 ;
        RECT 1974.135 1116.560 1974.465 1117.040 ;
        RECT 1974.635 1116.390 1974.805 1116.870 ;
      LAYER li1 ;
        RECT 1970.435 1116.220 1973.125 1116.390 ;
      LAYER li1 ;
        RECT 1973.385 1116.220 1974.805 1116.390 ;
        RECT 1975.065 1116.315 1975.355 1117.040 ;
        RECT 1975.915 1116.240 1976.245 1117.040 ;
      LAYER li1 ;
        RECT 1976.415 1116.390 1976.585 1116.870 ;
      LAYER li1 ;
        RECT 1976.755 1116.560 1977.085 1117.040 ;
      LAYER li1 ;
        RECT 1977.255 1116.390 1977.425 1116.870 ;
      LAYER li1 ;
        RECT 1977.595 1116.560 1977.925 1117.040 ;
      LAYER li1 ;
        RECT 1978.095 1116.390 1978.265 1116.870 ;
      LAYER li1 ;
        RECT 1978.435 1116.560 1978.765 1117.040 ;
      LAYER li1 ;
        RECT 1978.935 1116.390 1979.105 1116.870 ;
      LAYER li1 ;
        RECT 1979.275 1116.560 1979.605 1117.040 ;
        RECT 1979.775 1116.390 1979.945 1116.865 ;
        RECT 1980.115 1116.560 1980.445 1117.040 ;
        RECT 1980.615 1116.390 1980.785 1116.870 ;
      LAYER li1 ;
        RECT 1976.415 1116.220 1979.105 1116.390 ;
      LAYER li1 ;
        RECT 1979.365 1116.220 1980.785 1116.390 ;
        RECT 1981.045 1116.315 1981.335 1117.040 ;
        RECT 1981.895 1116.240 1982.225 1117.040 ;
      LAYER li1 ;
        RECT 1982.395 1116.390 1982.565 1116.870 ;
      LAYER li1 ;
        RECT 1982.735 1116.560 1983.065 1117.040 ;
      LAYER li1 ;
        RECT 1983.235 1116.390 1983.405 1116.870 ;
      LAYER li1 ;
        RECT 1983.575 1116.560 1983.905 1117.040 ;
      LAYER li1 ;
        RECT 1984.075 1116.390 1984.245 1116.870 ;
      LAYER li1 ;
        RECT 1984.415 1116.560 1984.745 1117.040 ;
      LAYER li1 ;
        RECT 1984.915 1116.390 1985.085 1116.870 ;
      LAYER li1 ;
        RECT 1985.255 1116.560 1985.585 1117.040 ;
        RECT 1985.755 1116.390 1985.925 1116.865 ;
        RECT 1986.095 1116.560 1986.425 1117.040 ;
        RECT 1986.595 1116.390 1986.765 1116.870 ;
      LAYER li1 ;
        RECT 1982.395 1116.220 1985.085 1116.390 ;
      LAYER li1 ;
        RECT 1985.345 1116.220 1986.765 1116.390 ;
        RECT 1987.025 1116.315 1987.315 1117.040 ;
        RECT 1987.875 1116.240 1988.205 1117.040 ;
      LAYER li1 ;
        RECT 1988.375 1116.390 1988.545 1116.870 ;
      LAYER li1 ;
        RECT 1988.715 1116.560 1989.045 1117.040 ;
      LAYER li1 ;
        RECT 1989.215 1116.390 1989.385 1116.870 ;
      LAYER li1 ;
        RECT 1989.555 1116.560 1989.885 1117.040 ;
      LAYER li1 ;
        RECT 1990.055 1116.390 1990.225 1116.870 ;
      LAYER li1 ;
        RECT 1990.395 1116.560 1990.725 1117.040 ;
      LAYER li1 ;
        RECT 1990.895 1116.390 1991.065 1116.870 ;
      LAYER li1 ;
        RECT 1991.235 1116.560 1991.565 1117.040 ;
        RECT 1991.735 1116.390 1991.905 1116.865 ;
        RECT 1992.075 1116.560 1992.405 1117.040 ;
        RECT 1992.575 1116.390 1992.745 1116.870 ;
      LAYER li1 ;
        RECT 1988.375 1116.220 1991.065 1116.390 ;
      LAYER li1 ;
        RECT 1991.325 1116.220 1992.745 1116.390 ;
        RECT 1993.005 1116.315 1993.295 1117.040 ;
        RECT 1993.855 1116.240 1994.185 1117.040 ;
      LAYER li1 ;
        RECT 1994.355 1116.390 1994.525 1116.870 ;
      LAYER li1 ;
        RECT 1994.695 1116.560 1995.025 1117.040 ;
      LAYER li1 ;
        RECT 1995.195 1116.390 1995.365 1116.870 ;
      LAYER li1 ;
        RECT 1995.535 1116.560 1995.865 1117.040 ;
      LAYER li1 ;
        RECT 1996.035 1116.390 1996.205 1116.870 ;
      LAYER li1 ;
        RECT 1996.375 1116.560 1996.705 1117.040 ;
      LAYER li1 ;
        RECT 1996.875 1116.390 1997.045 1116.870 ;
      LAYER li1 ;
        RECT 1997.215 1116.560 1997.545 1117.040 ;
        RECT 1997.715 1116.390 1997.885 1116.865 ;
        RECT 1998.055 1116.560 1998.385 1117.040 ;
        RECT 1998.555 1116.390 1998.725 1116.870 ;
      LAYER li1 ;
        RECT 1994.355 1116.220 1997.045 1116.390 ;
      LAYER li1 ;
        RECT 1997.305 1116.220 1998.725 1116.390 ;
        RECT 1998.985 1116.315 1999.275 1117.040 ;
        RECT 1999.835 1116.240 2000.165 1117.040 ;
      LAYER li1 ;
        RECT 2000.335 1116.390 2000.505 1116.870 ;
      LAYER li1 ;
        RECT 2000.675 1116.560 2001.005 1117.040 ;
      LAYER li1 ;
        RECT 2001.175 1116.390 2001.345 1116.870 ;
      LAYER li1 ;
        RECT 2001.515 1116.560 2001.845 1117.040 ;
      LAYER li1 ;
        RECT 2002.015 1116.390 2002.185 1116.870 ;
      LAYER li1 ;
        RECT 2002.355 1116.560 2002.685 1117.040 ;
      LAYER li1 ;
        RECT 2002.855 1116.390 2003.025 1116.870 ;
      LAYER li1 ;
        RECT 2003.195 1116.560 2003.525 1117.040 ;
        RECT 2003.695 1116.390 2003.865 1116.865 ;
        RECT 2004.035 1116.560 2004.365 1117.040 ;
        RECT 2004.535 1116.390 2004.705 1116.870 ;
      LAYER li1 ;
        RECT 2000.335 1116.220 2003.025 1116.390 ;
      LAYER li1 ;
        RECT 2003.285 1116.220 2004.705 1116.390 ;
        RECT 2004.965 1116.315 2005.255 1117.040 ;
        RECT 2005.815 1116.240 2006.145 1117.040 ;
      LAYER li1 ;
        RECT 2006.315 1116.390 2006.485 1116.870 ;
      LAYER li1 ;
        RECT 2006.655 1116.560 2006.985 1117.040 ;
      LAYER li1 ;
        RECT 2007.155 1116.390 2007.325 1116.870 ;
      LAYER li1 ;
        RECT 2007.495 1116.560 2007.825 1117.040 ;
      LAYER li1 ;
        RECT 2007.995 1116.390 2008.165 1116.870 ;
      LAYER li1 ;
        RECT 2008.335 1116.560 2008.665 1117.040 ;
      LAYER li1 ;
        RECT 2008.835 1116.390 2009.005 1116.870 ;
      LAYER li1 ;
        RECT 2009.175 1116.560 2009.505 1117.040 ;
        RECT 2009.675 1116.390 2009.845 1116.865 ;
        RECT 2010.015 1116.560 2010.345 1117.040 ;
        RECT 2010.515 1116.390 2010.685 1116.870 ;
      LAYER li1 ;
        RECT 2006.315 1116.220 2009.005 1116.390 ;
      LAYER li1 ;
        RECT 2009.265 1116.220 2010.685 1116.390 ;
        RECT 2010.945 1116.315 2011.235 1117.040 ;
        RECT 2011.795 1116.240 2012.125 1117.040 ;
      LAYER li1 ;
        RECT 2012.295 1116.390 2012.465 1116.870 ;
      LAYER li1 ;
        RECT 2012.635 1116.560 2012.965 1117.040 ;
      LAYER li1 ;
        RECT 2013.135 1116.390 2013.305 1116.870 ;
      LAYER li1 ;
        RECT 2013.475 1116.560 2013.805 1117.040 ;
      LAYER li1 ;
        RECT 2013.975 1116.390 2014.145 1116.870 ;
      LAYER li1 ;
        RECT 2014.315 1116.560 2014.645 1117.040 ;
      LAYER li1 ;
        RECT 2014.815 1116.390 2014.985 1116.870 ;
      LAYER li1 ;
        RECT 2015.155 1116.560 2015.485 1117.040 ;
        RECT 2015.655 1116.390 2015.825 1116.865 ;
        RECT 2015.995 1116.560 2016.325 1117.040 ;
        RECT 2016.495 1116.390 2016.665 1116.870 ;
      LAYER li1 ;
        RECT 2012.295 1116.220 2014.985 1116.390 ;
      LAYER li1 ;
        RECT 2015.245 1116.220 2016.665 1116.390 ;
        RECT 2016.925 1116.315 2017.215 1117.040 ;
        RECT 2017.775 1116.240 2018.105 1117.040 ;
      LAYER li1 ;
        RECT 2018.275 1116.390 2018.445 1116.870 ;
      LAYER li1 ;
        RECT 2018.615 1116.560 2018.945 1117.040 ;
      LAYER li1 ;
        RECT 2019.115 1116.390 2019.285 1116.870 ;
      LAYER li1 ;
        RECT 2019.455 1116.560 2019.785 1117.040 ;
      LAYER li1 ;
        RECT 2019.955 1116.390 2020.125 1116.870 ;
      LAYER li1 ;
        RECT 2020.295 1116.560 2020.625 1117.040 ;
      LAYER li1 ;
        RECT 2020.795 1116.390 2020.965 1116.870 ;
      LAYER li1 ;
        RECT 2021.135 1116.560 2021.465 1117.040 ;
        RECT 2021.635 1116.390 2021.805 1116.865 ;
        RECT 2021.975 1116.560 2022.305 1117.040 ;
        RECT 2022.475 1116.390 2022.645 1116.870 ;
      LAYER li1 ;
        RECT 2018.275 1116.220 2020.965 1116.390 ;
      LAYER li1 ;
        RECT 2021.225 1116.220 2022.645 1116.390 ;
        RECT 2022.905 1116.315 2023.195 1117.040 ;
        RECT 2023.755 1116.240 2024.085 1117.040 ;
      LAYER li1 ;
        RECT 2024.255 1116.390 2024.425 1116.870 ;
      LAYER li1 ;
        RECT 2024.595 1116.560 2024.925 1117.040 ;
      LAYER li1 ;
        RECT 2025.095 1116.390 2025.265 1116.870 ;
      LAYER li1 ;
        RECT 2025.435 1116.560 2025.765 1117.040 ;
      LAYER li1 ;
        RECT 2025.935 1116.390 2026.105 1116.870 ;
      LAYER li1 ;
        RECT 2026.275 1116.560 2026.605 1117.040 ;
      LAYER li1 ;
        RECT 2026.775 1116.390 2026.945 1116.870 ;
      LAYER li1 ;
        RECT 2027.115 1116.560 2027.445 1117.040 ;
        RECT 2027.615 1116.390 2027.785 1116.865 ;
        RECT 2027.955 1116.560 2028.285 1117.040 ;
        RECT 2028.455 1116.390 2028.625 1116.870 ;
      LAYER li1 ;
        RECT 2024.255 1116.220 2026.945 1116.390 ;
      LAYER li1 ;
        RECT 2027.205 1116.220 2028.625 1116.390 ;
        RECT 2028.885 1116.315 2029.175 1117.040 ;
        RECT 2029.735 1116.240 2030.065 1117.040 ;
      LAYER li1 ;
        RECT 2030.235 1116.390 2030.405 1116.870 ;
      LAYER li1 ;
        RECT 2030.575 1116.560 2030.905 1117.040 ;
      LAYER li1 ;
        RECT 2031.075 1116.390 2031.245 1116.870 ;
      LAYER li1 ;
        RECT 2031.415 1116.560 2031.745 1117.040 ;
      LAYER li1 ;
        RECT 2031.915 1116.390 2032.085 1116.870 ;
      LAYER li1 ;
        RECT 2032.255 1116.560 2032.585 1117.040 ;
      LAYER li1 ;
        RECT 2032.755 1116.390 2032.925 1116.870 ;
      LAYER li1 ;
        RECT 2033.095 1116.560 2033.425 1117.040 ;
        RECT 2033.595 1116.390 2033.765 1116.865 ;
        RECT 2033.935 1116.560 2034.265 1117.040 ;
        RECT 2034.435 1116.390 2034.605 1116.870 ;
      LAYER li1 ;
        RECT 2030.235 1116.220 2032.925 1116.390 ;
      LAYER li1 ;
        RECT 2033.185 1116.220 2034.605 1116.390 ;
        RECT 2034.865 1116.315 2035.155 1117.040 ;
        RECT 2035.715 1116.240 2036.045 1117.040 ;
      LAYER li1 ;
        RECT 2036.215 1116.390 2036.385 1116.870 ;
      LAYER li1 ;
        RECT 2036.555 1116.560 2036.885 1117.040 ;
      LAYER li1 ;
        RECT 2037.055 1116.390 2037.225 1116.870 ;
      LAYER li1 ;
        RECT 2037.395 1116.560 2037.725 1117.040 ;
      LAYER li1 ;
        RECT 2037.895 1116.390 2038.065 1116.870 ;
      LAYER li1 ;
        RECT 2038.235 1116.560 2038.565 1117.040 ;
      LAYER li1 ;
        RECT 2038.735 1116.390 2038.905 1116.870 ;
      LAYER li1 ;
        RECT 2039.075 1116.560 2039.405 1117.040 ;
        RECT 2039.575 1116.390 2039.745 1116.865 ;
        RECT 2039.915 1116.560 2040.245 1117.040 ;
        RECT 2040.415 1116.390 2040.585 1116.870 ;
      LAYER li1 ;
        RECT 2036.215 1116.220 2038.905 1116.390 ;
      LAYER li1 ;
        RECT 2039.165 1116.220 2040.585 1116.390 ;
        RECT 2040.845 1116.315 2041.135 1117.040 ;
        RECT 2041.695 1116.240 2042.025 1117.040 ;
      LAYER li1 ;
        RECT 2042.195 1116.390 2042.365 1116.870 ;
      LAYER li1 ;
        RECT 2042.535 1116.560 2042.865 1117.040 ;
      LAYER li1 ;
        RECT 2043.035 1116.390 2043.205 1116.870 ;
      LAYER li1 ;
        RECT 2043.375 1116.560 2043.705 1117.040 ;
      LAYER li1 ;
        RECT 2043.875 1116.390 2044.045 1116.870 ;
      LAYER li1 ;
        RECT 2044.215 1116.560 2044.545 1117.040 ;
      LAYER li1 ;
        RECT 2044.715 1116.390 2044.885 1116.870 ;
      LAYER li1 ;
        RECT 2045.055 1116.560 2045.385 1117.040 ;
        RECT 2045.555 1116.390 2045.725 1116.865 ;
        RECT 2045.895 1116.560 2046.225 1117.040 ;
        RECT 2046.395 1116.390 2046.565 1116.870 ;
      LAYER li1 ;
        RECT 2042.195 1116.220 2044.885 1116.390 ;
      LAYER li1 ;
        RECT 2045.145 1116.220 2046.565 1116.390 ;
        RECT 2046.825 1116.315 2047.115 1117.040 ;
        RECT 2047.675 1116.240 2048.005 1117.040 ;
      LAYER li1 ;
        RECT 2048.175 1116.390 2048.345 1116.870 ;
      LAYER li1 ;
        RECT 2048.515 1116.560 2048.845 1117.040 ;
      LAYER li1 ;
        RECT 2049.015 1116.390 2049.185 1116.870 ;
      LAYER li1 ;
        RECT 2049.355 1116.560 2049.685 1117.040 ;
      LAYER li1 ;
        RECT 2049.855 1116.390 2050.025 1116.870 ;
      LAYER li1 ;
        RECT 2050.195 1116.560 2050.525 1117.040 ;
      LAYER li1 ;
        RECT 2050.695 1116.390 2050.865 1116.870 ;
      LAYER li1 ;
        RECT 2051.035 1116.560 2051.365 1117.040 ;
        RECT 2051.535 1116.390 2051.705 1116.865 ;
        RECT 2051.875 1116.560 2052.205 1117.040 ;
        RECT 2052.375 1116.390 2052.545 1116.870 ;
      LAYER li1 ;
        RECT 2048.175 1116.220 2050.865 1116.390 ;
      LAYER li1 ;
        RECT 2051.125 1116.220 2052.545 1116.390 ;
        RECT 2052.805 1116.315 2053.095 1117.040 ;
        RECT 2053.655 1116.240 2053.985 1117.040 ;
      LAYER li1 ;
        RECT 2054.155 1116.390 2054.325 1116.870 ;
      LAYER li1 ;
        RECT 2054.495 1116.560 2054.825 1117.040 ;
      LAYER li1 ;
        RECT 2054.995 1116.390 2055.165 1116.870 ;
      LAYER li1 ;
        RECT 2055.335 1116.560 2055.665 1117.040 ;
      LAYER li1 ;
        RECT 2055.835 1116.390 2056.005 1116.870 ;
      LAYER li1 ;
        RECT 2056.175 1116.560 2056.505 1117.040 ;
      LAYER li1 ;
        RECT 2056.675 1116.390 2056.845 1116.870 ;
      LAYER li1 ;
        RECT 2057.015 1116.560 2057.345 1117.040 ;
        RECT 2057.515 1116.390 2057.685 1116.865 ;
        RECT 2057.855 1116.560 2058.185 1117.040 ;
        RECT 2058.355 1116.390 2058.525 1116.870 ;
      LAYER li1 ;
        RECT 2054.155 1116.220 2056.845 1116.390 ;
      LAYER li1 ;
        RECT 2057.105 1116.220 2058.525 1116.390 ;
        RECT 2058.785 1116.315 2059.075 1117.040 ;
        RECT 2059.635 1116.240 2059.965 1117.040 ;
      LAYER li1 ;
        RECT 2060.135 1116.390 2060.305 1116.870 ;
      LAYER li1 ;
        RECT 2060.475 1116.560 2060.805 1117.040 ;
      LAYER li1 ;
        RECT 2060.975 1116.390 2061.145 1116.870 ;
      LAYER li1 ;
        RECT 2061.315 1116.560 2061.645 1117.040 ;
      LAYER li1 ;
        RECT 2061.815 1116.390 2061.985 1116.870 ;
      LAYER li1 ;
        RECT 2062.155 1116.560 2062.485 1117.040 ;
      LAYER li1 ;
        RECT 2062.655 1116.390 2062.825 1116.870 ;
      LAYER li1 ;
        RECT 2062.995 1116.560 2063.325 1117.040 ;
        RECT 2063.495 1116.390 2063.665 1116.865 ;
        RECT 2063.835 1116.560 2064.165 1117.040 ;
        RECT 2064.335 1116.390 2064.505 1116.870 ;
      LAYER li1 ;
        RECT 2060.135 1116.220 2062.825 1116.390 ;
      LAYER li1 ;
        RECT 2063.085 1116.220 2064.505 1116.390 ;
        RECT 2064.765 1116.315 2065.055 1117.040 ;
        RECT 2065.615 1116.240 2065.945 1117.040 ;
      LAYER li1 ;
        RECT 2066.115 1116.390 2066.285 1116.870 ;
      LAYER li1 ;
        RECT 2066.455 1116.560 2066.785 1117.040 ;
      LAYER li1 ;
        RECT 2066.955 1116.390 2067.125 1116.870 ;
      LAYER li1 ;
        RECT 2067.295 1116.560 2067.625 1117.040 ;
      LAYER li1 ;
        RECT 2067.795 1116.390 2067.965 1116.870 ;
      LAYER li1 ;
        RECT 2068.135 1116.560 2068.465 1117.040 ;
      LAYER li1 ;
        RECT 2068.635 1116.390 2068.805 1116.870 ;
      LAYER li1 ;
        RECT 2068.975 1116.560 2069.305 1117.040 ;
        RECT 2069.475 1116.390 2069.645 1116.865 ;
        RECT 2069.815 1116.560 2070.145 1117.040 ;
        RECT 2070.315 1116.390 2070.485 1116.870 ;
      LAYER li1 ;
        RECT 2066.115 1116.220 2068.805 1116.390 ;
      LAYER li1 ;
        RECT 2069.065 1116.220 2070.485 1116.390 ;
        RECT 2070.745 1116.315 2071.035 1117.040 ;
        RECT 2071.595 1116.240 2071.925 1117.040 ;
      LAYER li1 ;
        RECT 2072.095 1116.390 2072.265 1116.870 ;
      LAYER li1 ;
        RECT 2072.435 1116.560 2072.765 1117.040 ;
      LAYER li1 ;
        RECT 2072.935 1116.390 2073.105 1116.870 ;
      LAYER li1 ;
        RECT 2073.275 1116.560 2073.605 1117.040 ;
      LAYER li1 ;
        RECT 2073.775 1116.390 2073.945 1116.870 ;
      LAYER li1 ;
        RECT 2074.115 1116.560 2074.445 1117.040 ;
      LAYER li1 ;
        RECT 2074.615 1116.390 2074.785 1116.870 ;
      LAYER li1 ;
        RECT 2074.955 1116.560 2075.285 1117.040 ;
        RECT 2075.455 1116.390 2075.625 1116.865 ;
        RECT 2075.795 1116.560 2076.125 1117.040 ;
        RECT 2076.295 1116.390 2076.465 1116.870 ;
      LAYER li1 ;
        RECT 2072.095 1116.220 2074.785 1116.390 ;
      LAYER li1 ;
        RECT 2075.045 1116.220 2076.465 1116.390 ;
        RECT 2076.725 1116.315 2077.015 1117.040 ;
        RECT 2077.575 1116.240 2077.905 1117.040 ;
      LAYER li1 ;
        RECT 2078.075 1116.390 2078.245 1116.870 ;
      LAYER li1 ;
        RECT 2078.415 1116.560 2078.745 1117.040 ;
      LAYER li1 ;
        RECT 2078.915 1116.390 2079.085 1116.870 ;
      LAYER li1 ;
        RECT 2079.255 1116.560 2079.585 1117.040 ;
      LAYER li1 ;
        RECT 2079.755 1116.390 2079.925 1116.870 ;
      LAYER li1 ;
        RECT 2080.095 1116.560 2080.425 1117.040 ;
      LAYER li1 ;
        RECT 2080.595 1116.390 2080.765 1116.870 ;
      LAYER li1 ;
        RECT 2080.935 1116.560 2081.265 1117.040 ;
        RECT 2081.435 1116.390 2081.605 1116.865 ;
        RECT 2081.775 1116.560 2082.105 1117.040 ;
        RECT 2082.275 1116.390 2082.445 1116.870 ;
      LAYER li1 ;
        RECT 2078.075 1116.220 2080.765 1116.390 ;
      LAYER li1 ;
        RECT 2081.025 1116.220 2082.445 1116.390 ;
        RECT 2082.705 1116.315 2082.995 1117.040 ;
        RECT 2083.555 1116.240 2083.885 1117.040 ;
      LAYER li1 ;
        RECT 2084.055 1116.390 2084.225 1116.870 ;
      LAYER li1 ;
        RECT 2084.395 1116.560 2084.725 1117.040 ;
      LAYER li1 ;
        RECT 2084.895 1116.390 2085.065 1116.870 ;
      LAYER li1 ;
        RECT 2085.235 1116.560 2085.565 1117.040 ;
      LAYER li1 ;
        RECT 2085.735 1116.390 2085.905 1116.870 ;
      LAYER li1 ;
        RECT 2086.075 1116.560 2086.405 1117.040 ;
      LAYER li1 ;
        RECT 2086.575 1116.390 2086.745 1116.870 ;
      LAYER li1 ;
        RECT 2086.915 1116.560 2087.245 1117.040 ;
        RECT 2087.415 1116.390 2087.585 1116.865 ;
        RECT 2087.755 1116.560 2088.085 1117.040 ;
        RECT 2088.255 1116.390 2088.425 1116.870 ;
      LAYER li1 ;
        RECT 2084.055 1116.220 2086.745 1116.390 ;
      LAYER li1 ;
        RECT 2087.005 1116.220 2088.425 1116.390 ;
        RECT 2088.685 1116.315 2088.975 1117.040 ;
        RECT 2089.535 1116.240 2089.865 1117.040 ;
      LAYER li1 ;
        RECT 2090.035 1116.390 2090.205 1116.870 ;
      LAYER li1 ;
        RECT 2090.375 1116.560 2090.705 1117.040 ;
      LAYER li1 ;
        RECT 2090.875 1116.390 2091.045 1116.870 ;
      LAYER li1 ;
        RECT 2091.215 1116.560 2091.545 1117.040 ;
      LAYER li1 ;
        RECT 2091.715 1116.390 2091.885 1116.870 ;
      LAYER li1 ;
        RECT 2092.055 1116.560 2092.385 1117.040 ;
      LAYER li1 ;
        RECT 2092.555 1116.390 2092.725 1116.870 ;
      LAYER li1 ;
        RECT 2092.895 1116.560 2093.225 1117.040 ;
        RECT 2093.395 1116.390 2093.565 1116.865 ;
        RECT 2093.735 1116.560 2094.065 1117.040 ;
        RECT 2094.235 1116.390 2094.405 1116.870 ;
      LAYER li1 ;
        RECT 2090.035 1116.220 2092.725 1116.390 ;
      LAYER li1 ;
        RECT 2092.985 1116.220 2094.405 1116.390 ;
        RECT 2094.665 1116.315 2094.955 1117.040 ;
      LAYER li1 ;
        RECT 670.435 1115.680 670.690 1116.220 ;
      LAYER li1 ;
        RECT 673.385 1116.050 673.560 1116.220 ;
        RECT 670.935 1115.880 673.560 1116.050 ;
        RECT 673.385 1115.680 673.560 1115.880 ;
      LAYER li1 ;
        RECT 673.740 1115.850 675.330 1116.050 ;
        RECT 676.415 1115.680 676.670 1116.220 ;
      LAYER li1 ;
        RECT 679.365 1116.050 679.540 1116.220 ;
        RECT 676.915 1115.880 679.540 1116.050 ;
        RECT 679.365 1115.680 679.540 1115.880 ;
      LAYER li1 ;
        RECT 679.720 1115.850 681.310 1116.050 ;
        RECT 682.395 1115.680 682.650 1116.220 ;
      LAYER li1 ;
        RECT 685.345 1116.050 685.520 1116.220 ;
        RECT 682.895 1115.880 685.520 1116.050 ;
        RECT 685.345 1115.680 685.520 1115.880 ;
      LAYER li1 ;
        RECT 685.700 1115.850 687.290 1116.050 ;
        RECT 688.375 1115.680 688.630 1116.220 ;
      LAYER li1 ;
        RECT 691.325 1116.050 691.500 1116.220 ;
        RECT 688.875 1115.880 691.500 1116.050 ;
        RECT 691.325 1115.680 691.500 1115.880 ;
      LAYER li1 ;
        RECT 691.680 1115.850 693.270 1116.050 ;
        RECT 694.355 1115.680 694.610 1116.220 ;
      LAYER li1 ;
        RECT 697.305 1116.050 697.480 1116.220 ;
        RECT 694.855 1115.880 697.480 1116.050 ;
        RECT 697.305 1115.680 697.480 1115.880 ;
      LAYER li1 ;
        RECT 697.660 1115.850 699.250 1116.050 ;
        RECT 700.335 1115.680 700.590 1116.220 ;
      LAYER li1 ;
        RECT 703.285 1116.050 703.460 1116.220 ;
        RECT 700.835 1115.880 703.460 1116.050 ;
        RECT 703.285 1115.680 703.460 1115.880 ;
      LAYER li1 ;
        RECT 703.640 1115.850 705.230 1116.050 ;
        RECT 706.315 1115.680 706.570 1116.220 ;
      LAYER li1 ;
        RECT 709.265 1116.050 709.440 1116.220 ;
        RECT 706.815 1115.880 709.440 1116.050 ;
        RECT 709.265 1115.680 709.440 1115.880 ;
      LAYER li1 ;
        RECT 709.620 1115.850 711.210 1116.050 ;
        RECT 712.295 1115.680 712.550 1116.220 ;
      LAYER li1 ;
        RECT 715.245 1116.050 715.420 1116.220 ;
        RECT 712.795 1115.880 715.420 1116.050 ;
        RECT 715.245 1115.680 715.420 1115.880 ;
      LAYER li1 ;
        RECT 715.600 1115.850 717.190 1116.050 ;
        RECT 718.275 1115.680 718.530 1116.220 ;
      LAYER li1 ;
        RECT 721.225 1116.050 721.400 1116.220 ;
        RECT 718.775 1115.880 721.400 1116.050 ;
        RECT 721.225 1115.680 721.400 1115.880 ;
      LAYER li1 ;
        RECT 721.580 1115.850 723.170 1116.050 ;
        RECT 724.255 1115.680 724.510 1116.220 ;
      LAYER li1 ;
        RECT 727.205 1116.050 727.380 1116.220 ;
        RECT 724.755 1115.880 727.380 1116.050 ;
        RECT 727.205 1115.680 727.380 1115.880 ;
      LAYER li1 ;
        RECT 727.560 1115.850 729.150 1116.050 ;
        RECT 730.235 1115.680 730.490 1116.220 ;
      LAYER li1 ;
        RECT 733.185 1116.050 733.360 1116.220 ;
        RECT 730.735 1115.880 733.360 1116.050 ;
        RECT 733.185 1115.680 733.360 1115.880 ;
      LAYER li1 ;
        RECT 733.540 1115.850 735.130 1116.050 ;
        RECT 736.215 1115.680 736.470 1116.220 ;
      LAYER li1 ;
        RECT 739.165 1116.050 739.340 1116.220 ;
        RECT 736.715 1115.880 739.340 1116.050 ;
        RECT 739.165 1115.680 739.340 1115.880 ;
      LAYER li1 ;
        RECT 739.520 1115.850 741.110 1116.050 ;
        RECT 742.195 1115.680 742.450 1116.220 ;
      LAYER li1 ;
        RECT 745.145 1116.050 745.320 1116.220 ;
        RECT 742.695 1115.880 745.320 1116.050 ;
        RECT 745.145 1115.680 745.320 1115.880 ;
      LAYER li1 ;
        RECT 745.500 1115.850 747.090 1116.050 ;
        RECT 748.175 1115.680 748.430 1116.220 ;
      LAYER li1 ;
        RECT 751.125 1116.050 751.300 1116.220 ;
        RECT 748.675 1115.880 751.300 1116.050 ;
        RECT 751.125 1115.680 751.300 1115.880 ;
      LAYER li1 ;
        RECT 751.480 1115.850 753.070 1116.050 ;
        RECT 754.155 1115.680 754.410 1116.220 ;
      LAYER li1 ;
        RECT 757.105 1116.050 757.280 1116.220 ;
        RECT 763.085 1116.050 763.260 1116.220 ;
        RECT 769.065 1116.050 769.240 1116.220 ;
        RECT 775.045 1116.050 775.220 1116.220 ;
        RECT 781.025 1116.050 781.200 1116.220 ;
        RECT 787.005 1116.050 787.180 1116.220 ;
        RECT 792.985 1116.050 793.160 1116.220 ;
        RECT 754.655 1115.880 757.280 1116.050 ;
        RECT 757.105 1115.680 757.280 1115.880 ;
      LAYER li1 ;
        RECT 757.460 1115.850 759.050 1116.050 ;
      LAYER li1 ;
        RECT 760.635 1115.880 763.260 1116.050 ;
        RECT 763.085 1115.680 763.260 1115.880 ;
      LAYER li1 ;
        RECT 763.440 1115.850 765.030 1116.050 ;
      LAYER li1 ;
        RECT 766.615 1115.880 769.240 1116.050 ;
        RECT 769.065 1115.680 769.240 1115.880 ;
      LAYER li1 ;
        RECT 769.420 1115.850 771.010 1116.050 ;
      LAYER li1 ;
        RECT 772.595 1115.880 775.220 1116.050 ;
        RECT 775.045 1115.680 775.220 1115.880 ;
      LAYER li1 ;
        RECT 775.400 1115.850 776.990 1116.050 ;
      LAYER li1 ;
        RECT 778.575 1115.880 781.200 1116.050 ;
        RECT 781.025 1115.680 781.200 1115.880 ;
      LAYER li1 ;
        RECT 781.380 1115.850 782.970 1116.050 ;
      LAYER li1 ;
        RECT 784.555 1115.880 787.180 1116.050 ;
        RECT 787.005 1115.680 787.180 1115.880 ;
      LAYER li1 ;
        RECT 787.360 1115.850 788.950 1116.050 ;
      LAYER li1 ;
        RECT 790.535 1115.880 793.160 1116.050 ;
        RECT 792.985 1115.680 793.160 1115.880 ;
      LAYER li1 ;
        RECT 793.340 1115.850 794.930 1116.050 ;
        RECT 1970.435 1115.680 1970.690 1116.220 ;
      LAYER li1 ;
        RECT 1973.385 1116.050 1973.560 1116.220 ;
        RECT 1970.935 1115.880 1973.560 1116.050 ;
        RECT 1973.385 1115.680 1973.560 1115.880 ;
      LAYER li1 ;
        RECT 1976.415 1115.680 1976.670 1116.220 ;
      LAYER li1 ;
        RECT 1979.365 1116.050 1979.540 1116.220 ;
        RECT 1976.915 1115.880 1979.540 1116.050 ;
        RECT 1979.365 1115.680 1979.540 1115.880 ;
      LAYER li1 ;
        RECT 1982.395 1115.680 1982.650 1116.220 ;
      LAYER li1 ;
        RECT 1985.345 1116.050 1985.520 1116.220 ;
        RECT 1982.895 1115.880 1985.520 1116.050 ;
        RECT 1985.345 1115.680 1985.520 1115.880 ;
      LAYER li1 ;
        RECT 1988.375 1115.680 1988.630 1116.220 ;
      LAYER li1 ;
        RECT 1991.325 1116.050 1991.500 1116.220 ;
        RECT 1988.875 1115.880 1991.500 1116.050 ;
        RECT 1991.325 1115.680 1991.500 1115.880 ;
      LAYER li1 ;
        RECT 1994.355 1115.680 1994.610 1116.220 ;
      LAYER li1 ;
        RECT 1997.305 1116.050 1997.480 1116.220 ;
        RECT 1994.855 1115.880 1997.480 1116.050 ;
        RECT 1997.305 1115.680 1997.480 1115.880 ;
      LAYER li1 ;
        RECT 2000.335 1115.680 2000.590 1116.220 ;
      LAYER li1 ;
        RECT 2003.285 1116.050 2003.460 1116.220 ;
        RECT 2000.835 1115.880 2003.460 1116.050 ;
        RECT 2003.285 1115.680 2003.460 1115.880 ;
      LAYER li1 ;
        RECT 2006.315 1115.680 2006.570 1116.220 ;
      LAYER li1 ;
        RECT 2009.265 1116.050 2009.440 1116.220 ;
        RECT 2006.815 1115.880 2009.440 1116.050 ;
        RECT 2009.265 1115.680 2009.440 1115.880 ;
      LAYER li1 ;
        RECT 2012.295 1115.680 2012.550 1116.220 ;
      LAYER li1 ;
        RECT 2015.245 1116.050 2015.420 1116.220 ;
        RECT 2012.795 1115.880 2015.420 1116.050 ;
        RECT 2015.245 1115.680 2015.420 1115.880 ;
      LAYER li1 ;
        RECT 2018.275 1115.680 2018.530 1116.220 ;
      LAYER li1 ;
        RECT 2021.225 1116.050 2021.400 1116.220 ;
        RECT 2018.775 1115.880 2021.400 1116.050 ;
        RECT 2021.225 1115.680 2021.400 1115.880 ;
      LAYER li1 ;
        RECT 2024.255 1115.680 2024.510 1116.220 ;
      LAYER li1 ;
        RECT 2027.205 1116.050 2027.380 1116.220 ;
        RECT 2024.755 1115.880 2027.380 1116.050 ;
        RECT 2027.205 1115.680 2027.380 1115.880 ;
      LAYER li1 ;
        RECT 2030.235 1115.680 2030.490 1116.220 ;
      LAYER li1 ;
        RECT 2033.185 1116.050 2033.360 1116.220 ;
        RECT 2030.735 1115.880 2033.360 1116.050 ;
        RECT 2033.185 1115.680 2033.360 1115.880 ;
      LAYER li1 ;
        RECT 2036.215 1115.680 2036.470 1116.220 ;
      LAYER li1 ;
        RECT 2039.165 1116.050 2039.340 1116.220 ;
        RECT 2036.715 1115.880 2039.340 1116.050 ;
        RECT 2039.165 1115.680 2039.340 1115.880 ;
      LAYER li1 ;
        RECT 2042.195 1115.680 2042.450 1116.220 ;
      LAYER li1 ;
        RECT 2045.145 1116.050 2045.320 1116.220 ;
        RECT 2042.695 1115.880 2045.320 1116.050 ;
        RECT 2045.145 1115.680 2045.320 1115.880 ;
      LAYER li1 ;
        RECT 2048.175 1115.680 2048.430 1116.220 ;
      LAYER li1 ;
        RECT 2051.125 1116.050 2051.300 1116.220 ;
        RECT 2048.675 1115.880 2051.300 1116.050 ;
        RECT 2051.125 1115.680 2051.300 1115.880 ;
      LAYER li1 ;
        RECT 2054.155 1115.680 2054.410 1116.220 ;
      LAYER li1 ;
        RECT 2057.105 1116.050 2057.280 1116.220 ;
        RECT 2054.655 1115.880 2057.280 1116.050 ;
        RECT 2057.105 1115.680 2057.280 1115.880 ;
      LAYER li1 ;
        RECT 2060.135 1115.680 2060.390 1116.220 ;
      LAYER li1 ;
        RECT 2063.085 1116.050 2063.260 1116.220 ;
        RECT 2060.635 1115.880 2063.260 1116.050 ;
        RECT 2063.085 1115.680 2063.260 1115.880 ;
      LAYER li1 ;
        RECT 2066.115 1115.680 2066.370 1116.220 ;
      LAYER li1 ;
        RECT 2069.065 1116.050 2069.240 1116.220 ;
        RECT 2066.615 1115.880 2069.240 1116.050 ;
        RECT 2069.065 1115.680 2069.240 1115.880 ;
      LAYER li1 ;
        RECT 2072.095 1115.680 2072.350 1116.220 ;
      LAYER li1 ;
        RECT 2075.045 1116.050 2075.220 1116.220 ;
        RECT 2072.595 1115.880 2075.220 1116.050 ;
        RECT 2075.045 1115.680 2075.220 1115.880 ;
      LAYER li1 ;
        RECT 2078.075 1115.680 2078.330 1116.220 ;
      LAYER li1 ;
        RECT 2081.025 1116.050 2081.200 1116.220 ;
        RECT 2078.575 1115.880 2081.200 1116.050 ;
        RECT 2081.025 1115.680 2081.200 1115.880 ;
      LAYER li1 ;
        RECT 2084.055 1115.680 2084.310 1116.220 ;
      LAYER li1 ;
        RECT 2087.005 1116.050 2087.180 1116.220 ;
        RECT 2084.555 1115.880 2087.180 1116.050 ;
        RECT 2087.005 1115.680 2087.180 1115.880 ;
      LAYER li1 ;
        RECT 2090.035 1115.680 2090.290 1116.220 ;
      LAYER li1 ;
        RECT 2092.985 1116.050 2093.160 1116.220 ;
        RECT 2090.535 1115.880 2093.160 1116.050 ;
        RECT 2092.985 1115.680 2093.160 1115.880 ;
        RECT 669.085 1114.490 669.375 1115.655 ;
        RECT 669.935 1114.490 670.265 1115.640 ;
      LAYER li1 ;
        RECT 670.435 1115.510 673.125 1115.680 ;
      LAYER li1 ;
        RECT 673.385 1115.510 674.885 1115.680 ;
      LAYER li1 ;
        RECT 670.435 1114.660 670.605 1115.510 ;
      LAYER li1 ;
        RECT 670.775 1114.490 671.105 1115.290 ;
      LAYER li1 ;
        RECT 671.275 1114.660 671.445 1115.510 ;
      LAYER li1 ;
        RECT 671.615 1114.490 671.945 1115.290 ;
      LAYER li1 ;
        RECT 672.115 1114.660 672.285 1115.510 ;
      LAYER li1 ;
        RECT 672.455 1114.490 672.785 1115.290 ;
      LAYER li1 ;
        RECT 672.955 1114.660 673.125 1115.510 ;
      LAYER li1 ;
        RECT 673.375 1114.490 673.545 1115.290 ;
        RECT 673.715 1114.660 674.045 1115.510 ;
        RECT 674.215 1114.490 674.385 1115.290 ;
        RECT 674.555 1114.660 674.885 1115.510 ;
        RECT 675.065 1114.490 675.355 1115.655 ;
        RECT 675.915 1114.490 676.245 1115.640 ;
      LAYER li1 ;
        RECT 676.415 1115.510 679.105 1115.680 ;
      LAYER li1 ;
        RECT 679.365 1115.510 680.865 1115.680 ;
      LAYER li1 ;
        RECT 676.415 1114.660 676.585 1115.510 ;
      LAYER li1 ;
        RECT 676.755 1114.490 677.085 1115.290 ;
      LAYER li1 ;
        RECT 677.255 1114.660 677.425 1115.510 ;
      LAYER li1 ;
        RECT 677.595 1114.490 677.925 1115.290 ;
      LAYER li1 ;
        RECT 678.095 1114.660 678.265 1115.510 ;
      LAYER li1 ;
        RECT 678.435 1114.490 678.765 1115.290 ;
      LAYER li1 ;
        RECT 678.935 1114.660 679.105 1115.510 ;
      LAYER li1 ;
        RECT 679.355 1114.490 679.525 1115.290 ;
        RECT 679.695 1114.660 680.025 1115.510 ;
        RECT 680.195 1114.490 680.365 1115.290 ;
        RECT 680.535 1114.660 680.865 1115.510 ;
        RECT 681.045 1114.490 681.335 1115.655 ;
        RECT 681.895 1114.490 682.225 1115.640 ;
      LAYER li1 ;
        RECT 682.395 1115.510 685.085 1115.680 ;
      LAYER li1 ;
        RECT 685.345 1115.510 686.845 1115.680 ;
      LAYER li1 ;
        RECT 682.395 1114.660 682.565 1115.510 ;
      LAYER li1 ;
        RECT 682.735 1114.490 683.065 1115.290 ;
      LAYER li1 ;
        RECT 683.235 1114.660 683.405 1115.510 ;
      LAYER li1 ;
        RECT 683.575 1114.490 683.905 1115.290 ;
      LAYER li1 ;
        RECT 684.075 1114.660 684.245 1115.510 ;
      LAYER li1 ;
        RECT 684.415 1114.490 684.745 1115.290 ;
      LAYER li1 ;
        RECT 684.915 1114.660 685.085 1115.510 ;
      LAYER li1 ;
        RECT 685.335 1114.490 685.505 1115.290 ;
        RECT 685.675 1114.660 686.005 1115.510 ;
        RECT 686.175 1114.490 686.345 1115.290 ;
        RECT 686.515 1114.660 686.845 1115.510 ;
        RECT 687.025 1114.490 687.315 1115.655 ;
        RECT 687.875 1114.490 688.205 1115.640 ;
      LAYER li1 ;
        RECT 688.375 1115.510 691.065 1115.680 ;
      LAYER li1 ;
        RECT 691.325 1115.510 692.825 1115.680 ;
      LAYER li1 ;
        RECT 688.375 1114.660 688.545 1115.510 ;
      LAYER li1 ;
        RECT 688.715 1114.490 689.045 1115.290 ;
      LAYER li1 ;
        RECT 689.215 1114.660 689.385 1115.510 ;
      LAYER li1 ;
        RECT 689.555 1114.490 689.885 1115.290 ;
      LAYER li1 ;
        RECT 690.055 1114.660 690.225 1115.510 ;
      LAYER li1 ;
        RECT 690.395 1114.490 690.725 1115.290 ;
      LAYER li1 ;
        RECT 690.895 1114.660 691.065 1115.510 ;
      LAYER li1 ;
        RECT 691.315 1114.490 691.485 1115.290 ;
        RECT 691.655 1114.660 691.985 1115.510 ;
        RECT 692.155 1114.490 692.325 1115.290 ;
        RECT 692.495 1114.660 692.825 1115.510 ;
        RECT 693.005 1114.490 693.295 1115.655 ;
        RECT 693.855 1114.490 694.185 1115.640 ;
      LAYER li1 ;
        RECT 694.355 1115.510 697.045 1115.680 ;
      LAYER li1 ;
        RECT 697.305 1115.510 698.805 1115.680 ;
      LAYER li1 ;
        RECT 694.355 1114.660 694.525 1115.510 ;
      LAYER li1 ;
        RECT 694.695 1114.490 695.025 1115.290 ;
      LAYER li1 ;
        RECT 695.195 1114.660 695.365 1115.510 ;
      LAYER li1 ;
        RECT 695.535 1114.490 695.865 1115.290 ;
      LAYER li1 ;
        RECT 696.035 1114.660 696.205 1115.510 ;
      LAYER li1 ;
        RECT 696.375 1114.490 696.705 1115.290 ;
      LAYER li1 ;
        RECT 696.875 1114.660 697.045 1115.510 ;
      LAYER li1 ;
        RECT 697.295 1114.490 697.465 1115.290 ;
        RECT 697.635 1114.660 697.965 1115.510 ;
        RECT 698.135 1114.490 698.305 1115.290 ;
        RECT 698.475 1114.660 698.805 1115.510 ;
        RECT 698.985 1114.490 699.275 1115.655 ;
        RECT 699.835 1114.490 700.165 1115.640 ;
      LAYER li1 ;
        RECT 700.335 1115.510 703.025 1115.680 ;
      LAYER li1 ;
        RECT 703.285 1115.510 704.785 1115.680 ;
      LAYER li1 ;
        RECT 700.335 1114.660 700.505 1115.510 ;
      LAYER li1 ;
        RECT 700.675 1114.490 701.005 1115.290 ;
      LAYER li1 ;
        RECT 701.175 1114.660 701.345 1115.510 ;
      LAYER li1 ;
        RECT 701.515 1114.490 701.845 1115.290 ;
      LAYER li1 ;
        RECT 702.015 1114.660 702.185 1115.510 ;
      LAYER li1 ;
        RECT 702.355 1114.490 702.685 1115.290 ;
      LAYER li1 ;
        RECT 702.855 1114.660 703.025 1115.510 ;
      LAYER li1 ;
        RECT 703.275 1114.490 703.445 1115.290 ;
        RECT 703.615 1114.660 703.945 1115.510 ;
        RECT 704.115 1114.490 704.285 1115.290 ;
        RECT 704.455 1114.660 704.785 1115.510 ;
        RECT 704.965 1114.490 705.255 1115.655 ;
        RECT 705.815 1114.490 706.145 1115.640 ;
      LAYER li1 ;
        RECT 706.315 1115.510 709.005 1115.680 ;
      LAYER li1 ;
        RECT 709.265 1115.510 710.765 1115.680 ;
      LAYER li1 ;
        RECT 706.315 1114.660 706.485 1115.510 ;
      LAYER li1 ;
        RECT 706.655 1114.490 706.985 1115.290 ;
      LAYER li1 ;
        RECT 707.155 1114.660 707.325 1115.510 ;
      LAYER li1 ;
        RECT 707.495 1114.490 707.825 1115.290 ;
      LAYER li1 ;
        RECT 707.995 1114.660 708.165 1115.510 ;
      LAYER li1 ;
        RECT 708.335 1114.490 708.665 1115.290 ;
      LAYER li1 ;
        RECT 708.835 1114.660 709.005 1115.510 ;
      LAYER li1 ;
        RECT 709.255 1114.490 709.425 1115.290 ;
        RECT 709.595 1114.660 709.925 1115.510 ;
        RECT 710.095 1114.490 710.265 1115.290 ;
        RECT 710.435 1114.660 710.765 1115.510 ;
        RECT 710.945 1114.490 711.235 1115.655 ;
        RECT 711.795 1114.490 712.125 1115.640 ;
      LAYER li1 ;
        RECT 712.295 1115.510 714.985 1115.680 ;
      LAYER li1 ;
        RECT 715.245 1115.510 716.745 1115.680 ;
      LAYER li1 ;
        RECT 712.295 1114.660 712.465 1115.510 ;
      LAYER li1 ;
        RECT 712.635 1114.490 712.965 1115.290 ;
      LAYER li1 ;
        RECT 713.135 1114.660 713.305 1115.510 ;
      LAYER li1 ;
        RECT 713.475 1114.490 713.805 1115.290 ;
      LAYER li1 ;
        RECT 713.975 1114.660 714.145 1115.510 ;
      LAYER li1 ;
        RECT 714.315 1114.490 714.645 1115.290 ;
      LAYER li1 ;
        RECT 714.815 1114.660 714.985 1115.510 ;
      LAYER li1 ;
        RECT 715.235 1114.490 715.405 1115.290 ;
        RECT 715.575 1114.660 715.905 1115.510 ;
        RECT 716.075 1114.490 716.245 1115.290 ;
        RECT 716.415 1114.660 716.745 1115.510 ;
        RECT 716.925 1114.490 717.215 1115.655 ;
        RECT 717.775 1114.490 718.105 1115.640 ;
      LAYER li1 ;
        RECT 718.275 1115.510 720.965 1115.680 ;
      LAYER li1 ;
        RECT 721.225 1115.510 722.725 1115.680 ;
      LAYER li1 ;
        RECT 718.275 1114.660 718.445 1115.510 ;
      LAYER li1 ;
        RECT 718.615 1114.490 718.945 1115.290 ;
      LAYER li1 ;
        RECT 719.115 1114.660 719.285 1115.510 ;
      LAYER li1 ;
        RECT 719.455 1114.490 719.785 1115.290 ;
      LAYER li1 ;
        RECT 719.955 1114.660 720.125 1115.510 ;
      LAYER li1 ;
        RECT 720.295 1114.490 720.625 1115.290 ;
      LAYER li1 ;
        RECT 720.795 1114.660 720.965 1115.510 ;
      LAYER li1 ;
        RECT 721.215 1114.490 721.385 1115.290 ;
        RECT 721.555 1114.660 721.885 1115.510 ;
        RECT 722.055 1114.490 722.225 1115.290 ;
        RECT 722.395 1114.660 722.725 1115.510 ;
        RECT 722.905 1114.490 723.195 1115.655 ;
        RECT 723.755 1114.490 724.085 1115.640 ;
      LAYER li1 ;
        RECT 724.255 1115.510 726.945 1115.680 ;
      LAYER li1 ;
        RECT 727.205 1115.510 728.705 1115.680 ;
      LAYER li1 ;
        RECT 724.255 1114.660 724.425 1115.510 ;
      LAYER li1 ;
        RECT 724.595 1114.490 724.925 1115.290 ;
      LAYER li1 ;
        RECT 725.095 1114.660 725.265 1115.510 ;
      LAYER li1 ;
        RECT 725.435 1114.490 725.765 1115.290 ;
      LAYER li1 ;
        RECT 725.935 1114.660 726.105 1115.510 ;
      LAYER li1 ;
        RECT 726.275 1114.490 726.605 1115.290 ;
      LAYER li1 ;
        RECT 726.775 1114.660 726.945 1115.510 ;
      LAYER li1 ;
        RECT 727.195 1114.490 727.365 1115.290 ;
        RECT 727.535 1114.660 727.865 1115.510 ;
        RECT 728.035 1114.490 728.205 1115.290 ;
        RECT 728.375 1114.660 728.705 1115.510 ;
        RECT 728.885 1114.490 729.175 1115.655 ;
        RECT 729.735 1114.490 730.065 1115.640 ;
      LAYER li1 ;
        RECT 730.235 1115.510 732.925 1115.680 ;
      LAYER li1 ;
        RECT 733.185 1115.510 734.685 1115.680 ;
      LAYER li1 ;
        RECT 730.235 1114.660 730.405 1115.510 ;
      LAYER li1 ;
        RECT 730.575 1114.490 730.905 1115.290 ;
      LAYER li1 ;
        RECT 731.075 1114.660 731.245 1115.510 ;
      LAYER li1 ;
        RECT 731.415 1114.490 731.745 1115.290 ;
      LAYER li1 ;
        RECT 731.915 1114.660 732.085 1115.510 ;
      LAYER li1 ;
        RECT 732.255 1114.490 732.585 1115.290 ;
      LAYER li1 ;
        RECT 732.755 1114.660 732.925 1115.510 ;
      LAYER li1 ;
        RECT 733.175 1114.490 733.345 1115.290 ;
        RECT 733.515 1114.660 733.845 1115.510 ;
        RECT 734.015 1114.490 734.185 1115.290 ;
        RECT 734.355 1114.660 734.685 1115.510 ;
        RECT 734.865 1114.490 735.155 1115.655 ;
        RECT 735.715 1114.490 736.045 1115.640 ;
      LAYER li1 ;
        RECT 736.215 1115.510 738.905 1115.680 ;
      LAYER li1 ;
        RECT 739.165 1115.510 740.665 1115.680 ;
      LAYER li1 ;
        RECT 736.215 1114.660 736.385 1115.510 ;
      LAYER li1 ;
        RECT 736.555 1114.490 736.885 1115.290 ;
      LAYER li1 ;
        RECT 737.055 1114.660 737.225 1115.510 ;
      LAYER li1 ;
        RECT 737.395 1114.490 737.725 1115.290 ;
      LAYER li1 ;
        RECT 737.895 1114.660 738.065 1115.510 ;
      LAYER li1 ;
        RECT 738.235 1114.490 738.565 1115.290 ;
      LAYER li1 ;
        RECT 738.735 1114.660 738.905 1115.510 ;
      LAYER li1 ;
        RECT 739.155 1114.490 739.325 1115.290 ;
        RECT 739.495 1114.660 739.825 1115.510 ;
        RECT 739.995 1114.490 740.165 1115.290 ;
        RECT 740.335 1114.660 740.665 1115.510 ;
        RECT 740.845 1114.490 741.135 1115.655 ;
        RECT 741.695 1114.490 742.025 1115.640 ;
      LAYER li1 ;
        RECT 742.195 1115.510 744.885 1115.680 ;
      LAYER li1 ;
        RECT 745.145 1115.510 746.645 1115.680 ;
      LAYER li1 ;
        RECT 742.195 1114.660 742.365 1115.510 ;
      LAYER li1 ;
        RECT 742.535 1114.490 742.865 1115.290 ;
      LAYER li1 ;
        RECT 743.035 1114.660 743.205 1115.510 ;
      LAYER li1 ;
        RECT 743.375 1114.490 743.705 1115.290 ;
      LAYER li1 ;
        RECT 743.875 1114.660 744.045 1115.510 ;
      LAYER li1 ;
        RECT 744.215 1114.490 744.545 1115.290 ;
      LAYER li1 ;
        RECT 744.715 1114.660 744.885 1115.510 ;
      LAYER li1 ;
        RECT 745.135 1114.490 745.305 1115.290 ;
        RECT 745.475 1114.660 745.805 1115.510 ;
        RECT 745.975 1114.490 746.145 1115.290 ;
        RECT 746.315 1114.660 746.645 1115.510 ;
        RECT 746.825 1114.490 747.115 1115.655 ;
        RECT 747.675 1114.490 748.005 1115.640 ;
      LAYER li1 ;
        RECT 748.175 1115.510 750.865 1115.680 ;
      LAYER li1 ;
        RECT 751.125 1115.510 752.625 1115.680 ;
      LAYER li1 ;
        RECT 748.175 1114.660 748.345 1115.510 ;
      LAYER li1 ;
        RECT 748.515 1114.490 748.845 1115.290 ;
      LAYER li1 ;
        RECT 749.015 1114.660 749.185 1115.510 ;
      LAYER li1 ;
        RECT 749.355 1114.490 749.685 1115.290 ;
      LAYER li1 ;
        RECT 749.855 1114.660 750.025 1115.510 ;
      LAYER li1 ;
        RECT 750.195 1114.490 750.525 1115.290 ;
      LAYER li1 ;
        RECT 750.695 1114.660 750.865 1115.510 ;
      LAYER li1 ;
        RECT 751.115 1114.490 751.285 1115.290 ;
        RECT 751.455 1114.660 751.785 1115.510 ;
        RECT 751.955 1114.490 752.125 1115.290 ;
        RECT 752.295 1114.660 752.625 1115.510 ;
        RECT 752.805 1114.490 753.095 1115.655 ;
        RECT 753.655 1114.490 753.985 1115.640 ;
      LAYER li1 ;
        RECT 754.155 1115.510 756.845 1115.680 ;
      LAYER li1 ;
        RECT 757.105 1115.510 758.605 1115.680 ;
      LAYER li1 ;
        RECT 754.155 1114.660 754.325 1115.510 ;
      LAYER li1 ;
        RECT 754.495 1114.490 754.825 1115.290 ;
      LAYER li1 ;
        RECT 754.995 1114.660 755.165 1115.510 ;
      LAYER li1 ;
        RECT 755.335 1114.490 755.665 1115.290 ;
      LAYER li1 ;
        RECT 755.835 1114.660 756.005 1115.510 ;
      LAYER li1 ;
        RECT 756.175 1114.490 756.505 1115.290 ;
      LAYER li1 ;
        RECT 756.675 1114.660 756.845 1115.510 ;
      LAYER li1 ;
        RECT 757.095 1114.490 757.265 1115.290 ;
        RECT 757.435 1114.660 757.765 1115.510 ;
        RECT 757.935 1114.490 758.105 1115.290 ;
        RECT 758.275 1114.660 758.605 1115.510 ;
        RECT 758.785 1114.490 759.075 1115.655 ;
        RECT 759.635 1114.490 759.965 1115.640 ;
        RECT 763.085 1115.510 764.585 1115.680 ;
        RECT 760.475 1114.490 760.805 1115.290 ;
        RECT 761.315 1114.490 761.645 1115.290 ;
        RECT 762.155 1114.490 762.485 1115.290 ;
        RECT 763.075 1114.490 763.245 1115.290 ;
        RECT 763.415 1114.660 763.745 1115.510 ;
        RECT 763.915 1114.490 764.085 1115.290 ;
        RECT 764.255 1114.660 764.585 1115.510 ;
        RECT 764.765 1114.490 765.055 1115.655 ;
        RECT 765.615 1114.490 765.945 1115.640 ;
        RECT 769.065 1115.510 770.565 1115.680 ;
        RECT 766.455 1114.490 766.785 1115.290 ;
        RECT 767.295 1114.490 767.625 1115.290 ;
        RECT 768.135 1114.490 768.465 1115.290 ;
        RECT 769.055 1114.490 769.225 1115.290 ;
        RECT 769.395 1114.660 769.725 1115.510 ;
        RECT 769.895 1114.490 770.065 1115.290 ;
        RECT 770.235 1114.660 770.565 1115.510 ;
        RECT 770.745 1114.490 771.035 1115.655 ;
        RECT 771.595 1114.490 771.925 1115.640 ;
        RECT 775.045 1115.510 776.545 1115.680 ;
        RECT 772.435 1114.490 772.765 1115.290 ;
        RECT 773.275 1114.490 773.605 1115.290 ;
        RECT 774.115 1114.490 774.445 1115.290 ;
        RECT 775.035 1114.490 775.205 1115.290 ;
        RECT 775.375 1114.660 775.705 1115.510 ;
        RECT 775.875 1114.490 776.045 1115.290 ;
        RECT 776.215 1114.660 776.545 1115.510 ;
        RECT 776.725 1114.490 777.015 1115.655 ;
        RECT 777.575 1114.490 777.905 1115.640 ;
        RECT 781.025 1115.510 782.525 1115.680 ;
        RECT 778.415 1114.490 778.745 1115.290 ;
        RECT 779.255 1114.490 779.585 1115.290 ;
        RECT 780.095 1114.490 780.425 1115.290 ;
        RECT 781.015 1114.490 781.185 1115.290 ;
        RECT 781.355 1114.660 781.685 1115.510 ;
        RECT 781.855 1114.490 782.025 1115.290 ;
        RECT 782.195 1114.660 782.525 1115.510 ;
        RECT 782.705 1114.490 782.995 1115.655 ;
        RECT 783.555 1114.490 783.885 1115.640 ;
        RECT 787.005 1115.510 788.505 1115.680 ;
        RECT 784.395 1114.490 784.725 1115.290 ;
        RECT 785.235 1114.490 785.565 1115.290 ;
        RECT 786.075 1114.490 786.405 1115.290 ;
        RECT 786.995 1114.490 787.165 1115.290 ;
        RECT 787.335 1114.660 787.665 1115.510 ;
        RECT 787.835 1114.490 788.005 1115.290 ;
        RECT 788.175 1114.660 788.505 1115.510 ;
        RECT 788.685 1114.490 788.975 1115.655 ;
        RECT 789.535 1114.490 789.865 1115.640 ;
        RECT 792.985 1115.510 794.485 1115.680 ;
        RECT 790.375 1114.490 790.705 1115.290 ;
        RECT 791.215 1114.490 791.545 1115.290 ;
        RECT 792.055 1114.490 792.385 1115.290 ;
        RECT 792.975 1114.490 793.145 1115.290 ;
        RECT 793.315 1114.660 793.645 1115.510 ;
        RECT 793.815 1114.490 793.985 1115.290 ;
        RECT 794.155 1114.660 794.485 1115.510 ;
        RECT 794.665 1114.490 794.955 1115.655 ;
        RECT 1969.085 1114.490 1969.375 1115.655 ;
        RECT 1969.935 1114.490 1970.265 1115.640 ;
      LAYER li1 ;
        RECT 1970.435 1115.510 1973.125 1115.680 ;
      LAYER li1 ;
        RECT 1973.385 1115.510 1974.885 1115.680 ;
      LAYER li1 ;
        RECT 1970.435 1114.660 1970.605 1115.510 ;
      LAYER li1 ;
        RECT 1970.775 1114.490 1971.105 1115.290 ;
      LAYER li1 ;
        RECT 1971.275 1114.660 1971.445 1115.510 ;
      LAYER li1 ;
        RECT 1971.615 1114.490 1971.945 1115.290 ;
      LAYER li1 ;
        RECT 1972.115 1114.660 1972.285 1115.510 ;
      LAYER li1 ;
        RECT 1972.455 1114.490 1972.785 1115.290 ;
      LAYER li1 ;
        RECT 1972.955 1114.660 1973.125 1115.510 ;
      LAYER li1 ;
        RECT 1973.375 1114.490 1973.545 1115.290 ;
        RECT 1973.715 1114.660 1974.045 1115.510 ;
        RECT 1974.215 1114.490 1974.385 1115.290 ;
        RECT 1974.555 1114.660 1974.885 1115.510 ;
        RECT 1975.065 1114.490 1975.355 1115.655 ;
        RECT 1975.915 1114.490 1976.245 1115.640 ;
      LAYER li1 ;
        RECT 1976.415 1115.510 1979.105 1115.680 ;
      LAYER li1 ;
        RECT 1979.365 1115.510 1980.865 1115.680 ;
      LAYER li1 ;
        RECT 1976.415 1114.660 1976.585 1115.510 ;
      LAYER li1 ;
        RECT 1976.755 1114.490 1977.085 1115.290 ;
      LAYER li1 ;
        RECT 1977.255 1114.660 1977.425 1115.510 ;
      LAYER li1 ;
        RECT 1977.595 1114.490 1977.925 1115.290 ;
      LAYER li1 ;
        RECT 1978.095 1114.660 1978.265 1115.510 ;
      LAYER li1 ;
        RECT 1978.435 1114.490 1978.765 1115.290 ;
      LAYER li1 ;
        RECT 1978.935 1114.660 1979.105 1115.510 ;
      LAYER li1 ;
        RECT 1979.355 1114.490 1979.525 1115.290 ;
        RECT 1979.695 1114.660 1980.025 1115.510 ;
        RECT 1980.195 1114.490 1980.365 1115.290 ;
        RECT 1980.535 1114.660 1980.865 1115.510 ;
        RECT 1981.045 1114.490 1981.335 1115.655 ;
        RECT 1981.895 1114.490 1982.225 1115.640 ;
      LAYER li1 ;
        RECT 1982.395 1115.510 1985.085 1115.680 ;
      LAYER li1 ;
        RECT 1985.345 1115.510 1986.845 1115.680 ;
      LAYER li1 ;
        RECT 1982.395 1114.660 1982.565 1115.510 ;
      LAYER li1 ;
        RECT 1982.735 1114.490 1983.065 1115.290 ;
      LAYER li1 ;
        RECT 1983.235 1114.660 1983.405 1115.510 ;
      LAYER li1 ;
        RECT 1983.575 1114.490 1983.905 1115.290 ;
      LAYER li1 ;
        RECT 1984.075 1114.660 1984.245 1115.510 ;
      LAYER li1 ;
        RECT 1984.415 1114.490 1984.745 1115.290 ;
      LAYER li1 ;
        RECT 1984.915 1114.660 1985.085 1115.510 ;
      LAYER li1 ;
        RECT 1985.335 1114.490 1985.505 1115.290 ;
        RECT 1985.675 1114.660 1986.005 1115.510 ;
        RECT 1986.175 1114.490 1986.345 1115.290 ;
        RECT 1986.515 1114.660 1986.845 1115.510 ;
        RECT 1987.025 1114.490 1987.315 1115.655 ;
        RECT 1987.875 1114.490 1988.205 1115.640 ;
      LAYER li1 ;
        RECT 1988.375 1115.510 1991.065 1115.680 ;
      LAYER li1 ;
        RECT 1991.325 1115.510 1992.825 1115.680 ;
      LAYER li1 ;
        RECT 1988.375 1114.660 1988.545 1115.510 ;
      LAYER li1 ;
        RECT 1988.715 1114.490 1989.045 1115.290 ;
      LAYER li1 ;
        RECT 1989.215 1114.660 1989.385 1115.510 ;
      LAYER li1 ;
        RECT 1989.555 1114.490 1989.885 1115.290 ;
      LAYER li1 ;
        RECT 1990.055 1114.660 1990.225 1115.510 ;
      LAYER li1 ;
        RECT 1990.395 1114.490 1990.725 1115.290 ;
      LAYER li1 ;
        RECT 1990.895 1114.660 1991.065 1115.510 ;
      LAYER li1 ;
        RECT 1991.315 1114.490 1991.485 1115.290 ;
        RECT 1991.655 1114.660 1991.985 1115.510 ;
        RECT 1992.155 1114.490 1992.325 1115.290 ;
        RECT 1992.495 1114.660 1992.825 1115.510 ;
        RECT 1993.005 1114.490 1993.295 1115.655 ;
        RECT 1993.855 1114.490 1994.185 1115.640 ;
      LAYER li1 ;
        RECT 1994.355 1115.510 1997.045 1115.680 ;
      LAYER li1 ;
        RECT 1997.305 1115.510 1998.805 1115.680 ;
      LAYER li1 ;
        RECT 1994.355 1114.660 1994.525 1115.510 ;
      LAYER li1 ;
        RECT 1994.695 1114.490 1995.025 1115.290 ;
      LAYER li1 ;
        RECT 1995.195 1114.660 1995.365 1115.510 ;
      LAYER li1 ;
        RECT 1995.535 1114.490 1995.865 1115.290 ;
      LAYER li1 ;
        RECT 1996.035 1114.660 1996.205 1115.510 ;
      LAYER li1 ;
        RECT 1996.375 1114.490 1996.705 1115.290 ;
      LAYER li1 ;
        RECT 1996.875 1114.660 1997.045 1115.510 ;
      LAYER li1 ;
        RECT 1997.295 1114.490 1997.465 1115.290 ;
        RECT 1997.635 1114.660 1997.965 1115.510 ;
        RECT 1998.135 1114.490 1998.305 1115.290 ;
        RECT 1998.475 1114.660 1998.805 1115.510 ;
        RECT 1998.985 1114.490 1999.275 1115.655 ;
        RECT 1999.835 1114.490 2000.165 1115.640 ;
      LAYER li1 ;
        RECT 2000.335 1115.510 2003.025 1115.680 ;
      LAYER li1 ;
        RECT 2003.285 1115.510 2004.785 1115.680 ;
      LAYER li1 ;
        RECT 2000.335 1114.660 2000.505 1115.510 ;
      LAYER li1 ;
        RECT 2000.675 1114.490 2001.005 1115.290 ;
      LAYER li1 ;
        RECT 2001.175 1114.660 2001.345 1115.510 ;
      LAYER li1 ;
        RECT 2001.515 1114.490 2001.845 1115.290 ;
      LAYER li1 ;
        RECT 2002.015 1114.660 2002.185 1115.510 ;
      LAYER li1 ;
        RECT 2002.355 1114.490 2002.685 1115.290 ;
      LAYER li1 ;
        RECT 2002.855 1114.660 2003.025 1115.510 ;
      LAYER li1 ;
        RECT 2003.275 1114.490 2003.445 1115.290 ;
        RECT 2003.615 1114.660 2003.945 1115.510 ;
        RECT 2004.115 1114.490 2004.285 1115.290 ;
        RECT 2004.455 1114.660 2004.785 1115.510 ;
        RECT 2004.965 1114.490 2005.255 1115.655 ;
        RECT 2005.815 1114.490 2006.145 1115.640 ;
      LAYER li1 ;
        RECT 2006.315 1115.510 2009.005 1115.680 ;
      LAYER li1 ;
        RECT 2009.265 1115.510 2010.765 1115.680 ;
      LAYER li1 ;
        RECT 2006.315 1114.660 2006.485 1115.510 ;
      LAYER li1 ;
        RECT 2006.655 1114.490 2006.985 1115.290 ;
      LAYER li1 ;
        RECT 2007.155 1114.660 2007.325 1115.510 ;
      LAYER li1 ;
        RECT 2007.495 1114.490 2007.825 1115.290 ;
      LAYER li1 ;
        RECT 2007.995 1114.660 2008.165 1115.510 ;
      LAYER li1 ;
        RECT 2008.335 1114.490 2008.665 1115.290 ;
      LAYER li1 ;
        RECT 2008.835 1114.660 2009.005 1115.510 ;
      LAYER li1 ;
        RECT 2009.255 1114.490 2009.425 1115.290 ;
        RECT 2009.595 1114.660 2009.925 1115.510 ;
        RECT 2010.095 1114.490 2010.265 1115.290 ;
        RECT 2010.435 1114.660 2010.765 1115.510 ;
        RECT 2010.945 1114.490 2011.235 1115.655 ;
        RECT 2011.795 1114.490 2012.125 1115.640 ;
      LAYER li1 ;
        RECT 2012.295 1115.510 2014.985 1115.680 ;
      LAYER li1 ;
        RECT 2015.245 1115.510 2016.745 1115.680 ;
      LAYER li1 ;
        RECT 2012.295 1114.660 2012.465 1115.510 ;
      LAYER li1 ;
        RECT 2012.635 1114.490 2012.965 1115.290 ;
      LAYER li1 ;
        RECT 2013.135 1114.660 2013.305 1115.510 ;
      LAYER li1 ;
        RECT 2013.475 1114.490 2013.805 1115.290 ;
      LAYER li1 ;
        RECT 2013.975 1114.660 2014.145 1115.510 ;
      LAYER li1 ;
        RECT 2014.315 1114.490 2014.645 1115.290 ;
      LAYER li1 ;
        RECT 2014.815 1114.660 2014.985 1115.510 ;
      LAYER li1 ;
        RECT 2015.235 1114.490 2015.405 1115.290 ;
        RECT 2015.575 1114.660 2015.905 1115.510 ;
        RECT 2016.075 1114.490 2016.245 1115.290 ;
        RECT 2016.415 1114.660 2016.745 1115.510 ;
        RECT 2016.925 1114.490 2017.215 1115.655 ;
        RECT 2017.775 1114.490 2018.105 1115.640 ;
      LAYER li1 ;
        RECT 2018.275 1115.510 2020.965 1115.680 ;
      LAYER li1 ;
        RECT 2021.225 1115.510 2022.725 1115.680 ;
      LAYER li1 ;
        RECT 2018.275 1114.660 2018.445 1115.510 ;
      LAYER li1 ;
        RECT 2018.615 1114.490 2018.945 1115.290 ;
      LAYER li1 ;
        RECT 2019.115 1114.660 2019.285 1115.510 ;
      LAYER li1 ;
        RECT 2019.455 1114.490 2019.785 1115.290 ;
      LAYER li1 ;
        RECT 2019.955 1114.660 2020.125 1115.510 ;
      LAYER li1 ;
        RECT 2020.295 1114.490 2020.625 1115.290 ;
      LAYER li1 ;
        RECT 2020.795 1114.660 2020.965 1115.510 ;
      LAYER li1 ;
        RECT 2021.215 1114.490 2021.385 1115.290 ;
        RECT 2021.555 1114.660 2021.885 1115.510 ;
        RECT 2022.055 1114.490 2022.225 1115.290 ;
        RECT 2022.395 1114.660 2022.725 1115.510 ;
        RECT 2022.905 1114.490 2023.195 1115.655 ;
        RECT 2023.755 1114.490 2024.085 1115.640 ;
      LAYER li1 ;
        RECT 2024.255 1115.510 2026.945 1115.680 ;
      LAYER li1 ;
        RECT 2027.205 1115.510 2028.705 1115.680 ;
      LAYER li1 ;
        RECT 2024.255 1114.660 2024.425 1115.510 ;
      LAYER li1 ;
        RECT 2024.595 1114.490 2024.925 1115.290 ;
      LAYER li1 ;
        RECT 2025.095 1114.660 2025.265 1115.510 ;
      LAYER li1 ;
        RECT 2025.435 1114.490 2025.765 1115.290 ;
      LAYER li1 ;
        RECT 2025.935 1114.660 2026.105 1115.510 ;
      LAYER li1 ;
        RECT 2026.275 1114.490 2026.605 1115.290 ;
      LAYER li1 ;
        RECT 2026.775 1114.660 2026.945 1115.510 ;
      LAYER li1 ;
        RECT 2027.195 1114.490 2027.365 1115.290 ;
        RECT 2027.535 1114.660 2027.865 1115.510 ;
        RECT 2028.035 1114.490 2028.205 1115.290 ;
        RECT 2028.375 1114.660 2028.705 1115.510 ;
        RECT 2028.885 1114.490 2029.175 1115.655 ;
        RECT 2029.735 1114.490 2030.065 1115.640 ;
      LAYER li1 ;
        RECT 2030.235 1115.510 2032.925 1115.680 ;
      LAYER li1 ;
        RECT 2033.185 1115.510 2034.685 1115.680 ;
      LAYER li1 ;
        RECT 2030.235 1114.660 2030.405 1115.510 ;
      LAYER li1 ;
        RECT 2030.575 1114.490 2030.905 1115.290 ;
      LAYER li1 ;
        RECT 2031.075 1114.660 2031.245 1115.510 ;
      LAYER li1 ;
        RECT 2031.415 1114.490 2031.745 1115.290 ;
      LAYER li1 ;
        RECT 2031.915 1114.660 2032.085 1115.510 ;
      LAYER li1 ;
        RECT 2032.255 1114.490 2032.585 1115.290 ;
      LAYER li1 ;
        RECT 2032.755 1114.660 2032.925 1115.510 ;
      LAYER li1 ;
        RECT 2033.175 1114.490 2033.345 1115.290 ;
        RECT 2033.515 1114.660 2033.845 1115.510 ;
        RECT 2034.015 1114.490 2034.185 1115.290 ;
        RECT 2034.355 1114.660 2034.685 1115.510 ;
        RECT 2034.865 1114.490 2035.155 1115.655 ;
        RECT 2035.715 1114.490 2036.045 1115.640 ;
      LAYER li1 ;
        RECT 2036.215 1115.510 2038.905 1115.680 ;
      LAYER li1 ;
        RECT 2039.165 1115.510 2040.665 1115.680 ;
      LAYER li1 ;
        RECT 2036.215 1114.660 2036.385 1115.510 ;
      LAYER li1 ;
        RECT 2036.555 1114.490 2036.885 1115.290 ;
      LAYER li1 ;
        RECT 2037.055 1114.660 2037.225 1115.510 ;
      LAYER li1 ;
        RECT 2037.395 1114.490 2037.725 1115.290 ;
      LAYER li1 ;
        RECT 2037.895 1114.660 2038.065 1115.510 ;
      LAYER li1 ;
        RECT 2038.235 1114.490 2038.565 1115.290 ;
      LAYER li1 ;
        RECT 2038.735 1114.660 2038.905 1115.510 ;
      LAYER li1 ;
        RECT 2039.155 1114.490 2039.325 1115.290 ;
        RECT 2039.495 1114.660 2039.825 1115.510 ;
        RECT 2039.995 1114.490 2040.165 1115.290 ;
        RECT 2040.335 1114.660 2040.665 1115.510 ;
        RECT 2040.845 1114.490 2041.135 1115.655 ;
        RECT 2041.695 1114.490 2042.025 1115.640 ;
      LAYER li1 ;
        RECT 2042.195 1115.510 2044.885 1115.680 ;
      LAYER li1 ;
        RECT 2045.145 1115.510 2046.645 1115.680 ;
      LAYER li1 ;
        RECT 2042.195 1114.660 2042.365 1115.510 ;
      LAYER li1 ;
        RECT 2042.535 1114.490 2042.865 1115.290 ;
      LAYER li1 ;
        RECT 2043.035 1114.660 2043.205 1115.510 ;
      LAYER li1 ;
        RECT 2043.375 1114.490 2043.705 1115.290 ;
      LAYER li1 ;
        RECT 2043.875 1114.660 2044.045 1115.510 ;
      LAYER li1 ;
        RECT 2044.215 1114.490 2044.545 1115.290 ;
      LAYER li1 ;
        RECT 2044.715 1114.660 2044.885 1115.510 ;
      LAYER li1 ;
        RECT 2045.135 1114.490 2045.305 1115.290 ;
        RECT 2045.475 1114.660 2045.805 1115.510 ;
        RECT 2045.975 1114.490 2046.145 1115.290 ;
        RECT 2046.315 1114.660 2046.645 1115.510 ;
        RECT 2046.825 1114.490 2047.115 1115.655 ;
        RECT 2047.675 1114.490 2048.005 1115.640 ;
      LAYER li1 ;
        RECT 2048.175 1115.510 2050.865 1115.680 ;
      LAYER li1 ;
        RECT 2051.125 1115.510 2052.625 1115.680 ;
      LAYER li1 ;
        RECT 2048.175 1114.660 2048.345 1115.510 ;
      LAYER li1 ;
        RECT 2048.515 1114.490 2048.845 1115.290 ;
      LAYER li1 ;
        RECT 2049.015 1114.660 2049.185 1115.510 ;
      LAYER li1 ;
        RECT 2049.355 1114.490 2049.685 1115.290 ;
      LAYER li1 ;
        RECT 2049.855 1114.660 2050.025 1115.510 ;
      LAYER li1 ;
        RECT 2050.195 1114.490 2050.525 1115.290 ;
      LAYER li1 ;
        RECT 2050.695 1114.660 2050.865 1115.510 ;
      LAYER li1 ;
        RECT 2051.115 1114.490 2051.285 1115.290 ;
        RECT 2051.455 1114.660 2051.785 1115.510 ;
        RECT 2051.955 1114.490 2052.125 1115.290 ;
        RECT 2052.295 1114.660 2052.625 1115.510 ;
        RECT 2052.805 1114.490 2053.095 1115.655 ;
        RECT 2053.655 1114.490 2053.985 1115.640 ;
      LAYER li1 ;
        RECT 2054.155 1115.510 2056.845 1115.680 ;
      LAYER li1 ;
        RECT 2057.105 1115.510 2058.605 1115.680 ;
      LAYER li1 ;
        RECT 2054.155 1114.660 2054.325 1115.510 ;
      LAYER li1 ;
        RECT 2054.495 1114.490 2054.825 1115.290 ;
      LAYER li1 ;
        RECT 2054.995 1114.660 2055.165 1115.510 ;
      LAYER li1 ;
        RECT 2055.335 1114.490 2055.665 1115.290 ;
      LAYER li1 ;
        RECT 2055.835 1114.660 2056.005 1115.510 ;
      LAYER li1 ;
        RECT 2056.175 1114.490 2056.505 1115.290 ;
      LAYER li1 ;
        RECT 2056.675 1114.660 2056.845 1115.510 ;
      LAYER li1 ;
        RECT 2057.095 1114.490 2057.265 1115.290 ;
        RECT 2057.435 1114.660 2057.765 1115.510 ;
        RECT 2057.935 1114.490 2058.105 1115.290 ;
        RECT 2058.275 1114.660 2058.605 1115.510 ;
        RECT 2058.785 1114.490 2059.075 1115.655 ;
        RECT 2059.635 1114.490 2059.965 1115.640 ;
      LAYER li1 ;
        RECT 2060.135 1115.510 2062.825 1115.680 ;
      LAYER li1 ;
        RECT 2063.085 1115.510 2064.585 1115.680 ;
      LAYER li1 ;
        RECT 2060.135 1114.660 2060.305 1115.510 ;
      LAYER li1 ;
        RECT 2060.475 1114.490 2060.805 1115.290 ;
      LAYER li1 ;
        RECT 2060.975 1114.660 2061.145 1115.510 ;
      LAYER li1 ;
        RECT 2061.315 1114.490 2061.645 1115.290 ;
      LAYER li1 ;
        RECT 2061.815 1114.660 2061.985 1115.510 ;
      LAYER li1 ;
        RECT 2062.155 1114.490 2062.485 1115.290 ;
      LAYER li1 ;
        RECT 2062.655 1114.660 2062.825 1115.510 ;
      LAYER li1 ;
        RECT 2063.075 1114.490 2063.245 1115.290 ;
        RECT 2063.415 1114.660 2063.745 1115.510 ;
        RECT 2063.915 1114.490 2064.085 1115.290 ;
        RECT 2064.255 1114.660 2064.585 1115.510 ;
        RECT 2064.765 1114.490 2065.055 1115.655 ;
        RECT 2065.615 1114.490 2065.945 1115.640 ;
      LAYER li1 ;
        RECT 2066.115 1115.510 2068.805 1115.680 ;
      LAYER li1 ;
        RECT 2069.065 1115.510 2070.565 1115.680 ;
      LAYER li1 ;
        RECT 2066.115 1114.660 2066.285 1115.510 ;
      LAYER li1 ;
        RECT 2066.455 1114.490 2066.785 1115.290 ;
      LAYER li1 ;
        RECT 2066.955 1114.660 2067.125 1115.510 ;
      LAYER li1 ;
        RECT 2067.295 1114.490 2067.625 1115.290 ;
      LAYER li1 ;
        RECT 2067.795 1114.660 2067.965 1115.510 ;
      LAYER li1 ;
        RECT 2068.135 1114.490 2068.465 1115.290 ;
      LAYER li1 ;
        RECT 2068.635 1114.660 2068.805 1115.510 ;
      LAYER li1 ;
        RECT 2069.055 1114.490 2069.225 1115.290 ;
        RECT 2069.395 1114.660 2069.725 1115.510 ;
        RECT 2069.895 1114.490 2070.065 1115.290 ;
        RECT 2070.235 1114.660 2070.565 1115.510 ;
        RECT 2070.745 1114.490 2071.035 1115.655 ;
        RECT 2071.595 1114.490 2071.925 1115.640 ;
      LAYER li1 ;
        RECT 2072.095 1115.510 2074.785 1115.680 ;
      LAYER li1 ;
        RECT 2075.045 1115.510 2076.545 1115.680 ;
      LAYER li1 ;
        RECT 2072.095 1114.660 2072.265 1115.510 ;
      LAYER li1 ;
        RECT 2072.435 1114.490 2072.765 1115.290 ;
      LAYER li1 ;
        RECT 2072.935 1114.660 2073.105 1115.510 ;
      LAYER li1 ;
        RECT 2073.275 1114.490 2073.605 1115.290 ;
      LAYER li1 ;
        RECT 2073.775 1114.660 2073.945 1115.510 ;
      LAYER li1 ;
        RECT 2074.115 1114.490 2074.445 1115.290 ;
      LAYER li1 ;
        RECT 2074.615 1114.660 2074.785 1115.510 ;
      LAYER li1 ;
        RECT 2075.035 1114.490 2075.205 1115.290 ;
        RECT 2075.375 1114.660 2075.705 1115.510 ;
        RECT 2075.875 1114.490 2076.045 1115.290 ;
        RECT 2076.215 1114.660 2076.545 1115.510 ;
        RECT 2076.725 1114.490 2077.015 1115.655 ;
        RECT 2077.575 1114.490 2077.905 1115.640 ;
      LAYER li1 ;
        RECT 2078.075 1115.510 2080.765 1115.680 ;
      LAYER li1 ;
        RECT 2081.025 1115.510 2082.525 1115.680 ;
      LAYER li1 ;
        RECT 2078.075 1114.660 2078.245 1115.510 ;
      LAYER li1 ;
        RECT 2078.415 1114.490 2078.745 1115.290 ;
      LAYER li1 ;
        RECT 2078.915 1114.660 2079.085 1115.510 ;
      LAYER li1 ;
        RECT 2079.255 1114.490 2079.585 1115.290 ;
      LAYER li1 ;
        RECT 2079.755 1114.660 2079.925 1115.510 ;
      LAYER li1 ;
        RECT 2080.095 1114.490 2080.425 1115.290 ;
      LAYER li1 ;
        RECT 2080.595 1114.660 2080.765 1115.510 ;
      LAYER li1 ;
        RECT 2081.015 1114.490 2081.185 1115.290 ;
        RECT 2081.355 1114.660 2081.685 1115.510 ;
        RECT 2081.855 1114.490 2082.025 1115.290 ;
        RECT 2082.195 1114.660 2082.525 1115.510 ;
        RECT 2082.705 1114.490 2082.995 1115.655 ;
        RECT 2083.555 1114.490 2083.885 1115.640 ;
      LAYER li1 ;
        RECT 2084.055 1115.510 2086.745 1115.680 ;
      LAYER li1 ;
        RECT 2087.005 1115.510 2088.505 1115.680 ;
      LAYER li1 ;
        RECT 2084.055 1114.660 2084.225 1115.510 ;
      LAYER li1 ;
        RECT 2084.395 1114.490 2084.725 1115.290 ;
      LAYER li1 ;
        RECT 2084.895 1114.660 2085.065 1115.510 ;
      LAYER li1 ;
        RECT 2085.235 1114.490 2085.565 1115.290 ;
      LAYER li1 ;
        RECT 2085.735 1114.660 2085.905 1115.510 ;
      LAYER li1 ;
        RECT 2086.075 1114.490 2086.405 1115.290 ;
      LAYER li1 ;
        RECT 2086.575 1114.660 2086.745 1115.510 ;
      LAYER li1 ;
        RECT 2086.995 1114.490 2087.165 1115.290 ;
        RECT 2087.335 1114.660 2087.665 1115.510 ;
        RECT 2087.835 1114.490 2088.005 1115.290 ;
        RECT 2088.175 1114.660 2088.505 1115.510 ;
        RECT 2088.685 1114.490 2088.975 1115.655 ;
        RECT 2089.535 1114.490 2089.865 1115.640 ;
      LAYER li1 ;
        RECT 2090.035 1115.510 2092.725 1115.680 ;
      LAYER li1 ;
        RECT 2092.985 1115.510 2094.485 1115.680 ;
      LAYER li1 ;
        RECT 2090.035 1114.660 2090.205 1115.510 ;
      LAYER li1 ;
        RECT 2090.375 1114.490 2090.705 1115.290 ;
      LAYER li1 ;
        RECT 2090.875 1114.660 2091.045 1115.510 ;
      LAYER li1 ;
        RECT 2091.215 1114.490 2091.545 1115.290 ;
      LAYER li1 ;
        RECT 2091.715 1114.660 2091.885 1115.510 ;
      LAYER li1 ;
        RECT 2092.055 1114.490 2092.385 1115.290 ;
      LAYER li1 ;
        RECT 2092.555 1114.660 2092.725 1115.510 ;
      LAYER li1 ;
        RECT 2092.975 1114.490 2093.145 1115.290 ;
        RECT 2093.315 1114.660 2093.645 1115.510 ;
        RECT 2093.815 1114.490 2093.985 1115.290 ;
        RECT 2094.155 1114.660 2094.485 1115.510 ;
        RECT 2094.665 1114.490 2094.955 1115.655 ;
        RECT 669.000 1114.320 669.145 1114.490 ;
        RECT 669.315 1114.320 669.605 1114.490 ;
        RECT 669.775 1114.320 670.065 1114.490 ;
        RECT 670.235 1114.320 670.525 1114.490 ;
        RECT 670.695 1114.320 670.985 1114.490 ;
        RECT 671.155 1114.320 671.445 1114.490 ;
        RECT 671.615 1114.320 671.905 1114.490 ;
        RECT 672.075 1114.320 672.365 1114.490 ;
        RECT 672.535 1114.320 672.825 1114.490 ;
        RECT 672.995 1114.320 673.285 1114.490 ;
        RECT 673.455 1114.320 673.745 1114.490 ;
        RECT 673.915 1114.320 674.205 1114.490 ;
        RECT 674.375 1114.320 674.665 1114.490 ;
        RECT 674.835 1114.320 675.125 1114.490 ;
        RECT 675.295 1114.320 675.585 1114.490 ;
        RECT 675.755 1114.320 676.045 1114.490 ;
        RECT 676.215 1114.320 676.505 1114.490 ;
        RECT 676.675 1114.320 676.965 1114.490 ;
        RECT 677.135 1114.320 677.425 1114.490 ;
        RECT 677.595 1114.320 677.885 1114.490 ;
        RECT 678.055 1114.320 678.345 1114.490 ;
        RECT 678.515 1114.320 678.805 1114.490 ;
        RECT 678.975 1114.320 679.265 1114.490 ;
        RECT 679.435 1114.320 679.725 1114.490 ;
        RECT 679.895 1114.320 680.185 1114.490 ;
        RECT 680.355 1114.320 680.645 1114.490 ;
        RECT 680.815 1114.320 681.105 1114.490 ;
        RECT 681.275 1114.320 681.565 1114.490 ;
        RECT 681.735 1114.320 682.025 1114.490 ;
        RECT 682.195 1114.320 682.485 1114.490 ;
        RECT 682.655 1114.320 682.945 1114.490 ;
        RECT 683.115 1114.320 683.405 1114.490 ;
        RECT 683.575 1114.320 683.865 1114.490 ;
        RECT 684.035 1114.320 684.325 1114.490 ;
        RECT 684.495 1114.320 684.785 1114.490 ;
        RECT 684.955 1114.320 685.245 1114.490 ;
        RECT 685.415 1114.320 685.705 1114.490 ;
        RECT 685.875 1114.320 686.165 1114.490 ;
        RECT 686.335 1114.320 686.625 1114.490 ;
        RECT 686.795 1114.320 687.085 1114.490 ;
        RECT 687.255 1114.320 687.545 1114.490 ;
        RECT 687.715 1114.320 688.005 1114.490 ;
        RECT 688.175 1114.320 688.465 1114.490 ;
        RECT 688.635 1114.320 688.925 1114.490 ;
        RECT 689.095 1114.320 689.385 1114.490 ;
        RECT 689.555 1114.320 689.845 1114.490 ;
        RECT 690.015 1114.320 690.305 1114.490 ;
        RECT 690.475 1114.320 690.765 1114.490 ;
        RECT 690.935 1114.320 691.225 1114.490 ;
        RECT 691.395 1114.320 691.685 1114.490 ;
        RECT 691.855 1114.320 692.145 1114.490 ;
        RECT 692.315 1114.320 692.605 1114.490 ;
        RECT 692.775 1114.320 693.065 1114.490 ;
        RECT 693.235 1114.320 693.525 1114.490 ;
        RECT 693.695 1114.320 693.985 1114.490 ;
        RECT 694.155 1114.320 694.445 1114.490 ;
        RECT 694.615 1114.320 694.905 1114.490 ;
        RECT 695.075 1114.320 695.365 1114.490 ;
        RECT 695.535 1114.320 695.825 1114.490 ;
        RECT 695.995 1114.320 696.285 1114.490 ;
        RECT 696.455 1114.320 696.745 1114.490 ;
        RECT 696.915 1114.320 697.205 1114.490 ;
        RECT 697.375 1114.320 697.665 1114.490 ;
        RECT 697.835 1114.320 698.125 1114.490 ;
        RECT 698.295 1114.320 698.585 1114.490 ;
        RECT 698.755 1114.320 699.045 1114.490 ;
        RECT 699.215 1114.320 699.505 1114.490 ;
        RECT 699.675 1114.320 699.965 1114.490 ;
        RECT 700.135 1114.320 700.425 1114.490 ;
        RECT 700.595 1114.320 700.885 1114.490 ;
        RECT 701.055 1114.320 701.345 1114.490 ;
        RECT 701.515 1114.320 701.805 1114.490 ;
        RECT 701.975 1114.320 702.265 1114.490 ;
        RECT 702.435 1114.320 702.725 1114.490 ;
        RECT 702.895 1114.320 703.185 1114.490 ;
        RECT 703.355 1114.320 703.645 1114.490 ;
        RECT 703.815 1114.320 704.105 1114.490 ;
        RECT 704.275 1114.320 704.565 1114.490 ;
        RECT 704.735 1114.320 705.025 1114.490 ;
        RECT 705.195 1114.320 705.485 1114.490 ;
        RECT 705.655 1114.320 705.945 1114.490 ;
        RECT 706.115 1114.320 706.405 1114.490 ;
        RECT 706.575 1114.320 706.865 1114.490 ;
        RECT 707.035 1114.320 707.325 1114.490 ;
        RECT 707.495 1114.320 707.785 1114.490 ;
        RECT 707.955 1114.320 708.245 1114.490 ;
        RECT 708.415 1114.320 708.705 1114.490 ;
        RECT 708.875 1114.320 709.165 1114.490 ;
        RECT 709.335 1114.320 709.625 1114.490 ;
        RECT 709.795 1114.320 710.085 1114.490 ;
        RECT 710.255 1114.320 710.545 1114.490 ;
        RECT 710.715 1114.320 711.005 1114.490 ;
        RECT 711.175 1114.320 711.465 1114.490 ;
        RECT 711.635 1114.320 711.925 1114.490 ;
        RECT 712.095 1114.320 712.385 1114.490 ;
        RECT 712.555 1114.320 712.845 1114.490 ;
        RECT 713.015 1114.320 713.305 1114.490 ;
        RECT 713.475 1114.320 713.765 1114.490 ;
        RECT 713.935 1114.320 714.225 1114.490 ;
        RECT 714.395 1114.320 714.685 1114.490 ;
        RECT 714.855 1114.320 715.145 1114.490 ;
        RECT 715.315 1114.320 715.605 1114.490 ;
        RECT 715.775 1114.320 716.065 1114.490 ;
        RECT 716.235 1114.320 716.525 1114.490 ;
        RECT 716.695 1114.320 716.985 1114.490 ;
        RECT 717.155 1114.320 717.445 1114.490 ;
        RECT 717.615 1114.320 717.905 1114.490 ;
        RECT 718.075 1114.320 718.365 1114.490 ;
        RECT 718.535 1114.320 718.825 1114.490 ;
        RECT 718.995 1114.320 719.285 1114.490 ;
        RECT 719.455 1114.320 719.745 1114.490 ;
        RECT 719.915 1114.320 720.205 1114.490 ;
        RECT 720.375 1114.320 720.665 1114.490 ;
        RECT 720.835 1114.320 721.125 1114.490 ;
        RECT 721.295 1114.320 721.585 1114.490 ;
        RECT 721.755 1114.320 722.045 1114.490 ;
        RECT 722.215 1114.320 722.505 1114.490 ;
        RECT 722.675 1114.320 722.965 1114.490 ;
        RECT 723.135 1114.320 723.425 1114.490 ;
        RECT 723.595 1114.320 723.885 1114.490 ;
        RECT 724.055 1114.320 724.345 1114.490 ;
        RECT 724.515 1114.320 724.805 1114.490 ;
        RECT 724.975 1114.320 725.265 1114.490 ;
        RECT 725.435 1114.320 725.725 1114.490 ;
        RECT 725.895 1114.320 726.185 1114.490 ;
        RECT 726.355 1114.320 726.645 1114.490 ;
        RECT 726.815 1114.320 727.105 1114.490 ;
        RECT 727.275 1114.320 727.565 1114.490 ;
        RECT 727.735 1114.320 728.025 1114.490 ;
        RECT 728.195 1114.320 728.485 1114.490 ;
        RECT 728.655 1114.320 728.945 1114.490 ;
        RECT 729.115 1114.320 729.405 1114.490 ;
        RECT 729.575 1114.320 729.865 1114.490 ;
        RECT 730.035 1114.320 730.325 1114.490 ;
        RECT 730.495 1114.320 730.785 1114.490 ;
        RECT 730.955 1114.320 731.245 1114.490 ;
        RECT 731.415 1114.320 731.705 1114.490 ;
        RECT 731.875 1114.320 732.165 1114.490 ;
        RECT 732.335 1114.320 732.625 1114.490 ;
        RECT 732.795 1114.320 733.085 1114.490 ;
        RECT 733.255 1114.320 733.545 1114.490 ;
        RECT 733.715 1114.320 734.005 1114.490 ;
        RECT 734.175 1114.320 734.465 1114.490 ;
        RECT 734.635 1114.320 734.925 1114.490 ;
        RECT 735.095 1114.320 735.385 1114.490 ;
        RECT 735.555 1114.320 735.845 1114.490 ;
        RECT 736.015 1114.320 736.305 1114.490 ;
        RECT 736.475 1114.320 736.765 1114.490 ;
        RECT 736.935 1114.320 737.225 1114.490 ;
        RECT 737.395 1114.320 737.685 1114.490 ;
        RECT 737.855 1114.320 738.145 1114.490 ;
        RECT 738.315 1114.320 738.605 1114.490 ;
        RECT 738.775 1114.320 739.065 1114.490 ;
        RECT 739.235 1114.320 739.525 1114.490 ;
        RECT 739.695 1114.320 739.985 1114.490 ;
        RECT 740.155 1114.320 740.445 1114.490 ;
        RECT 740.615 1114.320 740.905 1114.490 ;
        RECT 741.075 1114.320 741.365 1114.490 ;
        RECT 741.535 1114.320 741.825 1114.490 ;
        RECT 741.995 1114.320 742.285 1114.490 ;
        RECT 742.455 1114.320 742.745 1114.490 ;
        RECT 742.915 1114.320 743.205 1114.490 ;
        RECT 743.375 1114.320 743.665 1114.490 ;
        RECT 743.835 1114.320 744.125 1114.490 ;
        RECT 744.295 1114.320 744.585 1114.490 ;
        RECT 744.755 1114.320 745.045 1114.490 ;
        RECT 745.215 1114.320 745.505 1114.490 ;
        RECT 745.675 1114.320 745.965 1114.490 ;
        RECT 746.135 1114.320 746.425 1114.490 ;
        RECT 746.595 1114.320 746.885 1114.490 ;
        RECT 747.055 1114.320 747.345 1114.490 ;
        RECT 747.515 1114.320 747.805 1114.490 ;
        RECT 747.975 1114.320 748.265 1114.490 ;
        RECT 748.435 1114.320 748.725 1114.490 ;
        RECT 748.895 1114.320 749.185 1114.490 ;
        RECT 749.355 1114.320 749.645 1114.490 ;
        RECT 749.815 1114.320 750.105 1114.490 ;
        RECT 750.275 1114.320 750.565 1114.490 ;
        RECT 750.735 1114.320 751.025 1114.490 ;
        RECT 751.195 1114.320 751.485 1114.490 ;
        RECT 751.655 1114.320 751.945 1114.490 ;
        RECT 752.115 1114.320 752.405 1114.490 ;
        RECT 752.575 1114.320 752.865 1114.490 ;
        RECT 753.035 1114.320 753.325 1114.490 ;
        RECT 753.495 1114.320 753.785 1114.490 ;
        RECT 753.955 1114.320 754.245 1114.490 ;
        RECT 754.415 1114.320 754.705 1114.490 ;
        RECT 754.875 1114.320 755.165 1114.490 ;
        RECT 755.335 1114.320 755.625 1114.490 ;
        RECT 755.795 1114.320 756.085 1114.490 ;
        RECT 756.255 1114.320 756.545 1114.490 ;
        RECT 756.715 1114.320 757.005 1114.490 ;
        RECT 757.175 1114.320 757.465 1114.490 ;
        RECT 757.635 1114.320 757.925 1114.490 ;
        RECT 758.095 1114.320 758.385 1114.490 ;
        RECT 758.555 1114.320 758.845 1114.490 ;
        RECT 759.015 1114.320 759.305 1114.490 ;
        RECT 759.475 1114.320 759.765 1114.490 ;
        RECT 759.935 1114.320 760.225 1114.490 ;
        RECT 760.395 1114.320 760.685 1114.490 ;
        RECT 760.855 1114.320 761.145 1114.490 ;
        RECT 761.315 1114.320 761.605 1114.490 ;
        RECT 761.775 1114.320 762.065 1114.490 ;
        RECT 762.235 1114.320 762.525 1114.490 ;
        RECT 762.695 1114.320 762.985 1114.490 ;
        RECT 763.155 1114.320 763.445 1114.490 ;
        RECT 763.615 1114.320 763.905 1114.490 ;
        RECT 764.075 1114.320 764.365 1114.490 ;
        RECT 764.535 1114.320 764.825 1114.490 ;
        RECT 764.995 1114.320 765.285 1114.490 ;
        RECT 765.455 1114.320 765.745 1114.490 ;
        RECT 765.915 1114.320 766.205 1114.490 ;
        RECT 766.375 1114.320 766.665 1114.490 ;
        RECT 766.835 1114.320 767.125 1114.490 ;
        RECT 767.295 1114.320 767.585 1114.490 ;
        RECT 767.755 1114.320 768.045 1114.490 ;
        RECT 768.215 1114.320 768.505 1114.490 ;
        RECT 768.675 1114.320 768.965 1114.490 ;
        RECT 769.135 1114.320 769.425 1114.490 ;
        RECT 769.595 1114.320 769.885 1114.490 ;
        RECT 770.055 1114.320 770.345 1114.490 ;
        RECT 770.515 1114.320 770.805 1114.490 ;
        RECT 770.975 1114.320 771.265 1114.490 ;
        RECT 771.435 1114.320 771.725 1114.490 ;
        RECT 771.895 1114.320 772.185 1114.490 ;
        RECT 772.355 1114.320 772.645 1114.490 ;
        RECT 772.815 1114.320 773.105 1114.490 ;
        RECT 773.275 1114.320 773.565 1114.490 ;
        RECT 773.735 1114.320 774.025 1114.490 ;
        RECT 774.195 1114.320 774.485 1114.490 ;
        RECT 774.655 1114.320 774.945 1114.490 ;
        RECT 775.115 1114.320 775.405 1114.490 ;
        RECT 775.575 1114.320 775.865 1114.490 ;
        RECT 776.035 1114.320 776.325 1114.490 ;
        RECT 776.495 1114.320 776.785 1114.490 ;
        RECT 776.955 1114.320 777.245 1114.490 ;
        RECT 777.415 1114.320 777.705 1114.490 ;
        RECT 777.875 1114.320 778.165 1114.490 ;
        RECT 778.335 1114.320 778.625 1114.490 ;
        RECT 778.795 1114.320 779.085 1114.490 ;
        RECT 779.255 1114.320 779.545 1114.490 ;
        RECT 779.715 1114.320 780.005 1114.490 ;
        RECT 780.175 1114.320 780.465 1114.490 ;
        RECT 780.635 1114.320 780.925 1114.490 ;
        RECT 781.095 1114.320 781.385 1114.490 ;
        RECT 781.555 1114.320 781.845 1114.490 ;
        RECT 782.015 1114.320 782.305 1114.490 ;
        RECT 782.475 1114.320 782.765 1114.490 ;
        RECT 782.935 1114.320 783.225 1114.490 ;
        RECT 783.395 1114.320 783.685 1114.490 ;
        RECT 783.855 1114.320 784.145 1114.490 ;
        RECT 784.315 1114.320 784.605 1114.490 ;
        RECT 784.775 1114.320 785.065 1114.490 ;
        RECT 785.235 1114.320 785.525 1114.490 ;
        RECT 785.695 1114.320 785.985 1114.490 ;
        RECT 786.155 1114.320 786.445 1114.490 ;
        RECT 786.615 1114.320 786.905 1114.490 ;
        RECT 787.075 1114.320 787.365 1114.490 ;
        RECT 787.535 1114.320 787.825 1114.490 ;
        RECT 787.995 1114.320 788.285 1114.490 ;
        RECT 788.455 1114.320 788.745 1114.490 ;
        RECT 788.915 1114.320 789.205 1114.490 ;
        RECT 789.375 1114.320 789.665 1114.490 ;
        RECT 789.835 1114.320 790.125 1114.490 ;
        RECT 790.295 1114.320 790.585 1114.490 ;
        RECT 790.755 1114.320 791.045 1114.490 ;
        RECT 791.215 1114.320 791.505 1114.490 ;
        RECT 791.675 1114.320 791.965 1114.490 ;
        RECT 792.135 1114.320 792.425 1114.490 ;
        RECT 792.595 1114.320 792.885 1114.490 ;
        RECT 793.055 1114.320 793.345 1114.490 ;
        RECT 793.515 1114.320 793.805 1114.490 ;
        RECT 793.975 1114.320 794.265 1114.490 ;
        RECT 794.435 1114.320 794.725 1114.490 ;
        RECT 794.895 1114.320 795.040 1114.490 ;
        RECT 1969.000 1114.320 1969.145 1114.490 ;
        RECT 1969.315 1114.320 1969.605 1114.490 ;
        RECT 1969.775 1114.320 1970.065 1114.490 ;
        RECT 1970.235 1114.320 1970.525 1114.490 ;
        RECT 1970.695 1114.320 1970.985 1114.490 ;
        RECT 1971.155 1114.320 1971.445 1114.490 ;
        RECT 1971.615 1114.320 1971.905 1114.490 ;
        RECT 1972.075 1114.320 1972.365 1114.490 ;
        RECT 1972.535 1114.320 1972.825 1114.490 ;
        RECT 1972.995 1114.320 1973.285 1114.490 ;
        RECT 1973.455 1114.320 1973.745 1114.490 ;
        RECT 1973.915 1114.320 1974.205 1114.490 ;
        RECT 1974.375 1114.320 1974.665 1114.490 ;
        RECT 1974.835 1114.320 1975.125 1114.490 ;
        RECT 1975.295 1114.320 1975.585 1114.490 ;
        RECT 1975.755 1114.320 1976.045 1114.490 ;
        RECT 1976.215 1114.320 1976.505 1114.490 ;
        RECT 1976.675 1114.320 1976.965 1114.490 ;
        RECT 1977.135 1114.320 1977.425 1114.490 ;
        RECT 1977.595 1114.320 1977.885 1114.490 ;
        RECT 1978.055 1114.320 1978.345 1114.490 ;
        RECT 1978.515 1114.320 1978.805 1114.490 ;
        RECT 1978.975 1114.320 1979.265 1114.490 ;
        RECT 1979.435 1114.320 1979.725 1114.490 ;
        RECT 1979.895 1114.320 1980.185 1114.490 ;
        RECT 1980.355 1114.320 1980.645 1114.490 ;
        RECT 1980.815 1114.320 1981.105 1114.490 ;
        RECT 1981.275 1114.320 1981.565 1114.490 ;
        RECT 1981.735 1114.320 1982.025 1114.490 ;
        RECT 1982.195 1114.320 1982.485 1114.490 ;
        RECT 1982.655 1114.320 1982.945 1114.490 ;
        RECT 1983.115 1114.320 1983.405 1114.490 ;
        RECT 1983.575 1114.320 1983.865 1114.490 ;
        RECT 1984.035 1114.320 1984.325 1114.490 ;
        RECT 1984.495 1114.320 1984.785 1114.490 ;
        RECT 1984.955 1114.320 1985.245 1114.490 ;
        RECT 1985.415 1114.320 1985.705 1114.490 ;
        RECT 1985.875 1114.320 1986.165 1114.490 ;
        RECT 1986.335 1114.320 1986.625 1114.490 ;
        RECT 1986.795 1114.320 1987.085 1114.490 ;
        RECT 1987.255 1114.320 1987.545 1114.490 ;
        RECT 1987.715 1114.320 1988.005 1114.490 ;
        RECT 1988.175 1114.320 1988.465 1114.490 ;
        RECT 1988.635 1114.320 1988.925 1114.490 ;
        RECT 1989.095 1114.320 1989.385 1114.490 ;
        RECT 1989.555 1114.320 1989.845 1114.490 ;
        RECT 1990.015 1114.320 1990.305 1114.490 ;
        RECT 1990.475 1114.320 1990.765 1114.490 ;
        RECT 1990.935 1114.320 1991.225 1114.490 ;
        RECT 1991.395 1114.320 1991.685 1114.490 ;
        RECT 1991.855 1114.320 1992.145 1114.490 ;
        RECT 1992.315 1114.320 1992.605 1114.490 ;
        RECT 1992.775 1114.320 1993.065 1114.490 ;
        RECT 1993.235 1114.320 1993.525 1114.490 ;
        RECT 1993.695 1114.320 1993.985 1114.490 ;
        RECT 1994.155 1114.320 1994.445 1114.490 ;
        RECT 1994.615 1114.320 1994.905 1114.490 ;
        RECT 1995.075 1114.320 1995.365 1114.490 ;
        RECT 1995.535 1114.320 1995.825 1114.490 ;
        RECT 1995.995 1114.320 1996.285 1114.490 ;
        RECT 1996.455 1114.320 1996.745 1114.490 ;
        RECT 1996.915 1114.320 1997.205 1114.490 ;
        RECT 1997.375 1114.320 1997.665 1114.490 ;
        RECT 1997.835 1114.320 1998.125 1114.490 ;
        RECT 1998.295 1114.320 1998.585 1114.490 ;
        RECT 1998.755 1114.320 1999.045 1114.490 ;
        RECT 1999.215 1114.320 1999.505 1114.490 ;
        RECT 1999.675 1114.320 1999.965 1114.490 ;
        RECT 2000.135 1114.320 2000.425 1114.490 ;
        RECT 2000.595 1114.320 2000.885 1114.490 ;
        RECT 2001.055 1114.320 2001.345 1114.490 ;
        RECT 2001.515 1114.320 2001.805 1114.490 ;
        RECT 2001.975 1114.320 2002.265 1114.490 ;
        RECT 2002.435 1114.320 2002.725 1114.490 ;
        RECT 2002.895 1114.320 2003.185 1114.490 ;
        RECT 2003.355 1114.320 2003.645 1114.490 ;
        RECT 2003.815 1114.320 2004.105 1114.490 ;
        RECT 2004.275 1114.320 2004.565 1114.490 ;
        RECT 2004.735 1114.320 2005.025 1114.490 ;
        RECT 2005.195 1114.320 2005.485 1114.490 ;
        RECT 2005.655 1114.320 2005.945 1114.490 ;
        RECT 2006.115 1114.320 2006.405 1114.490 ;
        RECT 2006.575 1114.320 2006.865 1114.490 ;
        RECT 2007.035 1114.320 2007.325 1114.490 ;
        RECT 2007.495 1114.320 2007.785 1114.490 ;
        RECT 2007.955 1114.320 2008.245 1114.490 ;
        RECT 2008.415 1114.320 2008.705 1114.490 ;
        RECT 2008.875 1114.320 2009.165 1114.490 ;
        RECT 2009.335 1114.320 2009.625 1114.490 ;
        RECT 2009.795 1114.320 2010.085 1114.490 ;
        RECT 2010.255 1114.320 2010.545 1114.490 ;
        RECT 2010.715 1114.320 2011.005 1114.490 ;
        RECT 2011.175 1114.320 2011.465 1114.490 ;
        RECT 2011.635 1114.320 2011.925 1114.490 ;
        RECT 2012.095 1114.320 2012.385 1114.490 ;
        RECT 2012.555 1114.320 2012.845 1114.490 ;
        RECT 2013.015 1114.320 2013.305 1114.490 ;
        RECT 2013.475 1114.320 2013.765 1114.490 ;
        RECT 2013.935 1114.320 2014.225 1114.490 ;
        RECT 2014.395 1114.320 2014.685 1114.490 ;
        RECT 2014.855 1114.320 2015.145 1114.490 ;
        RECT 2015.315 1114.320 2015.605 1114.490 ;
        RECT 2015.775 1114.320 2016.065 1114.490 ;
        RECT 2016.235 1114.320 2016.525 1114.490 ;
        RECT 2016.695 1114.320 2016.985 1114.490 ;
        RECT 2017.155 1114.320 2017.445 1114.490 ;
        RECT 2017.615 1114.320 2017.905 1114.490 ;
        RECT 2018.075 1114.320 2018.365 1114.490 ;
        RECT 2018.535 1114.320 2018.825 1114.490 ;
        RECT 2018.995 1114.320 2019.285 1114.490 ;
        RECT 2019.455 1114.320 2019.745 1114.490 ;
        RECT 2019.915 1114.320 2020.205 1114.490 ;
        RECT 2020.375 1114.320 2020.665 1114.490 ;
        RECT 2020.835 1114.320 2021.125 1114.490 ;
        RECT 2021.295 1114.320 2021.585 1114.490 ;
        RECT 2021.755 1114.320 2022.045 1114.490 ;
        RECT 2022.215 1114.320 2022.505 1114.490 ;
        RECT 2022.675 1114.320 2022.965 1114.490 ;
        RECT 2023.135 1114.320 2023.425 1114.490 ;
        RECT 2023.595 1114.320 2023.885 1114.490 ;
        RECT 2024.055 1114.320 2024.345 1114.490 ;
        RECT 2024.515 1114.320 2024.805 1114.490 ;
        RECT 2024.975 1114.320 2025.265 1114.490 ;
        RECT 2025.435 1114.320 2025.725 1114.490 ;
        RECT 2025.895 1114.320 2026.185 1114.490 ;
        RECT 2026.355 1114.320 2026.645 1114.490 ;
        RECT 2026.815 1114.320 2027.105 1114.490 ;
        RECT 2027.275 1114.320 2027.565 1114.490 ;
        RECT 2027.735 1114.320 2028.025 1114.490 ;
        RECT 2028.195 1114.320 2028.485 1114.490 ;
        RECT 2028.655 1114.320 2028.945 1114.490 ;
        RECT 2029.115 1114.320 2029.405 1114.490 ;
        RECT 2029.575 1114.320 2029.865 1114.490 ;
        RECT 2030.035 1114.320 2030.325 1114.490 ;
        RECT 2030.495 1114.320 2030.785 1114.490 ;
        RECT 2030.955 1114.320 2031.245 1114.490 ;
        RECT 2031.415 1114.320 2031.705 1114.490 ;
        RECT 2031.875 1114.320 2032.165 1114.490 ;
        RECT 2032.335 1114.320 2032.625 1114.490 ;
        RECT 2032.795 1114.320 2033.085 1114.490 ;
        RECT 2033.255 1114.320 2033.545 1114.490 ;
        RECT 2033.715 1114.320 2034.005 1114.490 ;
        RECT 2034.175 1114.320 2034.465 1114.490 ;
        RECT 2034.635 1114.320 2034.925 1114.490 ;
        RECT 2035.095 1114.320 2035.385 1114.490 ;
        RECT 2035.555 1114.320 2035.845 1114.490 ;
        RECT 2036.015 1114.320 2036.305 1114.490 ;
        RECT 2036.475 1114.320 2036.765 1114.490 ;
        RECT 2036.935 1114.320 2037.225 1114.490 ;
        RECT 2037.395 1114.320 2037.685 1114.490 ;
        RECT 2037.855 1114.320 2038.145 1114.490 ;
        RECT 2038.315 1114.320 2038.605 1114.490 ;
        RECT 2038.775 1114.320 2039.065 1114.490 ;
        RECT 2039.235 1114.320 2039.525 1114.490 ;
        RECT 2039.695 1114.320 2039.985 1114.490 ;
        RECT 2040.155 1114.320 2040.445 1114.490 ;
        RECT 2040.615 1114.320 2040.905 1114.490 ;
        RECT 2041.075 1114.320 2041.365 1114.490 ;
        RECT 2041.535 1114.320 2041.825 1114.490 ;
        RECT 2041.995 1114.320 2042.285 1114.490 ;
        RECT 2042.455 1114.320 2042.745 1114.490 ;
        RECT 2042.915 1114.320 2043.205 1114.490 ;
        RECT 2043.375 1114.320 2043.665 1114.490 ;
        RECT 2043.835 1114.320 2044.125 1114.490 ;
        RECT 2044.295 1114.320 2044.585 1114.490 ;
        RECT 2044.755 1114.320 2045.045 1114.490 ;
        RECT 2045.215 1114.320 2045.505 1114.490 ;
        RECT 2045.675 1114.320 2045.965 1114.490 ;
        RECT 2046.135 1114.320 2046.425 1114.490 ;
        RECT 2046.595 1114.320 2046.885 1114.490 ;
        RECT 2047.055 1114.320 2047.345 1114.490 ;
        RECT 2047.515 1114.320 2047.805 1114.490 ;
        RECT 2047.975 1114.320 2048.265 1114.490 ;
        RECT 2048.435 1114.320 2048.725 1114.490 ;
        RECT 2048.895 1114.320 2049.185 1114.490 ;
        RECT 2049.355 1114.320 2049.645 1114.490 ;
        RECT 2049.815 1114.320 2050.105 1114.490 ;
        RECT 2050.275 1114.320 2050.565 1114.490 ;
        RECT 2050.735 1114.320 2051.025 1114.490 ;
        RECT 2051.195 1114.320 2051.485 1114.490 ;
        RECT 2051.655 1114.320 2051.945 1114.490 ;
        RECT 2052.115 1114.320 2052.405 1114.490 ;
        RECT 2052.575 1114.320 2052.865 1114.490 ;
        RECT 2053.035 1114.320 2053.325 1114.490 ;
        RECT 2053.495 1114.320 2053.785 1114.490 ;
        RECT 2053.955 1114.320 2054.245 1114.490 ;
        RECT 2054.415 1114.320 2054.705 1114.490 ;
        RECT 2054.875 1114.320 2055.165 1114.490 ;
        RECT 2055.335 1114.320 2055.625 1114.490 ;
        RECT 2055.795 1114.320 2056.085 1114.490 ;
        RECT 2056.255 1114.320 2056.545 1114.490 ;
        RECT 2056.715 1114.320 2057.005 1114.490 ;
        RECT 2057.175 1114.320 2057.465 1114.490 ;
        RECT 2057.635 1114.320 2057.925 1114.490 ;
        RECT 2058.095 1114.320 2058.385 1114.490 ;
        RECT 2058.555 1114.320 2058.845 1114.490 ;
        RECT 2059.015 1114.320 2059.305 1114.490 ;
        RECT 2059.475 1114.320 2059.765 1114.490 ;
        RECT 2059.935 1114.320 2060.225 1114.490 ;
        RECT 2060.395 1114.320 2060.685 1114.490 ;
        RECT 2060.855 1114.320 2061.145 1114.490 ;
        RECT 2061.315 1114.320 2061.605 1114.490 ;
        RECT 2061.775 1114.320 2062.065 1114.490 ;
        RECT 2062.235 1114.320 2062.525 1114.490 ;
        RECT 2062.695 1114.320 2062.985 1114.490 ;
        RECT 2063.155 1114.320 2063.445 1114.490 ;
        RECT 2063.615 1114.320 2063.905 1114.490 ;
        RECT 2064.075 1114.320 2064.365 1114.490 ;
        RECT 2064.535 1114.320 2064.825 1114.490 ;
        RECT 2064.995 1114.320 2065.285 1114.490 ;
        RECT 2065.455 1114.320 2065.745 1114.490 ;
        RECT 2065.915 1114.320 2066.205 1114.490 ;
        RECT 2066.375 1114.320 2066.665 1114.490 ;
        RECT 2066.835 1114.320 2067.125 1114.490 ;
        RECT 2067.295 1114.320 2067.585 1114.490 ;
        RECT 2067.755 1114.320 2068.045 1114.490 ;
        RECT 2068.215 1114.320 2068.505 1114.490 ;
        RECT 2068.675 1114.320 2068.965 1114.490 ;
        RECT 2069.135 1114.320 2069.425 1114.490 ;
        RECT 2069.595 1114.320 2069.885 1114.490 ;
        RECT 2070.055 1114.320 2070.345 1114.490 ;
        RECT 2070.515 1114.320 2070.805 1114.490 ;
        RECT 2070.975 1114.320 2071.265 1114.490 ;
        RECT 2071.435 1114.320 2071.725 1114.490 ;
        RECT 2071.895 1114.320 2072.185 1114.490 ;
        RECT 2072.355 1114.320 2072.645 1114.490 ;
        RECT 2072.815 1114.320 2073.105 1114.490 ;
        RECT 2073.275 1114.320 2073.565 1114.490 ;
        RECT 2073.735 1114.320 2074.025 1114.490 ;
        RECT 2074.195 1114.320 2074.485 1114.490 ;
        RECT 2074.655 1114.320 2074.945 1114.490 ;
        RECT 2075.115 1114.320 2075.405 1114.490 ;
        RECT 2075.575 1114.320 2075.865 1114.490 ;
        RECT 2076.035 1114.320 2076.325 1114.490 ;
        RECT 2076.495 1114.320 2076.785 1114.490 ;
        RECT 2076.955 1114.320 2077.245 1114.490 ;
        RECT 2077.415 1114.320 2077.705 1114.490 ;
        RECT 2077.875 1114.320 2078.165 1114.490 ;
        RECT 2078.335 1114.320 2078.625 1114.490 ;
        RECT 2078.795 1114.320 2079.085 1114.490 ;
        RECT 2079.255 1114.320 2079.545 1114.490 ;
        RECT 2079.715 1114.320 2080.005 1114.490 ;
        RECT 2080.175 1114.320 2080.465 1114.490 ;
        RECT 2080.635 1114.320 2080.925 1114.490 ;
        RECT 2081.095 1114.320 2081.385 1114.490 ;
        RECT 2081.555 1114.320 2081.845 1114.490 ;
        RECT 2082.015 1114.320 2082.305 1114.490 ;
        RECT 2082.475 1114.320 2082.765 1114.490 ;
        RECT 2082.935 1114.320 2083.225 1114.490 ;
        RECT 2083.395 1114.320 2083.685 1114.490 ;
        RECT 2083.855 1114.320 2084.145 1114.490 ;
        RECT 2084.315 1114.320 2084.605 1114.490 ;
        RECT 2084.775 1114.320 2085.065 1114.490 ;
        RECT 2085.235 1114.320 2085.525 1114.490 ;
        RECT 2085.695 1114.320 2085.985 1114.490 ;
        RECT 2086.155 1114.320 2086.445 1114.490 ;
        RECT 2086.615 1114.320 2086.905 1114.490 ;
        RECT 2087.075 1114.320 2087.365 1114.490 ;
        RECT 2087.535 1114.320 2087.825 1114.490 ;
        RECT 2087.995 1114.320 2088.285 1114.490 ;
        RECT 2088.455 1114.320 2088.745 1114.490 ;
        RECT 2088.915 1114.320 2089.205 1114.490 ;
        RECT 2089.375 1114.320 2089.665 1114.490 ;
        RECT 2089.835 1114.320 2090.125 1114.490 ;
        RECT 2090.295 1114.320 2090.585 1114.490 ;
        RECT 2090.755 1114.320 2091.045 1114.490 ;
        RECT 2091.215 1114.320 2091.505 1114.490 ;
        RECT 2091.675 1114.320 2091.965 1114.490 ;
        RECT 2092.135 1114.320 2092.425 1114.490 ;
        RECT 2092.595 1114.320 2092.885 1114.490 ;
        RECT 2093.055 1114.320 2093.345 1114.490 ;
        RECT 2093.515 1114.320 2093.805 1114.490 ;
        RECT 2093.975 1114.320 2094.265 1114.490 ;
        RECT 2094.435 1114.320 2094.725 1114.490 ;
        RECT 2094.895 1114.320 2095.040 1114.490 ;
        RECT 675.065 1113.155 675.355 1114.320 ;
        RECT 675.535 1113.300 675.865 1114.150 ;
        RECT 676.035 1113.520 676.205 1114.320 ;
        RECT 676.375 1113.300 676.705 1114.150 ;
        RECT 676.875 1113.520 677.045 1114.320 ;
      LAYER li1 ;
        RECT 677.295 1113.300 677.465 1114.150 ;
      LAYER li1 ;
        RECT 677.635 1113.520 677.965 1114.320 ;
      LAYER li1 ;
        RECT 678.135 1113.300 678.305 1114.150 ;
      LAYER li1 ;
        RECT 678.475 1113.520 678.805 1114.320 ;
      LAYER li1 ;
        RECT 678.975 1113.300 679.145 1114.150 ;
      LAYER li1 ;
        RECT 679.315 1113.520 679.645 1114.320 ;
      LAYER li1 ;
        RECT 679.815 1113.300 679.985 1114.150 ;
      LAYER li1 ;
        RECT 675.535 1113.130 677.035 1113.300 ;
      LAYER li1 ;
        RECT 677.295 1113.130 679.985 1113.300 ;
      LAYER li1 ;
        RECT 680.155 1113.170 680.485 1114.320 ;
        RECT 681.045 1113.155 681.335 1114.320 ;
        RECT 681.515 1113.300 681.845 1114.150 ;
        RECT 682.015 1113.520 682.185 1114.320 ;
        RECT 682.355 1113.300 682.685 1114.150 ;
        RECT 682.855 1113.520 683.025 1114.320 ;
      LAYER li1 ;
        RECT 683.275 1113.300 683.445 1114.150 ;
      LAYER li1 ;
        RECT 683.615 1113.520 683.945 1114.320 ;
      LAYER li1 ;
        RECT 684.115 1113.300 684.285 1114.150 ;
      LAYER li1 ;
        RECT 684.455 1113.520 684.785 1114.320 ;
      LAYER li1 ;
        RECT 684.955 1113.300 685.125 1114.150 ;
      LAYER li1 ;
        RECT 685.295 1113.520 685.625 1114.320 ;
      LAYER li1 ;
        RECT 685.795 1113.300 685.965 1114.150 ;
      LAYER li1 ;
        RECT 681.515 1113.130 683.015 1113.300 ;
      LAYER li1 ;
        RECT 683.275 1113.130 685.965 1113.300 ;
      LAYER li1 ;
        RECT 686.135 1113.170 686.465 1114.320 ;
        RECT 687.025 1113.155 687.315 1114.320 ;
        RECT 687.495 1113.300 687.825 1114.150 ;
        RECT 687.995 1113.520 688.165 1114.320 ;
        RECT 688.335 1113.300 688.665 1114.150 ;
        RECT 688.835 1113.520 689.005 1114.320 ;
      LAYER li1 ;
        RECT 689.255 1113.300 689.425 1114.150 ;
      LAYER li1 ;
        RECT 689.595 1113.520 689.925 1114.320 ;
      LAYER li1 ;
        RECT 690.095 1113.300 690.265 1114.150 ;
      LAYER li1 ;
        RECT 690.435 1113.520 690.765 1114.320 ;
      LAYER li1 ;
        RECT 690.935 1113.300 691.105 1114.150 ;
      LAYER li1 ;
        RECT 691.275 1113.520 691.605 1114.320 ;
      LAYER li1 ;
        RECT 691.775 1113.300 691.945 1114.150 ;
      LAYER li1 ;
        RECT 687.495 1113.130 688.995 1113.300 ;
      LAYER li1 ;
        RECT 689.255 1113.130 691.945 1113.300 ;
      LAYER li1 ;
        RECT 692.115 1113.170 692.445 1114.320 ;
        RECT 693.005 1113.155 693.295 1114.320 ;
        RECT 693.475 1113.300 693.805 1114.150 ;
        RECT 693.975 1113.520 694.145 1114.320 ;
        RECT 694.315 1113.300 694.645 1114.150 ;
        RECT 694.815 1113.520 694.985 1114.320 ;
      LAYER li1 ;
        RECT 695.235 1113.300 695.405 1114.150 ;
      LAYER li1 ;
        RECT 695.575 1113.520 695.905 1114.320 ;
      LAYER li1 ;
        RECT 696.075 1113.300 696.245 1114.150 ;
      LAYER li1 ;
        RECT 696.415 1113.520 696.745 1114.320 ;
      LAYER li1 ;
        RECT 696.915 1113.300 697.085 1114.150 ;
      LAYER li1 ;
        RECT 697.255 1113.520 697.585 1114.320 ;
      LAYER li1 ;
        RECT 697.755 1113.300 697.925 1114.150 ;
      LAYER li1 ;
        RECT 693.475 1113.130 694.975 1113.300 ;
      LAYER li1 ;
        RECT 695.235 1113.130 697.925 1113.300 ;
      LAYER li1 ;
        RECT 698.095 1113.170 698.425 1114.320 ;
        RECT 698.985 1113.155 699.275 1114.320 ;
        RECT 699.455 1113.300 699.785 1114.150 ;
        RECT 699.955 1113.520 700.125 1114.320 ;
        RECT 700.295 1113.300 700.625 1114.150 ;
        RECT 700.795 1113.520 700.965 1114.320 ;
      LAYER li1 ;
        RECT 701.215 1113.300 701.385 1114.150 ;
      LAYER li1 ;
        RECT 701.555 1113.520 701.885 1114.320 ;
      LAYER li1 ;
        RECT 702.055 1113.300 702.225 1114.150 ;
      LAYER li1 ;
        RECT 702.395 1113.520 702.725 1114.320 ;
      LAYER li1 ;
        RECT 702.895 1113.300 703.065 1114.150 ;
      LAYER li1 ;
        RECT 703.235 1113.520 703.565 1114.320 ;
      LAYER li1 ;
        RECT 703.735 1113.300 703.905 1114.150 ;
      LAYER li1 ;
        RECT 699.455 1113.130 700.955 1113.300 ;
      LAYER li1 ;
        RECT 701.215 1113.130 703.905 1113.300 ;
      LAYER li1 ;
        RECT 704.075 1113.170 704.405 1114.320 ;
        RECT 704.965 1113.155 705.255 1114.320 ;
        RECT 705.435 1113.300 705.765 1114.150 ;
        RECT 705.935 1113.520 706.105 1114.320 ;
        RECT 706.275 1113.300 706.605 1114.150 ;
        RECT 706.775 1113.520 706.945 1114.320 ;
      LAYER li1 ;
        RECT 707.195 1113.300 707.365 1114.150 ;
      LAYER li1 ;
        RECT 707.535 1113.520 707.865 1114.320 ;
      LAYER li1 ;
        RECT 708.035 1113.300 708.205 1114.150 ;
      LAYER li1 ;
        RECT 708.375 1113.520 708.705 1114.320 ;
      LAYER li1 ;
        RECT 708.875 1113.300 709.045 1114.150 ;
      LAYER li1 ;
        RECT 709.215 1113.520 709.545 1114.320 ;
      LAYER li1 ;
        RECT 709.715 1113.300 709.885 1114.150 ;
      LAYER li1 ;
        RECT 705.435 1113.130 706.935 1113.300 ;
      LAYER li1 ;
        RECT 707.195 1113.130 709.885 1113.300 ;
      LAYER li1 ;
        RECT 710.055 1113.170 710.385 1114.320 ;
        RECT 710.945 1113.155 711.235 1114.320 ;
        RECT 711.415 1113.300 711.745 1114.150 ;
        RECT 711.915 1113.520 712.085 1114.320 ;
        RECT 712.255 1113.300 712.585 1114.150 ;
        RECT 712.755 1113.520 712.925 1114.320 ;
      LAYER li1 ;
        RECT 713.175 1113.300 713.345 1114.150 ;
      LAYER li1 ;
        RECT 713.515 1113.520 713.845 1114.320 ;
      LAYER li1 ;
        RECT 714.015 1113.300 714.185 1114.150 ;
      LAYER li1 ;
        RECT 714.355 1113.520 714.685 1114.320 ;
      LAYER li1 ;
        RECT 714.855 1113.300 715.025 1114.150 ;
      LAYER li1 ;
        RECT 715.195 1113.520 715.525 1114.320 ;
      LAYER li1 ;
        RECT 715.695 1113.300 715.865 1114.150 ;
      LAYER li1 ;
        RECT 711.415 1113.130 712.915 1113.300 ;
      LAYER li1 ;
        RECT 713.175 1113.130 715.865 1113.300 ;
      LAYER li1 ;
        RECT 716.035 1113.170 716.365 1114.320 ;
        RECT 716.925 1113.155 717.215 1114.320 ;
        RECT 717.395 1113.300 717.725 1114.150 ;
        RECT 717.895 1113.520 718.065 1114.320 ;
        RECT 718.235 1113.300 718.565 1114.150 ;
        RECT 718.735 1113.520 718.905 1114.320 ;
      LAYER li1 ;
        RECT 719.155 1113.300 719.325 1114.150 ;
      LAYER li1 ;
        RECT 719.495 1113.520 719.825 1114.320 ;
      LAYER li1 ;
        RECT 719.995 1113.300 720.165 1114.150 ;
      LAYER li1 ;
        RECT 720.335 1113.520 720.665 1114.320 ;
      LAYER li1 ;
        RECT 720.835 1113.300 721.005 1114.150 ;
      LAYER li1 ;
        RECT 721.175 1113.520 721.505 1114.320 ;
      LAYER li1 ;
        RECT 721.675 1113.300 721.845 1114.150 ;
      LAYER li1 ;
        RECT 717.395 1113.130 718.895 1113.300 ;
      LAYER li1 ;
        RECT 719.155 1113.130 721.845 1113.300 ;
      LAYER li1 ;
        RECT 722.015 1113.170 722.345 1114.320 ;
        RECT 722.905 1113.155 723.195 1114.320 ;
        RECT 723.375 1113.300 723.705 1114.150 ;
        RECT 723.875 1113.520 724.045 1114.320 ;
        RECT 724.215 1113.300 724.545 1114.150 ;
        RECT 724.715 1113.520 724.885 1114.320 ;
      LAYER li1 ;
        RECT 725.135 1113.300 725.305 1114.150 ;
      LAYER li1 ;
        RECT 725.475 1113.520 725.805 1114.320 ;
      LAYER li1 ;
        RECT 725.975 1113.300 726.145 1114.150 ;
      LAYER li1 ;
        RECT 726.315 1113.520 726.645 1114.320 ;
      LAYER li1 ;
        RECT 726.815 1113.300 726.985 1114.150 ;
      LAYER li1 ;
        RECT 727.155 1113.520 727.485 1114.320 ;
      LAYER li1 ;
        RECT 727.655 1113.300 727.825 1114.150 ;
      LAYER li1 ;
        RECT 723.375 1113.130 724.875 1113.300 ;
      LAYER li1 ;
        RECT 725.135 1113.130 727.825 1113.300 ;
      LAYER li1 ;
        RECT 727.995 1113.170 728.325 1114.320 ;
        RECT 728.885 1113.155 729.175 1114.320 ;
        RECT 729.355 1113.300 729.685 1114.150 ;
        RECT 729.855 1113.520 730.025 1114.320 ;
        RECT 730.195 1113.300 730.525 1114.150 ;
        RECT 730.695 1113.520 730.865 1114.320 ;
      LAYER li1 ;
        RECT 731.115 1113.300 731.285 1114.150 ;
      LAYER li1 ;
        RECT 731.455 1113.520 731.785 1114.320 ;
      LAYER li1 ;
        RECT 731.955 1113.300 732.125 1114.150 ;
      LAYER li1 ;
        RECT 732.295 1113.520 732.625 1114.320 ;
      LAYER li1 ;
        RECT 732.795 1113.300 732.965 1114.150 ;
      LAYER li1 ;
        RECT 733.135 1113.520 733.465 1114.320 ;
      LAYER li1 ;
        RECT 733.635 1113.300 733.805 1114.150 ;
      LAYER li1 ;
        RECT 729.355 1113.130 730.855 1113.300 ;
      LAYER li1 ;
        RECT 731.115 1113.130 733.805 1113.300 ;
      LAYER li1 ;
        RECT 733.975 1113.170 734.305 1114.320 ;
        RECT 734.865 1113.155 735.155 1114.320 ;
        RECT 735.335 1113.300 735.665 1114.150 ;
        RECT 735.835 1113.520 736.005 1114.320 ;
        RECT 736.175 1113.300 736.505 1114.150 ;
        RECT 736.675 1113.520 736.845 1114.320 ;
      LAYER li1 ;
        RECT 737.095 1113.300 737.265 1114.150 ;
      LAYER li1 ;
        RECT 737.435 1113.520 737.765 1114.320 ;
      LAYER li1 ;
        RECT 737.935 1113.300 738.105 1114.150 ;
      LAYER li1 ;
        RECT 738.275 1113.520 738.605 1114.320 ;
      LAYER li1 ;
        RECT 738.775 1113.300 738.945 1114.150 ;
      LAYER li1 ;
        RECT 739.115 1113.520 739.445 1114.320 ;
      LAYER li1 ;
        RECT 739.615 1113.300 739.785 1114.150 ;
      LAYER li1 ;
        RECT 735.335 1113.130 736.835 1113.300 ;
      LAYER li1 ;
        RECT 737.095 1113.130 739.785 1113.300 ;
      LAYER li1 ;
        RECT 739.955 1113.170 740.285 1114.320 ;
        RECT 740.845 1113.155 741.135 1114.320 ;
        RECT 741.315 1113.300 741.645 1114.150 ;
        RECT 741.815 1113.520 741.985 1114.320 ;
        RECT 742.155 1113.300 742.485 1114.150 ;
        RECT 742.655 1113.520 742.825 1114.320 ;
      LAYER li1 ;
        RECT 743.075 1113.300 743.245 1114.150 ;
      LAYER li1 ;
        RECT 743.415 1113.520 743.745 1114.320 ;
      LAYER li1 ;
        RECT 743.915 1113.300 744.085 1114.150 ;
      LAYER li1 ;
        RECT 744.255 1113.520 744.585 1114.320 ;
      LAYER li1 ;
        RECT 744.755 1113.300 744.925 1114.150 ;
      LAYER li1 ;
        RECT 745.095 1113.520 745.425 1114.320 ;
      LAYER li1 ;
        RECT 745.595 1113.300 745.765 1114.150 ;
      LAYER li1 ;
        RECT 741.315 1113.130 742.815 1113.300 ;
      LAYER li1 ;
        RECT 743.075 1113.130 745.765 1113.300 ;
      LAYER li1 ;
        RECT 745.935 1113.170 746.265 1114.320 ;
        RECT 746.825 1113.155 747.115 1114.320 ;
        RECT 747.295 1113.300 747.625 1114.150 ;
        RECT 747.795 1113.520 747.965 1114.320 ;
        RECT 748.135 1113.300 748.465 1114.150 ;
        RECT 748.635 1113.520 748.805 1114.320 ;
      LAYER li1 ;
        RECT 749.055 1113.300 749.225 1114.150 ;
      LAYER li1 ;
        RECT 749.395 1113.520 749.725 1114.320 ;
      LAYER li1 ;
        RECT 749.895 1113.300 750.065 1114.150 ;
      LAYER li1 ;
        RECT 750.235 1113.520 750.565 1114.320 ;
      LAYER li1 ;
        RECT 750.735 1113.300 750.905 1114.150 ;
      LAYER li1 ;
        RECT 751.075 1113.520 751.405 1114.320 ;
      LAYER li1 ;
        RECT 751.575 1113.300 751.745 1114.150 ;
      LAYER li1 ;
        RECT 747.295 1113.130 748.795 1113.300 ;
      LAYER li1 ;
        RECT 749.055 1113.130 751.745 1113.300 ;
      LAYER li1 ;
        RECT 751.915 1113.170 752.245 1114.320 ;
        RECT 752.805 1113.155 753.095 1114.320 ;
        RECT 753.275 1113.300 753.605 1114.150 ;
        RECT 753.775 1113.520 753.945 1114.320 ;
        RECT 754.115 1113.300 754.445 1114.150 ;
        RECT 754.615 1113.520 754.785 1114.320 ;
      LAYER li1 ;
        RECT 755.035 1113.300 755.205 1114.150 ;
      LAYER li1 ;
        RECT 755.375 1113.520 755.705 1114.320 ;
      LAYER li1 ;
        RECT 755.875 1113.300 756.045 1114.150 ;
      LAYER li1 ;
        RECT 756.215 1113.520 756.545 1114.320 ;
      LAYER li1 ;
        RECT 756.715 1113.300 756.885 1114.150 ;
      LAYER li1 ;
        RECT 757.055 1113.520 757.385 1114.320 ;
      LAYER li1 ;
        RECT 757.555 1113.300 757.725 1114.150 ;
      LAYER li1 ;
        RECT 753.275 1113.130 754.775 1113.300 ;
      LAYER li1 ;
        RECT 755.035 1113.130 757.725 1113.300 ;
      LAYER li1 ;
        RECT 757.895 1113.170 758.225 1114.320 ;
        RECT 758.785 1113.155 759.075 1114.320 ;
        RECT 759.255 1113.300 759.585 1114.150 ;
        RECT 759.755 1113.520 759.925 1114.320 ;
        RECT 760.095 1113.300 760.425 1114.150 ;
        RECT 760.595 1113.520 760.765 1114.320 ;
      LAYER li1 ;
        RECT 761.015 1113.300 761.185 1114.150 ;
      LAYER li1 ;
        RECT 761.355 1113.520 761.685 1114.320 ;
      LAYER li1 ;
        RECT 761.855 1113.300 762.025 1114.150 ;
      LAYER li1 ;
        RECT 762.195 1113.520 762.525 1114.320 ;
      LAYER li1 ;
        RECT 762.695 1113.300 762.865 1114.150 ;
      LAYER li1 ;
        RECT 763.035 1113.520 763.365 1114.320 ;
      LAYER li1 ;
        RECT 763.535 1113.300 763.705 1114.150 ;
      LAYER li1 ;
        RECT 759.255 1113.130 760.755 1113.300 ;
      LAYER li1 ;
        RECT 761.015 1113.130 763.705 1113.300 ;
      LAYER li1 ;
        RECT 763.875 1113.170 764.205 1114.320 ;
        RECT 764.765 1113.155 765.055 1114.320 ;
        RECT 765.235 1113.300 765.565 1114.150 ;
        RECT 765.735 1113.520 765.905 1114.320 ;
        RECT 766.075 1113.300 766.405 1114.150 ;
        RECT 766.575 1113.520 766.745 1114.320 ;
      LAYER li1 ;
        RECT 766.995 1113.300 767.165 1114.150 ;
      LAYER li1 ;
        RECT 767.335 1113.520 767.665 1114.320 ;
      LAYER li1 ;
        RECT 767.835 1113.300 768.005 1114.150 ;
      LAYER li1 ;
        RECT 768.175 1113.520 768.505 1114.320 ;
      LAYER li1 ;
        RECT 768.675 1113.300 768.845 1114.150 ;
      LAYER li1 ;
        RECT 769.015 1113.520 769.345 1114.320 ;
      LAYER li1 ;
        RECT 769.515 1113.300 769.685 1114.150 ;
      LAYER li1 ;
        RECT 765.235 1113.130 766.735 1113.300 ;
      LAYER li1 ;
        RECT 766.995 1113.130 769.685 1113.300 ;
      LAYER li1 ;
        RECT 769.855 1113.170 770.185 1114.320 ;
        RECT 770.745 1113.155 771.035 1114.320 ;
        RECT 771.215 1113.300 771.545 1114.150 ;
        RECT 771.715 1113.520 771.885 1114.320 ;
        RECT 772.055 1113.300 772.385 1114.150 ;
        RECT 772.555 1113.520 772.725 1114.320 ;
      LAYER li1 ;
        RECT 772.975 1113.300 773.145 1114.150 ;
      LAYER li1 ;
        RECT 773.315 1113.520 773.645 1114.320 ;
      LAYER li1 ;
        RECT 773.815 1113.300 773.985 1114.150 ;
      LAYER li1 ;
        RECT 774.155 1113.520 774.485 1114.320 ;
      LAYER li1 ;
        RECT 774.655 1113.300 774.825 1114.150 ;
      LAYER li1 ;
        RECT 774.995 1113.520 775.325 1114.320 ;
      LAYER li1 ;
        RECT 775.495 1113.300 775.665 1114.150 ;
      LAYER li1 ;
        RECT 771.215 1113.130 772.715 1113.300 ;
      LAYER li1 ;
        RECT 772.975 1113.130 775.665 1113.300 ;
      LAYER li1 ;
        RECT 775.835 1113.170 776.165 1114.320 ;
        RECT 776.725 1113.155 777.015 1114.320 ;
        RECT 777.195 1113.300 777.525 1114.150 ;
        RECT 777.695 1113.520 777.865 1114.320 ;
        RECT 778.035 1113.300 778.365 1114.150 ;
        RECT 778.535 1113.520 778.705 1114.320 ;
      LAYER li1 ;
        RECT 778.955 1113.300 779.125 1114.150 ;
      LAYER li1 ;
        RECT 779.295 1113.520 779.625 1114.320 ;
      LAYER li1 ;
        RECT 779.795 1113.300 779.965 1114.150 ;
      LAYER li1 ;
        RECT 780.135 1113.520 780.465 1114.320 ;
      LAYER li1 ;
        RECT 780.635 1113.300 780.805 1114.150 ;
      LAYER li1 ;
        RECT 780.975 1113.520 781.305 1114.320 ;
      LAYER li1 ;
        RECT 781.475 1113.300 781.645 1114.150 ;
      LAYER li1 ;
        RECT 777.195 1113.130 778.695 1113.300 ;
      LAYER li1 ;
        RECT 778.955 1113.130 781.645 1113.300 ;
      LAYER li1 ;
        RECT 781.815 1113.170 782.145 1114.320 ;
        RECT 782.705 1113.155 782.995 1114.320 ;
        RECT 783.175 1113.300 783.505 1114.150 ;
        RECT 783.675 1113.520 783.845 1114.320 ;
        RECT 784.015 1113.300 784.345 1114.150 ;
        RECT 784.515 1113.520 784.685 1114.320 ;
      LAYER li1 ;
        RECT 784.935 1113.300 785.105 1114.150 ;
      LAYER li1 ;
        RECT 785.275 1113.520 785.605 1114.320 ;
      LAYER li1 ;
        RECT 785.775 1113.300 785.945 1114.150 ;
      LAYER li1 ;
        RECT 786.115 1113.520 786.445 1114.320 ;
      LAYER li1 ;
        RECT 786.615 1113.300 786.785 1114.150 ;
      LAYER li1 ;
        RECT 786.955 1113.520 787.285 1114.320 ;
      LAYER li1 ;
        RECT 787.455 1113.300 787.625 1114.150 ;
      LAYER li1 ;
        RECT 783.175 1113.130 784.675 1113.300 ;
      LAYER li1 ;
        RECT 784.935 1113.130 787.625 1113.300 ;
      LAYER li1 ;
        RECT 787.795 1113.170 788.125 1114.320 ;
        RECT 788.685 1113.155 788.975 1114.320 ;
        RECT 789.535 1113.170 789.865 1114.320 ;
        RECT 790.375 1113.520 790.705 1114.320 ;
        RECT 791.215 1113.520 791.545 1114.320 ;
        RECT 792.055 1113.520 792.385 1114.320 ;
        RECT 792.975 1113.520 793.145 1114.320 ;
        RECT 793.315 1113.300 793.645 1114.150 ;
        RECT 793.815 1113.520 793.985 1114.320 ;
        RECT 794.155 1113.300 794.485 1114.150 ;
      LAYER li1 ;
        RECT 675.580 1112.760 676.680 1112.960 ;
      LAYER li1 ;
        RECT 676.860 1112.930 677.035 1113.130 ;
        RECT 676.860 1112.760 679.485 1112.930 ;
        RECT 676.860 1112.590 677.035 1112.760 ;
      LAYER li1 ;
        RECT 679.730 1112.590 679.985 1113.130 ;
        RECT 681.560 1112.760 682.660 1112.960 ;
      LAYER li1 ;
        RECT 682.840 1112.930 683.015 1113.130 ;
        RECT 682.840 1112.760 685.465 1112.930 ;
        RECT 682.840 1112.590 683.015 1112.760 ;
      LAYER li1 ;
        RECT 685.710 1112.590 685.965 1113.130 ;
        RECT 687.540 1112.760 688.640 1112.960 ;
      LAYER li1 ;
        RECT 688.820 1112.930 688.995 1113.130 ;
        RECT 688.820 1112.760 691.445 1112.930 ;
        RECT 688.820 1112.590 688.995 1112.760 ;
      LAYER li1 ;
        RECT 691.690 1112.590 691.945 1113.130 ;
        RECT 693.520 1112.760 694.620 1112.960 ;
      LAYER li1 ;
        RECT 694.800 1112.930 694.975 1113.130 ;
        RECT 694.800 1112.760 697.425 1112.930 ;
        RECT 694.800 1112.590 694.975 1112.760 ;
      LAYER li1 ;
        RECT 697.670 1112.590 697.925 1113.130 ;
        RECT 699.500 1112.760 700.600 1112.960 ;
      LAYER li1 ;
        RECT 700.780 1112.930 700.955 1113.130 ;
        RECT 700.780 1112.760 703.405 1112.930 ;
        RECT 700.780 1112.590 700.955 1112.760 ;
      LAYER li1 ;
        RECT 703.650 1112.590 703.905 1113.130 ;
        RECT 705.480 1112.760 706.580 1112.960 ;
      LAYER li1 ;
        RECT 706.760 1112.930 706.935 1113.130 ;
        RECT 706.760 1112.760 709.385 1112.930 ;
        RECT 706.760 1112.590 706.935 1112.760 ;
      LAYER li1 ;
        RECT 709.630 1112.590 709.885 1113.130 ;
        RECT 711.460 1112.760 712.560 1112.960 ;
      LAYER li1 ;
        RECT 712.740 1112.930 712.915 1113.130 ;
        RECT 712.740 1112.760 715.365 1112.930 ;
        RECT 712.740 1112.590 712.915 1112.760 ;
      LAYER li1 ;
        RECT 715.610 1112.590 715.865 1113.130 ;
        RECT 717.440 1112.760 718.540 1112.960 ;
      LAYER li1 ;
        RECT 718.720 1112.930 718.895 1113.130 ;
        RECT 718.720 1112.760 721.345 1112.930 ;
        RECT 718.720 1112.590 718.895 1112.760 ;
      LAYER li1 ;
        RECT 721.590 1112.590 721.845 1113.130 ;
        RECT 723.420 1112.760 724.520 1112.960 ;
      LAYER li1 ;
        RECT 724.700 1112.930 724.875 1113.130 ;
        RECT 724.700 1112.760 727.325 1112.930 ;
        RECT 724.700 1112.590 724.875 1112.760 ;
      LAYER li1 ;
        RECT 727.570 1112.590 727.825 1113.130 ;
        RECT 729.400 1112.760 730.500 1112.960 ;
      LAYER li1 ;
        RECT 730.680 1112.930 730.855 1113.130 ;
        RECT 730.680 1112.760 733.305 1112.930 ;
        RECT 730.680 1112.590 730.855 1112.760 ;
      LAYER li1 ;
        RECT 733.550 1112.590 733.805 1113.130 ;
        RECT 735.380 1112.760 736.480 1112.960 ;
      LAYER li1 ;
        RECT 736.660 1112.930 736.835 1113.130 ;
        RECT 736.660 1112.760 739.285 1112.930 ;
        RECT 736.660 1112.590 736.835 1112.760 ;
      LAYER li1 ;
        RECT 739.530 1112.590 739.785 1113.130 ;
        RECT 741.360 1112.760 742.460 1112.960 ;
      LAYER li1 ;
        RECT 742.640 1112.930 742.815 1113.130 ;
        RECT 742.640 1112.760 745.265 1112.930 ;
        RECT 742.640 1112.590 742.815 1112.760 ;
      LAYER li1 ;
        RECT 745.510 1112.590 745.765 1113.130 ;
        RECT 747.340 1112.760 748.440 1112.960 ;
      LAYER li1 ;
        RECT 748.620 1112.930 748.795 1113.130 ;
        RECT 748.620 1112.760 751.245 1112.930 ;
        RECT 748.620 1112.590 748.795 1112.760 ;
      LAYER li1 ;
        RECT 751.490 1112.590 751.745 1113.130 ;
        RECT 753.320 1112.760 754.420 1112.960 ;
      LAYER li1 ;
        RECT 754.600 1112.930 754.775 1113.130 ;
        RECT 754.600 1112.760 757.225 1112.930 ;
        RECT 754.600 1112.590 754.775 1112.760 ;
      LAYER li1 ;
        RECT 757.470 1112.590 757.725 1113.130 ;
        RECT 759.300 1112.760 760.400 1112.960 ;
      LAYER li1 ;
        RECT 760.580 1112.930 760.755 1113.130 ;
        RECT 760.580 1112.760 763.205 1112.930 ;
        RECT 760.580 1112.590 760.755 1112.760 ;
      LAYER li1 ;
        RECT 763.450 1112.590 763.705 1113.130 ;
      LAYER li1 ;
        RECT 766.560 1112.930 766.735 1113.130 ;
        RECT 766.560 1112.760 769.185 1112.930 ;
        RECT 766.560 1112.590 766.735 1112.760 ;
      LAYER li1 ;
        RECT 769.430 1112.590 769.685 1113.130 ;
      LAYER li1 ;
        RECT 772.540 1112.930 772.715 1113.130 ;
        RECT 772.540 1112.760 775.165 1112.930 ;
        RECT 772.540 1112.590 772.715 1112.760 ;
      LAYER li1 ;
        RECT 775.410 1112.590 775.665 1113.130 ;
      LAYER li1 ;
        RECT 778.520 1112.930 778.695 1113.130 ;
        RECT 778.520 1112.760 781.145 1112.930 ;
        RECT 778.520 1112.590 778.695 1112.760 ;
      LAYER li1 ;
        RECT 781.390 1112.590 781.645 1113.130 ;
      LAYER li1 ;
        RECT 784.500 1112.930 784.675 1113.130 ;
        RECT 784.500 1112.760 787.125 1112.930 ;
        RECT 784.500 1112.590 784.675 1112.760 ;
      LAYER li1 ;
        RECT 787.370 1112.590 787.625 1113.130 ;
      LAYER li1 ;
        RECT 792.985 1113.130 794.485 1113.300 ;
        RECT 794.665 1113.155 794.955 1114.320 ;
        RECT 1975.065 1113.155 1975.355 1114.320 ;
        RECT 1975.535 1113.300 1975.865 1114.150 ;
        RECT 1976.035 1113.520 1976.205 1114.320 ;
        RECT 1976.375 1113.300 1976.705 1114.150 ;
        RECT 1976.875 1113.520 1977.045 1114.320 ;
        RECT 1977.635 1113.520 1977.965 1114.320 ;
        RECT 1978.475 1113.520 1978.805 1114.320 ;
        RECT 1979.315 1113.520 1979.645 1114.320 ;
        RECT 1975.535 1113.130 1977.035 1113.300 ;
        RECT 1980.155 1113.170 1980.485 1114.320 ;
        RECT 1981.045 1113.155 1981.335 1114.320 ;
        RECT 1981.515 1113.300 1981.845 1114.150 ;
        RECT 1982.015 1113.520 1982.185 1114.320 ;
        RECT 1982.355 1113.300 1982.685 1114.150 ;
        RECT 1982.855 1113.520 1983.025 1114.320 ;
        RECT 1983.615 1113.520 1983.945 1114.320 ;
        RECT 1984.455 1113.520 1984.785 1114.320 ;
        RECT 1985.295 1113.520 1985.625 1114.320 ;
        RECT 1981.515 1113.130 1983.015 1113.300 ;
        RECT 1986.135 1113.170 1986.465 1114.320 ;
        RECT 1987.025 1113.155 1987.315 1114.320 ;
        RECT 1987.495 1113.300 1987.825 1114.150 ;
        RECT 1987.995 1113.520 1988.165 1114.320 ;
        RECT 1988.335 1113.300 1988.665 1114.150 ;
        RECT 1988.835 1113.520 1989.005 1114.320 ;
        RECT 1989.595 1113.520 1989.925 1114.320 ;
        RECT 1990.435 1113.520 1990.765 1114.320 ;
        RECT 1991.275 1113.520 1991.605 1114.320 ;
        RECT 1987.495 1113.130 1988.995 1113.300 ;
        RECT 1992.115 1113.170 1992.445 1114.320 ;
        RECT 1993.005 1113.155 1993.295 1114.320 ;
        RECT 1993.475 1113.300 1993.805 1114.150 ;
        RECT 1993.975 1113.520 1994.145 1114.320 ;
        RECT 1994.315 1113.300 1994.645 1114.150 ;
        RECT 1994.815 1113.520 1994.985 1114.320 ;
        RECT 1995.575 1113.520 1995.905 1114.320 ;
        RECT 1996.415 1113.520 1996.745 1114.320 ;
        RECT 1997.255 1113.520 1997.585 1114.320 ;
        RECT 1993.475 1113.130 1994.975 1113.300 ;
        RECT 1998.095 1113.170 1998.425 1114.320 ;
        RECT 1998.985 1113.155 1999.275 1114.320 ;
        RECT 1999.455 1113.300 1999.785 1114.150 ;
        RECT 1999.955 1113.520 2000.125 1114.320 ;
        RECT 2000.295 1113.300 2000.625 1114.150 ;
        RECT 2000.795 1113.520 2000.965 1114.320 ;
        RECT 2001.555 1113.520 2001.885 1114.320 ;
        RECT 2002.395 1113.520 2002.725 1114.320 ;
        RECT 2003.235 1113.520 2003.565 1114.320 ;
        RECT 1999.455 1113.130 2000.955 1113.300 ;
        RECT 2004.075 1113.170 2004.405 1114.320 ;
        RECT 2004.965 1113.155 2005.255 1114.320 ;
        RECT 2005.435 1113.300 2005.765 1114.150 ;
        RECT 2005.935 1113.520 2006.105 1114.320 ;
        RECT 2006.275 1113.300 2006.605 1114.150 ;
        RECT 2006.775 1113.520 2006.945 1114.320 ;
        RECT 2007.535 1113.520 2007.865 1114.320 ;
        RECT 2008.375 1113.520 2008.705 1114.320 ;
        RECT 2009.215 1113.520 2009.545 1114.320 ;
        RECT 2005.435 1113.130 2006.935 1113.300 ;
        RECT 2010.055 1113.170 2010.385 1114.320 ;
        RECT 2010.945 1113.155 2011.235 1114.320 ;
        RECT 2011.415 1113.300 2011.745 1114.150 ;
        RECT 2011.915 1113.520 2012.085 1114.320 ;
        RECT 2012.255 1113.300 2012.585 1114.150 ;
        RECT 2012.755 1113.520 2012.925 1114.320 ;
        RECT 2013.515 1113.520 2013.845 1114.320 ;
        RECT 2014.355 1113.520 2014.685 1114.320 ;
        RECT 2015.195 1113.520 2015.525 1114.320 ;
        RECT 2011.415 1113.130 2012.915 1113.300 ;
        RECT 2016.035 1113.170 2016.365 1114.320 ;
        RECT 2016.925 1113.155 2017.215 1114.320 ;
        RECT 2017.395 1113.300 2017.725 1114.150 ;
        RECT 2017.895 1113.520 2018.065 1114.320 ;
        RECT 2018.235 1113.300 2018.565 1114.150 ;
        RECT 2018.735 1113.520 2018.905 1114.320 ;
        RECT 2019.495 1113.520 2019.825 1114.320 ;
        RECT 2020.335 1113.520 2020.665 1114.320 ;
        RECT 2021.175 1113.520 2021.505 1114.320 ;
        RECT 2017.395 1113.130 2018.895 1113.300 ;
        RECT 2022.015 1113.170 2022.345 1114.320 ;
        RECT 2022.905 1113.155 2023.195 1114.320 ;
        RECT 2023.375 1113.300 2023.705 1114.150 ;
        RECT 2023.875 1113.520 2024.045 1114.320 ;
        RECT 2024.215 1113.300 2024.545 1114.150 ;
        RECT 2024.715 1113.520 2024.885 1114.320 ;
        RECT 2025.475 1113.520 2025.805 1114.320 ;
        RECT 2026.315 1113.520 2026.645 1114.320 ;
        RECT 2027.155 1113.520 2027.485 1114.320 ;
        RECT 2023.375 1113.130 2024.875 1113.300 ;
        RECT 2027.995 1113.170 2028.325 1114.320 ;
        RECT 2028.885 1113.155 2029.175 1114.320 ;
        RECT 2029.355 1113.300 2029.685 1114.150 ;
        RECT 2029.855 1113.520 2030.025 1114.320 ;
        RECT 2030.195 1113.300 2030.525 1114.150 ;
        RECT 2030.695 1113.520 2030.865 1114.320 ;
        RECT 2031.455 1113.520 2031.785 1114.320 ;
        RECT 2032.295 1113.520 2032.625 1114.320 ;
        RECT 2033.135 1113.520 2033.465 1114.320 ;
        RECT 2029.355 1113.130 2030.855 1113.300 ;
        RECT 2033.975 1113.170 2034.305 1114.320 ;
        RECT 2034.865 1113.155 2035.155 1114.320 ;
        RECT 2035.335 1113.300 2035.665 1114.150 ;
        RECT 2035.835 1113.520 2036.005 1114.320 ;
        RECT 2036.175 1113.300 2036.505 1114.150 ;
        RECT 2036.675 1113.520 2036.845 1114.320 ;
        RECT 2037.435 1113.520 2037.765 1114.320 ;
        RECT 2038.275 1113.520 2038.605 1114.320 ;
        RECT 2039.115 1113.520 2039.445 1114.320 ;
        RECT 2035.335 1113.130 2036.835 1113.300 ;
        RECT 2039.955 1113.170 2040.285 1114.320 ;
        RECT 2040.845 1113.155 2041.135 1114.320 ;
        RECT 2041.315 1113.300 2041.645 1114.150 ;
        RECT 2041.815 1113.520 2041.985 1114.320 ;
        RECT 2042.155 1113.300 2042.485 1114.150 ;
        RECT 2042.655 1113.520 2042.825 1114.320 ;
        RECT 2043.415 1113.520 2043.745 1114.320 ;
        RECT 2044.255 1113.520 2044.585 1114.320 ;
        RECT 2045.095 1113.520 2045.425 1114.320 ;
        RECT 2041.315 1113.130 2042.815 1113.300 ;
        RECT 2045.935 1113.170 2046.265 1114.320 ;
        RECT 2046.825 1113.155 2047.115 1114.320 ;
        RECT 2047.295 1113.300 2047.625 1114.150 ;
        RECT 2047.795 1113.520 2047.965 1114.320 ;
        RECT 2048.135 1113.300 2048.465 1114.150 ;
        RECT 2048.635 1113.520 2048.805 1114.320 ;
        RECT 2049.395 1113.520 2049.725 1114.320 ;
        RECT 2050.235 1113.520 2050.565 1114.320 ;
        RECT 2051.075 1113.520 2051.405 1114.320 ;
        RECT 2047.295 1113.130 2048.795 1113.300 ;
        RECT 2051.915 1113.170 2052.245 1114.320 ;
        RECT 2052.805 1113.155 2053.095 1114.320 ;
        RECT 2053.275 1113.300 2053.605 1114.150 ;
        RECT 2053.775 1113.520 2053.945 1114.320 ;
        RECT 2054.115 1113.300 2054.445 1114.150 ;
        RECT 2054.615 1113.520 2054.785 1114.320 ;
        RECT 2055.375 1113.520 2055.705 1114.320 ;
        RECT 2056.215 1113.520 2056.545 1114.320 ;
        RECT 2057.055 1113.520 2057.385 1114.320 ;
        RECT 2053.275 1113.130 2054.775 1113.300 ;
        RECT 2057.895 1113.170 2058.225 1114.320 ;
        RECT 2058.785 1113.155 2059.075 1114.320 ;
        RECT 2059.255 1113.300 2059.585 1114.150 ;
        RECT 2059.755 1113.520 2059.925 1114.320 ;
        RECT 2060.095 1113.300 2060.425 1114.150 ;
        RECT 2060.595 1113.520 2060.765 1114.320 ;
        RECT 2061.355 1113.520 2061.685 1114.320 ;
        RECT 2062.195 1113.520 2062.525 1114.320 ;
        RECT 2063.035 1113.520 2063.365 1114.320 ;
        RECT 2059.255 1113.130 2060.755 1113.300 ;
        RECT 2063.875 1113.170 2064.205 1114.320 ;
        RECT 2064.765 1113.155 2065.055 1114.320 ;
        RECT 2065.235 1113.300 2065.565 1114.150 ;
        RECT 2065.735 1113.520 2065.905 1114.320 ;
        RECT 2066.075 1113.300 2066.405 1114.150 ;
        RECT 2066.575 1113.520 2066.745 1114.320 ;
        RECT 2067.335 1113.520 2067.665 1114.320 ;
        RECT 2068.175 1113.520 2068.505 1114.320 ;
        RECT 2069.015 1113.520 2069.345 1114.320 ;
        RECT 2065.235 1113.130 2066.735 1113.300 ;
        RECT 2069.855 1113.170 2070.185 1114.320 ;
        RECT 2070.745 1113.155 2071.035 1114.320 ;
        RECT 2071.215 1113.300 2071.545 1114.150 ;
        RECT 2071.715 1113.520 2071.885 1114.320 ;
        RECT 2072.055 1113.300 2072.385 1114.150 ;
        RECT 2072.555 1113.520 2072.725 1114.320 ;
        RECT 2073.315 1113.520 2073.645 1114.320 ;
        RECT 2074.155 1113.520 2074.485 1114.320 ;
        RECT 2074.995 1113.520 2075.325 1114.320 ;
        RECT 2071.215 1113.130 2072.715 1113.300 ;
        RECT 2075.835 1113.170 2076.165 1114.320 ;
        RECT 2076.725 1113.155 2077.015 1114.320 ;
        RECT 2077.195 1113.300 2077.525 1114.150 ;
        RECT 2077.695 1113.520 2077.865 1114.320 ;
        RECT 2078.035 1113.300 2078.365 1114.150 ;
        RECT 2078.535 1113.520 2078.705 1114.320 ;
        RECT 2079.295 1113.520 2079.625 1114.320 ;
        RECT 2080.135 1113.520 2080.465 1114.320 ;
        RECT 2080.975 1113.520 2081.305 1114.320 ;
        RECT 2077.195 1113.130 2078.695 1113.300 ;
        RECT 2081.815 1113.170 2082.145 1114.320 ;
        RECT 2082.705 1113.155 2082.995 1114.320 ;
        RECT 2083.175 1113.300 2083.505 1114.150 ;
        RECT 2083.675 1113.520 2083.845 1114.320 ;
        RECT 2084.015 1113.300 2084.345 1114.150 ;
        RECT 2084.515 1113.520 2084.685 1114.320 ;
        RECT 2085.275 1113.520 2085.605 1114.320 ;
        RECT 2086.115 1113.520 2086.445 1114.320 ;
        RECT 2086.955 1113.520 2087.285 1114.320 ;
        RECT 2083.175 1113.130 2084.675 1113.300 ;
        RECT 2087.795 1113.170 2088.125 1114.320 ;
        RECT 2088.685 1113.155 2088.975 1114.320 ;
        RECT 2089.535 1113.170 2089.865 1114.320 ;
      LAYER li1 ;
        RECT 2090.035 1113.300 2090.205 1114.150 ;
      LAYER li1 ;
        RECT 2090.375 1113.520 2090.705 1114.320 ;
      LAYER li1 ;
        RECT 2090.875 1113.300 2091.045 1114.150 ;
      LAYER li1 ;
        RECT 2091.215 1113.520 2091.545 1114.320 ;
      LAYER li1 ;
        RECT 2091.715 1113.300 2091.885 1114.150 ;
      LAYER li1 ;
        RECT 2092.055 1113.520 2092.385 1114.320 ;
      LAYER li1 ;
        RECT 2092.555 1113.300 2092.725 1114.150 ;
      LAYER li1 ;
        RECT 2092.975 1113.520 2093.145 1114.320 ;
        RECT 2093.315 1113.300 2093.645 1114.150 ;
        RECT 2093.815 1113.520 2093.985 1114.320 ;
        RECT 2094.155 1113.300 2094.485 1114.150 ;
        RECT 792.985 1112.930 793.160 1113.130 ;
        RECT 790.535 1112.760 793.160 1112.930 ;
      LAYER li1 ;
        RECT 793.340 1112.760 794.440 1112.960 ;
        RECT 1975.580 1112.760 1976.680 1112.960 ;
      LAYER li1 ;
        RECT 1976.860 1112.930 1977.035 1113.130 ;
        RECT 1976.860 1112.760 1979.485 1112.930 ;
      LAYER li1 ;
        RECT 1981.560 1112.760 1982.660 1112.960 ;
      LAYER li1 ;
        RECT 1982.840 1112.930 1983.015 1113.130 ;
        RECT 1982.840 1112.760 1985.465 1112.930 ;
      LAYER li1 ;
        RECT 1987.540 1112.760 1988.640 1112.960 ;
      LAYER li1 ;
        RECT 1988.820 1112.930 1988.995 1113.130 ;
        RECT 1988.820 1112.760 1991.445 1112.930 ;
      LAYER li1 ;
        RECT 1993.520 1112.760 1994.620 1112.960 ;
      LAYER li1 ;
        RECT 1994.800 1112.930 1994.975 1113.130 ;
        RECT 1994.800 1112.760 1997.425 1112.930 ;
      LAYER li1 ;
        RECT 1999.500 1112.760 2000.600 1112.960 ;
      LAYER li1 ;
        RECT 2000.780 1112.930 2000.955 1113.130 ;
        RECT 2000.780 1112.760 2003.405 1112.930 ;
      LAYER li1 ;
        RECT 2005.480 1112.760 2006.580 1112.960 ;
      LAYER li1 ;
        RECT 2006.760 1112.930 2006.935 1113.130 ;
        RECT 2006.760 1112.760 2009.385 1112.930 ;
      LAYER li1 ;
        RECT 2011.460 1112.760 2012.560 1112.960 ;
      LAYER li1 ;
        RECT 2012.740 1112.930 2012.915 1113.130 ;
        RECT 2012.740 1112.760 2015.365 1112.930 ;
      LAYER li1 ;
        RECT 2017.440 1112.760 2018.540 1112.960 ;
      LAYER li1 ;
        RECT 2018.720 1112.930 2018.895 1113.130 ;
        RECT 2018.720 1112.760 2021.345 1112.930 ;
      LAYER li1 ;
        RECT 2023.420 1112.760 2024.520 1112.960 ;
      LAYER li1 ;
        RECT 2024.700 1112.930 2024.875 1113.130 ;
        RECT 2024.700 1112.760 2027.325 1112.930 ;
      LAYER li1 ;
        RECT 2029.400 1112.760 2030.500 1112.960 ;
      LAYER li1 ;
        RECT 2030.680 1112.930 2030.855 1113.130 ;
        RECT 2030.680 1112.760 2033.305 1112.930 ;
      LAYER li1 ;
        RECT 2035.380 1112.760 2036.480 1112.960 ;
      LAYER li1 ;
        RECT 2036.660 1112.930 2036.835 1113.130 ;
        RECT 2036.660 1112.760 2039.285 1112.930 ;
      LAYER li1 ;
        RECT 2041.360 1112.760 2042.460 1112.960 ;
      LAYER li1 ;
        RECT 2042.640 1112.930 2042.815 1113.130 ;
        RECT 2042.640 1112.760 2045.265 1112.930 ;
      LAYER li1 ;
        RECT 2047.340 1112.760 2048.440 1112.960 ;
      LAYER li1 ;
        RECT 2048.620 1112.930 2048.795 1113.130 ;
        RECT 2048.620 1112.760 2051.245 1112.930 ;
      LAYER li1 ;
        RECT 2053.320 1112.760 2054.420 1112.960 ;
      LAYER li1 ;
        RECT 2054.600 1112.930 2054.775 1113.130 ;
        RECT 2054.600 1112.760 2057.225 1112.930 ;
      LAYER li1 ;
        RECT 2059.300 1112.760 2060.400 1112.960 ;
      LAYER li1 ;
        RECT 2060.580 1112.930 2060.755 1113.130 ;
        RECT 2060.580 1112.760 2063.205 1112.930 ;
      LAYER li1 ;
        RECT 2065.280 1112.760 2066.380 1112.960 ;
      LAYER li1 ;
        RECT 2066.560 1112.930 2066.735 1113.130 ;
        RECT 2066.560 1112.760 2069.185 1112.930 ;
      LAYER li1 ;
        RECT 2071.260 1112.760 2072.360 1112.960 ;
      LAYER li1 ;
        RECT 2072.540 1112.930 2072.715 1113.130 ;
        RECT 2072.540 1112.760 2075.165 1112.930 ;
      LAYER li1 ;
        RECT 2077.240 1112.760 2078.340 1112.960 ;
      LAYER li1 ;
        RECT 2078.520 1112.930 2078.695 1113.130 ;
        RECT 2078.520 1112.760 2081.145 1112.930 ;
      LAYER li1 ;
        RECT 2083.220 1112.760 2084.320 1112.960 ;
      LAYER li1 ;
        RECT 2084.500 1112.930 2084.675 1113.130 ;
      LAYER li1 ;
        RECT 2090.035 1113.130 2092.725 1113.300 ;
      LAYER li1 ;
        RECT 2092.985 1113.130 2094.485 1113.300 ;
        RECT 2094.665 1113.155 2094.955 1114.320 ;
        RECT 2084.500 1112.760 2087.125 1112.930 ;
        RECT 675.065 1111.770 675.355 1112.495 ;
        RECT 675.615 1112.420 677.035 1112.590 ;
      LAYER li1 ;
        RECT 677.295 1112.420 679.985 1112.590 ;
      LAYER li1 ;
        RECT 675.615 1111.940 675.785 1112.420 ;
        RECT 675.955 1111.770 676.285 1112.250 ;
        RECT 676.455 1111.945 676.625 1112.420 ;
        RECT 676.795 1111.770 677.125 1112.250 ;
      LAYER li1 ;
        RECT 677.295 1111.940 677.465 1112.420 ;
      LAYER li1 ;
        RECT 677.635 1111.770 677.965 1112.250 ;
      LAYER li1 ;
        RECT 678.135 1111.940 678.305 1112.420 ;
      LAYER li1 ;
        RECT 678.475 1111.770 678.805 1112.250 ;
      LAYER li1 ;
        RECT 678.975 1111.940 679.145 1112.420 ;
      LAYER li1 ;
        RECT 679.315 1111.770 679.645 1112.250 ;
      LAYER li1 ;
        RECT 679.815 1111.940 679.985 1112.420 ;
      LAYER li1 ;
        RECT 680.155 1111.770 680.485 1112.570 ;
        RECT 681.045 1111.770 681.335 1112.495 ;
        RECT 681.595 1112.420 683.015 1112.590 ;
      LAYER li1 ;
        RECT 683.275 1112.420 685.965 1112.590 ;
      LAYER li1 ;
        RECT 681.595 1111.940 681.765 1112.420 ;
        RECT 681.935 1111.770 682.265 1112.250 ;
        RECT 682.435 1111.945 682.605 1112.420 ;
        RECT 682.775 1111.770 683.105 1112.250 ;
      LAYER li1 ;
        RECT 683.275 1111.940 683.445 1112.420 ;
      LAYER li1 ;
        RECT 683.615 1111.770 683.945 1112.250 ;
      LAYER li1 ;
        RECT 684.115 1111.940 684.285 1112.420 ;
      LAYER li1 ;
        RECT 684.455 1111.770 684.785 1112.250 ;
      LAYER li1 ;
        RECT 684.955 1111.940 685.125 1112.420 ;
      LAYER li1 ;
        RECT 685.295 1111.770 685.625 1112.250 ;
      LAYER li1 ;
        RECT 685.795 1111.940 685.965 1112.420 ;
      LAYER li1 ;
        RECT 686.135 1111.770 686.465 1112.570 ;
        RECT 687.025 1111.770 687.315 1112.495 ;
        RECT 687.575 1112.420 688.995 1112.590 ;
      LAYER li1 ;
        RECT 689.255 1112.420 691.945 1112.590 ;
      LAYER li1 ;
        RECT 687.575 1111.940 687.745 1112.420 ;
        RECT 687.915 1111.770 688.245 1112.250 ;
        RECT 688.415 1111.945 688.585 1112.420 ;
        RECT 688.755 1111.770 689.085 1112.250 ;
      LAYER li1 ;
        RECT 689.255 1111.940 689.425 1112.420 ;
      LAYER li1 ;
        RECT 689.595 1111.770 689.925 1112.250 ;
      LAYER li1 ;
        RECT 690.095 1111.940 690.265 1112.420 ;
      LAYER li1 ;
        RECT 690.435 1111.770 690.765 1112.250 ;
      LAYER li1 ;
        RECT 690.935 1111.940 691.105 1112.420 ;
      LAYER li1 ;
        RECT 691.275 1111.770 691.605 1112.250 ;
      LAYER li1 ;
        RECT 691.775 1111.940 691.945 1112.420 ;
      LAYER li1 ;
        RECT 692.115 1111.770 692.445 1112.570 ;
        RECT 693.005 1111.770 693.295 1112.495 ;
        RECT 693.555 1112.420 694.975 1112.590 ;
      LAYER li1 ;
        RECT 695.235 1112.420 697.925 1112.590 ;
      LAYER li1 ;
        RECT 693.555 1111.940 693.725 1112.420 ;
        RECT 693.895 1111.770 694.225 1112.250 ;
        RECT 694.395 1111.945 694.565 1112.420 ;
        RECT 694.735 1111.770 695.065 1112.250 ;
      LAYER li1 ;
        RECT 695.235 1111.940 695.405 1112.420 ;
      LAYER li1 ;
        RECT 695.575 1111.770 695.905 1112.250 ;
      LAYER li1 ;
        RECT 696.075 1111.940 696.245 1112.420 ;
      LAYER li1 ;
        RECT 696.415 1111.770 696.745 1112.250 ;
      LAYER li1 ;
        RECT 696.915 1111.940 697.085 1112.420 ;
      LAYER li1 ;
        RECT 697.255 1111.770 697.585 1112.250 ;
      LAYER li1 ;
        RECT 697.755 1111.940 697.925 1112.420 ;
      LAYER li1 ;
        RECT 698.095 1111.770 698.425 1112.570 ;
        RECT 698.985 1111.770 699.275 1112.495 ;
        RECT 699.535 1112.420 700.955 1112.590 ;
      LAYER li1 ;
        RECT 701.215 1112.420 703.905 1112.590 ;
      LAYER li1 ;
        RECT 699.535 1111.940 699.705 1112.420 ;
        RECT 699.875 1111.770 700.205 1112.250 ;
        RECT 700.375 1111.945 700.545 1112.420 ;
        RECT 700.715 1111.770 701.045 1112.250 ;
      LAYER li1 ;
        RECT 701.215 1111.940 701.385 1112.420 ;
      LAYER li1 ;
        RECT 701.555 1111.770 701.885 1112.250 ;
      LAYER li1 ;
        RECT 702.055 1111.940 702.225 1112.420 ;
      LAYER li1 ;
        RECT 702.395 1111.770 702.725 1112.250 ;
      LAYER li1 ;
        RECT 702.895 1111.940 703.065 1112.420 ;
      LAYER li1 ;
        RECT 703.235 1111.770 703.565 1112.250 ;
      LAYER li1 ;
        RECT 703.735 1111.940 703.905 1112.420 ;
      LAYER li1 ;
        RECT 704.075 1111.770 704.405 1112.570 ;
        RECT 704.965 1111.770 705.255 1112.495 ;
        RECT 705.515 1112.420 706.935 1112.590 ;
      LAYER li1 ;
        RECT 707.195 1112.420 709.885 1112.590 ;
      LAYER li1 ;
        RECT 705.515 1111.940 705.685 1112.420 ;
        RECT 705.855 1111.770 706.185 1112.250 ;
        RECT 706.355 1111.945 706.525 1112.420 ;
        RECT 706.695 1111.770 707.025 1112.250 ;
      LAYER li1 ;
        RECT 707.195 1111.940 707.365 1112.420 ;
      LAYER li1 ;
        RECT 707.535 1111.770 707.865 1112.250 ;
      LAYER li1 ;
        RECT 708.035 1111.940 708.205 1112.420 ;
      LAYER li1 ;
        RECT 708.375 1111.770 708.705 1112.250 ;
      LAYER li1 ;
        RECT 708.875 1111.940 709.045 1112.420 ;
      LAYER li1 ;
        RECT 709.215 1111.770 709.545 1112.250 ;
      LAYER li1 ;
        RECT 709.715 1111.940 709.885 1112.420 ;
      LAYER li1 ;
        RECT 710.055 1111.770 710.385 1112.570 ;
        RECT 710.945 1111.770 711.235 1112.495 ;
        RECT 711.495 1112.420 712.915 1112.590 ;
      LAYER li1 ;
        RECT 713.175 1112.420 715.865 1112.590 ;
      LAYER li1 ;
        RECT 711.495 1111.940 711.665 1112.420 ;
        RECT 711.835 1111.770 712.165 1112.250 ;
        RECT 712.335 1111.945 712.505 1112.420 ;
        RECT 712.675 1111.770 713.005 1112.250 ;
      LAYER li1 ;
        RECT 713.175 1111.940 713.345 1112.420 ;
      LAYER li1 ;
        RECT 713.515 1111.770 713.845 1112.250 ;
      LAYER li1 ;
        RECT 714.015 1111.940 714.185 1112.420 ;
      LAYER li1 ;
        RECT 714.355 1111.770 714.685 1112.250 ;
      LAYER li1 ;
        RECT 714.855 1111.940 715.025 1112.420 ;
      LAYER li1 ;
        RECT 715.195 1111.770 715.525 1112.250 ;
      LAYER li1 ;
        RECT 715.695 1111.940 715.865 1112.420 ;
      LAYER li1 ;
        RECT 716.035 1111.770 716.365 1112.570 ;
        RECT 716.925 1111.770 717.215 1112.495 ;
        RECT 717.475 1112.420 718.895 1112.590 ;
      LAYER li1 ;
        RECT 719.155 1112.420 721.845 1112.590 ;
      LAYER li1 ;
        RECT 717.475 1111.940 717.645 1112.420 ;
        RECT 717.815 1111.770 718.145 1112.250 ;
        RECT 718.315 1111.945 718.485 1112.420 ;
        RECT 718.655 1111.770 718.985 1112.250 ;
      LAYER li1 ;
        RECT 719.155 1111.940 719.325 1112.420 ;
      LAYER li1 ;
        RECT 719.495 1111.770 719.825 1112.250 ;
      LAYER li1 ;
        RECT 719.995 1111.940 720.165 1112.420 ;
      LAYER li1 ;
        RECT 720.335 1111.770 720.665 1112.250 ;
      LAYER li1 ;
        RECT 720.835 1111.940 721.005 1112.420 ;
      LAYER li1 ;
        RECT 721.175 1111.770 721.505 1112.250 ;
      LAYER li1 ;
        RECT 721.675 1111.940 721.845 1112.420 ;
      LAYER li1 ;
        RECT 722.015 1111.770 722.345 1112.570 ;
        RECT 722.905 1111.770 723.195 1112.495 ;
        RECT 723.455 1112.420 724.875 1112.590 ;
      LAYER li1 ;
        RECT 725.135 1112.420 727.825 1112.590 ;
      LAYER li1 ;
        RECT 723.455 1111.940 723.625 1112.420 ;
        RECT 723.795 1111.770 724.125 1112.250 ;
        RECT 724.295 1111.945 724.465 1112.420 ;
        RECT 724.635 1111.770 724.965 1112.250 ;
      LAYER li1 ;
        RECT 725.135 1111.940 725.305 1112.420 ;
      LAYER li1 ;
        RECT 725.475 1111.770 725.805 1112.250 ;
      LAYER li1 ;
        RECT 725.975 1111.940 726.145 1112.420 ;
      LAYER li1 ;
        RECT 726.315 1111.770 726.645 1112.250 ;
      LAYER li1 ;
        RECT 726.815 1111.940 726.985 1112.420 ;
      LAYER li1 ;
        RECT 727.155 1111.770 727.485 1112.250 ;
      LAYER li1 ;
        RECT 727.655 1111.940 727.825 1112.420 ;
      LAYER li1 ;
        RECT 727.995 1111.770 728.325 1112.570 ;
        RECT 728.885 1111.770 729.175 1112.495 ;
        RECT 729.435 1112.420 730.855 1112.590 ;
      LAYER li1 ;
        RECT 731.115 1112.420 733.805 1112.590 ;
      LAYER li1 ;
        RECT 729.435 1111.940 729.605 1112.420 ;
        RECT 729.775 1111.770 730.105 1112.250 ;
        RECT 730.275 1111.945 730.445 1112.420 ;
        RECT 730.615 1111.770 730.945 1112.250 ;
      LAYER li1 ;
        RECT 731.115 1111.940 731.285 1112.420 ;
      LAYER li1 ;
        RECT 731.455 1111.770 731.785 1112.250 ;
      LAYER li1 ;
        RECT 731.955 1111.940 732.125 1112.420 ;
      LAYER li1 ;
        RECT 732.295 1111.770 732.625 1112.250 ;
      LAYER li1 ;
        RECT 732.795 1111.940 732.965 1112.420 ;
      LAYER li1 ;
        RECT 733.135 1111.770 733.465 1112.250 ;
      LAYER li1 ;
        RECT 733.635 1111.940 733.805 1112.420 ;
      LAYER li1 ;
        RECT 733.975 1111.770 734.305 1112.570 ;
        RECT 734.865 1111.770 735.155 1112.495 ;
        RECT 735.415 1112.420 736.835 1112.590 ;
      LAYER li1 ;
        RECT 737.095 1112.420 739.785 1112.590 ;
      LAYER li1 ;
        RECT 735.415 1111.940 735.585 1112.420 ;
        RECT 735.755 1111.770 736.085 1112.250 ;
        RECT 736.255 1111.945 736.425 1112.420 ;
        RECT 736.595 1111.770 736.925 1112.250 ;
      LAYER li1 ;
        RECT 737.095 1111.940 737.265 1112.420 ;
      LAYER li1 ;
        RECT 737.435 1111.770 737.765 1112.250 ;
      LAYER li1 ;
        RECT 737.935 1111.940 738.105 1112.420 ;
      LAYER li1 ;
        RECT 738.275 1111.770 738.605 1112.250 ;
      LAYER li1 ;
        RECT 738.775 1111.940 738.945 1112.420 ;
      LAYER li1 ;
        RECT 739.115 1111.770 739.445 1112.250 ;
      LAYER li1 ;
        RECT 739.615 1111.940 739.785 1112.420 ;
      LAYER li1 ;
        RECT 739.955 1111.770 740.285 1112.570 ;
        RECT 740.845 1111.770 741.135 1112.495 ;
        RECT 741.395 1112.420 742.815 1112.590 ;
      LAYER li1 ;
        RECT 743.075 1112.420 745.765 1112.590 ;
      LAYER li1 ;
        RECT 741.395 1111.940 741.565 1112.420 ;
        RECT 741.735 1111.770 742.065 1112.250 ;
        RECT 742.235 1111.945 742.405 1112.420 ;
        RECT 742.575 1111.770 742.905 1112.250 ;
      LAYER li1 ;
        RECT 743.075 1111.940 743.245 1112.420 ;
      LAYER li1 ;
        RECT 743.415 1111.770 743.745 1112.250 ;
      LAYER li1 ;
        RECT 743.915 1111.940 744.085 1112.420 ;
      LAYER li1 ;
        RECT 744.255 1111.770 744.585 1112.250 ;
      LAYER li1 ;
        RECT 744.755 1111.940 744.925 1112.420 ;
      LAYER li1 ;
        RECT 745.095 1111.770 745.425 1112.250 ;
      LAYER li1 ;
        RECT 745.595 1111.940 745.765 1112.420 ;
      LAYER li1 ;
        RECT 745.935 1111.770 746.265 1112.570 ;
        RECT 746.825 1111.770 747.115 1112.495 ;
        RECT 747.375 1112.420 748.795 1112.590 ;
      LAYER li1 ;
        RECT 749.055 1112.420 751.745 1112.590 ;
      LAYER li1 ;
        RECT 747.375 1111.940 747.545 1112.420 ;
        RECT 747.715 1111.770 748.045 1112.250 ;
        RECT 748.215 1111.945 748.385 1112.420 ;
        RECT 748.555 1111.770 748.885 1112.250 ;
      LAYER li1 ;
        RECT 749.055 1111.940 749.225 1112.420 ;
      LAYER li1 ;
        RECT 749.395 1111.770 749.725 1112.250 ;
      LAYER li1 ;
        RECT 749.895 1111.940 750.065 1112.420 ;
      LAYER li1 ;
        RECT 750.235 1111.770 750.565 1112.250 ;
      LAYER li1 ;
        RECT 750.735 1111.940 750.905 1112.420 ;
      LAYER li1 ;
        RECT 751.075 1111.770 751.405 1112.250 ;
      LAYER li1 ;
        RECT 751.575 1111.940 751.745 1112.420 ;
      LAYER li1 ;
        RECT 751.915 1111.770 752.245 1112.570 ;
        RECT 752.805 1111.770 753.095 1112.495 ;
        RECT 753.355 1112.420 754.775 1112.590 ;
      LAYER li1 ;
        RECT 755.035 1112.420 757.725 1112.590 ;
      LAYER li1 ;
        RECT 753.355 1111.940 753.525 1112.420 ;
        RECT 753.695 1111.770 754.025 1112.250 ;
        RECT 754.195 1111.945 754.365 1112.420 ;
        RECT 754.535 1111.770 754.865 1112.250 ;
      LAYER li1 ;
        RECT 755.035 1111.940 755.205 1112.420 ;
      LAYER li1 ;
        RECT 755.375 1111.770 755.705 1112.250 ;
      LAYER li1 ;
        RECT 755.875 1111.940 756.045 1112.420 ;
      LAYER li1 ;
        RECT 756.215 1111.770 756.545 1112.250 ;
      LAYER li1 ;
        RECT 756.715 1111.940 756.885 1112.420 ;
      LAYER li1 ;
        RECT 757.055 1111.770 757.385 1112.250 ;
      LAYER li1 ;
        RECT 757.555 1111.940 757.725 1112.420 ;
      LAYER li1 ;
        RECT 757.895 1111.770 758.225 1112.570 ;
        RECT 758.785 1111.770 759.075 1112.495 ;
        RECT 759.335 1112.420 760.755 1112.590 ;
      LAYER li1 ;
        RECT 761.015 1112.420 763.705 1112.590 ;
      LAYER li1 ;
        RECT 759.335 1111.940 759.505 1112.420 ;
        RECT 759.675 1111.770 760.005 1112.250 ;
        RECT 760.175 1111.945 760.345 1112.420 ;
        RECT 760.515 1111.770 760.845 1112.250 ;
      LAYER li1 ;
        RECT 761.015 1111.940 761.185 1112.420 ;
      LAYER li1 ;
        RECT 761.355 1111.770 761.685 1112.250 ;
      LAYER li1 ;
        RECT 761.855 1111.940 762.025 1112.420 ;
      LAYER li1 ;
        RECT 762.195 1111.770 762.525 1112.250 ;
      LAYER li1 ;
        RECT 762.695 1111.940 762.865 1112.420 ;
      LAYER li1 ;
        RECT 763.035 1111.770 763.365 1112.250 ;
      LAYER li1 ;
        RECT 763.535 1111.940 763.705 1112.420 ;
      LAYER li1 ;
        RECT 763.875 1111.770 764.205 1112.570 ;
        RECT 764.765 1111.770 765.055 1112.495 ;
        RECT 765.315 1112.420 766.735 1112.590 ;
      LAYER li1 ;
        RECT 766.995 1112.420 769.685 1112.590 ;
      LAYER li1 ;
        RECT 765.315 1111.940 765.485 1112.420 ;
        RECT 765.655 1111.770 765.985 1112.250 ;
        RECT 766.155 1111.945 766.325 1112.420 ;
        RECT 766.495 1111.770 766.825 1112.250 ;
      LAYER li1 ;
        RECT 766.995 1111.940 767.165 1112.420 ;
      LAYER li1 ;
        RECT 767.335 1111.770 767.665 1112.250 ;
      LAYER li1 ;
        RECT 767.835 1111.940 768.005 1112.420 ;
      LAYER li1 ;
        RECT 768.175 1111.770 768.505 1112.250 ;
      LAYER li1 ;
        RECT 768.675 1111.940 768.845 1112.420 ;
      LAYER li1 ;
        RECT 769.015 1111.770 769.345 1112.250 ;
      LAYER li1 ;
        RECT 769.515 1111.940 769.685 1112.420 ;
      LAYER li1 ;
        RECT 769.855 1111.770 770.185 1112.570 ;
        RECT 770.745 1111.770 771.035 1112.495 ;
        RECT 771.295 1112.420 772.715 1112.590 ;
      LAYER li1 ;
        RECT 772.975 1112.420 775.665 1112.590 ;
      LAYER li1 ;
        RECT 771.295 1111.940 771.465 1112.420 ;
        RECT 771.635 1111.770 771.965 1112.250 ;
        RECT 772.135 1111.945 772.305 1112.420 ;
        RECT 772.475 1111.770 772.805 1112.250 ;
      LAYER li1 ;
        RECT 772.975 1111.940 773.145 1112.420 ;
      LAYER li1 ;
        RECT 773.315 1111.770 773.645 1112.250 ;
      LAYER li1 ;
        RECT 773.815 1111.940 773.985 1112.420 ;
      LAYER li1 ;
        RECT 774.155 1111.770 774.485 1112.250 ;
      LAYER li1 ;
        RECT 774.655 1111.940 774.825 1112.420 ;
      LAYER li1 ;
        RECT 774.995 1111.770 775.325 1112.250 ;
      LAYER li1 ;
        RECT 775.495 1111.940 775.665 1112.420 ;
      LAYER li1 ;
        RECT 775.835 1111.770 776.165 1112.570 ;
        RECT 776.725 1111.770 777.015 1112.495 ;
        RECT 777.275 1112.420 778.695 1112.590 ;
      LAYER li1 ;
        RECT 778.955 1112.420 781.645 1112.590 ;
      LAYER li1 ;
        RECT 777.275 1111.940 777.445 1112.420 ;
        RECT 777.615 1111.770 777.945 1112.250 ;
        RECT 778.115 1111.945 778.285 1112.420 ;
        RECT 778.455 1111.770 778.785 1112.250 ;
      LAYER li1 ;
        RECT 778.955 1111.940 779.125 1112.420 ;
      LAYER li1 ;
        RECT 779.295 1111.770 779.625 1112.250 ;
      LAYER li1 ;
        RECT 779.795 1111.940 779.965 1112.420 ;
      LAYER li1 ;
        RECT 780.135 1111.770 780.465 1112.250 ;
      LAYER li1 ;
        RECT 780.635 1111.940 780.805 1112.420 ;
      LAYER li1 ;
        RECT 780.975 1111.770 781.305 1112.250 ;
      LAYER li1 ;
        RECT 781.475 1111.940 781.645 1112.420 ;
      LAYER li1 ;
        RECT 781.815 1111.770 782.145 1112.570 ;
        RECT 782.705 1111.770 782.995 1112.495 ;
        RECT 783.255 1112.420 784.675 1112.590 ;
      LAYER li1 ;
        RECT 784.935 1112.420 787.625 1112.590 ;
      LAYER li1 ;
        RECT 792.985 1112.590 793.160 1112.760 ;
        RECT 1976.860 1112.590 1977.035 1112.760 ;
        RECT 1982.840 1112.590 1983.015 1112.760 ;
        RECT 1988.820 1112.590 1988.995 1112.760 ;
        RECT 1994.800 1112.590 1994.975 1112.760 ;
        RECT 2000.780 1112.590 2000.955 1112.760 ;
        RECT 2006.760 1112.590 2006.935 1112.760 ;
        RECT 2012.740 1112.590 2012.915 1112.760 ;
        RECT 2018.720 1112.590 2018.895 1112.760 ;
        RECT 2024.700 1112.590 2024.875 1112.760 ;
        RECT 2030.680 1112.590 2030.855 1112.760 ;
        RECT 2036.660 1112.590 2036.835 1112.760 ;
        RECT 2042.640 1112.590 2042.815 1112.760 ;
        RECT 2048.620 1112.590 2048.795 1112.760 ;
        RECT 2054.600 1112.590 2054.775 1112.760 ;
        RECT 2060.580 1112.590 2060.755 1112.760 ;
        RECT 2066.560 1112.590 2066.735 1112.760 ;
        RECT 2072.540 1112.590 2072.715 1112.760 ;
        RECT 2078.520 1112.590 2078.695 1112.760 ;
        RECT 2084.500 1112.590 2084.675 1112.760 ;
        RECT 783.255 1111.940 783.425 1112.420 ;
        RECT 783.595 1111.770 783.925 1112.250 ;
        RECT 784.095 1111.945 784.265 1112.420 ;
        RECT 784.435 1111.770 784.765 1112.250 ;
      LAYER li1 ;
        RECT 784.935 1111.940 785.105 1112.420 ;
      LAYER li1 ;
        RECT 785.275 1111.770 785.605 1112.250 ;
      LAYER li1 ;
        RECT 785.775 1111.940 785.945 1112.420 ;
      LAYER li1 ;
        RECT 786.115 1111.770 786.445 1112.250 ;
      LAYER li1 ;
        RECT 786.615 1111.940 786.785 1112.420 ;
      LAYER li1 ;
        RECT 786.955 1111.770 787.285 1112.250 ;
      LAYER li1 ;
        RECT 787.455 1111.940 787.625 1112.420 ;
      LAYER li1 ;
        RECT 787.795 1111.770 788.125 1112.570 ;
        RECT 788.685 1111.770 788.975 1112.495 ;
        RECT 789.535 1111.770 789.865 1112.570 ;
        RECT 792.985 1112.420 794.405 1112.590 ;
        RECT 790.375 1111.770 790.705 1112.250 ;
        RECT 791.215 1111.770 791.545 1112.250 ;
        RECT 792.055 1111.770 792.385 1112.250 ;
        RECT 792.895 1111.770 793.225 1112.250 ;
        RECT 793.395 1111.945 793.565 1112.420 ;
        RECT 793.735 1111.770 794.065 1112.250 ;
        RECT 794.235 1111.940 794.405 1112.420 ;
        RECT 794.665 1111.770 794.955 1112.495 ;
        RECT 1975.065 1111.770 1975.355 1112.495 ;
        RECT 1975.615 1112.420 1977.035 1112.590 ;
        RECT 1975.615 1111.940 1975.785 1112.420 ;
        RECT 1975.955 1111.770 1976.285 1112.250 ;
        RECT 1976.455 1111.945 1976.625 1112.420 ;
        RECT 1976.795 1111.770 1977.125 1112.250 ;
        RECT 1977.635 1111.770 1977.965 1112.250 ;
        RECT 1978.475 1111.770 1978.805 1112.250 ;
        RECT 1979.315 1111.770 1979.645 1112.250 ;
        RECT 1980.155 1111.770 1980.485 1112.570 ;
        RECT 1981.045 1111.770 1981.335 1112.495 ;
        RECT 1981.595 1112.420 1983.015 1112.590 ;
        RECT 1981.595 1111.940 1981.765 1112.420 ;
        RECT 1981.935 1111.770 1982.265 1112.250 ;
        RECT 1982.435 1111.945 1982.605 1112.420 ;
        RECT 1982.775 1111.770 1983.105 1112.250 ;
        RECT 1983.615 1111.770 1983.945 1112.250 ;
        RECT 1984.455 1111.770 1984.785 1112.250 ;
        RECT 1985.295 1111.770 1985.625 1112.250 ;
        RECT 1986.135 1111.770 1986.465 1112.570 ;
        RECT 1987.025 1111.770 1987.315 1112.495 ;
        RECT 1987.575 1112.420 1988.995 1112.590 ;
        RECT 1987.575 1111.940 1987.745 1112.420 ;
        RECT 1987.915 1111.770 1988.245 1112.250 ;
        RECT 1988.415 1111.945 1988.585 1112.420 ;
        RECT 1988.755 1111.770 1989.085 1112.250 ;
        RECT 1989.595 1111.770 1989.925 1112.250 ;
        RECT 1990.435 1111.770 1990.765 1112.250 ;
        RECT 1991.275 1111.770 1991.605 1112.250 ;
        RECT 1992.115 1111.770 1992.445 1112.570 ;
        RECT 1993.005 1111.770 1993.295 1112.495 ;
        RECT 1993.555 1112.420 1994.975 1112.590 ;
        RECT 1993.555 1111.940 1993.725 1112.420 ;
        RECT 1993.895 1111.770 1994.225 1112.250 ;
        RECT 1994.395 1111.945 1994.565 1112.420 ;
        RECT 1994.735 1111.770 1995.065 1112.250 ;
        RECT 1995.575 1111.770 1995.905 1112.250 ;
        RECT 1996.415 1111.770 1996.745 1112.250 ;
        RECT 1997.255 1111.770 1997.585 1112.250 ;
        RECT 1998.095 1111.770 1998.425 1112.570 ;
        RECT 1998.985 1111.770 1999.275 1112.495 ;
        RECT 1999.535 1112.420 2000.955 1112.590 ;
        RECT 1999.535 1111.940 1999.705 1112.420 ;
        RECT 1999.875 1111.770 2000.205 1112.250 ;
        RECT 2000.375 1111.945 2000.545 1112.420 ;
        RECT 2000.715 1111.770 2001.045 1112.250 ;
        RECT 2001.555 1111.770 2001.885 1112.250 ;
        RECT 2002.395 1111.770 2002.725 1112.250 ;
        RECT 2003.235 1111.770 2003.565 1112.250 ;
        RECT 2004.075 1111.770 2004.405 1112.570 ;
        RECT 2004.965 1111.770 2005.255 1112.495 ;
        RECT 2005.515 1112.420 2006.935 1112.590 ;
        RECT 2005.515 1111.940 2005.685 1112.420 ;
        RECT 2005.855 1111.770 2006.185 1112.250 ;
        RECT 2006.355 1111.945 2006.525 1112.420 ;
        RECT 2006.695 1111.770 2007.025 1112.250 ;
        RECT 2007.535 1111.770 2007.865 1112.250 ;
        RECT 2008.375 1111.770 2008.705 1112.250 ;
        RECT 2009.215 1111.770 2009.545 1112.250 ;
        RECT 2010.055 1111.770 2010.385 1112.570 ;
        RECT 2010.945 1111.770 2011.235 1112.495 ;
        RECT 2011.495 1112.420 2012.915 1112.590 ;
        RECT 2011.495 1111.940 2011.665 1112.420 ;
        RECT 2011.835 1111.770 2012.165 1112.250 ;
        RECT 2012.335 1111.945 2012.505 1112.420 ;
        RECT 2012.675 1111.770 2013.005 1112.250 ;
        RECT 2013.515 1111.770 2013.845 1112.250 ;
        RECT 2014.355 1111.770 2014.685 1112.250 ;
        RECT 2015.195 1111.770 2015.525 1112.250 ;
        RECT 2016.035 1111.770 2016.365 1112.570 ;
        RECT 2016.925 1111.770 2017.215 1112.495 ;
        RECT 2017.475 1112.420 2018.895 1112.590 ;
        RECT 2017.475 1111.940 2017.645 1112.420 ;
        RECT 2017.815 1111.770 2018.145 1112.250 ;
        RECT 2018.315 1111.945 2018.485 1112.420 ;
        RECT 2018.655 1111.770 2018.985 1112.250 ;
        RECT 2019.495 1111.770 2019.825 1112.250 ;
        RECT 2020.335 1111.770 2020.665 1112.250 ;
        RECT 2021.175 1111.770 2021.505 1112.250 ;
        RECT 2022.015 1111.770 2022.345 1112.570 ;
        RECT 2022.905 1111.770 2023.195 1112.495 ;
        RECT 2023.455 1112.420 2024.875 1112.590 ;
        RECT 2023.455 1111.940 2023.625 1112.420 ;
        RECT 2023.795 1111.770 2024.125 1112.250 ;
        RECT 2024.295 1111.945 2024.465 1112.420 ;
        RECT 2024.635 1111.770 2024.965 1112.250 ;
        RECT 2025.475 1111.770 2025.805 1112.250 ;
        RECT 2026.315 1111.770 2026.645 1112.250 ;
        RECT 2027.155 1111.770 2027.485 1112.250 ;
        RECT 2027.995 1111.770 2028.325 1112.570 ;
        RECT 2028.885 1111.770 2029.175 1112.495 ;
        RECT 2029.435 1112.420 2030.855 1112.590 ;
        RECT 2029.435 1111.940 2029.605 1112.420 ;
        RECT 2029.775 1111.770 2030.105 1112.250 ;
        RECT 2030.275 1111.945 2030.445 1112.420 ;
        RECT 2030.615 1111.770 2030.945 1112.250 ;
        RECT 2031.455 1111.770 2031.785 1112.250 ;
        RECT 2032.295 1111.770 2032.625 1112.250 ;
        RECT 2033.135 1111.770 2033.465 1112.250 ;
        RECT 2033.975 1111.770 2034.305 1112.570 ;
        RECT 2034.865 1111.770 2035.155 1112.495 ;
        RECT 2035.415 1112.420 2036.835 1112.590 ;
        RECT 2035.415 1111.940 2035.585 1112.420 ;
        RECT 2035.755 1111.770 2036.085 1112.250 ;
        RECT 2036.255 1111.945 2036.425 1112.420 ;
        RECT 2036.595 1111.770 2036.925 1112.250 ;
        RECT 2037.435 1111.770 2037.765 1112.250 ;
        RECT 2038.275 1111.770 2038.605 1112.250 ;
        RECT 2039.115 1111.770 2039.445 1112.250 ;
        RECT 2039.955 1111.770 2040.285 1112.570 ;
        RECT 2040.845 1111.770 2041.135 1112.495 ;
        RECT 2041.395 1112.420 2042.815 1112.590 ;
        RECT 2041.395 1111.940 2041.565 1112.420 ;
        RECT 2041.735 1111.770 2042.065 1112.250 ;
        RECT 2042.235 1111.945 2042.405 1112.420 ;
        RECT 2042.575 1111.770 2042.905 1112.250 ;
        RECT 2043.415 1111.770 2043.745 1112.250 ;
        RECT 2044.255 1111.770 2044.585 1112.250 ;
        RECT 2045.095 1111.770 2045.425 1112.250 ;
        RECT 2045.935 1111.770 2046.265 1112.570 ;
        RECT 2046.825 1111.770 2047.115 1112.495 ;
        RECT 2047.375 1112.420 2048.795 1112.590 ;
        RECT 2047.375 1111.940 2047.545 1112.420 ;
        RECT 2047.715 1111.770 2048.045 1112.250 ;
        RECT 2048.215 1111.945 2048.385 1112.420 ;
        RECT 2048.555 1111.770 2048.885 1112.250 ;
        RECT 2049.395 1111.770 2049.725 1112.250 ;
        RECT 2050.235 1111.770 2050.565 1112.250 ;
        RECT 2051.075 1111.770 2051.405 1112.250 ;
        RECT 2051.915 1111.770 2052.245 1112.570 ;
        RECT 2052.805 1111.770 2053.095 1112.495 ;
        RECT 2053.355 1112.420 2054.775 1112.590 ;
        RECT 2053.355 1111.940 2053.525 1112.420 ;
        RECT 2053.695 1111.770 2054.025 1112.250 ;
        RECT 2054.195 1111.945 2054.365 1112.420 ;
        RECT 2054.535 1111.770 2054.865 1112.250 ;
        RECT 2055.375 1111.770 2055.705 1112.250 ;
        RECT 2056.215 1111.770 2056.545 1112.250 ;
        RECT 2057.055 1111.770 2057.385 1112.250 ;
        RECT 2057.895 1111.770 2058.225 1112.570 ;
        RECT 2058.785 1111.770 2059.075 1112.495 ;
        RECT 2059.335 1112.420 2060.755 1112.590 ;
        RECT 2059.335 1111.940 2059.505 1112.420 ;
        RECT 2059.675 1111.770 2060.005 1112.250 ;
        RECT 2060.175 1111.945 2060.345 1112.420 ;
        RECT 2060.515 1111.770 2060.845 1112.250 ;
        RECT 2061.355 1111.770 2061.685 1112.250 ;
        RECT 2062.195 1111.770 2062.525 1112.250 ;
        RECT 2063.035 1111.770 2063.365 1112.250 ;
        RECT 2063.875 1111.770 2064.205 1112.570 ;
        RECT 2064.765 1111.770 2065.055 1112.495 ;
        RECT 2065.315 1112.420 2066.735 1112.590 ;
        RECT 2065.315 1111.940 2065.485 1112.420 ;
        RECT 2065.655 1111.770 2065.985 1112.250 ;
        RECT 2066.155 1111.945 2066.325 1112.420 ;
        RECT 2066.495 1111.770 2066.825 1112.250 ;
        RECT 2067.335 1111.770 2067.665 1112.250 ;
        RECT 2068.175 1111.770 2068.505 1112.250 ;
        RECT 2069.015 1111.770 2069.345 1112.250 ;
        RECT 2069.855 1111.770 2070.185 1112.570 ;
        RECT 2070.745 1111.770 2071.035 1112.495 ;
        RECT 2071.295 1112.420 2072.715 1112.590 ;
        RECT 2071.295 1111.940 2071.465 1112.420 ;
        RECT 2071.635 1111.770 2071.965 1112.250 ;
        RECT 2072.135 1111.945 2072.305 1112.420 ;
        RECT 2072.475 1111.770 2072.805 1112.250 ;
        RECT 2073.315 1111.770 2073.645 1112.250 ;
        RECT 2074.155 1111.770 2074.485 1112.250 ;
        RECT 2074.995 1111.770 2075.325 1112.250 ;
        RECT 2075.835 1111.770 2076.165 1112.570 ;
        RECT 2076.725 1111.770 2077.015 1112.495 ;
        RECT 2077.275 1112.420 2078.695 1112.590 ;
        RECT 2077.275 1111.940 2077.445 1112.420 ;
        RECT 2077.615 1111.770 2077.945 1112.250 ;
        RECT 2078.115 1111.945 2078.285 1112.420 ;
        RECT 2078.455 1111.770 2078.785 1112.250 ;
        RECT 2079.295 1111.770 2079.625 1112.250 ;
        RECT 2080.135 1111.770 2080.465 1112.250 ;
        RECT 2080.975 1111.770 2081.305 1112.250 ;
        RECT 2081.815 1111.770 2082.145 1112.570 ;
        RECT 2082.705 1111.770 2082.995 1112.495 ;
        RECT 2083.255 1112.420 2084.675 1112.590 ;
      LAYER li1 ;
        RECT 2090.035 1112.590 2090.290 1113.130 ;
      LAYER li1 ;
        RECT 2092.985 1112.930 2093.160 1113.130 ;
        RECT 2090.535 1112.760 2093.160 1112.930 ;
        RECT 2092.985 1112.590 2093.160 1112.760 ;
        RECT 2083.255 1111.940 2083.425 1112.420 ;
        RECT 2083.595 1111.770 2083.925 1112.250 ;
        RECT 2084.095 1111.945 2084.265 1112.420 ;
        RECT 2084.435 1111.770 2084.765 1112.250 ;
        RECT 2085.275 1111.770 2085.605 1112.250 ;
        RECT 2086.115 1111.770 2086.445 1112.250 ;
        RECT 2086.955 1111.770 2087.285 1112.250 ;
        RECT 2087.795 1111.770 2088.125 1112.570 ;
        RECT 2088.685 1111.770 2088.975 1112.495 ;
        RECT 2089.535 1111.770 2089.865 1112.570 ;
      LAYER li1 ;
        RECT 2090.035 1112.420 2092.725 1112.590 ;
      LAYER li1 ;
        RECT 2092.985 1112.420 2094.405 1112.590 ;
      LAYER li1 ;
        RECT 2090.035 1111.940 2090.205 1112.420 ;
      LAYER li1 ;
        RECT 2090.375 1111.770 2090.705 1112.250 ;
      LAYER li1 ;
        RECT 2090.875 1111.940 2091.045 1112.420 ;
      LAYER li1 ;
        RECT 2091.215 1111.770 2091.545 1112.250 ;
      LAYER li1 ;
        RECT 2091.715 1111.940 2091.885 1112.420 ;
      LAYER li1 ;
        RECT 2092.055 1111.770 2092.385 1112.250 ;
      LAYER li1 ;
        RECT 2092.555 1111.940 2092.725 1112.420 ;
      LAYER li1 ;
        RECT 2092.895 1111.770 2093.225 1112.250 ;
        RECT 2093.395 1111.945 2093.565 1112.420 ;
        RECT 2093.735 1111.770 2094.065 1112.250 ;
        RECT 2094.235 1111.940 2094.405 1112.420 ;
        RECT 2094.665 1111.770 2094.955 1112.495 ;
        RECT 674.980 1111.600 675.125 1111.770 ;
        RECT 675.295 1111.600 675.585 1111.770 ;
        RECT 675.755 1111.600 676.045 1111.770 ;
        RECT 676.215 1111.600 676.505 1111.770 ;
        RECT 676.675 1111.600 676.965 1111.770 ;
        RECT 677.135 1111.600 677.425 1111.770 ;
        RECT 677.595 1111.600 677.885 1111.770 ;
        RECT 678.055 1111.600 678.345 1111.770 ;
        RECT 678.515 1111.600 678.805 1111.770 ;
        RECT 678.975 1111.600 679.265 1111.770 ;
        RECT 679.435 1111.600 679.725 1111.770 ;
        RECT 679.895 1111.600 680.185 1111.770 ;
        RECT 680.355 1111.600 680.645 1111.770 ;
        RECT 680.815 1111.600 681.105 1111.770 ;
        RECT 681.275 1111.600 681.565 1111.770 ;
        RECT 681.735 1111.600 682.025 1111.770 ;
        RECT 682.195 1111.600 682.485 1111.770 ;
        RECT 682.655 1111.600 682.945 1111.770 ;
        RECT 683.115 1111.600 683.405 1111.770 ;
        RECT 683.575 1111.600 683.865 1111.770 ;
        RECT 684.035 1111.600 684.325 1111.770 ;
        RECT 684.495 1111.600 684.785 1111.770 ;
        RECT 684.955 1111.600 685.245 1111.770 ;
        RECT 685.415 1111.600 685.705 1111.770 ;
        RECT 685.875 1111.600 686.165 1111.770 ;
        RECT 686.335 1111.600 686.625 1111.770 ;
        RECT 686.795 1111.600 687.085 1111.770 ;
        RECT 687.255 1111.600 687.545 1111.770 ;
        RECT 687.715 1111.600 688.005 1111.770 ;
        RECT 688.175 1111.600 688.465 1111.770 ;
        RECT 688.635 1111.600 688.925 1111.770 ;
        RECT 689.095 1111.600 689.385 1111.770 ;
        RECT 689.555 1111.600 689.845 1111.770 ;
        RECT 690.015 1111.600 690.305 1111.770 ;
        RECT 690.475 1111.600 690.765 1111.770 ;
        RECT 690.935 1111.600 691.225 1111.770 ;
        RECT 691.395 1111.600 691.685 1111.770 ;
        RECT 691.855 1111.600 692.145 1111.770 ;
        RECT 692.315 1111.600 692.605 1111.770 ;
        RECT 692.775 1111.600 693.065 1111.770 ;
        RECT 693.235 1111.600 693.525 1111.770 ;
        RECT 693.695 1111.600 693.985 1111.770 ;
        RECT 694.155 1111.600 694.445 1111.770 ;
        RECT 694.615 1111.600 694.905 1111.770 ;
        RECT 695.075 1111.600 695.365 1111.770 ;
        RECT 695.535 1111.600 695.825 1111.770 ;
        RECT 695.995 1111.600 696.285 1111.770 ;
        RECT 696.455 1111.600 696.745 1111.770 ;
        RECT 696.915 1111.600 697.205 1111.770 ;
        RECT 697.375 1111.600 697.665 1111.770 ;
        RECT 697.835 1111.600 698.125 1111.770 ;
        RECT 698.295 1111.600 698.585 1111.770 ;
        RECT 698.755 1111.600 699.045 1111.770 ;
        RECT 699.215 1111.600 699.505 1111.770 ;
        RECT 699.675 1111.600 699.965 1111.770 ;
        RECT 700.135 1111.600 700.425 1111.770 ;
        RECT 700.595 1111.600 700.885 1111.770 ;
        RECT 701.055 1111.600 701.345 1111.770 ;
        RECT 701.515 1111.600 701.805 1111.770 ;
        RECT 701.975 1111.600 702.265 1111.770 ;
        RECT 702.435 1111.600 702.725 1111.770 ;
        RECT 702.895 1111.600 703.185 1111.770 ;
        RECT 703.355 1111.600 703.645 1111.770 ;
        RECT 703.815 1111.600 704.105 1111.770 ;
        RECT 704.275 1111.600 704.565 1111.770 ;
        RECT 704.735 1111.600 705.025 1111.770 ;
        RECT 705.195 1111.600 705.485 1111.770 ;
        RECT 705.655 1111.600 705.945 1111.770 ;
        RECT 706.115 1111.600 706.405 1111.770 ;
        RECT 706.575 1111.600 706.865 1111.770 ;
        RECT 707.035 1111.600 707.325 1111.770 ;
        RECT 707.495 1111.600 707.785 1111.770 ;
        RECT 707.955 1111.600 708.245 1111.770 ;
        RECT 708.415 1111.600 708.705 1111.770 ;
        RECT 708.875 1111.600 709.165 1111.770 ;
        RECT 709.335 1111.600 709.625 1111.770 ;
        RECT 709.795 1111.600 710.085 1111.770 ;
        RECT 710.255 1111.600 710.545 1111.770 ;
        RECT 710.715 1111.600 711.005 1111.770 ;
        RECT 711.175 1111.600 711.465 1111.770 ;
        RECT 711.635 1111.600 711.925 1111.770 ;
        RECT 712.095 1111.600 712.385 1111.770 ;
        RECT 712.555 1111.600 712.845 1111.770 ;
        RECT 713.015 1111.600 713.305 1111.770 ;
        RECT 713.475 1111.600 713.765 1111.770 ;
        RECT 713.935 1111.600 714.225 1111.770 ;
        RECT 714.395 1111.600 714.685 1111.770 ;
        RECT 714.855 1111.600 715.145 1111.770 ;
        RECT 715.315 1111.600 715.605 1111.770 ;
        RECT 715.775 1111.600 716.065 1111.770 ;
        RECT 716.235 1111.600 716.525 1111.770 ;
        RECT 716.695 1111.600 716.985 1111.770 ;
        RECT 717.155 1111.600 717.445 1111.770 ;
        RECT 717.615 1111.600 717.905 1111.770 ;
        RECT 718.075 1111.600 718.365 1111.770 ;
        RECT 718.535 1111.600 718.825 1111.770 ;
        RECT 718.995 1111.600 719.285 1111.770 ;
        RECT 719.455 1111.600 719.745 1111.770 ;
        RECT 719.915 1111.600 720.205 1111.770 ;
        RECT 720.375 1111.600 720.665 1111.770 ;
        RECT 720.835 1111.600 721.125 1111.770 ;
        RECT 721.295 1111.600 721.585 1111.770 ;
        RECT 721.755 1111.600 722.045 1111.770 ;
        RECT 722.215 1111.600 722.505 1111.770 ;
        RECT 722.675 1111.600 722.965 1111.770 ;
        RECT 723.135 1111.600 723.425 1111.770 ;
        RECT 723.595 1111.600 723.885 1111.770 ;
        RECT 724.055 1111.600 724.345 1111.770 ;
        RECT 724.515 1111.600 724.805 1111.770 ;
        RECT 724.975 1111.600 725.265 1111.770 ;
        RECT 725.435 1111.600 725.725 1111.770 ;
        RECT 725.895 1111.600 726.185 1111.770 ;
        RECT 726.355 1111.600 726.645 1111.770 ;
        RECT 726.815 1111.600 727.105 1111.770 ;
        RECT 727.275 1111.600 727.565 1111.770 ;
        RECT 727.735 1111.600 728.025 1111.770 ;
        RECT 728.195 1111.600 728.485 1111.770 ;
        RECT 728.655 1111.600 728.945 1111.770 ;
        RECT 729.115 1111.600 729.405 1111.770 ;
        RECT 729.575 1111.600 729.865 1111.770 ;
        RECT 730.035 1111.600 730.325 1111.770 ;
        RECT 730.495 1111.600 730.785 1111.770 ;
        RECT 730.955 1111.600 731.245 1111.770 ;
        RECT 731.415 1111.600 731.705 1111.770 ;
        RECT 731.875 1111.600 732.165 1111.770 ;
        RECT 732.335 1111.600 732.625 1111.770 ;
        RECT 732.795 1111.600 733.085 1111.770 ;
        RECT 733.255 1111.600 733.545 1111.770 ;
        RECT 733.715 1111.600 734.005 1111.770 ;
        RECT 734.175 1111.600 734.465 1111.770 ;
        RECT 734.635 1111.600 734.925 1111.770 ;
        RECT 735.095 1111.600 735.385 1111.770 ;
        RECT 735.555 1111.600 735.845 1111.770 ;
        RECT 736.015 1111.600 736.305 1111.770 ;
        RECT 736.475 1111.600 736.765 1111.770 ;
        RECT 736.935 1111.600 737.225 1111.770 ;
        RECT 737.395 1111.600 737.685 1111.770 ;
        RECT 737.855 1111.600 738.145 1111.770 ;
        RECT 738.315 1111.600 738.605 1111.770 ;
        RECT 738.775 1111.600 739.065 1111.770 ;
        RECT 739.235 1111.600 739.525 1111.770 ;
        RECT 739.695 1111.600 739.985 1111.770 ;
        RECT 740.155 1111.600 740.445 1111.770 ;
        RECT 740.615 1111.600 740.905 1111.770 ;
        RECT 741.075 1111.600 741.365 1111.770 ;
        RECT 741.535 1111.600 741.825 1111.770 ;
        RECT 741.995 1111.600 742.285 1111.770 ;
        RECT 742.455 1111.600 742.745 1111.770 ;
        RECT 742.915 1111.600 743.205 1111.770 ;
        RECT 743.375 1111.600 743.665 1111.770 ;
        RECT 743.835 1111.600 744.125 1111.770 ;
        RECT 744.295 1111.600 744.585 1111.770 ;
        RECT 744.755 1111.600 745.045 1111.770 ;
        RECT 745.215 1111.600 745.505 1111.770 ;
        RECT 745.675 1111.600 745.965 1111.770 ;
        RECT 746.135 1111.600 746.425 1111.770 ;
        RECT 746.595 1111.600 746.885 1111.770 ;
        RECT 747.055 1111.600 747.345 1111.770 ;
        RECT 747.515 1111.600 747.805 1111.770 ;
        RECT 747.975 1111.600 748.265 1111.770 ;
        RECT 748.435 1111.600 748.725 1111.770 ;
        RECT 748.895 1111.600 749.185 1111.770 ;
        RECT 749.355 1111.600 749.645 1111.770 ;
        RECT 749.815 1111.600 750.105 1111.770 ;
        RECT 750.275 1111.600 750.565 1111.770 ;
        RECT 750.735 1111.600 751.025 1111.770 ;
        RECT 751.195 1111.600 751.485 1111.770 ;
        RECT 751.655 1111.600 751.945 1111.770 ;
        RECT 752.115 1111.600 752.405 1111.770 ;
        RECT 752.575 1111.600 752.865 1111.770 ;
        RECT 753.035 1111.600 753.325 1111.770 ;
        RECT 753.495 1111.600 753.785 1111.770 ;
        RECT 753.955 1111.600 754.245 1111.770 ;
        RECT 754.415 1111.600 754.705 1111.770 ;
        RECT 754.875 1111.600 755.165 1111.770 ;
        RECT 755.335 1111.600 755.625 1111.770 ;
        RECT 755.795 1111.600 756.085 1111.770 ;
        RECT 756.255 1111.600 756.545 1111.770 ;
        RECT 756.715 1111.600 757.005 1111.770 ;
        RECT 757.175 1111.600 757.465 1111.770 ;
        RECT 757.635 1111.600 757.925 1111.770 ;
        RECT 758.095 1111.600 758.385 1111.770 ;
        RECT 758.555 1111.600 758.845 1111.770 ;
        RECT 759.015 1111.600 759.305 1111.770 ;
        RECT 759.475 1111.600 759.765 1111.770 ;
        RECT 759.935 1111.600 760.225 1111.770 ;
        RECT 760.395 1111.600 760.685 1111.770 ;
        RECT 760.855 1111.600 761.145 1111.770 ;
        RECT 761.315 1111.600 761.605 1111.770 ;
        RECT 761.775 1111.600 762.065 1111.770 ;
        RECT 762.235 1111.600 762.525 1111.770 ;
        RECT 762.695 1111.600 762.985 1111.770 ;
        RECT 763.155 1111.600 763.445 1111.770 ;
        RECT 763.615 1111.600 763.905 1111.770 ;
        RECT 764.075 1111.600 764.365 1111.770 ;
        RECT 764.535 1111.600 764.825 1111.770 ;
        RECT 764.995 1111.600 765.285 1111.770 ;
        RECT 765.455 1111.600 765.745 1111.770 ;
        RECT 765.915 1111.600 766.205 1111.770 ;
        RECT 766.375 1111.600 766.665 1111.770 ;
        RECT 766.835 1111.600 767.125 1111.770 ;
        RECT 767.295 1111.600 767.585 1111.770 ;
        RECT 767.755 1111.600 768.045 1111.770 ;
        RECT 768.215 1111.600 768.505 1111.770 ;
        RECT 768.675 1111.600 768.965 1111.770 ;
        RECT 769.135 1111.600 769.425 1111.770 ;
        RECT 769.595 1111.600 769.885 1111.770 ;
        RECT 770.055 1111.600 770.345 1111.770 ;
        RECT 770.515 1111.600 770.805 1111.770 ;
        RECT 770.975 1111.600 771.265 1111.770 ;
        RECT 771.435 1111.600 771.725 1111.770 ;
        RECT 771.895 1111.600 772.185 1111.770 ;
        RECT 772.355 1111.600 772.645 1111.770 ;
        RECT 772.815 1111.600 773.105 1111.770 ;
        RECT 773.275 1111.600 773.565 1111.770 ;
        RECT 773.735 1111.600 774.025 1111.770 ;
        RECT 774.195 1111.600 774.485 1111.770 ;
        RECT 774.655 1111.600 774.945 1111.770 ;
        RECT 775.115 1111.600 775.405 1111.770 ;
        RECT 775.575 1111.600 775.865 1111.770 ;
        RECT 776.035 1111.600 776.325 1111.770 ;
        RECT 776.495 1111.600 776.785 1111.770 ;
        RECT 776.955 1111.600 777.245 1111.770 ;
        RECT 777.415 1111.600 777.705 1111.770 ;
        RECT 777.875 1111.600 778.165 1111.770 ;
        RECT 778.335 1111.600 778.625 1111.770 ;
        RECT 778.795 1111.600 779.085 1111.770 ;
        RECT 779.255 1111.600 779.545 1111.770 ;
        RECT 779.715 1111.600 780.005 1111.770 ;
        RECT 780.175 1111.600 780.465 1111.770 ;
        RECT 780.635 1111.600 780.925 1111.770 ;
        RECT 781.095 1111.600 781.385 1111.770 ;
        RECT 781.555 1111.600 781.845 1111.770 ;
        RECT 782.015 1111.600 782.305 1111.770 ;
        RECT 782.475 1111.600 782.765 1111.770 ;
        RECT 782.935 1111.600 783.225 1111.770 ;
        RECT 783.395 1111.600 783.685 1111.770 ;
        RECT 783.855 1111.600 784.145 1111.770 ;
        RECT 784.315 1111.600 784.605 1111.770 ;
        RECT 784.775 1111.600 785.065 1111.770 ;
        RECT 785.235 1111.600 785.525 1111.770 ;
        RECT 785.695 1111.600 785.985 1111.770 ;
        RECT 786.155 1111.600 786.445 1111.770 ;
        RECT 786.615 1111.600 786.905 1111.770 ;
        RECT 787.075 1111.600 787.365 1111.770 ;
        RECT 787.535 1111.600 787.825 1111.770 ;
        RECT 787.995 1111.600 788.285 1111.770 ;
        RECT 788.455 1111.600 788.745 1111.770 ;
        RECT 788.915 1111.600 789.205 1111.770 ;
        RECT 789.375 1111.600 789.665 1111.770 ;
        RECT 789.835 1111.600 790.125 1111.770 ;
        RECT 790.295 1111.600 790.585 1111.770 ;
        RECT 790.755 1111.600 791.045 1111.770 ;
        RECT 791.215 1111.600 791.505 1111.770 ;
        RECT 791.675 1111.600 791.965 1111.770 ;
        RECT 792.135 1111.600 792.425 1111.770 ;
        RECT 792.595 1111.600 792.885 1111.770 ;
        RECT 793.055 1111.600 793.345 1111.770 ;
        RECT 793.515 1111.600 793.805 1111.770 ;
        RECT 793.975 1111.600 794.265 1111.770 ;
        RECT 794.435 1111.600 794.725 1111.770 ;
        RECT 794.895 1111.600 795.040 1111.770 ;
        RECT 1974.980 1111.600 1975.125 1111.770 ;
        RECT 1975.295 1111.600 1975.585 1111.770 ;
        RECT 1975.755 1111.600 1976.045 1111.770 ;
        RECT 1976.215 1111.600 1976.505 1111.770 ;
        RECT 1976.675 1111.600 1976.965 1111.770 ;
        RECT 1977.135 1111.600 1977.425 1111.770 ;
        RECT 1977.595 1111.600 1977.885 1111.770 ;
        RECT 1978.055 1111.600 1978.345 1111.770 ;
        RECT 1978.515 1111.600 1978.805 1111.770 ;
        RECT 1978.975 1111.600 1979.265 1111.770 ;
        RECT 1979.435 1111.600 1979.725 1111.770 ;
        RECT 1979.895 1111.600 1980.185 1111.770 ;
        RECT 1980.355 1111.600 1980.645 1111.770 ;
        RECT 1980.815 1111.600 1981.105 1111.770 ;
        RECT 1981.275 1111.600 1981.565 1111.770 ;
        RECT 1981.735 1111.600 1982.025 1111.770 ;
        RECT 1982.195 1111.600 1982.485 1111.770 ;
        RECT 1982.655 1111.600 1982.945 1111.770 ;
        RECT 1983.115 1111.600 1983.405 1111.770 ;
        RECT 1983.575 1111.600 1983.865 1111.770 ;
        RECT 1984.035 1111.600 1984.325 1111.770 ;
        RECT 1984.495 1111.600 1984.785 1111.770 ;
        RECT 1984.955 1111.600 1985.245 1111.770 ;
        RECT 1985.415 1111.600 1985.705 1111.770 ;
        RECT 1985.875 1111.600 1986.165 1111.770 ;
        RECT 1986.335 1111.600 1986.625 1111.770 ;
        RECT 1986.795 1111.600 1987.085 1111.770 ;
        RECT 1987.255 1111.600 1987.545 1111.770 ;
        RECT 1987.715 1111.600 1988.005 1111.770 ;
        RECT 1988.175 1111.600 1988.465 1111.770 ;
        RECT 1988.635 1111.600 1988.925 1111.770 ;
        RECT 1989.095 1111.600 1989.385 1111.770 ;
        RECT 1989.555 1111.600 1989.845 1111.770 ;
        RECT 1990.015 1111.600 1990.305 1111.770 ;
        RECT 1990.475 1111.600 1990.765 1111.770 ;
        RECT 1990.935 1111.600 1991.225 1111.770 ;
        RECT 1991.395 1111.600 1991.685 1111.770 ;
        RECT 1991.855 1111.600 1992.145 1111.770 ;
        RECT 1992.315 1111.600 1992.605 1111.770 ;
        RECT 1992.775 1111.600 1993.065 1111.770 ;
        RECT 1993.235 1111.600 1993.525 1111.770 ;
        RECT 1993.695 1111.600 1993.985 1111.770 ;
        RECT 1994.155 1111.600 1994.445 1111.770 ;
        RECT 1994.615 1111.600 1994.905 1111.770 ;
        RECT 1995.075 1111.600 1995.365 1111.770 ;
        RECT 1995.535 1111.600 1995.825 1111.770 ;
        RECT 1995.995 1111.600 1996.285 1111.770 ;
        RECT 1996.455 1111.600 1996.745 1111.770 ;
        RECT 1996.915 1111.600 1997.205 1111.770 ;
        RECT 1997.375 1111.600 1997.665 1111.770 ;
        RECT 1997.835 1111.600 1998.125 1111.770 ;
        RECT 1998.295 1111.600 1998.585 1111.770 ;
        RECT 1998.755 1111.600 1999.045 1111.770 ;
        RECT 1999.215 1111.600 1999.505 1111.770 ;
        RECT 1999.675 1111.600 1999.965 1111.770 ;
        RECT 2000.135 1111.600 2000.425 1111.770 ;
        RECT 2000.595 1111.600 2000.885 1111.770 ;
        RECT 2001.055 1111.600 2001.345 1111.770 ;
        RECT 2001.515 1111.600 2001.805 1111.770 ;
        RECT 2001.975 1111.600 2002.265 1111.770 ;
        RECT 2002.435 1111.600 2002.725 1111.770 ;
        RECT 2002.895 1111.600 2003.185 1111.770 ;
        RECT 2003.355 1111.600 2003.645 1111.770 ;
        RECT 2003.815 1111.600 2004.105 1111.770 ;
        RECT 2004.275 1111.600 2004.565 1111.770 ;
        RECT 2004.735 1111.600 2005.025 1111.770 ;
        RECT 2005.195 1111.600 2005.485 1111.770 ;
        RECT 2005.655 1111.600 2005.945 1111.770 ;
        RECT 2006.115 1111.600 2006.405 1111.770 ;
        RECT 2006.575 1111.600 2006.865 1111.770 ;
        RECT 2007.035 1111.600 2007.325 1111.770 ;
        RECT 2007.495 1111.600 2007.785 1111.770 ;
        RECT 2007.955 1111.600 2008.245 1111.770 ;
        RECT 2008.415 1111.600 2008.705 1111.770 ;
        RECT 2008.875 1111.600 2009.165 1111.770 ;
        RECT 2009.335 1111.600 2009.625 1111.770 ;
        RECT 2009.795 1111.600 2010.085 1111.770 ;
        RECT 2010.255 1111.600 2010.545 1111.770 ;
        RECT 2010.715 1111.600 2011.005 1111.770 ;
        RECT 2011.175 1111.600 2011.465 1111.770 ;
        RECT 2011.635 1111.600 2011.925 1111.770 ;
        RECT 2012.095 1111.600 2012.385 1111.770 ;
        RECT 2012.555 1111.600 2012.845 1111.770 ;
        RECT 2013.015 1111.600 2013.305 1111.770 ;
        RECT 2013.475 1111.600 2013.765 1111.770 ;
        RECT 2013.935 1111.600 2014.225 1111.770 ;
        RECT 2014.395 1111.600 2014.685 1111.770 ;
        RECT 2014.855 1111.600 2015.145 1111.770 ;
        RECT 2015.315 1111.600 2015.605 1111.770 ;
        RECT 2015.775 1111.600 2016.065 1111.770 ;
        RECT 2016.235 1111.600 2016.525 1111.770 ;
        RECT 2016.695 1111.600 2016.985 1111.770 ;
        RECT 2017.155 1111.600 2017.445 1111.770 ;
        RECT 2017.615 1111.600 2017.905 1111.770 ;
        RECT 2018.075 1111.600 2018.365 1111.770 ;
        RECT 2018.535 1111.600 2018.825 1111.770 ;
        RECT 2018.995 1111.600 2019.285 1111.770 ;
        RECT 2019.455 1111.600 2019.745 1111.770 ;
        RECT 2019.915 1111.600 2020.205 1111.770 ;
        RECT 2020.375 1111.600 2020.665 1111.770 ;
        RECT 2020.835 1111.600 2021.125 1111.770 ;
        RECT 2021.295 1111.600 2021.585 1111.770 ;
        RECT 2021.755 1111.600 2022.045 1111.770 ;
        RECT 2022.215 1111.600 2022.505 1111.770 ;
        RECT 2022.675 1111.600 2022.965 1111.770 ;
        RECT 2023.135 1111.600 2023.425 1111.770 ;
        RECT 2023.595 1111.600 2023.885 1111.770 ;
        RECT 2024.055 1111.600 2024.345 1111.770 ;
        RECT 2024.515 1111.600 2024.805 1111.770 ;
        RECT 2024.975 1111.600 2025.265 1111.770 ;
        RECT 2025.435 1111.600 2025.725 1111.770 ;
        RECT 2025.895 1111.600 2026.185 1111.770 ;
        RECT 2026.355 1111.600 2026.645 1111.770 ;
        RECT 2026.815 1111.600 2027.105 1111.770 ;
        RECT 2027.275 1111.600 2027.565 1111.770 ;
        RECT 2027.735 1111.600 2028.025 1111.770 ;
        RECT 2028.195 1111.600 2028.485 1111.770 ;
        RECT 2028.655 1111.600 2028.945 1111.770 ;
        RECT 2029.115 1111.600 2029.405 1111.770 ;
        RECT 2029.575 1111.600 2029.865 1111.770 ;
        RECT 2030.035 1111.600 2030.325 1111.770 ;
        RECT 2030.495 1111.600 2030.785 1111.770 ;
        RECT 2030.955 1111.600 2031.245 1111.770 ;
        RECT 2031.415 1111.600 2031.705 1111.770 ;
        RECT 2031.875 1111.600 2032.165 1111.770 ;
        RECT 2032.335 1111.600 2032.625 1111.770 ;
        RECT 2032.795 1111.600 2033.085 1111.770 ;
        RECT 2033.255 1111.600 2033.545 1111.770 ;
        RECT 2033.715 1111.600 2034.005 1111.770 ;
        RECT 2034.175 1111.600 2034.465 1111.770 ;
        RECT 2034.635 1111.600 2034.925 1111.770 ;
        RECT 2035.095 1111.600 2035.385 1111.770 ;
        RECT 2035.555 1111.600 2035.845 1111.770 ;
        RECT 2036.015 1111.600 2036.305 1111.770 ;
        RECT 2036.475 1111.600 2036.765 1111.770 ;
        RECT 2036.935 1111.600 2037.225 1111.770 ;
        RECT 2037.395 1111.600 2037.685 1111.770 ;
        RECT 2037.855 1111.600 2038.145 1111.770 ;
        RECT 2038.315 1111.600 2038.605 1111.770 ;
        RECT 2038.775 1111.600 2039.065 1111.770 ;
        RECT 2039.235 1111.600 2039.525 1111.770 ;
        RECT 2039.695 1111.600 2039.985 1111.770 ;
        RECT 2040.155 1111.600 2040.445 1111.770 ;
        RECT 2040.615 1111.600 2040.905 1111.770 ;
        RECT 2041.075 1111.600 2041.365 1111.770 ;
        RECT 2041.535 1111.600 2041.825 1111.770 ;
        RECT 2041.995 1111.600 2042.285 1111.770 ;
        RECT 2042.455 1111.600 2042.745 1111.770 ;
        RECT 2042.915 1111.600 2043.205 1111.770 ;
        RECT 2043.375 1111.600 2043.665 1111.770 ;
        RECT 2043.835 1111.600 2044.125 1111.770 ;
        RECT 2044.295 1111.600 2044.585 1111.770 ;
        RECT 2044.755 1111.600 2045.045 1111.770 ;
        RECT 2045.215 1111.600 2045.505 1111.770 ;
        RECT 2045.675 1111.600 2045.965 1111.770 ;
        RECT 2046.135 1111.600 2046.425 1111.770 ;
        RECT 2046.595 1111.600 2046.885 1111.770 ;
        RECT 2047.055 1111.600 2047.345 1111.770 ;
        RECT 2047.515 1111.600 2047.805 1111.770 ;
        RECT 2047.975 1111.600 2048.265 1111.770 ;
        RECT 2048.435 1111.600 2048.725 1111.770 ;
        RECT 2048.895 1111.600 2049.185 1111.770 ;
        RECT 2049.355 1111.600 2049.645 1111.770 ;
        RECT 2049.815 1111.600 2050.105 1111.770 ;
        RECT 2050.275 1111.600 2050.565 1111.770 ;
        RECT 2050.735 1111.600 2051.025 1111.770 ;
        RECT 2051.195 1111.600 2051.485 1111.770 ;
        RECT 2051.655 1111.600 2051.945 1111.770 ;
        RECT 2052.115 1111.600 2052.405 1111.770 ;
        RECT 2052.575 1111.600 2052.865 1111.770 ;
        RECT 2053.035 1111.600 2053.325 1111.770 ;
        RECT 2053.495 1111.600 2053.785 1111.770 ;
        RECT 2053.955 1111.600 2054.245 1111.770 ;
        RECT 2054.415 1111.600 2054.705 1111.770 ;
        RECT 2054.875 1111.600 2055.165 1111.770 ;
        RECT 2055.335 1111.600 2055.625 1111.770 ;
        RECT 2055.795 1111.600 2056.085 1111.770 ;
        RECT 2056.255 1111.600 2056.545 1111.770 ;
        RECT 2056.715 1111.600 2057.005 1111.770 ;
        RECT 2057.175 1111.600 2057.465 1111.770 ;
        RECT 2057.635 1111.600 2057.925 1111.770 ;
        RECT 2058.095 1111.600 2058.385 1111.770 ;
        RECT 2058.555 1111.600 2058.845 1111.770 ;
        RECT 2059.015 1111.600 2059.305 1111.770 ;
        RECT 2059.475 1111.600 2059.765 1111.770 ;
        RECT 2059.935 1111.600 2060.225 1111.770 ;
        RECT 2060.395 1111.600 2060.685 1111.770 ;
        RECT 2060.855 1111.600 2061.145 1111.770 ;
        RECT 2061.315 1111.600 2061.605 1111.770 ;
        RECT 2061.775 1111.600 2062.065 1111.770 ;
        RECT 2062.235 1111.600 2062.525 1111.770 ;
        RECT 2062.695 1111.600 2062.985 1111.770 ;
        RECT 2063.155 1111.600 2063.445 1111.770 ;
        RECT 2063.615 1111.600 2063.905 1111.770 ;
        RECT 2064.075 1111.600 2064.365 1111.770 ;
        RECT 2064.535 1111.600 2064.825 1111.770 ;
        RECT 2064.995 1111.600 2065.285 1111.770 ;
        RECT 2065.455 1111.600 2065.745 1111.770 ;
        RECT 2065.915 1111.600 2066.205 1111.770 ;
        RECT 2066.375 1111.600 2066.665 1111.770 ;
        RECT 2066.835 1111.600 2067.125 1111.770 ;
        RECT 2067.295 1111.600 2067.585 1111.770 ;
        RECT 2067.755 1111.600 2068.045 1111.770 ;
        RECT 2068.215 1111.600 2068.505 1111.770 ;
        RECT 2068.675 1111.600 2068.965 1111.770 ;
        RECT 2069.135 1111.600 2069.425 1111.770 ;
        RECT 2069.595 1111.600 2069.885 1111.770 ;
        RECT 2070.055 1111.600 2070.345 1111.770 ;
        RECT 2070.515 1111.600 2070.805 1111.770 ;
        RECT 2070.975 1111.600 2071.265 1111.770 ;
        RECT 2071.435 1111.600 2071.725 1111.770 ;
        RECT 2071.895 1111.600 2072.185 1111.770 ;
        RECT 2072.355 1111.600 2072.645 1111.770 ;
        RECT 2072.815 1111.600 2073.105 1111.770 ;
        RECT 2073.275 1111.600 2073.565 1111.770 ;
        RECT 2073.735 1111.600 2074.025 1111.770 ;
        RECT 2074.195 1111.600 2074.485 1111.770 ;
        RECT 2074.655 1111.600 2074.945 1111.770 ;
        RECT 2075.115 1111.600 2075.405 1111.770 ;
        RECT 2075.575 1111.600 2075.865 1111.770 ;
        RECT 2076.035 1111.600 2076.325 1111.770 ;
        RECT 2076.495 1111.600 2076.785 1111.770 ;
        RECT 2076.955 1111.600 2077.245 1111.770 ;
        RECT 2077.415 1111.600 2077.705 1111.770 ;
        RECT 2077.875 1111.600 2078.165 1111.770 ;
        RECT 2078.335 1111.600 2078.625 1111.770 ;
        RECT 2078.795 1111.600 2079.085 1111.770 ;
        RECT 2079.255 1111.600 2079.545 1111.770 ;
        RECT 2079.715 1111.600 2080.005 1111.770 ;
        RECT 2080.175 1111.600 2080.465 1111.770 ;
        RECT 2080.635 1111.600 2080.925 1111.770 ;
        RECT 2081.095 1111.600 2081.385 1111.770 ;
        RECT 2081.555 1111.600 2081.845 1111.770 ;
        RECT 2082.015 1111.600 2082.305 1111.770 ;
        RECT 2082.475 1111.600 2082.765 1111.770 ;
        RECT 2082.935 1111.600 2083.225 1111.770 ;
        RECT 2083.395 1111.600 2083.685 1111.770 ;
        RECT 2083.855 1111.600 2084.145 1111.770 ;
        RECT 2084.315 1111.600 2084.605 1111.770 ;
        RECT 2084.775 1111.600 2085.065 1111.770 ;
        RECT 2085.235 1111.600 2085.525 1111.770 ;
        RECT 2085.695 1111.600 2085.985 1111.770 ;
        RECT 2086.155 1111.600 2086.445 1111.770 ;
        RECT 2086.615 1111.600 2086.905 1111.770 ;
        RECT 2087.075 1111.600 2087.365 1111.770 ;
        RECT 2087.535 1111.600 2087.825 1111.770 ;
        RECT 2087.995 1111.600 2088.285 1111.770 ;
        RECT 2088.455 1111.600 2088.745 1111.770 ;
        RECT 2088.915 1111.600 2089.205 1111.770 ;
        RECT 2089.375 1111.600 2089.665 1111.770 ;
        RECT 2089.835 1111.600 2090.125 1111.770 ;
        RECT 2090.295 1111.600 2090.585 1111.770 ;
        RECT 2090.755 1111.600 2091.045 1111.770 ;
        RECT 2091.215 1111.600 2091.505 1111.770 ;
        RECT 2091.675 1111.600 2091.965 1111.770 ;
        RECT 2092.135 1111.600 2092.425 1111.770 ;
        RECT 2092.595 1111.600 2092.885 1111.770 ;
        RECT 2093.055 1111.600 2093.345 1111.770 ;
        RECT 2093.515 1111.600 2093.805 1111.770 ;
        RECT 2093.975 1111.600 2094.265 1111.770 ;
        RECT 2094.435 1111.600 2094.725 1111.770 ;
        RECT 2094.895 1111.600 2095.040 1111.770 ;
      LAYER mcon ;
        RECT 835.260 4984.800 836.350 4984.970 ;
        RECT 841.240 4984.800 842.330 4984.970 ;
        RECT 847.220 4984.800 848.310 4984.970 ;
        RECT 836.170 4981.400 836.340 4982.250 ;
        RECT 842.150 4981.400 842.320 4982.250 ;
        RECT 848.130 4981.400 848.300 4982.250 ;
        RECT 2087.580 4983.025 2087.750 4983.875 ;
        RECT 3314.355 4985.675 3314.525 4986.525 ;
        RECT 3312.945 4982.955 3314.035 4983.125 ;
        RECT 3317.585 4982.615 3317.755 4983.465 ;
        RECT 3323.565 4982.615 3323.735 4983.465 ;
        RECT 3329.545 4982.615 3329.715 4983.465 ;
        RECT 3335.525 4982.615 3335.695 4983.465 ;
        RECT 199.410 4455.510 200.260 4455.680 ;
        RECT 202.810 4456.000 202.980 4457.090 ;
        RECT 199.750 4451.370 199.920 4452.460 ;
        RECT 202.470 4452.280 203.320 4452.450 ;
        RECT 199.410 4449.530 200.260 4449.700 ;
        RECT 202.810 4450.020 202.980 4451.110 ;
        RECT 199.750 4445.390 199.920 4446.480 ;
        RECT 202.470 4446.300 203.320 4446.470 ;
        RECT 199.410 4443.550 200.260 4443.720 ;
        RECT 202.810 4444.040 202.980 4445.130 ;
        RECT 199.750 4439.410 199.920 4440.500 ;
        RECT 202.470 4440.320 203.320 4440.490 ;
        RECT 199.750 4433.430 199.920 4434.520 ;
        RECT 202.470 4434.340 203.320 4434.510 ;
        RECT 199.750 4427.450 199.920 4428.540 ;
        RECT 202.470 4428.360 203.320 4428.530 ;
        RECT 3384.690 3571.200 3384.860 3572.290 ;
        RECT 3384.350 3567.480 3385.200 3567.650 ;
        RECT 3387.750 3566.570 3387.920 3567.660 ;
        RECT 3384.690 3565.220 3384.860 3566.310 ;
        RECT 3384.350 3561.500 3385.200 3561.670 ;
        RECT 3387.750 3560.590 3387.920 3561.680 ;
        RECT 3384.690 3559.240 3384.860 3560.330 ;
        RECT 3384.350 3555.520 3385.200 3555.690 ;
        RECT 3387.750 3554.610 3387.920 3555.700 ;
        RECT 3384.690 3553.260 3384.860 3554.350 ;
        RECT 3384.350 3549.540 3385.200 3549.710 ;
        RECT 3387.750 3548.630 3387.920 3549.720 ;
        RECT 3384.350 3543.560 3385.200 3543.730 ;
        RECT 3387.750 3542.650 3387.920 3543.740 ;
        RECT 3384.350 3537.580 3385.200 3537.750 ;
        RECT 3387.750 3536.670 3387.920 3537.760 ;
        RECT 199.535 3052.280 200.385 3052.450 ;
        RECT 202.935 3052.770 203.105 3053.860 ;
        RECT 199.875 3048.140 200.045 3049.230 ;
        RECT 202.595 3049.050 203.445 3049.220 ;
        RECT 199.535 3046.300 200.385 3046.470 ;
        RECT 202.935 3046.790 203.105 3047.880 ;
        RECT 199.875 3042.160 200.045 3043.250 ;
        RECT 202.595 3043.070 203.445 3043.240 ;
        RECT 199.535 3040.320 200.385 3040.490 ;
        RECT 202.935 3040.810 203.105 3041.900 ;
        RECT 199.875 3036.180 200.045 3037.270 ;
        RECT 202.595 3037.090 203.445 3037.260 ;
        RECT 199.535 3034.340 200.385 3034.510 ;
        RECT 202.935 3034.830 203.105 3035.920 ;
        RECT 199.875 3030.200 200.045 3031.290 ;
        RECT 202.595 3031.110 203.445 3031.280 ;
        RECT 199.535 3028.360 200.385 3028.530 ;
        RECT 202.935 3028.850 203.105 3029.940 ;
        RECT 199.875 3024.220 200.045 3025.310 ;
        RECT 202.595 3025.130 203.445 3025.300 ;
        RECT 199.875 3018.240 200.045 3019.330 ;
        RECT 202.595 3019.150 203.445 3019.320 ;
        RECT 199.875 3012.260 200.045 3013.350 ;
        RECT 202.595 3013.170 203.445 3013.340 ;
        RECT 199.875 3006.280 200.045 3007.370 ;
        RECT 202.595 3007.190 203.445 3007.360 ;
        RECT 199.875 3000.300 200.045 3001.390 ;
        RECT 202.595 3001.210 203.445 3001.380 ;
        RECT 199.875 2994.320 200.045 2995.410 ;
        RECT 202.595 2995.230 203.445 2995.400 ;
        RECT 199.875 2988.340 200.045 2989.430 ;
        RECT 202.595 2989.250 203.445 2989.420 ;
        RECT 3384.690 2267.080 3384.860 2268.170 ;
        RECT 3384.690 2261.100 3384.860 2262.190 ;
        RECT 3384.690 2255.120 3384.860 2256.210 ;
        RECT 3384.690 2249.140 3384.860 2250.230 ;
        RECT 3384.690 2243.160 3384.860 2244.250 ;
        RECT 3384.690 2237.180 3384.860 2238.270 ;
        RECT 199.645 1761.375 200.495 1761.545 ;
        RECT 203.045 1761.865 203.215 1762.955 ;
        RECT 199.985 1757.235 200.155 1758.325 ;
        RECT 202.705 1758.145 203.555 1758.315 ;
        RECT 199.645 1755.395 200.495 1755.565 ;
        RECT 203.045 1755.885 203.215 1756.975 ;
        RECT 199.985 1751.255 200.155 1752.345 ;
        RECT 202.705 1752.165 203.555 1752.335 ;
        RECT 199.645 1749.415 200.495 1749.585 ;
        RECT 203.045 1749.905 203.215 1750.995 ;
        RECT 199.985 1745.275 200.155 1746.365 ;
        RECT 202.705 1746.185 203.555 1746.355 ;
        RECT 199.645 1743.435 200.495 1743.605 ;
        RECT 203.045 1743.925 203.215 1745.015 ;
        RECT 199.985 1739.295 200.155 1740.385 ;
        RECT 202.705 1740.205 203.555 1740.375 ;
        RECT 199.645 1737.455 200.495 1737.625 ;
        RECT 203.045 1737.945 203.215 1739.035 ;
        RECT 199.985 1733.315 200.155 1734.405 ;
        RECT 202.705 1734.225 203.555 1734.395 ;
        RECT 199.645 1731.475 200.495 1731.645 ;
        RECT 203.045 1731.965 203.215 1733.055 ;
        RECT 199.985 1727.335 200.155 1728.425 ;
        RECT 202.705 1728.245 203.555 1728.415 ;
        RECT 199.645 1725.495 200.495 1725.665 ;
        RECT 203.045 1725.985 203.215 1727.075 ;
        RECT 199.985 1721.355 200.155 1722.445 ;
        RECT 202.705 1722.265 203.555 1722.435 ;
        RECT 199.645 1719.515 200.495 1719.685 ;
        RECT 203.045 1720.005 203.215 1721.095 ;
        RECT 199.985 1715.375 200.155 1716.465 ;
        RECT 202.705 1716.285 203.555 1716.455 ;
        RECT 199.645 1713.535 200.495 1713.705 ;
        RECT 203.045 1714.025 203.215 1715.115 ;
        RECT 199.985 1709.395 200.155 1710.485 ;
        RECT 202.705 1710.305 203.555 1710.475 ;
        RECT 199.645 1707.555 200.495 1707.725 ;
        RECT 203.045 1708.045 203.215 1709.135 ;
        RECT 199.985 1703.415 200.155 1704.505 ;
        RECT 202.705 1704.325 203.555 1704.495 ;
        RECT 199.645 1701.575 200.495 1701.745 ;
        RECT 203.045 1702.065 203.215 1703.155 ;
        RECT 199.985 1697.435 200.155 1698.525 ;
        RECT 202.705 1698.345 203.555 1698.515 ;
        RECT 199.985 1691.455 200.155 1692.545 ;
        RECT 202.705 1692.365 203.555 1692.535 ;
        RECT 199.985 1685.475 200.155 1686.565 ;
        RECT 202.705 1686.385 203.555 1686.555 ;
        RECT 199.985 1679.495 200.155 1680.585 ;
        RECT 202.705 1680.405 203.555 1680.575 ;
        RECT 199.985 1673.515 200.155 1674.605 ;
        RECT 202.705 1674.425 203.555 1674.595 ;
        RECT 670.520 1115.510 670.690 1116.360 ;
        RECT 674.240 1115.850 675.330 1116.020 ;
        RECT 676.500 1115.510 676.670 1116.360 ;
        RECT 680.220 1115.850 681.310 1116.020 ;
        RECT 682.480 1115.510 682.650 1116.360 ;
        RECT 686.200 1115.850 687.290 1116.020 ;
        RECT 688.460 1115.510 688.630 1116.360 ;
        RECT 692.180 1115.850 693.270 1116.020 ;
        RECT 694.440 1115.510 694.610 1116.360 ;
        RECT 698.160 1115.850 699.250 1116.020 ;
        RECT 700.420 1115.510 700.590 1116.360 ;
        RECT 704.140 1115.850 705.230 1116.020 ;
        RECT 706.400 1115.510 706.570 1116.360 ;
        RECT 710.120 1115.850 711.210 1116.020 ;
        RECT 712.380 1115.510 712.550 1116.360 ;
        RECT 716.100 1115.850 717.190 1116.020 ;
        RECT 718.360 1115.510 718.530 1116.360 ;
        RECT 722.080 1115.850 723.170 1116.020 ;
        RECT 724.340 1115.510 724.510 1116.360 ;
        RECT 728.060 1115.850 729.150 1116.020 ;
        RECT 730.320 1115.510 730.490 1116.360 ;
        RECT 734.040 1115.850 735.130 1116.020 ;
        RECT 736.300 1115.510 736.470 1116.360 ;
        RECT 740.020 1115.850 741.110 1116.020 ;
        RECT 742.280 1115.510 742.450 1116.360 ;
        RECT 746.000 1115.850 747.090 1116.020 ;
        RECT 748.260 1115.510 748.430 1116.360 ;
        RECT 751.980 1115.850 753.070 1116.020 ;
        RECT 754.240 1115.510 754.410 1116.360 ;
        RECT 757.960 1115.850 759.050 1116.020 ;
        RECT 763.940 1115.850 765.030 1116.020 ;
        RECT 769.920 1115.850 771.010 1116.020 ;
        RECT 775.900 1115.850 776.990 1116.020 ;
        RECT 781.880 1115.850 782.970 1116.020 ;
        RECT 787.860 1115.850 788.950 1116.020 ;
        RECT 793.840 1115.850 794.930 1116.020 ;
        RECT 1970.520 1115.510 1970.690 1116.360 ;
        RECT 1976.500 1115.510 1976.670 1116.360 ;
        RECT 1982.480 1115.510 1982.650 1116.360 ;
        RECT 1988.460 1115.510 1988.630 1116.360 ;
        RECT 1994.440 1115.510 1994.610 1116.360 ;
        RECT 2000.420 1115.510 2000.590 1116.360 ;
        RECT 2006.400 1115.510 2006.570 1116.360 ;
        RECT 2012.380 1115.510 2012.550 1116.360 ;
        RECT 2018.360 1115.510 2018.530 1116.360 ;
        RECT 2024.340 1115.510 2024.510 1116.360 ;
        RECT 2030.320 1115.510 2030.490 1116.360 ;
        RECT 2036.300 1115.510 2036.470 1116.360 ;
        RECT 2042.280 1115.510 2042.450 1116.360 ;
        RECT 2048.260 1115.510 2048.430 1116.360 ;
        RECT 2054.240 1115.510 2054.410 1116.360 ;
        RECT 2060.220 1115.510 2060.390 1116.360 ;
        RECT 2066.200 1115.510 2066.370 1116.360 ;
        RECT 2072.180 1115.510 2072.350 1116.360 ;
        RECT 2078.160 1115.510 2078.330 1116.360 ;
        RECT 2084.140 1115.510 2084.310 1116.360 ;
        RECT 2090.120 1115.510 2090.290 1116.360 ;
        RECT 675.590 1112.790 676.680 1112.960 ;
        RECT 679.730 1112.450 679.900 1113.300 ;
        RECT 681.570 1112.790 682.660 1112.960 ;
        RECT 685.710 1112.450 685.880 1113.300 ;
        RECT 687.550 1112.790 688.640 1112.960 ;
        RECT 691.690 1112.450 691.860 1113.300 ;
        RECT 693.530 1112.790 694.620 1112.960 ;
        RECT 697.670 1112.450 697.840 1113.300 ;
        RECT 699.510 1112.790 700.600 1112.960 ;
        RECT 703.650 1112.450 703.820 1113.300 ;
        RECT 705.490 1112.790 706.580 1112.960 ;
        RECT 709.630 1112.450 709.800 1113.300 ;
        RECT 711.470 1112.790 712.560 1112.960 ;
        RECT 715.610 1112.450 715.780 1113.300 ;
        RECT 717.450 1112.790 718.540 1112.960 ;
        RECT 721.590 1112.450 721.760 1113.300 ;
        RECT 723.430 1112.790 724.520 1112.960 ;
        RECT 727.570 1112.450 727.740 1113.300 ;
        RECT 729.410 1112.790 730.500 1112.960 ;
        RECT 733.550 1112.450 733.720 1113.300 ;
        RECT 735.390 1112.790 736.480 1112.960 ;
        RECT 739.530 1112.450 739.700 1113.300 ;
        RECT 741.370 1112.790 742.460 1112.960 ;
        RECT 745.510 1112.450 745.680 1113.300 ;
        RECT 747.350 1112.790 748.440 1112.960 ;
        RECT 751.490 1112.450 751.660 1113.300 ;
        RECT 753.330 1112.790 754.420 1112.960 ;
        RECT 757.470 1112.450 757.640 1113.300 ;
        RECT 759.310 1112.790 760.400 1112.960 ;
        RECT 763.450 1112.450 763.620 1113.300 ;
        RECT 769.430 1112.450 769.600 1113.300 ;
        RECT 775.410 1112.450 775.580 1113.300 ;
        RECT 781.390 1112.450 781.560 1113.300 ;
        RECT 787.370 1112.450 787.540 1113.300 ;
        RECT 793.340 1112.790 794.430 1112.960 ;
        RECT 1975.590 1112.790 1976.680 1112.960 ;
        RECT 1981.570 1112.790 1982.660 1112.960 ;
        RECT 1987.550 1112.790 1988.640 1112.960 ;
        RECT 1993.530 1112.790 1994.620 1112.960 ;
        RECT 1999.510 1112.790 2000.600 1112.960 ;
        RECT 2005.490 1112.790 2006.580 1112.960 ;
        RECT 2011.470 1112.790 2012.560 1112.960 ;
        RECT 2017.450 1112.790 2018.540 1112.960 ;
        RECT 2023.430 1112.790 2024.520 1112.960 ;
        RECT 2029.410 1112.790 2030.500 1112.960 ;
        RECT 2035.390 1112.790 2036.480 1112.960 ;
        RECT 2041.370 1112.790 2042.460 1112.960 ;
        RECT 2047.350 1112.790 2048.440 1112.960 ;
        RECT 2053.330 1112.790 2054.420 1112.960 ;
        RECT 2059.310 1112.790 2060.400 1112.960 ;
        RECT 2065.290 1112.790 2066.380 1112.960 ;
        RECT 2071.270 1112.790 2072.360 1112.960 ;
        RECT 2077.250 1112.790 2078.340 1112.960 ;
        RECT 2083.230 1112.790 2084.320 1112.960 ;
        RECT 2090.120 1112.450 2090.290 1113.300 ;
      LAYER met1 ;
        RECT 2087.510 4986.375 2088.720 4986.635 ;
        RECT 3314.315 4985.615 3314.575 4986.585 ;
        RECT 3317.515 4985.965 3318.725 4986.225 ;
        RECT 3323.495 4985.965 3324.705 4986.225 ;
        RECT 3329.475 4985.965 3330.685 4986.225 ;
        RECT 3335.455 4985.965 3336.665 4986.225 ;
        RECT 835.200 4984.750 836.410 4985.010 ;
        RECT 841.180 4984.750 842.390 4985.010 ;
        RECT 847.160 4984.750 848.370 4985.010 ;
        RECT 2087.540 4982.965 2087.800 4983.935 ;
        RECT 3312.885 4982.905 3314.095 4983.165 ;
        RECT 3317.545 4982.555 3317.805 4983.525 ;
        RECT 3323.525 4982.555 3323.785 4983.525 ;
        RECT 3329.505 4982.555 3329.765 4983.525 ;
        RECT 3335.485 4982.555 3335.745 4983.525 ;
        RECT 836.120 4981.340 836.380 4982.310 ;
        RECT 842.100 4981.340 842.360 4982.310 ;
        RECT 848.080 4981.340 848.340 4982.310 ;
        RECT 212.455 4977.145 848.420 4977.285 ;
        RECT 202.770 4455.940 203.030 4457.150 ;
        RECT 212.455 4456.785 212.595 4977.145 ;
        RECT 848.100 4977.025 848.420 4977.145 ;
        RECT 212.335 4456.465 212.595 4456.785 ;
        RECT 212.735 4976.865 847.800 4977.005 ;
        RECT 212.735 4455.815 212.875 4976.865 ;
        RECT 847.480 4976.745 847.800 4976.865 ;
        RECT 199.350 4455.460 200.320 4455.720 ;
        RECT 212.615 4455.495 212.875 4455.815 ;
        RECT 213.015 4976.585 842.440 4976.725 ;
        RECT 199.710 4451.310 199.970 4452.520 ;
        RECT 202.410 4452.230 203.380 4452.490 ;
        RECT 212.315 4452.250 212.575 4452.570 ;
        RECT 202.770 4449.960 203.030 4451.170 ;
        RECT 199.350 4449.480 200.320 4449.740 ;
        RECT 199.710 4445.330 199.970 4446.540 ;
        RECT 202.410 4446.250 203.380 4446.510 ;
        RECT 202.770 4443.980 203.030 4445.190 ;
        RECT 199.350 4443.500 200.320 4443.760 ;
        RECT 199.710 4439.350 199.970 4440.560 ;
        RECT 202.410 4440.270 203.380 4440.530 ;
        RECT 199.710 4433.370 199.970 4434.580 ;
        RECT 202.410 4434.290 203.380 4434.550 ;
        RECT 199.710 4427.390 199.970 4428.600 ;
        RECT 202.410 4428.310 203.380 4428.570 ;
        RECT 202.895 3052.710 203.155 3053.920 ;
        RECT 212.315 3053.555 212.455 4452.250 ;
        RECT 212.195 3053.235 212.455 3053.555 ;
        RECT 212.595 4451.630 212.855 4451.950 ;
        RECT 212.595 3052.585 212.735 4451.630 ;
        RECT 213.015 4450.685 213.155 4976.585 ;
        RECT 842.120 4976.465 842.440 4976.585 ;
        RECT 212.895 4450.365 213.155 4450.685 ;
        RECT 213.295 4976.305 841.820 4976.445 ;
        RECT 213.295 4449.835 213.435 4976.305 ;
        RECT 841.500 4976.185 841.820 4976.305 ;
        RECT 2087.460 4976.235 3309.400 4976.375 ;
        RECT 3313.250 4976.235 3313.570 4976.355 ;
        RECT 213.175 4449.515 213.435 4449.835 ;
        RECT 213.575 4976.025 836.460 4976.165 ;
        RECT 2087.460 4976.115 2087.780 4976.235 ;
        RECT 3309.210 4976.095 3313.570 4976.235 ;
        RECT 3317.465 4976.235 3375.740 4976.375 ;
        RECT 3317.465 4976.115 3317.785 4976.235 ;
        RECT 199.475 3052.230 200.445 3052.490 ;
        RECT 212.475 3052.265 212.735 3052.585 ;
        RECT 212.875 4446.270 213.135 4446.590 ;
        RECT 199.835 3048.080 200.095 3049.290 ;
        RECT 202.535 3049.000 203.505 3049.260 ;
        RECT 212.175 3049.020 212.435 3049.340 ;
        RECT 202.895 3046.730 203.155 3047.940 ;
        RECT 199.475 3046.250 200.445 3046.510 ;
        RECT 199.835 3042.100 200.095 3043.310 ;
        RECT 202.535 3043.020 203.505 3043.280 ;
        RECT 202.895 3040.750 203.155 3041.960 ;
        RECT 199.475 3040.270 200.445 3040.530 ;
        RECT 199.835 3036.120 200.095 3037.330 ;
        RECT 202.535 3037.040 203.505 3037.300 ;
        RECT 202.895 3034.770 203.155 3035.980 ;
        RECT 199.475 3034.290 200.445 3034.550 ;
        RECT 199.835 3030.140 200.095 3031.350 ;
        RECT 202.535 3031.060 203.505 3031.320 ;
        RECT 202.895 3028.790 203.155 3030.000 ;
        RECT 199.475 3028.310 200.445 3028.570 ;
        RECT 199.835 3024.160 200.095 3025.370 ;
        RECT 202.535 3025.080 203.505 3025.340 ;
        RECT 199.835 3018.180 200.095 3019.390 ;
        RECT 202.535 3019.100 203.505 3019.360 ;
        RECT 199.835 3012.200 200.095 3013.410 ;
        RECT 202.535 3013.120 203.505 3013.380 ;
        RECT 199.835 3006.220 200.095 3007.430 ;
        RECT 202.535 3007.140 203.505 3007.400 ;
        RECT 199.835 3000.240 200.095 3001.450 ;
        RECT 202.535 3001.160 203.505 3001.420 ;
        RECT 199.835 2994.260 200.095 2995.470 ;
        RECT 202.535 2995.180 203.505 2995.440 ;
        RECT 199.835 2988.280 200.095 2989.490 ;
        RECT 202.535 2989.200 203.505 2989.460 ;
        RECT 203.005 1761.805 203.265 1763.015 ;
        RECT 212.175 1762.650 212.315 3049.020 ;
        RECT 212.055 1762.330 212.315 1762.650 ;
        RECT 212.455 3048.400 212.715 3048.720 ;
        RECT 212.455 1761.680 212.595 3048.400 ;
        RECT 212.875 3047.455 213.015 4446.270 ;
        RECT 212.755 3047.135 213.015 3047.455 ;
        RECT 213.155 4445.650 213.415 4445.970 ;
        RECT 213.155 3046.605 213.295 4445.650 ;
        RECT 213.575 4444.825 213.715 4976.025 ;
        RECT 836.140 4975.905 836.460 4976.025 ;
        RECT 2088.055 4975.955 3308.810 4976.095 ;
        RECT 3314.220 4975.955 3314.540 4976.075 ;
        RECT 213.455 4444.505 213.715 4444.825 ;
        RECT 213.855 4975.745 835.840 4975.885 ;
        RECT 2088.080 4975.835 2088.400 4975.955 ;
        RECT 3308.625 4975.815 3314.540 4975.955 ;
        RECT 3318.085 4975.955 3375.460 4976.095 ;
        RECT 3318.085 4975.835 3318.405 4975.955 ;
        RECT 213.855 4443.855 213.995 4975.745 ;
        RECT 835.520 4975.625 835.840 4975.745 ;
        RECT 3323.445 4975.675 3375.180 4975.815 ;
        RECT 3323.445 4975.555 3323.765 4975.675 ;
        RECT 3324.065 4975.395 3374.900 4975.535 ;
        RECT 3324.065 4975.275 3324.385 4975.395 ;
        RECT 3329.425 4975.115 3374.620 4975.255 ;
        RECT 3329.425 4974.995 3329.745 4975.115 ;
        RECT 3330.045 4974.835 3374.340 4974.975 ;
        RECT 3330.045 4974.715 3330.365 4974.835 ;
        RECT 3335.405 4974.555 3374.060 4974.695 ;
        RECT 3335.405 4974.435 3335.725 4974.555 ;
        RECT 3336.000 4974.275 3373.780 4974.415 ;
        RECT 3336.025 4974.155 3336.345 4974.275 ;
        RECT 213.735 4443.535 213.995 4443.855 ;
        RECT 213.035 3046.285 213.295 3046.605 ;
        RECT 213.435 4440.290 213.695 4440.610 ;
        RECT 199.585 1761.325 200.555 1761.585 ;
        RECT 212.335 1761.360 212.595 1761.680 ;
        RECT 212.735 3043.040 212.995 3043.360 ;
        RECT 199.945 1757.175 200.205 1758.385 ;
        RECT 202.645 1758.095 203.615 1758.355 ;
        RECT 212.035 1758.115 212.295 1758.435 ;
        RECT 203.005 1755.825 203.265 1757.035 ;
        RECT 199.585 1755.345 200.555 1755.605 ;
        RECT 199.945 1751.195 200.205 1752.405 ;
        RECT 202.645 1752.115 203.615 1752.375 ;
        RECT 203.005 1749.845 203.265 1751.055 ;
        RECT 199.585 1749.365 200.555 1749.625 ;
        RECT 199.945 1745.215 200.205 1746.425 ;
        RECT 202.645 1746.135 203.615 1746.395 ;
        RECT 203.005 1743.865 203.265 1745.075 ;
        RECT 199.585 1743.385 200.555 1743.645 ;
        RECT 199.945 1739.235 200.205 1740.445 ;
        RECT 202.645 1740.155 203.615 1740.415 ;
        RECT 203.005 1737.885 203.265 1739.095 ;
        RECT 199.585 1737.405 200.555 1737.665 ;
        RECT 199.945 1733.255 200.205 1734.465 ;
        RECT 202.645 1734.175 203.615 1734.435 ;
        RECT 203.005 1731.905 203.265 1733.115 ;
        RECT 199.585 1731.425 200.555 1731.685 ;
        RECT 199.945 1727.275 200.205 1728.485 ;
        RECT 202.645 1728.195 203.615 1728.455 ;
        RECT 203.005 1725.925 203.265 1727.135 ;
        RECT 199.585 1725.445 200.555 1725.705 ;
        RECT 199.945 1721.295 200.205 1722.505 ;
        RECT 202.645 1722.215 203.615 1722.475 ;
        RECT 203.005 1719.945 203.265 1721.155 ;
        RECT 199.585 1719.465 200.555 1719.725 ;
        RECT 199.945 1715.315 200.205 1716.525 ;
        RECT 202.645 1716.235 203.615 1716.495 ;
        RECT 203.005 1713.965 203.265 1715.175 ;
        RECT 199.585 1713.485 200.555 1713.745 ;
        RECT 199.945 1709.335 200.205 1710.545 ;
        RECT 202.645 1710.255 203.615 1710.515 ;
        RECT 203.005 1707.985 203.265 1709.195 ;
        RECT 199.585 1707.505 200.555 1707.765 ;
        RECT 199.945 1703.355 200.205 1704.565 ;
        RECT 202.645 1704.275 203.615 1704.535 ;
        RECT 203.005 1702.005 203.265 1703.215 ;
        RECT 199.585 1701.525 200.555 1701.785 ;
        RECT 199.945 1697.375 200.205 1698.585 ;
        RECT 202.645 1698.295 203.615 1698.555 ;
        RECT 199.945 1691.395 200.205 1692.605 ;
        RECT 202.645 1692.315 203.615 1692.575 ;
        RECT 199.945 1685.415 200.205 1686.625 ;
        RECT 202.645 1686.335 203.615 1686.595 ;
        RECT 199.945 1679.435 200.205 1680.645 ;
        RECT 202.645 1680.355 203.615 1680.615 ;
        RECT 199.945 1673.455 200.205 1674.665 ;
        RECT 202.645 1674.375 203.615 1674.635 ;
        RECT 212.035 1121.260 212.175 1758.115 ;
        RECT 212.315 1757.495 212.575 1757.815 ;
        RECT 212.315 1121.540 212.455 1757.495 ;
        RECT 212.735 1756.550 212.875 3043.040 ;
        RECT 212.615 1756.230 212.875 1756.550 ;
        RECT 213.015 3042.420 213.275 3042.740 ;
        RECT 213.015 1755.700 213.155 3042.420 ;
        RECT 213.435 3041.595 213.575 4440.290 ;
        RECT 213.315 3041.275 213.575 3041.595 ;
        RECT 213.715 4439.670 213.975 4439.990 ;
        RECT 213.715 3040.625 213.855 4439.670 ;
        RECT 213.595 3040.305 213.855 3040.625 ;
        RECT 213.995 4434.310 214.255 4434.630 ;
        RECT 212.895 1755.380 213.155 1755.700 ;
        RECT 213.295 3037.060 213.555 3037.380 ;
        RECT 212.595 1752.135 212.855 1752.455 ;
        RECT 212.595 1121.820 212.735 1752.135 ;
        RECT 212.875 1751.515 213.135 1751.835 ;
        RECT 212.875 1122.100 213.015 1751.515 ;
        RECT 213.295 1750.690 213.435 3037.060 ;
        RECT 213.175 1750.370 213.435 1750.690 ;
        RECT 213.575 3036.440 213.835 3036.760 ;
        RECT 213.575 1749.720 213.715 3036.440 ;
        RECT 213.995 3035.495 214.135 4434.310 ;
        RECT 213.875 3035.175 214.135 3035.495 ;
        RECT 214.275 4433.690 214.535 4434.010 ;
        RECT 214.275 3034.645 214.415 4433.690 ;
        RECT 214.155 3034.325 214.415 3034.645 ;
        RECT 214.555 4428.330 214.815 4428.650 ;
        RECT 213.455 1749.400 213.715 1749.720 ;
        RECT 213.855 3031.080 214.115 3031.400 ;
        RECT 213.155 1746.155 213.415 1746.475 ;
        RECT 213.155 1122.380 213.295 1746.155 ;
        RECT 213.435 1745.535 213.695 1745.855 ;
        RECT 213.435 1122.660 213.575 1745.535 ;
        RECT 213.855 1744.590 213.995 3031.080 ;
        RECT 213.735 1744.270 213.995 1744.590 ;
        RECT 214.135 3030.460 214.395 3030.780 ;
        RECT 214.135 1743.740 214.275 3030.460 ;
        RECT 214.555 3029.635 214.695 4428.330 ;
        RECT 214.435 3029.315 214.695 3029.635 ;
        RECT 214.835 4427.710 215.095 4428.030 ;
        RECT 214.835 3028.665 214.975 4427.710 ;
        RECT 3373.640 3579.995 3373.780 4974.275 ;
        RECT 3373.500 3579.815 3373.780 3579.995 ;
        RECT 3373.500 3553.075 3373.640 3579.815 ;
        RECT 3373.920 3579.360 3374.060 4974.555 ;
        RECT 3373.780 3579.180 3374.060 3579.360 ;
        RECT 3373.780 3554.045 3373.920 3579.180 ;
        RECT 3374.200 3578.690 3374.340 4974.835 ;
        RECT 3374.060 3578.515 3374.340 3578.690 ;
        RECT 3374.060 3559.055 3374.200 3578.515 ;
        RECT 3374.480 3577.990 3374.620 4975.115 ;
        RECT 3374.340 3577.810 3374.620 3577.990 ;
        RECT 3374.340 3560.025 3374.480 3577.810 ;
        RECT 3374.760 3577.305 3374.900 4975.395 ;
        RECT 3374.620 3577.125 3374.900 3577.305 ;
        RECT 3374.620 3565.035 3374.760 3577.125 ;
        RECT 3375.040 3576.575 3375.180 4975.675 ;
        RECT 3374.900 3576.390 3375.180 3576.575 ;
        RECT 3374.900 3566.005 3375.040 3576.390 ;
        RECT 3375.320 3575.930 3375.460 4975.955 ;
        RECT 3375.180 3575.755 3375.460 3575.930 ;
        RECT 3375.180 3571.015 3375.320 3575.755 ;
        RECT 3375.600 3575.385 3375.740 4976.235 ;
        RECT 3375.460 3575.210 3375.740 3575.385 ;
        RECT 3375.460 3571.865 3375.600 3575.210 ;
        RECT 3375.460 3571.545 3375.720 3571.865 ;
        RECT 3384.640 3571.140 3384.900 3572.350 ;
        RECT 3375.180 3570.695 3375.440 3571.015 ;
        RECT 3387.350 3570.660 3388.320 3570.920 ;
        RECT 3375.480 3567.450 3375.740 3567.770 ;
        RECT 3375.200 3566.830 3375.460 3567.150 ;
        RECT 3374.900 3565.685 3375.160 3566.005 ;
        RECT 3374.620 3564.715 3374.880 3565.035 ;
        RECT 3374.920 3561.470 3375.180 3561.790 ;
        RECT 3374.640 3560.850 3374.900 3561.170 ;
        RECT 3374.340 3559.705 3374.600 3560.025 ;
        RECT 3374.060 3558.735 3374.320 3559.055 ;
        RECT 3374.360 3555.490 3374.620 3555.810 ;
        RECT 3374.080 3554.870 3374.340 3555.190 ;
        RECT 3373.780 3553.725 3374.040 3554.045 ;
        RECT 3373.500 3552.755 3373.760 3553.075 ;
        RECT 3373.800 3549.510 3374.060 3549.830 ;
        RECT 3373.520 3548.890 3373.780 3549.210 ;
        RECT 3373.240 3543.530 3373.500 3543.850 ;
        RECT 3372.960 3542.910 3373.220 3543.230 ;
        RECT 3372.680 3537.550 3372.940 3537.870 ;
        RECT 3372.520 3537.250 3372.660 3537.275 ;
        RECT 3372.400 3536.930 3372.660 3537.250 ;
        RECT 214.715 3028.345 214.975 3028.665 ;
        RECT 214.015 1743.420 214.275 1743.740 ;
        RECT 214.415 3025.100 214.675 3025.420 ;
        RECT 213.715 1740.175 213.975 1740.495 ;
        RECT 213.715 1122.940 213.855 1740.175 ;
        RECT 213.995 1739.555 214.255 1739.875 ;
        RECT 213.995 1123.220 214.135 1739.555 ;
        RECT 214.415 1738.730 214.555 3025.100 ;
        RECT 214.295 1738.410 214.555 1738.730 ;
        RECT 214.695 3024.480 214.955 3024.800 ;
        RECT 214.695 1737.760 214.835 3024.480 ;
        RECT 214.575 1737.440 214.835 1737.760 ;
        RECT 214.975 3019.120 215.235 3019.440 ;
        RECT 214.275 1734.195 214.535 1734.515 ;
        RECT 214.275 1123.500 214.415 1734.195 ;
        RECT 214.555 1733.575 214.815 1733.895 ;
        RECT 214.555 1123.780 214.695 1733.575 ;
        RECT 214.975 1732.750 215.115 3019.120 ;
        RECT 214.855 1732.430 215.115 1732.750 ;
        RECT 215.255 3018.500 215.515 3018.820 ;
        RECT 215.255 1731.780 215.395 3018.500 ;
        RECT 215.135 1731.460 215.395 1731.780 ;
        RECT 215.535 3013.140 215.795 3013.460 ;
        RECT 214.835 1728.215 215.095 1728.535 ;
        RECT 214.835 1124.060 214.975 1728.215 ;
        RECT 215.115 1727.595 215.375 1727.915 ;
        RECT 215.115 1124.340 215.255 1727.595 ;
        RECT 215.535 1726.770 215.675 3013.140 ;
        RECT 215.415 1726.450 215.675 1726.770 ;
        RECT 215.815 3012.520 216.075 3012.840 ;
        RECT 215.815 1725.800 215.955 3012.520 ;
        RECT 215.695 1725.480 215.955 1725.800 ;
        RECT 216.095 3007.160 216.355 3007.480 ;
        RECT 215.395 1722.235 215.655 1722.555 ;
        RECT 215.395 1124.620 215.535 1722.235 ;
        RECT 215.675 1721.615 215.935 1721.935 ;
        RECT 215.675 1124.900 215.815 1721.615 ;
        RECT 216.095 1720.790 216.235 3007.160 ;
        RECT 215.975 1720.470 216.235 1720.790 ;
        RECT 216.375 3006.540 216.635 3006.860 ;
        RECT 216.375 1719.820 216.515 3006.540 ;
        RECT 216.255 1719.500 216.515 1719.820 ;
        RECT 216.655 3001.180 216.915 3001.500 ;
        RECT 215.955 1716.255 216.215 1716.575 ;
        RECT 215.955 1125.180 216.095 1716.255 ;
        RECT 216.235 1715.635 216.495 1715.955 ;
        RECT 216.235 1125.460 216.375 1715.635 ;
        RECT 216.655 1714.810 216.795 3001.180 ;
        RECT 216.535 1714.490 216.795 1714.810 ;
        RECT 216.935 3000.560 217.195 3000.880 ;
        RECT 216.935 1713.840 217.075 3000.560 ;
        RECT 216.815 1713.520 217.075 1713.840 ;
        RECT 217.215 2995.200 217.475 2995.520 ;
        RECT 216.515 1710.275 216.775 1710.595 ;
        RECT 216.515 1125.740 216.655 1710.275 ;
        RECT 216.795 1709.655 217.055 1709.975 ;
        RECT 216.795 1126.020 216.935 1709.655 ;
        RECT 217.215 1708.830 217.355 2995.200 ;
        RECT 217.095 1708.510 217.355 1708.830 ;
        RECT 217.495 2994.580 217.755 2994.900 ;
        RECT 217.495 1707.860 217.635 2994.580 ;
        RECT 217.375 1707.540 217.635 1707.860 ;
        RECT 217.775 2989.220 218.035 2989.540 ;
        RECT 217.075 1704.295 217.335 1704.615 ;
        RECT 217.075 1126.300 217.215 1704.295 ;
        RECT 217.355 1703.675 217.615 1703.995 ;
        RECT 217.355 1126.580 217.495 1703.675 ;
        RECT 217.775 1702.850 217.915 2989.220 ;
        RECT 217.655 1702.530 217.915 1702.850 ;
        RECT 218.055 2988.600 218.315 2988.920 ;
        RECT 218.055 1701.880 218.195 2988.600 ;
        RECT 3372.520 2275.540 3372.660 3536.930 ;
        RECT 3372.380 2275.395 3372.660 2275.540 ;
        RECT 3372.380 2236.995 3372.520 2275.395 ;
        RECT 3372.800 2275.250 3372.940 3537.550 ;
        RECT 3372.660 2275.100 3372.940 2275.250 ;
        RECT 3372.660 2237.965 3372.800 2275.100 ;
        RECT 3373.080 2274.955 3373.220 3542.910 ;
        RECT 3372.940 2274.815 3373.220 2274.955 ;
        RECT 3372.940 2242.975 3373.080 2274.815 ;
        RECT 3373.360 2274.655 3373.500 3543.530 ;
        RECT 3373.220 2274.490 3373.500 2274.655 ;
        RECT 3373.220 2243.945 3373.360 2274.490 ;
        RECT 3373.640 2274.330 3373.780 3548.890 ;
        RECT 3373.500 2274.180 3373.780 2274.330 ;
        RECT 3373.500 2248.955 3373.640 2274.180 ;
        RECT 3373.920 2274.025 3374.060 3549.510 ;
        RECT 3373.780 2273.845 3374.060 2274.025 ;
        RECT 3373.780 2249.805 3373.920 2273.845 ;
        RECT 3374.200 2273.665 3374.340 3554.870 ;
        RECT 3374.060 2273.495 3374.340 2273.665 ;
        RECT 3374.060 2254.935 3374.200 2273.495 ;
        RECT 3374.480 2273.330 3374.620 3555.490 ;
        RECT 3374.340 2273.175 3374.620 2273.330 ;
        RECT 3374.340 2255.905 3374.480 2273.175 ;
        RECT 3374.760 2273.030 3374.900 3560.850 ;
        RECT 3374.620 2272.865 3374.900 2273.030 ;
        RECT 3374.620 2260.915 3374.760 2272.865 ;
        RECT 3375.040 2272.720 3375.180 3561.470 ;
        RECT 3374.900 2272.505 3375.180 2272.720 ;
        RECT 3374.900 2261.765 3375.040 2272.505 ;
        RECT 3375.320 2272.360 3375.460 3566.830 ;
        RECT 3375.180 2272.160 3375.460 2272.360 ;
        RECT 3375.180 2266.895 3375.320 2272.160 ;
        RECT 3375.600 2272.015 3375.740 3567.450 ;
        RECT 3384.290 3567.430 3385.260 3567.690 ;
        RECT 3387.700 3566.510 3387.960 3567.720 ;
        RECT 3384.640 3565.160 3384.900 3566.370 ;
        RECT 3387.350 3564.680 3388.320 3564.940 ;
        RECT 3384.290 3561.450 3385.260 3561.710 ;
        RECT 3387.700 3560.530 3387.960 3561.740 ;
        RECT 3384.640 3559.180 3384.900 3560.390 ;
        RECT 3387.350 3558.700 3388.320 3558.960 ;
        RECT 3384.290 3555.470 3385.260 3555.730 ;
        RECT 3387.700 3554.550 3387.960 3555.760 ;
        RECT 3384.640 3553.200 3384.900 3554.410 ;
        RECT 3387.350 3552.720 3388.320 3552.980 ;
        RECT 3384.290 3549.490 3385.260 3549.750 ;
        RECT 3387.700 3548.570 3387.960 3549.780 ;
        RECT 3384.290 3543.510 3385.260 3543.770 ;
        RECT 3387.700 3542.590 3387.960 3543.800 ;
        RECT 3384.290 3537.530 3385.260 3537.790 ;
        RECT 3387.700 3536.610 3387.960 3537.820 ;
        RECT 3375.460 2271.825 3375.740 2272.015 ;
        RECT 3375.460 2267.865 3375.600 2271.825 ;
        RECT 3375.460 2267.545 3375.720 2267.865 ;
        RECT 3384.640 2267.020 3384.900 2268.230 ;
        RECT 3375.180 2266.575 3375.440 2266.895 ;
        RECT 3387.350 2266.540 3388.320 2266.800 ;
        RECT 3374.900 2261.445 3375.160 2261.765 ;
        RECT 3384.640 2261.040 3384.900 2262.250 ;
        RECT 3374.620 2260.595 3374.880 2260.915 ;
        RECT 3387.350 2260.560 3388.320 2260.820 ;
        RECT 3374.340 2255.585 3374.600 2255.905 ;
        RECT 3384.640 2255.060 3384.900 2256.270 ;
        RECT 3374.060 2254.615 3374.320 2254.935 ;
        RECT 3387.350 2254.580 3388.320 2254.840 ;
        RECT 3373.780 2249.485 3374.040 2249.805 ;
        RECT 3384.640 2249.080 3384.900 2250.290 ;
        RECT 3373.500 2248.635 3373.760 2248.955 ;
        RECT 3387.350 2248.600 3388.320 2248.860 ;
        RECT 3373.220 2243.625 3373.480 2243.945 ;
        RECT 3384.640 2243.100 3384.900 2244.310 ;
        RECT 3372.940 2242.655 3373.200 2242.975 ;
        RECT 3387.350 2242.620 3388.320 2242.880 ;
        RECT 3372.660 2237.645 3372.920 2237.965 ;
        RECT 3384.640 2237.120 3384.900 2238.330 ;
        RECT 3372.380 2236.675 3372.640 2236.995 ;
        RECT 3387.350 2236.640 3388.320 2236.900 ;
        RECT 217.935 1701.560 218.195 1701.880 ;
        RECT 217.635 1698.315 217.895 1698.635 ;
        RECT 217.635 1126.860 217.775 1698.315 ;
        RECT 217.915 1697.695 218.175 1698.015 ;
        RECT 217.915 1127.140 218.055 1697.695 ;
        RECT 218.195 1692.335 218.455 1692.655 ;
        RECT 218.195 1127.420 218.335 1692.335 ;
        RECT 218.475 1691.715 218.735 1692.035 ;
        RECT 218.475 1127.700 218.615 1691.715 ;
        RECT 218.755 1686.355 219.015 1686.675 ;
        RECT 218.755 1127.980 218.895 1686.355 ;
        RECT 219.035 1685.735 219.295 1686.055 ;
        RECT 219.035 1128.260 219.175 1685.735 ;
        RECT 219.315 1680.375 219.575 1680.695 ;
        RECT 219.315 1128.540 219.455 1680.375 ;
        RECT 219.595 1679.755 219.855 1680.075 ;
        RECT 219.595 1128.820 219.735 1679.755 ;
        RECT 219.875 1674.395 220.135 1674.715 ;
        RECT 219.875 1129.100 220.015 1674.395 ;
        RECT 220.155 1673.775 220.415 1674.095 ;
        RECT 220.155 1129.380 220.295 1673.775 ;
        RECT 1970.490 1129.520 1970.810 1129.640 ;
        RECT 670.490 1129.380 670.810 1129.500 ;
        RECT 220.155 1129.240 670.810 1129.380 ;
        RECT 674.705 1129.380 1970.810 1129.520 ;
        RECT 674.705 1129.260 675.025 1129.380 ;
        RECT 1975.850 1129.240 1976.170 1129.360 ;
        RECT 675.850 1129.100 676.170 1129.220 ;
        RECT 219.875 1128.960 676.170 1129.100 ;
        RECT 679.715 1129.100 1976.170 1129.240 ;
        RECT 679.715 1128.980 680.035 1129.100 ;
        RECT 1976.470 1128.960 1976.790 1129.080 ;
        RECT 676.470 1128.820 676.790 1128.940 ;
        RECT 219.595 1128.680 676.790 1128.820 ;
        RECT 680.685 1128.820 1976.790 1128.960 ;
        RECT 680.685 1128.700 681.005 1128.820 ;
        RECT 1981.830 1128.680 1982.150 1128.800 ;
        RECT 681.830 1128.540 682.150 1128.660 ;
        RECT 219.315 1128.400 682.150 1128.540 ;
        RECT 685.695 1128.540 1982.150 1128.680 ;
        RECT 685.695 1128.420 686.015 1128.540 ;
        RECT 1982.450 1128.400 1982.770 1128.520 ;
        RECT 682.450 1128.260 682.770 1128.380 ;
        RECT 219.035 1128.120 682.770 1128.260 ;
        RECT 686.665 1128.260 1982.770 1128.400 ;
        RECT 686.665 1128.140 686.985 1128.260 ;
        RECT 1987.810 1128.120 1988.130 1128.240 ;
        RECT 687.810 1127.980 688.130 1128.100 ;
        RECT 218.755 1127.840 688.130 1127.980 ;
        RECT 691.675 1127.980 1988.130 1128.120 ;
        RECT 691.675 1127.860 691.995 1127.980 ;
        RECT 1988.430 1127.840 1988.750 1127.960 ;
        RECT 688.430 1127.700 688.750 1127.820 ;
        RECT 218.475 1127.560 688.750 1127.700 ;
        RECT 692.645 1127.700 1988.750 1127.840 ;
        RECT 692.645 1127.580 692.965 1127.700 ;
        RECT 1993.790 1127.560 1994.110 1127.680 ;
        RECT 693.790 1127.420 694.110 1127.540 ;
        RECT 218.195 1127.280 694.110 1127.420 ;
        RECT 697.655 1127.420 1994.110 1127.560 ;
        RECT 697.655 1127.300 697.975 1127.420 ;
        RECT 1994.410 1127.280 1994.730 1127.400 ;
        RECT 694.410 1127.140 694.730 1127.260 ;
        RECT 217.915 1127.000 694.730 1127.140 ;
        RECT 698.625 1127.140 1994.730 1127.280 ;
        RECT 698.625 1127.020 698.945 1127.140 ;
        RECT 1999.770 1127.000 2000.090 1127.120 ;
        RECT 699.770 1126.860 700.090 1126.980 ;
        RECT 217.635 1126.720 700.090 1126.860 ;
        RECT 703.635 1126.860 2000.090 1127.000 ;
        RECT 703.635 1126.740 703.955 1126.860 ;
        RECT 2000.390 1126.720 2000.710 1126.840 ;
        RECT 700.390 1126.580 700.710 1126.700 ;
        RECT 217.355 1126.440 700.710 1126.580 ;
        RECT 704.485 1126.580 2000.710 1126.720 ;
        RECT 704.485 1126.460 704.805 1126.580 ;
        RECT 2005.750 1126.440 2006.070 1126.560 ;
        RECT 705.750 1126.300 706.070 1126.420 ;
        RECT 217.075 1126.160 706.070 1126.300 ;
        RECT 709.615 1126.300 2006.070 1126.440 ;
        RECT 709.615 1126.180 709.935 1126.300 ;
        RECT 2006.370 1126.160 2006.690 1126.280 ;
        RECT 706.370 1126.020 706.690 1126.140 ;
        RECT 216.795 1125.880 706.690 1126.020 ;
        RECT 710.585 1126.020 2006.690 1126.160 ;
        RECT 710.585 1125.900 710.905 1126.020 ;
        RECT 2011.730 1125.880 2012.050 1126.000 ;
        RECT 711.730 1125.740 712.050 1125.860 ;
        RECT 216.515 1125.600 712.050 1125.740 ;
        RECT 715.595 1125.740 2012.050 1125.880 ;
        RECT 715.595 1125.620 715.915 1125.740 ;
        RECT 2012.350 1125.600 2012.670 1125.720 ;
        RECT 712.350 1125.460 712.670 1125.580 ;
        RECT 216.235 1125.320 712.670 1125.460 ;
        RECT 716.445 1125.460 2012.670 1125.600 ;
        RECT 716.445 1125.340 716.765 1125.460 ;
        RECT 2017.710 1125.320 2018.030 1125.440 ;
        RECT 717.710 1125.180 718.030 1125.300 ;
        RECT 215.955 1125.040 718.030 1125.180 ;
        RECT 721.575 1125.180 2018.030 1125.320 ;
        RECT 721.575 1125.060 721.895 1125.180 ;
        RECT 2018.330 1125.040 2018.650 1125.160 ;
        RECT 718.330 1124.900 718.650 1125.020 ;
        RECT 215.675 1124.760 718.650 1124.900 ;
        RECT 722.545 1124.900 2018.650 1125.040 ;
        RECT 722.545 1124.780 722.865 1124.900 ;
        RECT 2023.690 1124.760 2024.010 1124.880 ;
        RECT 723.690 1124.620 724.010 1124.740 ;
        RECT 215.395 1124.480 724.010 1124.620 ;
        RECT 727.555 1124.620 2024.010 1124.760 ;
        RECT 727.555 1124.500 727.875 1124.620 ;
        RECT 2024.310 1124.480 2024.630 1124.600 ;
        RECT 724.310 1124.340 724.630 1124.460 ;
        RECT 215.115 1124.200 724.630 1124.340 ;
        RECT 728.525 1124.340 2024.630 1124.480 ;
        RECT 728.525 1124.220 728.845 1124.340 ;
        RECT 2029.670 1124.200 2029.990 1124.320 ;
        RECT 729.670 1124.060 729.990 1124.180 ;
        RECT 214.835 1123.920 729.990 1124.060 ;
        RECT 733.535 1124.060 2029.990 1124.200 ;
        RECT 733.535 1123.940 733.855 1124.060 ;
        RECT 2030.290 1123.920 2030.610 1124.040 ;
        RECT 730.290 1123.780 730.610 1123.900 ;
        RECT 214.555 1123.640 730.610 1123.780 ;
        RECT 734.505 1123.780 2030.610 1123.920 ;
        RECT 734.505 1123.660 734.825 1123.780 ;
        RECT 2035.650 1123.640 2035.970 1123.760 ;
        RECT 735.650 1123.500 735.970 1123.620 ;
        RECT 214.275 1123.360 735.970 1123.500 ;
        RECT 739.515 1123.500 2035.970 1123.640 ;
        RECT 739.515 1123.380 739.835 1123.500 ;
        RECT 2036.270 1123.360 2036.590 1123.480 ;
        RECT 736.270 1123.220 736.590 1123.340 ;
        RECT 213.995 1123.080 736.590 1123.220 ;
        RECT 740.485 1123.220 2036.590 1123.360 ;
        RECT 740.485 1123.100 740.805 1123.220 ;
        RECT 2041.630 1123.080 2041.950 1123.200 ;
        RECT 741.630 1122.940 741.950 1123.060 ;
        RECT 213.715 1122.800 741.950 1122.940 ;
        RECT 745.495 1122.940 2041.950 1123.080 ;
        RECT 745.495 1122.820 745.815 1122.940 ;
        RECT 2042.250 1122.800 2042.570 1122.920 ;
        RECT 742.250 1122.660 742.570 1122.780 ;
        RECT 213.435 1122.520 742.570 1122.660 ;
        RECT 746.465 1122.660 2042.570 1122.800 ;
        RECT 746.465 1122.540 746.785 1122.660 ;
        RECT 2047.610 1122.520 2047.930 1122.640 ;
        RECT 747.610 1122.380 747.930 1122.500 ;
        RECT 213.155 1122.240 747.930 1122.380 ;
        RECT 751.475 1122.380 2047.930 1122.520 ;
        RECT 751.475 1122.260 751.795 1122.380 ;
        RECT 2048.230 1122.240 2048.550 1122.360 ;
        RECT 748.230 1122.100 748.550 1122.220 ;
        RECT 212.875 1121.960 748.550 1122.100 ;
        RECT 752.445 1122.100 2048.550 1122.240 ;
        RECT 752.445 1121.980 752.765 1122.100 ;
        RECT 2053.590 1121.960 2053.910 1122.080 ;
        RECT 753.590 1121.820 753.910 1121.940 ;
        RECT 212.595 1121.680 753.910 1121.820 ;
        RECT 757.455 1121.820 2053.910 1121.960 ;
        RECT 757.455 1121.700 757.775 1121.820 ;
        RECT 2054.210 1121.680 2054.530 1121.800 ;
        RECT 754.210 1121.540 754.530 1121.660 ;
        RECT 212.315 1121.400 754.530 1121.540 ;
        RECT 758.425 1121.540 2054.530 1121.680 ;
        RECT 758.425 1121.420 758.745 1121.540 ;
        RECT 2059.570 1121.400 2059.890 1121.520 ;
        RECT 759.570 1121.260 759.890 1121.380 ;
        RECT 212.035 1121.120 759.890 1121.260 ;
        RECT 763.435 1121.260 2059.890 1121.400 ;
        RECT 763.435 1121.140 763.755 1121.260 ;
        RECT 2060.190 1121.120 2060.510 1121.240 ;
        RECT 764.405 1120.980 2060.510 1121.120 ;
        RECT 764.405 1120.860 764.725 1120.980 ;
        RECT 2065.550 1120.840 2065.870 1120.960 ;
        RECT 769.415 1120.700 2065.870 1120.840 ;
        RECT 769.415 1120.580 769.735 1120.700 ;
        RECT 2066.170 1120.560 2066.490 1120.680 ;
        RECT 770.385 1120.420 2066.490 1120.560 ;
        RECT 770.385 1120.300 770.705 1120.420 ;
        RECT 2071.530 1120.280 2071.850 1120.400 ;
        RECT 775.395 1120.140 2071.850 1120.280 ;
        RECT 775.395 1120.020 775.715 1120.140 ;
        RECT 2072.150 1120.000 2072.470 1120.120 ;
        RECT 776.245 1119.860 2072.470 1120.000 ;
        RECT 776.245 1119.740 776.565 1119.860 ;
        RECT 2077.510 1119.720 2077.830 1119.840 ;
        RECT 781.375 1119.580 2077.830 1119.720 ;
        RECT 781.375 1119.460 781.695 1119.580 ;
        RECT 2078.130 1119.440 2078.450 1119.560 ;
        RECT 782.345 1119.300 2078.450 1119.440 ;
        RECT 782.345 1119.180 782.665 1119.300 ;
        RECT 2083.490 1119.160 2083.810 1119.280 ;
        RECT 787.355 1119.020 2083.810 1119.160 ;
        RECT 787.355 1118.900 787.675 1119.020 ;
        RECT 2084.110 1118.880 2084.430 1119.000 ;
        RECT 788.205 1118.740 2084.430 1118.880 ;
        RECT 788.205 1118.620 788.525 1118.740 ;
        RECT 2089.470 1118.600 2089.790 1118.720 ;
        RECT 793.335 1118.460 2089.790 1118.600 ;
        RECT 793.335 1118.340 793.655 1118.460 ;
        RECT 2090.090 1118.320 2090.410 1118.440 ;
        RECT 794.305 1118.180 2090.410 1118.320 ;
        RECT 794.305 1118.060 794.625 1118.180 ;
        RECT 670.470 1115.450 670.730 1116.420 ;
        RECT 674.180 1115.810 675.390 1116.070 ;
        RECT 676.450 1115.450 676.710 1116.420 ;
        RECT 680.160 1115.810 681.370 1116.070 ;
        RECT 682.430 1115.450 682.690 1116.420 ;
        RECT 686.140 1115.810 687.350 1116.070 ;
        RECT 688.410 1115.450 688.670 1116.420 ;
        RECT 692.120 1115.810 693.330 1116.070 ;
        RECT 694.390 1115.450 694.650 1116.420 ;
        RECT 698.100 1115.810 699.310 1116.070 ;
        RECT 700.370 1115.450 700.630 1116.420 ;
        RECT 704.080 1115.810 705.290 1116.070 ;
        RECT 706.350 1115.450 706.610 1116.420 ;
        RECT 710.060 1115.810 711.270 1116.070 ;
        RECT 712.330 1115.450 712.590 1116.420 ;
        RECT 716.040 1115.810 717.250 1116.070 ;
        RECT 718.310 1115.450 718.570 1116.420 ;
        RECT 722.020 1115.810 723.230 1116.070 ;
        RECT 724.290 1115.450 724.550 1116.420 ;
        RECT 728.000 1115.810 729.210 1116.070 ;
        RECT 730.270 1115.450 730.530 1116.420 ;
        RECT 733.980 1115.810 735.190 1116.070 ;
        RECT 736.250 1115.450 736.510 1116.420 ;
        RECT 739.960 1115.810 741.170 1116.070 ;
        RECT 742.230 1115.450 742.490 1116.420 ;
        RECT 745.940 1115.810 747.150 1116.070 ;
        RECT 748.210 1115.450 748.470 1116.420 ;
        RECT 751.920 1115.810 753.130 1116.070 ;
        RECT 754.190 1115.450 754.450 1116.420 ;
        RECT 757.900 1115.810 759.110 1116.070 ;
        RECT 763.880 1115.810 765.090 1116.070 ;
        RECT 769.860 1115.810 771.070 1116.070 ;
        RECT 775.840 1115.810 777.050 1116.070 ;
        RECT 781.820 1115.810 783.030 1116.070 ;
        RECT 787.800 1115.810 789.010 1116.070 ;
        RECT 793.780 1115.810 794.990 1116.070 ;
        RECT 1970.470 1115.450 1970.730 1116.420 ;
        RECT 1976.450 1115.450 1976.710 1116.420 ;
        RECT 1982.430 1115.450 1982.690 1116.420 ;
        RECT 1988.410 1115.450 1988.670 1116.420 ;
        RECT 1994.390 1115.450 1994.650 1116.420 ;
        RECT 2000.370 1115.450 2000.630 1116.420 ;
        RECT 2006.350 1115.450 2006.610 1116.420 ;
        RECT 2012.330 1115.450 2012.590 1116.420 ;
        RECT 2018.310 1115.450 2018.570 1116.420 ;
        RECT 2024.290 1115.450 2024.550 1116.420 ;
        RECT 2030.270 1115.450 2030.530 1116.420 ;
        RECT 2036.250 1115.450 2036.510 1116.420 ;
        RECT 2042.230 1115.450 2042.490 1116.420 ;
        RECT 2048.210 1115.450 2048.470 1116.420 ;
        RECT 2054.190 1115.450 2054.450 1116.420 ;
        RECT 2060.170 1115.450 2060.430 1116.420 ;
        RECT 2066.150 1115.450 2066.410 1116.420 ;
        RECT 2072.130 1115.450 2072.390 1116.420 ;
        RECT 2078.110 1115.450 2078.370 1116.420 ;
        RECT 2084.090 1115.450 2084.350 1116.420 ;
        RECT 2090.070 1115.450 2090.330 1116.420 ;
        RECT 675.530 1112.750 676.740 1113.010 ;
        RECT 679.680 1112.390 679.940 1113.360 ;
        RECT 681.510 1112.750 682.720 1113.010 ;
        RECT 685.660 1112.390 685.920 1113.360 ;
        RECT 687.490 1112.750 688.700 1113.010 ;
        RECT 691.640 1112.390 691.900 1113.360 ;
        RECT 693.470 1112.750 694.680 1113.010 ;
        RECT 697.620 1112.390 697.880 1113.360 ;
        RECT 699.450 1112.750 700.660 1113.010 ;
        RECT 703.600 1112.390 703.860 1113.360 ;
        RECT 705.430 1112.750 706.640 1113.010 ;
        RECT 709.580 1112.390 709.840 1113.360 ;
        RECT 711.410 1112.750 712.620 1113.010 ;
        RECT 715.560 1112.390 715.820 1113.360 ;
        RECT 717.390 1112.750 718.600 1113.010 ;
        RECT 721.540 1112.390 721.800 1113.360 ;
        RECT 723.370 1112.750 724.580 1113.010 ;
        RECT 727.520 1112.390 727.780 1113.360 ;
        RECT 729.350 1112.750 730.560 1113.010 ;
        RECT 733.500 1112.390 733.760 1113.360 ;
        RECT 735.330 1112.750 736.540 1113.010 ;
        RECT 739.480 1112.390 739.740 1113.360 ;
        RECT 741.310 1112.750 742.520 1113.010 ;
        RECT 745.460 1112.390 745.720 1113.360 ;
        RECT 747.290 1112.750 748.500 1113.010 ;
        RECT 751.440 1112.390 751.700 1113.360 ;
        RECT 753.270 1112.750 754.480 1113.010 ;
        RECT 757.420 1112.390 757.680 1113.360 ;
        RECT 759.250 1112.750 760.460 1113.010 ;
        RECT 763.400 1112.390 763.660 1113.360 ;
        RECT 769.380 1112.390 769.640 1113.360 ;
        RECT 775.360 1112.390 775.620 1113.360 ;
        RECT 781.340 1112.390 781.600 1113.360 ;
        RECT 787.320 1112.390 787.580 1113.360 ;
        RECT 793.280 1112.750 794.490 1113.010 ;
        RECT 1975.530 1112.750 1976.740 1113.010 ;
        RECT 1981.510 1112.750 1982.720 1113.010 ;
        RECT 1987.490 1112.750 1988.700 1113.010 ;
        RECT 1993.470 1112.750 1994.680 1113.010 ;
        RECT 1999.450 1112.750 2000.660 1113.010 ;
        RECT 2005.430 1112.750 2006.640 1113.010 ;
        RECT 2011.410 1112.750 2012.620 1113.010 ;
        RECT 2017.390 1112.750 2018.600 1113.010 ;
        RECT 2023.370 1112.750 2024.580 1113.010 ;
        RECT 2029.350 1112.750 2030.560 1113.010 ;
        RECT 2035.330 1112.750 2036.540 1113.010 ;
        RECT 2041.310 1112.750 2042.520 1113.010 ;
        RECT 2047.290 1112.750 2048.500 1113.010 ;
        RECT 2053.270 1112.750 2054.480 1113.010 ;
        RECT 2059.250 1112.750 2060.460 1113.010 ;
        RECT 2065.230 1112.750 2066.440 1113.010 ;
        RECT 2071.210 1112.750 2072.420 1113.010 ;
        RECT 2077.190 1112.750 2078.400 1113.010 ;
        RECT 2083.170 1112.750 2084.380 1113.010 ;
        RECT 2090.080 1112.390 2090.340 1113.360 ;
      LAYER via ;
        RECT 2087.570 4986.375 2088.660 4986.635 ;
        RECT 3314.315 4985.675 3314.575 4986.525 ;
        RECT 3317.575 4985.965 3318.665 4986.225 ;
        RECT 3323.555 4985.965 3324.645 4986.225 ;
        RECT 3329.535 4985.965 3330.625 4986.225 ;
        RECT 3335.515 4985.965 3336.605 4986.225 ;
        RECT 835.260 4984.750 836.350 4985.010 ;
        RECT 841.240 4984.750 842.330 4985.010 ;
        RECT 847.220 4984.750 848.310 4985.010 ;
        RECT 2087.540 4983.025 2087.800 4983.875 ;
        RECT 3312.945 4982.905 3314.035 4983.165 ;
        RECT 3317.545 4982.615 3317.805 4983.465 ;
        RECT 3323.525 4982.615 3323.785 4983.465 ;
        RECT 3329.505 4982.615 3329.765 4983.465 ;
        RECT 3335.485 4982.615 3335.745 4983.465 ;
        RECT 836.120 4981.400 836.380 4982.250 ;
        RECT 842.100 4981.400 842.360 4982.250 ;
        RECT 848.080 4981.400 848.340 4982.250 ;
        RECT 202.770 4456.000 203.030 4457.090 ;
        RECT 848.130 4977.025 848.390 4977.285 ;
        RECT 212.335 4456.495 212.595 4456.755 ;
        RECT 847.510 4976.745 847.770 4977.005 ;
        RECT 199.410 4455.460 200.260 4455.720 ;
        RECT 212.615 4455.525 212.875 4455.785 ;
        RECT 199.710 4451.370 199.970 4452.460 ;
        RECT 202.470 4452.230 203.320 4452.490 ;
        RECT 212.315 4452.280 212.575 4452.540 ;
        RECT 202.770 4450.020 203.030 4451.110 ;
        RECT 199.410 4449.480 200.260 4449.740 ;
        RECT 199.710 4445.390 199.970 4446.480 ;
        RECT 202.470 4446.250 203.320 4446.510 ;
        RECT 202.770 4444.040 203.030 4445.130 ;
        RECT 199.410 4443.500 200.260 4443.760 ;
        RECT 199.710 4439.410 199.970 4440.500 ;
        RECT 202.470 4440.270 203.320 4440.530 ;
        RECT 199.710 4433.430 199.970 4434.520 ;
        RECT 202.470 4434.290 203.320 4434.550 ;
        RECT 199.710 4427.450 199.970 4428.540 ;
        RECT 202.470 4428.310 203.320 4428.570 ;
        RECT 202.895 3052.770 203.155 3053.860 ;
        RECT 212.195 3053.265 212.455 3053.525 ;
        RECT 212.595 4451.660 212.855 4451.920 ;
        RECT 842.150 4976.465 842.410 4976.725 ;
        RECT 212.895 4450.395 213.155 4450.655 ;
        RECT 841.530 4976.185 841.790 4976.445 ;
        RECT 213.175 4449.545 213.435 4449.805 ;
        RECT 199.535 3052.230 200.385 3052.490 ;
        RECT 212.475 3052.295 212.735 3052.555 ;
        RECT 212.875 4446.300 213.135 4446.560 ;
        RECT 199.835 3048.140 200.095 3049.230 ;
        RECT 202.595 3049.000 203.445 3049.260 ;
        RECT 212.175 3049.050 212.435 3049.310 ;
        RECT 202.895 3046.790 203.155 3047.880 ;
        RECT 199.535 3046.250 200.385 3046.510 ;
        RECT 199.835 3042.160 200.095 3043.250 ;
        RECT 202.595 3043.020 203.445 3043.280 ;
        RECT 202.895 3040.810 203.155 3041.900 ;
        RECT 199.535 3040.270 200.385 3040.530 ;
        RECT 199.835 3036.180 200.095 3037.270 ;
        RECT 202.595 3037.040 203.445 3037.300 ;
        RECT 202.895 3034.830 203.155 3035.920 ;
        RECT 199.535 3034.290 200.385 3034.550 ;
        RECT 199.835 3030.200 200.095 3031.290 ;
        RECT 202.595 3031.060 203.445 3031.320 ;
        RECT 202.895 3028.850 203.155 3029.940 ;
        RECT 199.535 3028.310 200.385 3028.570 ;
        RECT 199.835 3024.220 200.095 3025.310 ;
        RECT 202.595 3025.080 203.445 3025.340 ;
        RECT 199.835 3018.240 200.095 3019.330 ;
        RECT 202.595 3019.100 203.445 3019.360 ;
        RECT 199.835 3012.260 200.095 3013.350 ;
        RECT 202.595 3013.120 203.445 3013.380 ;
        RECT 199.835 3006.280 200.095 3007.370 ;
        RECT 202.595 3007.140 203.445 3007.400 ;
        RECT 199.835 3000.300 200.095 3001.390 ;
        RECT 202.595 3001.160 203.445 3001.420 ;
        RECT 199.835 2994.320 200.095 2995.410 ;
        RECT 202.595 2995.180 203.445 2995.440 ;
        RECT 199.835 2988.340 200.095 2989.430 ;
        RECT 202.595 2989.200 203.445 2989.460 ;
        RECT 203.005 1761.865 203.265 1762.955 ;
        RECT 212.055 1762.360 212.315 1762.620 ;
        RECT 212.455 3048.430 212.715 3048.690 ;
        RECT 212.755 3047.165 213.015 3047.425 ;
        RECT 213.155 4445.680 213.415 4445.940 ;
        RECT 836.170 4975.905 836.430 4976.165 ;
        RECT 2087.490 4976.115 2087.750 4976.375 ;
        RECT 3313.280 4976.095 3313.540 4976.355 ;
        RECT 3317.495 4976.115 3317.755 4976.375 ;
        RECT 213.455 4444.535 213.715 4444.795 ;
        RECT 835.550 4975.625 835.810 4975.885 ;
        RECT 2088.110 4975.835 2088.370 4976.095 ;
        RECT 3314.250 4975.815 3314.510 4976.075 ;
        RECT 3318.115 4975.835 3318.375 4976.095 ;
        RECT 3323.475 4975.555 3323.735 4975.815 ;
        RECT 3324.095 4975.275 3324.355 4975.535 ;
        RECT 3329.455 4974.995 3329.715 4975.255 ;
        RECT 3330.075 4974.715 3330.335 4974.975 ;
        RECT 3335.435 4974.435 3335.695 4974.695 ;
        RECT 3336.055 4974.155 3336.315 4974.415 ;
        RECT 213.735 4443.565 213.995 4443.825 ;
        RECT 213.035 3046.315 213.295 3046.575 ;
        RECT 213.435 4440.320 213.695 4440.580 ;
        RECT 199.645 1761.325 200.495 1761.585 ;
        RECT 212.335 1761.390 212.595 1761.650 ;
        RECT 212.735 3043.070 212.995 3043.330 ;
        RECT 199.945 1757.235 200.205 1758.325 ;
        RECT 202.705 1758.095 203.555 1758.355 ;
        RECT 212.035 1758.145 212.295 1758.405 ;
        RECT 203.005 1755.885 203.265 1756.975 ;
        RECT 199.645 1755.345 200.495 1755.605 ;
        RECT 199.945 1751.255 200.205 1752.345 ;
        RECT 202.705 1752.115 203.555 1752.375 ;
        RECT 203.005 1749.905 203.265 1750.995 ;
        RECT 199.645 1749.365 200.495 1749.625 ;
        RECT 199.945 1745.275 200.205 1746.365 ;
        RECT 202.705 1746.135 203.555 1746.395 ;
        RECT 203.005 1743.925 203.265 1745.015 ;
        RECT 199.645 1743.385 200.495 1743.645 ;
        RECT 199.945 1739.295 200.205 1740.385 ;
        RECT 202.705 1740.155 203.555 1740.415 ;
        RECT 203.005 1737.945 203.265 1739.035 ;
        RECT 199.645 1737.405 200.495 1737.665 ;
        RECT 199.945 1733.315 200.205 1734.405 ;
        RECT 202.705 1734.175 203.555 1734.435 ;
        RECT 203.005 1731.965 203.265 1733.055 ;
        RECT 199.645 1731.425 200.495 1731.685 ;
        RECT 199.945 1727.335 200.205 1728.425 ;
        RECT 202.705 1728.195 203.555 1728.455 ;
        RECT 203.005 1725.985 203.265 1727.075 ;
        RECT 199.645 1725.445 200.495 1725.705 ;
        RECT 199.945 1721.355 200.205 1722.445 ;
        RECT 202.705 1722.215 203.555 1722.475 ;
        RECT 203.005 1720.005 203.265 1721.095 ;
        RECT 199.645 1719.465 200.495 1719.725 ;
        RECT 199.945 1715.375 200.205 1716.465 ;
        RECT 202.705 1716.235 203.555 1716.495 ;
        RECT 203.005 1714.025 203.265 1715.115 ;
        RECT 199.645 1713.485 200.495 1713.745 ;
        RECT 199.945 1709.395 200.205 1710.485 ;
        RECT 202.705 1710.255 203.555 1710.515 ;
        RECT 203.005 1708.045 203.265 1709.135 ;
        RECT 199.645 1707.505 200.495 1707.765 ;
        RECT 199.945 1703.415 200.205 1704.505 ;
        RECT 202.705 1704.275 203.555 1704.535 ;
        RECT 203.005 1702.065 203.265 1703.155 ;
        RECT 199.645 1701.525 200.495 1701.785 ;
        RECT 199.945 1697.435 200.205 1698.525 ;
        RECT 202.705 1698.295 203.555 1698.555 ;
        RECT 199.945 1691.455 200.205 1692.545 ;
        RECT 202.705 1692.315 203.555 1692.575 ;
        RECT 199.945 1685.475 200.205 1686.565 ;
        RECT 202.705 1686.335 203.555 1686.595 ;
        RECT 199.945 1679.495 200.205 1680.585 ;
        RECT 202.705 1680.355 203.555 1680.615 ;
        RECT 199.945 1673.515 200.205 1674.605 ;
        RECT 202.705 1674.375 203.555 1674.635 ;
        RECT 212.315 1757.525 212.575 1757.785 ;
        RECT 212.615 1756.260 212.875 1756.520 ;
        RECT 213.015 3042.450 213.275 3042.710 ;
        RECT 213.315 3041.305 213.575 3041.565 ;
        RECT 213.715 4439.700 213.975 4439.960 ;
        RECT 213.595 3040.335 213.855 3040.595 ;
        RECT 213.995 4434.340 214.255 4434.600 ;
        RECT 212.895 1755.410 213.155 1755.670 ;
        RECT 213.295 3037.090 213.555 3037.350 ;
        RECT 212.595 1752.165 212.855 1752.425 ;
        RECT 212.875 1751.545 213.135 1751.805 ;
        RECT 213.175 1750.400 213.435 1750.660 ;
        RECT 213.575 3036.470 213.835 3036.730 ;
        RECT 213.875 3035.205 214.135 3035.465 ;
        RECT 214.275 4433.720 214.535 4433.980 ;
        RECT 214.155 3034.355 214.415 3034.615 ;
        RECT 214.555 4428.360 214.815 4428.620 ;
        RECT 213.455 1749.430 213.715 1749.690 ;
        RECT 213.855 3031.110 214.115 3031.370 ;
        RECT 213.155 1746.185 213.415 1746.445 ;
        RECT 213.435 1745.565 213.695 1745.825 ;
        RECT 213.735 1744.300 213.995 1744.560 ;
        RECT 214.135 3030.490 214.395 3030.750 ;
        RECT 214.435 3029.345 214.695 3029.605 ;
        RECT 214.835 4427.740 215.095 4428.000 ;
        RECT 3375.460 3571.575 3375.720 3571.835 ;
        RECT 3384.640 3571.200 3384.900 3572.290 ;
        RECT 3375.180 3570.725 3375.440 3570.985 ;
        RECT 3387.410 3570.660 3388.260 3570.920 ;
        RECT 3375.480 3567.480 3375.740 3567.740 ;
        RECT 3375.200 3566.860 3375.460 3567.120 ;
        RECT 3374.900 3565.715 3375.160 3565.975 ;
        RECT 3374.620 3564.745 3374.880 3565.005 ;
        RECT 3374.920 3561.500 3375.180 3561.760 ;
        RECT 3374.640 3560.880 3374.900 3561.140 ;
        RECT 3374.340 3559.735 3374.600 3559.995 ;
        RECT 3374.060 3558.765 3374.320 3559.025 ;
        RECT 3374.360 3555.520 3374.620 3555.780 ;
        RECT 3374.080 3554.900 3374.340 3555.160 ;
        RECT 3373.780 3553.755 3374.040 3554.015 ;
        RECT 3373.500 3552.785 3373.760 3553.045 ;
        RECT 3373.800 3549.540 3374.060 3549.800 ;
        RECT 3373.520 3548.920 3373.780 3549.180 ;
        RECT 3373.240 3543.560 3373.500 3543.820 ;
        RECT 3372.960 3542.940 3373.220 3543.200 ;
        RECT 3372.680 3537.580 3372.940 3537.840 ;
        RECT 3372.400 3536.960 3372.660 3537.220 ;
        RECT 214.715 3028.375 214.975 3028.635 ;
        RECT 214.015 1743.450 214.275 1743.710 ;
        RECT 214.415 3025.130 214.675 3025.390 ;
        RECT 213.715 1740.205 213.975 1740.465 ;
        RECT 213.995 1739.585 214.255 1739.845 ;
        RECT 214.295 1738.440 214.555 1738.700 ;
        RECT 214.695 3024.510 214.955 3024.770 ;
        RECT 214.575 1737.470 214.835 1737.730 ;
        RECT 214.975 3019.150 215.235 3019.410 ;
        RECT 214.275 1734.225 214.535 1734.485 ;
        RECT 214.555 1733.605 214.815 1733.865 ;
        RECT 214.855 1732.460 215.115 1732.720 ;
        RECT 215.255 3018.530 215.515 3018.790 ;
        RECT 215.135 1731.490 215.395 1731.750 ;
        RECT 215.535 3013.170 215.795 3013.430 ;
        RECT 214.835 1728.245 215.095 1728.505 ;
        RECT 215.115 1727.625 215.375 1727.885 ;
        RECT 215.415 1726.480 215.675 1726.740 ;
        RECT 215.815 3012.550 216.075 3012.810 ;
        RECT 215.695 1725.510 215.955 1725.770 ;
        RECT 216.095 3007.190 216.355 3007.450 ;
        RECT 215.395 1722.265 215.655 1722.525 ;
        RECT 215.675 1721.645 215.935 1721.905 ;
        RECT 215.975 1720.500 216.235 1720.760 ;
        RECT 216.375 3006.570 216.635 3006.830 ;
        RECT 216.255 1719.530 216.515 1719.790 ;
        RECT 216.655 3001.210 216.915 3001.470 ;
        RECT 215.955 1716.285 216.215 1716.545 ;
        RECT 216.235 1715.665 216.495 1715.925 ;
        RECT 216.535 1714.520 216.795 1714.780 ;
        RECT 216.935 3000.590 217.195 3000.850 ;
        RECT 216.815 1713.550 217.075 1713.810 ;
        RECT 217.215 2995.230 217.475 2995.490 ;
        RECT 216.515 1710.305 216.775 1710.565 ;
        RECT 216.795 1709.685 217.055 1709.945 ;
        RECT 217.095 1708.540 217.355 1708.800 ;
        RECT 217.495 2994.610 217.755 2994.870 ;
        RECT 217.375 1707.570 217.635 1707.830 ;
        RECT 217.775 2989.250 218.035 2989.510 ;
        RECT 217.075 1704.325 217.335 1704.585 ;
        RECT 217.355 1703.705 217.615 1703.965 ;
        RECT 217.655 1702.560 217.915 1702.820 ;
        RECT 218.055 2988.630 218.315 2988.890 ;
        RECT 3384.350 3567.430 3385.200 3567.690 ;
        RECT 3387.700 3566.570 3387.960 3567.660 ;
        RECT 3384.640 3565.220 3384.900 3566.310 ;
        RECT 3387.410 3564.680 3388.260 3564.940 ;
        RECT 3384.350 3561.450 3385.200 3561.710 ;
        RECT 3387.700 3560.590 3387.960 3561.680 ;
        RECT 3384.640 3559.240 3384.900 3560.330 ;
        RECT 3387.410 3558.700 3388.260 3558.960 ;
        RECT 3384.350 3555.470 3385.200 3555.730 ;
        RECT 3387.700 3554.610 3387.960 3555.700 ;
        RECT 3384.640 3553.260 3384.900 3554.350 ;
        RECT 3387.410 3552.720 3388.260 3552.980 ;
        RECT 3384.350 3549.490 3385.200 3549.750 ;
        RECT 3387.700 3548.630 3387.960 3549.720 ;
        RECT 3384.350 3543.510 3385.200 3543.770 ;
        RECT 3387.700 3542.650 3387.960 3543.740 ;
        RECT 3384.350 3537.530 3385.200 3537.790 ;
        RECT 3387.700 3536.670 3387.960 3537.760 ;
        RECT 3375.460 2267.575 3375.720 2267.835 ;
        RECT 3384.640 2267.080 3384.900 2268.170 ;
        RECT 3375.180 2266.605 3375.440 2266.865 ;
        RECT 3387.410 2266.540 3388.260 2266.800 ;
        RECT 3374.900 2261.475 3375.160 2261.735 ;
        RECT 3384.640 2261.100 3384.900 2262.190 ;
        RECT 3374.620 2260.625 3374.880 2260.885 ;
        RECT 3387.410 2260.560 3388.260 2260.820 ;
        RECT 3374.340 2255.615 3374.600 2255.875 ;
        RECT 3384.640 2255.120 3384.900 2256.210 ;
        RECT 3374.060 2254.645 3374.320 2254.905 ;
        RECT 3387.410 2254.580 3388.260 2254.840 ;
        RECT 3373.780 2249.515 3374.040 2249.775 ;
        RECT 3384.640 2249.140 3384.900 2250.230 ;
        RECT 3373.500 2248.665 3373.760 2248.925 ;
        RECT 3387.410 2248.600 3388.260 2248.860 ;
        RECT 3373.220 2243.655 3373.480 2243.915 ;
        RECT 3384.640 2243.160 3384.900 2244.250 ;
        RECT 3372.940 2242.685 3373.200 2242.945 ;
        RECT 3387.410 2242.620 3388.260 2242.880 ;
        RECT 3372.660 2237.675 3372.920 2237.935 ;
        RECT 3384.640 2237.180 3384.900 2238.270 ;
        RECT 3372.380 2236.705 3372.640 2236.965 ;
        RECT 3387.410 2236.640 3388.260 2236.900 ;
        RECT 217.935 1701.590 218.195 1701.850 ;
        RECT 217.635 1698.345 217.895 1698.605 ;
        RECT 217.915 1697.725 218.175 1697.985 ;
        RECT 218.195 1692.365 218.455 1692.625 ;
        RECT 218.475 1691.745 218.735 1692.005 ;
        RECT 218.755 1686.385 219.015 1686.645 ;
        RECT 219.035 1685.765 219.295 1686.025 ;
        RECT 219.315 1680.405 219.575 1680.665 ;
        RECT 219.595 1679.785 219.855 1680.045 ;
        RECT 219.875 1674.425 220.135 1674.685 ;
        RECT 220.155 1673.805 220.415 1674.065 ;
        RECT 670.520 1129.240 670.780 1129.500 ;
        RECT 674.735 1129.260 674.995 1129.520 ;
        RECT 1970.520 1129.380 1970.780 1129.640 ;
        RECT 675.880 1128.960 676.140 1129.220 ;
        RECT 679.745 1128.980 680.005 1129.240 ;
        RECT 1975.880 1129.100 1976.140 1129.360 ;
        RECT 676.500 1128.680 676.760 1128.940 ;
        RECT 680.715 1128.700 680.975 1128.960 ;
        RECT 1976.500 1128.820 1976.760 1129.080 ;
        RECT 681.860 1128.400 682.120 1128.660 ;
        RECT 685.725 1128.420 685.985 1128.680 ;
        RECT 1981.860 1128.540 1982.120 1128.800 ;
        RECT 682.480 1128.120 682.740 1128.380 ;
        RECT 686.695 1128.140 686.955 1128.400 ;
        RECT 1982.480 1128.260 1982.740 1128.520 ;
        RECT 687.840 1127.840 688.100 1128.100 ;
        RECT 691.705 1127.860 691.965 1128.120 ;
        RECT 1987.840 1127.980 1988.100 1128.240 ;
        RECT 688.460 1127.560 688.720 1127.820 ;
        RECT 692.675 1127.580 692.935 1127.840 ;
        RECT 1988.460 1127.700 1988.720 1127.960 ;
        RECT 693.820 1127.280 694.080 1127.540 ;
        RECT 697.685 1127.300 697.945 1127.560 ;
        RECT 1993.820 1127.420 1994.080 1127.680 ;
        RECT 694.440 1127.000 694.700 1127.260 ;
        RECT 698.655 1127.020 698.915 1127.280 ;
        RECT 1994.440 1127.140 1994.700 1127.400 ;
        RECT 699.800 1126.720 700.060 1126.980 ;
        RECT 703.665 1126.740 703.925 1127.000 ;
        RECT 1999.800 1126.860 2000.060 1127.120 ;
        RECT 700.420 1126.440 700.680 1126.700 ;
        RECT 704.515 1126.460 704.775 1126.720 ;
        RECT 2000.420 1126.580 2000.680 1126.840 ;
        RECT 705.780 1126.160 706.040 1126.420 ;
        RECT 709.645 1126.180 709.905 1126.440 ;
        RECT 2005.780 1126.300 2006.040 1126.560 ;
        RECT 706.400 1125.880 706.660 1126.140 ;
        RECT 710.615 1125.900 710.875 1126.160 ;
        RECT 2006.400 1126.020 2006.660 1126.280 ;
        RECT 711.760 1125.600 712.020 1125.860 ;
        RECT 715.625 1125.620 715.885 1125.880 ;
        RECT 2011.760 1125.740 2012.020 1126.000 ;
        RECT 712.380 1125.320 712.640 1125.580 ;
        RECT 716.475 1125.340 716.735 1125.600 ;
        RECT 2012.380 1125.460 2012.640 1125.720 ;
        RECT 717.740 1125.040 718.000 1125.300 ;
        RECT 721.605 1125.060 721.865 1125.320 ;
        RECT 2017.740 1125.180 2018.000 1125.440 ;
        RECT 718.360 1124.760 718.620 1125.020 ;
        RECT 722.575 1124.780 722.835 1125.040 ;
        RECT 2018.360 1124.900 2018.620 1125.160 ;
        RECT 723.720 1124.480 723.980 1124.740 ;
        RECT 727.585 1124.500 727.845 1124.760 ;
        RECT 2023.720 1124.620 2023.980 1124.880 ;
        RECT 724.340 1124.200 724.600 1124.460 ;
        RECT 728.555 1124.220 728.815 1124.480 ;
        RECT 2024.340 1124.340 2024.600 1124.600 ;
        RECT 729.700 1123.920 729.960 1124.180 ;
        RECT 733.565 1123.940 733.825 1124.200 ;
        RECT 2029.700 1124.060 2029.960 1124.320 ;
        RECT 730.320 1123.640 730.580 1123.900 ;
        RECT 734.535 1123.660 734.795 1123.920 ;
        RECT 2030.320 1123.780 2030.580 1124.040 ;
        RECT 735.680 1123.360 735.940 1123.620 ;
        RECT 739.545 1123.380 739.805 1123.640 ;
        RECT 2035.680 1123.500 2035.940 1123.760 ;
        RECT 736.300 1123.080 736.560 1123.340 ;
        RECT 740.515 1123.100 740.775 1123.360 ;
        RECT 2036.300 1123.220 2036.560 1123.480 ;
        RECT 741.660 1122.800 741.920 1123.060 ;
        RECT 745.525 1122.820 745.785 1123.080 ;
        RECT 2041.660 1122.940 2041.920 1123.200 ;
        RECT 742.280 1122.520 742.540 1122.780 ;
        RECT 746.495 1122.540 746.755 1122.800 ;
        RECT 2042.280 1122.660 2042.540 1122.920 ;
        RECT 747.640 1122.240 747.900 1122.500 ;
        RECT 751.505 1122.260 751.765 1122.520 ;
        RECT 2047.640 1122.380 2047.900 1122.640 ;
        RECT 748.260 1121.960 748.520 1122.220 ;
        RECT 752.475 1121.980 752.735 1122.240 ;
        RECT 2048.260 1122.100 2048.520 1122.360 ;
        RECT 753.620 1121.680 753.880 1121.940 ;
        RECT 757.485 1121.700 757.745 1121.960 ;
        RECT 2053.620 1121.820 2053.880 1122.080 ;
        RECT 754.240 1121.400 754.500 1121.660 ;
        RECT 758.455 1121.420 758.715 1121.680 ;
        RECT 2054.240 1121.540 2054.500 1121.800 ;
        RECT 759.600 1121.120 759.860 1121.380 ;
        RECT 763.465 1121.140 763.725 1121.400 ;
        RECT 2059.600 1121.260 2059.860 1121.520 ;
        RECT 764.435 1120.860 764.695 1121.120 ;
        RECT 2060.220 1120.980 2060.480 1121.240 ;
        RECT 769.445 1120.580 769.705 1120.840 ;
        RECT 2065.580 1120.700 2065.840 1120.960 ;
        RECT 770.415 1120.300 770.675 1120.560 ;
        RECT 2066.200 1120.420 2066.460 1120.680 ;
        RECT 775.425 1120.020 775.685 1120.280 ;
        RECT 2071.560 1120.140 2071.820 1120.400 ;
        RECT 776.275 1119.740 776.535 1120.000 ;
        RECT 2072.180 1119.860 2072.440 1120.120 ;
        RECT 781.405 1119.460 781.665 1119.720 ;
        RECT 2077.540 1119.580 2077.800 1119.840 ;
        RECT 782.375 1119.180 782.635 1119.440 ;
        RECT 2078.160 1119.300 2078.420 1119.560 ;
        RECT 787.385 1118.900 787.645 1119.160 ;
        RECT 2083.520 1119.020 2083.780 1119.280 ;
        RECT 788.235 1118.620 788.495 1118.880 ;
        RECT 2084.140 1118.740 2084.400 1119.000 ;
        RECT 793.365 1118.340 793.625 1118.600 ;
        RECT 2089.500 1118.460 2089.760 1118.720 ;
        RECT 794.335 1118.060 794.595 1118.320 ;
        RECT 2090.120 1118.180 2090.380 1118.440 ;
        RECT 670.470 1115.510 670.730 1116.360 ;
        RECT 674.240 1115.810 675.330 1116.070 ;
        RECT 676.450 1115.510 676.710 1116.360 ;
        RECT 680.220 1115.810 681.310 1116.070 ;
        RECT 682.430 1115.510 682.690 1116.360 ;
        RECT 686.200 1115.810 687.290 1116.070 ;
        RECT 688.410 1115.510 688.670 1116.360 ;
        RECT 692.180 1115.810 693.270 1116.070 ;
        RECT 694.390 1115.510 694.650 1116.360 ;
        RECT 698.160 1115.810 699.250 1116.070 ;
        RECT 700.370 1115.510 700.630 1116.360 ;
        RECT 704.140 1115.810 705.230 1116.070 ;
        RECT 706.350 1115.510 706.610 1116.360 ;
        RECT 710.120 1115.810 711.210 1116.070 ;
        RECT 712.330 1115.510 712.590 1116.360 ;
        RECT 716.100 1115.810 717.190 1116.070 ;
        RECT 718.310 1115.510 718.570 1116.360 ;
        RECT 722.080 1115.810 723.170 1116.070 ;
        RECT 724.290 1115.510 724.550 1116.360 ;
        RECT 728.060 1115.810 729.150 1116.070 ;
        RECT 730.270 1115.510 730.530 1116.360 ;
        RECT 734.040 1115.810 735.130 1116.070 ;
        RECT 736.250 1115.510 736.510 1116.360 ;
        RECT 740.020 1115.810 741.110 1116.070 ;
        RECT 742.230 1115.510 742.490 1116.360 ;
        RECT 746.000 1115.810 747.090 1116.070 ;
        RECT 748.210 1115.510 748.470 1116.360 ;
        RECT 751.980 1115.810 753.070 1116.070 ;
        RECT 754.190 1115.510 754.450 1116.360 ;
        RECT 757.960 1115.810 759.050 1116.070 ;
        RECT 763.940 1115.810 765.030 1116.070 ;
        RECT 769.920 1115.810 771.010 1116.070 ;
        RECT 775.900 1115.810 776.990 1116.070 ;
        RECT 781.880 1115.810 782.970 1116.070 ;
        RECT 787.860 1115.810 788.950 1116.070 ;
        RECT 793.840 1115.810 794.930 1116.070 ;
        RECT 1970.470 1115.510 1970.730 1116.360 ;
        RECT 1976.450 1115.510 1976.710 1116.360 ;
        RECT 1982.430 1115.510 1982.690 1116.360 ;
        RECT 1988.410 1115.510 1988.670 1116.360 ;
        RECT 1994.390 1115.510 1994.650 1116.360 ;
        RECT 2000.370 1115.510 2000.630 1116.360 ;
        RECT 2006.350 1115.510 2006.610 1116.360 ;
        RECT 2012.330 1115.510 2012.590 1116.360 ;
        RECT 2018.310 1115.510 2018.570 1116.360 ;
        RECT 2024.290 1115.510 2024.550 1116.360 ;
        RECT 2030.270 1115.510 2030.530 1116.360 ;
        RECT 2036.250 1115.510 2036.510 1116.360 ;
        RECT 2042.230 1115.510 2042.490 1116.360 ;
        RECT 2048.210 1115.510 2048.470 1116.360 ;
        RECT 2054.190 1115.510 2054.450 1116.360 ;
        RECT 2060.170 1115.510 2060.430 1116.360 ;
        RECT 2066.150 1115.510 2066.410 1116.360 ;
        RECT 2072.130 1115.510 2072.390 1116.360 ;
        RECT 2078.110 1115.510 2078.370 1116.360 ;
        RECT 2084.090 1115.510 2084.350 1116.360 ;
        RECT 2090.070 1115.510 2090.330 1116.360 ;
        RECT 675.590 1112.750 676.680 1113.010 ;
        RECT 679.680 1112.450 679.940 1113.300 ;
        RECT 681.570 1112.750 682.660 1113.010 ;
        RECT 685.660 1112.450 685.920 1113.300 ;
        RECT 687.550 1112.750 688.640 1113.010 ;
        RECT 691.640 1112.450 691.900 1113.300 ;
        RECT 693.530 1112.750 694.620 1113.010 ;
        RECT 697.620 1112.450 697.880 1113.300 ;
        RECT 699.510 1112.750 700.600 1113.010 ;
        RECT 703.600 1112.450 703.860 1113.300 ;
        RECT 705.490 1112.750 706.580 1113.010 ;
        RECT 709.580 1112.450 709.840 1113.300 ;
        RECT 711.470 1112.750 712.560 1113.010 ;
        RECT 715.560 1112.450 715.820 1113.300 ;
        RECT 717.450 1112.750 718.540 1113.010 ;
        RECT 721.540 1112.450 721.800 1113.300 ;
        RECT 723.430 1112.750 724.520 1113.010 ;
        RECT 727.520 1112.450 727.780 1113.300 ;
        RECT 729.410 1112.750 730.500 1113.010 ;
        RECT 733.500 1112.450 733.760 1113.300 ;
        RECT 735.390 1112.750 736.480 1113.010 ;
        RECT 739.480 1112.450 739.740 1113.300 ;
        RECT 741.370 1112.750 742.460 1113.010 ;
        RECT 745.460 1112.450 745.720 1113.300 ;
        RECT 747.350 1112.750 748.440 1113.010 ;
        RECT 751.440 1112.450 751.700 1113.300 ;
        RECT 753.330 1112.750 754.420 1113.010 ;
        RECT 757.420 1112.450 757.680 1113.300 ;
        RECT 759.310 1112.750 760.400 1113.010 ;
        RECT 763.400 1112.450 763.660 1113.300 ;
        RECT 769.380 1112.450 769.640 1113.300 ;
        RECT 775.360 1112.450 775.620 1113.300 ;
        RECT 781.340 1112.450 781.600 1113.300 ;
        RECT 787.320 1112.450 787.580 1113.300 ;
        RECT 793.340 1112.750 794.430 1113.010 ;
        RECT 1975.590 1112.750 1976.680 1113.010 ;
        RECT 1981.570 1112.750 1982.660 1113.010 ;
        RECT 1987.550 1112.750 1988.640 1113.010 ;
        RECT 1993.530 1112.750 1994.620 1113.010 ;
        RECT 1999.510 1112.750 2000.600 1113.010 ;
        RECT 2005.490 1112.750 2006.580 1113.010 ;
        RECT 2011.470 1112.750 2012.560 1113.010 ;
        RECT 2017.450 1112.750 2018.540 1113.010 ;
        RECT 2023.430 1112.750 2024.520 1113.010 ;
        RECT 2029.410 1112.750 2030.500 1113.010 ;
        RECT 2035.390 1112.750 2036.480 1113.010 ;
        RECT 2041.370 1112.750 2042.460 1113.010 ;
        RECT 2047.350 1112.750 2048.440 1113.010 ;
        RECT 2053.330 1112.750 2054.420 1113.010 ;
        RECT 2059.310 1112.750 2060.400 1113.010 ;
        RECT 2065.290 1112.750 2066.380 1113.010 ;
        RECT 2071.270 1112.750 2072.360 1113.010 ;
        RECT 2077.250 1112.750 2078.340 1113.010 ;
        RECT 2083.230 1112.750 2084.320 1113.010 ;
        RECT 2090.080 1112.450 2090.340 1113.300 ;
      LAYER met2 ;
        RECT 2087.570 4986.345 2088.660 4986.665 ;
        RECT 835.260 4984.720 836.350 4985.040 ;
        RECT 841.240 4984.720 842.330 4985.040 ;
        RECT 847.220 4984.720 848.310 4985.040 ;
        RECT 835.550 4975.915 835.690 4984.720 ;
        RECT 836.090 4981.400 836.410 4982.250 ;
        RECT 836.170 4976.195 836.310 4981.400 ;
        RECT 841.530 4976.475 841.670 4984.720 ;
        RECT 842.070 4981.400 842.390 4982.250 ;
        RECT 842.150 4976.755 842.290 4981.400 ;
        RECT 847.510 4977.035 847.650 4984.720 ;
        RECT 2087.510 4983.025 2087.830 4983.875 ;
        RECT 848.050 4981.400 848.370 4982.250 ;
        RECT 848.130 4977.315 848.270 4981.400 ;
        RECT 835.550 4975.595 835.810 4975.915 ;
        RECT 836.170 4975.875 836.430 4976.195 ;
        RECT 841.530 4976.155 841.790 4976.475 ;
        RECT 842.150 4976.435 842.410 4976.755 ;
        RECT 847.510 4976.715 847.770 4977.035 ;
        RECT 848.130 4976.995 848.390 4977.315 ;
        RECT 835.550 4975.520 835.690 4975.595 ;
        RECT 836.170 4975.520 836.310 4975.875 ;
        RECT 841.530 4975.520 841.670 4976.155 ;
        RECT 842.150 4975.520 842.290 4976.435 ;
        RECT 847.510 4975.520 847.650 4976.715 ;
        RECT 848.130 4975.520 848.270 4976.995 ;
        RECT 2087.610 4976.405 2087.750 4983.025 ;
        RECT 2087.490 4976.085 2087.750 4976.405 ;
        RECT 2088.230 4976.125 2088.370 4986.345 ;
        RECT 3314.285 4985.675 3314.605 4986.525 ;
        RECT 3317.575 4985.935 3318.665 4986.255 ;
        RECT 3323.555 4985.935 3324.645 4986.255 ;
        RECT 3329.535 4985.935 3330.625 4986.255 ;
        RECT 3335.515 4985.935 3336.605 4986.255 ;
        RECT 3312.945 4982.875 3314.035 4983.195 ;
        RECT 3313.400 4976.385 3313.540 4982.875 ;
        RECT 2087.610 4975.645 2087.750 4976.085 ;
        RECT 2088.110 4975.805 2088.370 4976.125 ;
        RECT 3313.280 4976.065 3313.540 4976.385 ;
        RECT 3314.370 4976.105 3314.510 4985.675 ;
        RECT 3317.515 4982.615 3317.835 4983.465 ;
        RECT 3317.615 4976.405 3317.755 4982.615 ;
        RECT 2088.230 4975.645 2088.370 4975.805 ;
        RECT 3313.400 4973.965 3313.540 4976.065 ;
        RECT 3314.250 4975.785 3314.510 4976.105 ;
        RECT 3317.495 4976.085 3317.755 4976.405 ;
        RECT 3318.235 4976.125 3318.375 4985.935 ;
        RECT 3323.495 4982.615 3323.815 4983.465 ;
        RECT 3314.370 4973.965 3314.510 4975.785 ;
        RECT 3317.615 4973.965 3317.755 4976.085 ;
        RECT 3318.115 4975.805 3318.375 4976.125 ;
        RECT 3323.595 4975.845 3323.735 4982.615 ;
        RECT 3318.235 4973.965 3318.375 4975.805 ;
        RECT 3323.475 4975.525 3323.735 4975.845 ;
        RECT 3324.215 4975.565 3324.355 4985.935 ;
        RECT 3329.475 4982.615 3329.795 4983.465 ;
        RECT 3323.595 4973.965 3323.735 4975.525 ;
        RECT 3324.095 4975.245 3324.355 4975.565 ;
        RECT 3329.575 4975.285 3329.715 4982.615 ;
        RECT 3324.215 4973.965 3324.355 4975.245 ;
        RECT 3329.455 4974.965 3329.715 4975.285 ;
        RECT 3330.195 4975.005 3330.335 4985.935 ;
        RECT 3335.455 4982.615 3335.775 4983.465 ;
        RECT 3329.575 4973.965 3329.715 4974.965 ;
        RECT 3330.075 4974.685 3330.335 4975.005 ;
        RECT 3335.555 4974.725 3335.695 4982.615 ;
        RECT 3330.195 4973.965 3330.335 4974.685 ;
        RECT 3335.435 4974.405 3335.695 4974.725 ;
        RECT 3336.175 4974.445 3336.315 4985.935 ;
        RECT 3335.555 4973.965 3335.695 4974.405 ;
        RECT 3336.055 4974.125 3336.315 4974.445 ;
        RECT 3336.175 4973.965 3336.315 4974.125 ;
        RECT 202.740 4456.635 203.060 4457.090 ;
        RECT 212.305 4456.635 212.625 4456.755 ;
        RECT 202.740 4456.495 215.175 4456.635 ;
        RECT 202.740 4456.000 203.060 4456.495 ;
        RECT 199.410 4455.665 200.260 4455.750 ;
        RECT 212.585 4455.665 212.905 4455.785 ;
        RECT 199.410 4455.525 215.175 4455.665 ;
        RECT 199.410 4455.430 200.260 4455.525 ;
        RECT 199.680 4451.800 200.000 4452.460 ;
        RECT 202.470 4452.420 203.320 4452.520 ;
        RECT 212.285 4452.420 212.605 4452.540 ;
        RECT 202.470 4452.280 215.175 4452.420 ;
        RECT 202.470 4452.200 203.320 4452.280 ;
        RECT 212.565 4451.800 212.885 4451.920 ;
        RECT 199.680 4451.660 215.175 4451.800 ;
        RECT 199.680 4451.370 200.000 4451.660 ;
        RECT 202.740 4450.655 203.060 4451.110 ;
        RECT 202.740 4450.515 215.175 4450.655 ;
        RECT 202.740 4450.020 203.060 4450.515 ;
        RECT 212.865 4450.395 213.185 4450.515 ;
        RECT 199.410 4449.685 200.260 4449.770 ;
        RECT 213.145 4449.685 213.465 4449.805 ;
        RECT 199.410 4449.545 215.175 4449.685 ;
        RECT 199.410 4449.450 200.260 4449.545 ;
        RECT 199.680 4445.820 200.000 4446.480 ;
        RECT 202.470 4446.440 203.320 4446.540 ;
        RECT 212.845 4446.440 213.165 4446.560 ;
        RECT 202.470 4446.300 215.175 4446.440 ;
        RECT 202.470 4446.220 203.320 4446.300 ;
        RECT 213.125 4445.820 213.445 4445.940 ;
        RECT 199.680 4445.680 215.175 4445.820 ;
        RECT 199.680 4445.390 200.000 4445.680 ;
        RECT 202.740 4444.675 203.060 4445.130 ;
        RECT 213.425 4444.675 213.745 4444.795 ;
        RECT 202.740 4444.535 215.175 4444.675 ;
        RECT 202.740 4444.040 203.060 4444.535 ;
        RECT 199.410 4443.705 200.260 4443.790 ;
        RECT 213.705 4443.705 214.025 4443.825 ;
        RECT 199.410 4443.565 215.175 4443.705 ;
        RECT 199.410 4443.470 200.260 4443.565 ;
        RECT 199.680 4439.840 200.000 4440.500 ;
        RECT 202.470 4440.460 203.320 4440.560 ;
        RECT 213.405 4440.460 213.725 4440.580 ;
        RECT 202.470 4440.320 215.175 4440.460 ;
        RECT 202.470 4440.240 203.320 4440.320 ;
        RECT 213.685 4439.840 214.005 4439.960 ;
        RECT 199.680 4439.700 215.175 4439.840 ;
        RECT 199.680 4439.410 200.000 4439.700 ;
        RECT 199.680 4433.860 200.000 4434.520 ;
        RECT 202.470 4434.480 203.320 4434.580 ;
        RECT 213.965 4434.480 214.285 4434.600 ;
        RECT 202.470 4434.340 215.175 4434.480 ;
        RECT 202.470 4434.260 203.320 4434.340 ;
        RECT 214.245 4433.860 214.565 4433.980 ;
        RECT 199.680 4433.720 215.175 4433.860 ;
        RECT 199.680 4433.430 200.000 4433.720 ;
        RECT 199.680 4427.880 200.000 4428.540 ;
        RECT 202.470 4428.500 203.320 4428.600 ;
        RECT 214.525 4428.500 214.845 4428.620 ;
        RECT 202.470 4428.360 215.175 4428.500 ;
        RECT 202.470 4428.280 203.320 4428.360 ;
        RECT 214.805 4427.880 215.125 4428.000 ;
        RECT 199.680 4427.740 215.175 4427.880 ;
        RECT 199.680 4427.450 200.000 4427.740 ;
        RECT 3384.610 3571.835 3384.930 3572.290 ;
        RECT 3375.090 3571.695 3384.930 3571.835 ;
        RECT 3375.430 3571.575 3375.750 3571.695 ;
        RECT 3384.610 3571.200 3384.930 3571.695 ;
        RECT 3375.150 3570.865 3375.470 3570.985 ;
        RECT 3387.410 3570.865 3388.260 3570.950 ;
        RECT 3375.090 3570.725 3388.260 3570.865 ;
        RECT 3387.410 3570.630 3388.260 3570.725 ;
        RECT 3375.450 3567.620 3375.770 3567.740 ;
        RECT 3384.350 3567.620 3385.200 3567.720 ;
        RECT 3375.205 3567.480 3385.200 3567.620 ;
        RECT 3384.350 3567.400 3385.200 3567.480 ;
        RECT 3375.170 3567.000 3375.490 3567.120 ;
        RECT 3387.670 3567.000 3387.990 3567.660 ;
        RECT 3375.170 3566.860 3387.990 3567.000 ;
        RECT 3387.670 3566.570 3387.990 3566.860 ;
        RECT 3374.870 3565.855 3375.190 3565.975 ;
        RECT 3384.610 3565.855 3384.930 3566.310 ;
        RECT 3372.210 3565.715 3384.930 3565.855 ;
        RECT 3384.610 3565.220 3384.930 3565.715 ;
        RECT 3374.590 3564.885 3374.910 3565.005 ;
        RECT 3387.410 3564.885 3388.260 3564.970 ;
        RECT 3372.210 3564.745 3388.260 3564.885 ;
        RECT 3387.410 3564.650 3388.260 3564.745 ;
        RECT 3374.890 3561.640 3375.210 3561.760 ;
        RECT 3384.350 3561.640 3385.200 3561.740 ;
        RECT 3372.210 3561.500 3385.200 3561.640 ;
        RECT 3384.350 3561.420 3385.200 3561.500 ;
        RECT 3374.610 3561.020 3374.930 3561.140 ;
        RECT 3387.670 3561.020 3387.990 3561.680 ;
        RECT 3372.210 3560.880 3387.990 3561.020 ;
        RECT 3387.670 3560.590 3387.990 3560.880 ;
        RECT 3374.310 3559.875 3374.630 3559.995 ;
        RECT 3384.610 3559.875 3384.930 3560.330 ;
        RECT 3372.210 3559.735 3384.930 3559.875 ;
        RECT 3384.610 3559.240 3384.930 3559.735 ;
        RECT 3374.030 3558.905 3374.350 3559.025 ;
        RECT 3387.410 3558.905 3388.260 3558.990 ;
        RECT 3372.210 3558.765 3388.260 3558.905 ;
        RECT 3387.410 3558.670 3388.260 3558.765 ;
        RECT 3374.330 3555.660 3374.650 3555.780 ;
        RECT 3384.350 3555.660 3385.200 3555.760 ;
        RECT 3372.210 3555.520 3385.200 3555.660 ;
        RECT 3384.350 3555.440 3385.200 3555.520 ;
        RECT 3374.050 3555.040 3374.370 3555.160 ;
        RECT 3387.670 3555.040 3387.990 3555.700 ;
        RECT 3372.210 3554.900 3387.990 3555.040 ;
        RECT 3387.670 3554.610 3387.990 3554.900 ;
        RECT 3373.750 3553.895 3374.070 3554.015 ;
        RECT 3384.610 3553.895 3384.930 3554.350 ;
        RECT 3372.210 3553.755 3384.930 3553.895 ;
        RECT 3384.610 3553.260 3384.930 3553.755 ;
        RECT 3373.470 3552.925 3373.790 3553.045 ;
        RECT 3387.410 3552.925 3388.260 3553.010 ;
        RECT 3372.210 3552.785 3388.260 3552.925 ;
        RECT 3387.410 3552.690 3388.260 3552.785 ;
        RECT 3373.770 3549.680 3374.090 3549.800 ;
        RECT 3384.350 3549.680 3385.200 3549.780 ;
        RECT 3372.210 3549.540 3385.200 3549.680 ;
        RECT 3384.350 3549.460 3385.200 3549.540 ;
        RECT 3373.490 3549.060 3373.810 3549.180 ;
        RECT 3387.670 3549.060 3387.990 3549.720 ;
        RECT 3372.210 3548.920 3387.990 3549.060 ;
        RECT 3387.670 3548.630 3387.990 3548.920 ;
        RECT 3373.210 3543.700 3373.530 3543.820 ;
        RECT 3384.350 3543.700 3385.200 3543.800 ;
        RECT 3372.210 3543.560 3385.200 3543.700 ;
        RECT 3384.350 3543.480 3385.200 3543.560 ;
        RECT 3372.930 3543.080 3373.250 3543.200 ;
        RECT 3387.670 3543.080 3387.990 3543.740 ;
        RECT 3372.210 3542.940 3387.990 3543.080 ;
        RECT 3387.670 3542.650 3387.990 3542.940 ;
        RECT 3372.650 3537.720 3372.970 3537.840 ;
        RECT 3384.350 3537.720 3385.200 3537.820 ;
        RECT 3372.210 3537.580 3385.200 3537.720 ;
        RECT 3384.350 3537.500 3385.200 3537.580 ;
        RECT 3372.370 3537.100 3372.690 3537.220 ;
        RECT 3387.670 3537.100 3387.990 3537.760 ;
        RECT 3372.210 3536.960 3387.990 3537.100 ;
        RECT 3387.670 3536.670 3387.990 3536.960 ;
        RECT 202.865 3053.405 203.185 3053.860 ;
        RECT 212.165 3053.405 212.485 3053.525 ;
        RECT 202.865 3053.265 218.400 3053.405 ;
        RECT 202.865 3052.770 203.185 3053.265 ;
        RECT 199.535 3052.435 200.385 3052.520 ;
        RECT 212.445 3052.435 212.765 3052.555 ;
        RECT 199.535 3052.295 218.400 3052.435 ;
        RECT 199.535 3052.200 200.385 3052.295 ;
        RECT 199.805 3048.570 200.125 3049.230 ;
        RECT 202.595 3049.190 203.445 3049.290 ;
        RECT 212.145 3049.190 212.465 3049.310 ;
        RECT 202.595 3049.050 218.400 3049.190 ;
        RECT 202.595 3048.970 203.445 3049.050 ;
        RECT 212.425 3048.570 212.745 3048.690 ;
        RECT 199.805 3048.430 218.400 3048.570 ;
        RECT 199.805 3048.140 200.125 3048.430 ;
        RECT 202.865 3047.425 203.185 3047.880 ;
        RECT 202.865 3047.285 218.400 3047.425 ;
        RECT 202.865 3046.790 203.185 3047.285 ;
        RECT 212.725 3047.165 213.045 3047.285 ;
        RECT 199.535 3046.455 200.385 3046.540 ;
        RECT 213.005 3046.455 213.325 3046.575 ;
        RECT 199.535 3046.315 218.400 3046.455 ;
        RECT 199.535 3046.220 200.385 3046.315 ;
        RECT 199.805 3042.590 200.125 3043.250 ;
        RECT 202.595 3043.210 203.445 3043.310 ;
        RECT 212.705 3043.210 213.025 3043.330 ;
        RECT 202.595 3043.070 218.400 3043.210 ;
        RECT 202.595 3042.990 203.445 3043.070 ;
        RECT 212.985 3042.590 213.305 3042.710 ;
        RECT 199.805 3042.450 218.400 3042.590 ;
        RECT 199.805 3042.160 200.125 3042.450 ;
        RECT 202.865 3041.445 203.185 3041.900 ;
        RECT 213.285 3041.445 213.605 3041.565 ;
        RECT 202.865 3041.305 218.400 3041.445 ;
        RECT 202.865 3040.810 203.185 3041.305 ;
        RECT 199.535 3040.475 200.385 3040.560 ;
        RECT 213.565 3040.475 213.885 3040.595 ;
        RECT 199.535 3040.335 218.400 3040.475 ;
        RECT 199.535 3040.240 200.385 3040.335 ;
        RECT 199.805 3036.610 200.125 3037.270 ;
        RECT 202.595 3037.230 203.445 3037.330 ;
        RECT 213.265 3037.230 213.585 3037.350 ;
        RECT 202.595 3037.090 218.400 3037.230 ;
        RECT 202.595 3037.010 203.445 3037.090 ;
        RECT 213.545 3036.610 213.865 3036.730 ;
        RECT 199.805 3036.470 218.400 3036.610 ;
        RECT 199.805 3036.180 200.125 3036.470 ;
        RECT 202.865 3035.465 203.185 3035.920 ;
        RECT 202.865 3035.325 218.400 3035.465 ;
        RECT 202.865 3034.830 203.185 3035.325 ;
        RECT 213.845 3035.205 214.165 3035.325 ;
        RECT 199.535 3034.495 200.385 3034.580 ;
        RECT 214.125 3034.495 214.445 3034.615 ;
        RECT 199.535 3034.355 218.400 3034.495 ;
        RECT 199.535 3034.260 200.385 3034.355 ;
        RECT 199.805 3030.630 200.125 3031.290 ;
        RECT 202.595 3031.250 203.445 3031.350 ;
        RECT 213.825 3031.250 214.145 3031.370 ;
        RECT 202.595 3031.110 218.400 3031.250 ;
        RECT 202.595 3031.030 203.445 3031.110 ;
        RECT 214.105 3030.630 214.425 3030.750 ;
        RECT 199.805 3030.490 218.400 3030.630 ;
        RECT 199.805 3030.200 200.125 3030.490 ;
        RECT 202.865 3029.485 203.185 3029.940 ;
        RECT 214.405 3029.485 214.725 3029.605 ;
        RECT 202.865 3029.345 218.400 3029.485 ;
        RECT 202.865 3028.850 203.185 3029.345 ;
        RECT 199.535 3028.515 200.385 3028.600 ;
        RECT 214.685 3028.515 215.005 3028.635 ;
        RECT 199.535 3028.375 218.400 3028.515 ;
        RECT 199.535 3028.280 200.385 3028.375 ;
        RECT 199.805 3024.650 200.125 3025.310 ;
        RECT 202.595 3025.270 203.445 3025.370 ;
        RECT 214.385 3025.270 214.705 3025.390 ;
        RECT 202.595 3025.130 218.400 3025.270 ;
        RECT 202.595 3025.050 203.445 3025.130 ;
        RECT 214.665 3024.650 214.985 3024.770 ;
        RECT 199.805 3024.510 218.400 3024.650 ;
        RECT 199.805 3024.220 200.125 3024.510 ;
        RECT 199.805 3018.670 200.125 3019.330 ;
        RECT 202.595 3019.290 203.445 3019.390 ;
        RECT 214.945 3019.290 215.265 3019.410 ;
        RECT 202.595 3019.150 218.400 3019.290 ;
        RECT 202.595 3019.070 203.445 3019.150 ;
        RECT 215.225 3018.670 215.545 3018.790 ;
        RECT 199.805 3018.530 218.400 3018.670 ;
        RECT 199.805 3018.240 200.125 3018.530 ;
        RECT 199.805 3012.690 200.125 3013.350 ;
        RECT 202.595 3013.310 203.445 3013.410 ;
        RECT 215.505 3013.310 215.825 3013.430 ;
        RECT 202.595 3013.170 218.400 3013.310 ;
        RECT 202.595 3013.090 203.445 3013.170 ;
        RECT 215.785 3012.690 216.105 3012.810 ;
        RECT 199.805 3012.550 218.400 3012.690 ;
        RECT 199.805 3012.260 200.125 3012.550 ;
        RECT 199.805 3006.710 200.125 3007.370 ;
        RECT 202.595 3007.330 203.445 3007.430 ;
        RECT 216.065 3007.330 216.385 3007.450 ;
        RECT 202.595 3007.190 218.400 3007.330 ;
        RECT 202.595 3007.110 203.445 3007.190 ;
        RECT 216.345 3006.710 216.665 3006.830 ;
        RECT 199.805 3006.570 218.400 3006.710 ;
        RECT 199.805 3006.280 200.125 3006.570 ;
        RECT 199.805 3000.730 200.125 3001.390 ;
        RECT 202.595 3001.350 203.445 3001.450 ;
        RECT 216.625 3001.350 216.945 3001.470 ;
        RECT 202.595 3001.210 218.400 3001.350 ;
        RECT 202.595 3001.130 203.445 3001.210 ;
        RECT 216.905 3000.730 217.225 3000.850 ;
        RECT 199.805 3000.590 218.400 3000.730 ;
        RECT 199.805 3000.300 200.125 3000.590 ;
        RECT 199.805 2994.750 200.125 2995.410 ;
        RECT 202.595 2995.370 203.445 2995.470 ;
        RECT 217.185 2995.370 217.505 2995.490 ;
        RECT 202.595 2995.230 218.400 2995.370 ;
        RECT 202.595 2995.150 203.445 2995.230 ;
        RECT 217.465 2994.750 217.785 2994.870 ;
        RECT 199.805 2994.610 218.400 2994.750 ;
        RECT 199.805 2994.320 200.125 2994.610 ;
        RECT 199.805 2988.770 200.125 2989.430 ;
        RECT 202.595 2989.390 203.445 2989.490 ;
        RECT 217.745 2989.390 218.065 2989.510 ;
        RECT 202.595 2989.250 218.400 2989.390 ;
        RECT 202.595 2989.170 203.445 2989.250 ;
        RECT 218.025 2988.770 218.345 2988.890 ;
        RECT 199.805 2988.630 218.400 2988.770 ;
        RECT 199.805 2988.340 200.125 2988.630 ;
        RECT 3375.430 2267.715 3375.750 2267.835 ;
        RECT 3384.610 2267.715 3384.930 2268.170 ;
        RECT 3368.850 2267.575 3384.930 2267.715 ;
        RECT 3384.610 2267.080 3384.930 2267.575 ;
        RECT 3375.150 2266.745 3375.470 2266.865 ;
        RECT 3387.410 2266.745 3388.260 2266.830 ;
        RECT 3368.850 2266.605 3388.260 2266.745 ;
        RECT 3387.410 2266.510 3388.260 2266.605 ;
        RECT 3384.610 2261.735 3384.930 2262.190 ;
        RECT 3368.850 2261.595 3384.930 2261.735 ;
        RECT 3374.870 2261.475 3375.190 2261.595 ;
        RECT 3384.610 2261.100 3384.930 2261.595 ;
        RECT 3374.590 2260.765 3374.910 2260.885 ;
        RECT 3387.410 2260.765 3388.260 2260.850 ;
        RECT 3368.850 2260.625 3388.260 2260.765 ;
        RECT 3387.410 2260.530 3388.260 2260.625 ;
        RECT 3374.310 2255.755 3374.630 2255.875 ;
        RECT 3384.610 2255.755 3384.930 2256.210 ;
        RECT 3368.850 2255.615 3384.930 2255.755 ;
        RECT 3384.610 2255.120 3384.930 2255.615 ;
        RECT 3374.030 2254.785 3374.350 2254.905 ;
        RECT 3387.410 2254.785 3388.260 2254.870 ;
        RECT 3368.850 2254.645 3388.260 2254.785 ;
        RECT 3387.410 2254.550 3388.260 2254.645 ;
        RECT 3384.610 2249.775 3384.930 2250.230 ;
        RECT 3368.850 2249.635 3384.930 2249.775 ;
        RECT 3373.750 2249.515 3374.070 2249.635 ;
        RECT 3384.610 2249.140 3384.930 2249.635 ;
        RECT 3373.470 2248.805 3373.790 2248.925 ;
        RECT 3387.410 2248.805 3388.260 2248.890 ;
        RECT 3368.850 2248.665 3388.260 2248.805 ;
        RECT 3387.410 2248.570 3388.260 2248.665 ;
        RECT 3373.190 2243.795 3373.510 2243.915 ;
        RECT 3384.610 2243.795 3384.930 2244.250 ;
        RECT 3368.850 2243.655 3384.930 2243.795 ;
        RECT 3384.610 2243.160 3384.930 2243.655 ;
        RECT 3372.910 2242.825 3373.230 2242.945 ;
        RECT 3387.410 2242.825 3388.260 2242.910 ;
        RECT 3368.850 2242.685 3388.260 2242.825 ;
        RECT 3387.410 2242.590 3388.260 2242.685 ;
        RECT 3372.630 2237.815 3372.950 2237.935 ;
        RECT 3384.610 2237.815 3384.930 2238.270 ;
        RECT 3368.850 2237.675 3384.930 2237.815 ;
        RECT 3384.610 2237.180 3384.930 2237.675 ;
        RECT 3372.350 2236.845 3372.670 2236.965 ;
        RECT 3387.410 2236.845 3388.260 2236.930 ;
        RECT 3368.850 2236.705 3388.260 2236.845 ;
        RECT 3387.410 2236.610 3388.260 2236.705 ;
        RECT 202.975 1762.500 203.295 1762.955 ;
        RECT 212.025 1762.500 212.345 1762.620 ;
        RECT 202.975 1762.360 220.540 1762.500 ;
        RECT 202.975 1761.865 203.295 1762.360 ;
        RECT 199.645 1761.530 200.495 1761.615 ;
        RECT 212.305 1761.530 212.625 1761.650 ;
        RECT 199.645 1761.390 220.540 1761.530 ;
        RECT 199.645 1761.295 200.495 1761.390 ;
        RECT 199.915 1757.665 200.235 1758.325 ;
        RECT 202.705 1758.285 203.555 1758.385 ;
        RECT 212.005 1758.285 212.325 1758.405 ;
        RECT 202.705 1758.145 220.540 1758.285 ;
        RECT 202.705 1758.065 203.555 1758.145 ;
        RECT 212.285 1757.665 212.605 1757.785 ;
        RECT 199.915 1757.525 220.540 1757.665 ;
        RECT 199.915 1757.235 200.235 1757.525 ;
        RECT 202.975 1756.520 203.295 1756.975 ;
        RECT 202.975 1756.380 220.540 1756.520 ;
        RECT 202.975 1755.885 203.295 1756.380 ;
        RECT 212.585 1756.260 212.905 1756.380 ;
        RECT 199.645 1755.550 200.495 1755.635 ;
        RECT 212.865 1755.550 213.185 1755.670 ;
        RECT 199.645 1755.410 220.540 1755.550 ;
        RECT 199.645 1755.315 200.495 1755.410 ;
        RECT 199.915 1751.685 200.235 1752.345 ;
        RECT 202.705 1752.305 203.555 1752.405 ;
        RECT 212.565 1752.305 212.885 1752.425 ;
        RECT 202.705 1752.165 220.540 1752.305 ;
        RECT 202.705 1752.085 203.555 1752.165 ;
        RECT 212.845 1751.685 213.165 1751.805 ;
        RECT 199.915 1751.545 220.540 1751.685 ;
        RECT 199.915 1751.255 200.235 1751.545 ;
        RECT 202.975 1750.540 203.295 1750.995 ;
        RECT 213.145 1750.540 213.465 1750.660 ;
        RECT 202.975 1750.400 220.540 1750.540 ;
        RECT 202.975 1749.905 203.295 1750.400 ;
        RECT 199.645 1749.570 200.495 1749.655 ;
        RECT 213.425 1749.570 213.745 1749.690 ;
        RECT 199.645 1749.430 220.540 1749.570 ;
        RECT 199.645 1749.335 200.495 1749.430 ;
        RECT 199.915 1745.705 200.235 1746.365 ;
        RECT 202.705 1746.325 203.555 1746.425 ;
        RECT 213.125 1746.325 213.445 1746.445 ;
        RECT 202.705 1746.185 220.540 1746.325 ;
        RECT 202.705 1746.105 203.555 1746.185 ;
        RECT 213.405 1745.705 213.725 1745.825 ;
        RECT 199.915 1745.565 220.540 1745.705 ;
        RECT 199.915 1745.275 200.235 1745.565 ;
        RECT 202.975 1744.560 203.295 1745.015 ;
        RECT 202.975 1744.420 220.540 1744.560 ;
        RECT 202.975 1743.925 203.295 1744.420 ;
        RECT 213.705 1744.300 214.025 1744.420 ;
        RECT 199.645 1743.590 200.495 1743.675 ;
        RECT 213.985 1743.590 214.305 1743.710 ;
        RECT 199.645 1743.450 220.540 1743.590 ;
        RECT 199.645 1743.355 200.495 1743.450 ;
        RECT 199.915 1739.725 200.235 1740.385 ;
        RECT 202.705 1740.345 203.555 1740.445 ;
        RECT 213.685 1740.345 214.005 1740.465 ;
        RECT 202.705 1740.205 220.540 1740.345 ;
        RECT 202.705 1740.125 203.555 1740.205 ;
        RECT 213.965 1739.725 214.285 1739.845 ;
        RECT 199.915 1739.585 220.540 1739.725 ;
        RECT 199.915 1739.295 200.235 1739.585 ;
        RECT 202.975 1738.580 203.295 1739.035 ;
        RECT 214.265 1738.580 214.585 1738.700 ;
        RECT 202.975 1738.440 220.540 1738.580 ;
        RECT 202.975 1737.945 203.295 1738.440 ;
        RECT 199.645 1737.610 200.495 1737.695 ;
        RECT 214.545 1737.610 214.865 1737.730 ;
        RECT 199.645 1737.470 220.540 1737.610 ;
        RECT 199.645 1737.375 200.495 1737.470 ;
        RECT 199.915 1733.745 200.235 1734.405 ;
        RECT 202.705 1734.365 203.555 1734.465 ;
        RECT 214.245 1734.365 214.565 1734.485 ;
        RECT 202.705 1734.225 220.540 1734.365 ;
        RECT 202.705 1734.145 203.555 1734.225 ;
        RECT 214.525 1733.745 214.845 1733.865 ;
        RECT 199.915 1733.605 220.540 1733.745 ;
        RECT 199.915 1733.315 200.235 1733.605 ;
        RECT 202.975 1732.600 203.295 1733.055 ;
        RECT 214.825 1732.600 215.145 1732.720 ;
        RECT 202.975 1732.460 220.540 1732.600 ;
        RECT 202.975 1731.965 203.295 1732.460 ;
        RECT 199.645 1731.630 200.495 1731.715 ;
        RECT 215.105 1731.630 215.425 1731.750 ;
        RECT 199.645 1731.490 220.540 1731.630 ;
        RECT 199.645 1731.395 200.495 1731.490 ;
        RECT 199.915 1727.765 200.235 1728.425 ;
        RECT 202.705 1728.385 203.555 1728.485 ;
        RECT 214.805 1728.385 215.125 1728.505 ;
        RECT 202.705 1728.245 220.540 1728.385 ;
        RECT 202.705 1728.165 203.555 1728.245 ;
        RECT 215.085 1727.765 215.405 1727.885 ;
        RECT 199.915 1727.625 220.540 1727.765 ;
        RECT 199.915 1727.335 200.235 1727.625 ;
        RECT 202.975 1726.620 203.295 1727.075 ;
        RECT 215.385 1726.620 215.705 1726.740 ;
        RECT 202.975 1726.480 220.540 1726.620 ;
        RECT 202.975 1725.985 203.295 1726.480 ;
        RECT 199.645 1725.650 200.495 1725.735 ;
        RECT 215.665 1725.650 215.985 1725.770 ;
        RECT 199.645 1725.510 220.540 1725.650 ;
        RECT 199.645 1725.415 200.495 1725.510 ;
        RECT 199.915 1721.785 200.235 1722.445 ;
        RECT 202.705 1722.405 203.555 1722.505 ;
        RECT 215.365 1722.405 215.685 1722.525 ;
        RECT 202.705 1722.265 220.540 1722.405 ;
        RECT 202.705 1722.185 203.555 1722.265 ;
        RECT 215.645 1721.785 215.965 1721.905 ;
        RECT 199.915 1721.645 220.540 1721.785 ;
        RECT 199.915 1721.355 200.235 1721.645 ;
        RECT 202.975 1720.640 203.295 1721.095 ;
        RECT 215.945 1720.640 216.265 1720.760 ;
        RECT 202.975 1720.500 220.540 1720.640 ;
        RECT 202.975 1720.005 203.295 1720.500 ;
        RECT 199.645 1719.670 200.495 1719.755 ;
        RECT 216.225 1719.670 216.545 1719.790 ;
        RECT 199.645 1719.530 220.540 1719.670 ;
        RECT 199.645 1719.435 200.495 1719.530 ;
        RECT 199.915 1715.805 200.235 1716.465 ;
        RECT 202.705 1716.425 203.555 1716.525 ;
        RECT 215.925 1716.425 216.245 1716.545 ;
        RECT 202.705 1716.285 220.540 1716.425 ;
        RECT 202.705 1716.205 203.555 1716.285 ;
        RECT 216.205 1715.805 216.525 1715.925 ;
        RECT 199.915 1715.665 220.540 1715.805 ;
        RECT 199.915 1715.375 200.235 1715.665 ;
        RECT 202.975 1714.660 203.295 1715.115 ;
        RECT 216.505 1714.660 216.825 1714.780 ;
        RECT 202.975 1714.520 220.540 1714.660 ;
        RECT 202.975 1714.025 203.295 1714.520 ;
        RECT 199.645 1713.690 200.495 1713.775 ;
        RECT 216.785 1713.690 217.105 1713.810 ;
        RECT 199.645 1713.550 220.540 1713.690 ;
        RECT 199.645 1713.455 200.495 1713.550 ;
        RECT 199.915 1709.825 200.235 1710.485 ;
        RECT 202.705 1710.445 203.555 1710.545 ;
        RECT 216.485 1710.445 216.805 1710.565 ;
        RECT 202.705 1710.305 220.540 1710.445 ;
        RECT 202.705 1710.225 203.555 1710.305 ;
        RECT 216.765 1709.825 217.085 1709.945 ;
        RECT 199.915 1709.685 220.540 1709.825 ;
        RECT 199.915 1709.395 200.235 1709.685 ;
        RECT 202.975 1708.680 203.295 1709.135 ;
        RECT 217.065 1708.680 217.385 1708.800 ;
        RECT 202.975 1708.540 220.540 1708.680 ;
        RECT 202.975 1708.045 203.295 1708.540 ;
        RECT 199.645 1707.710 200.495 1707.795 ;
        RECT 217.345 1707.710 217.665 1707.830 ;
        RECT 199.645 1707.570 220.540 1707.710 ;
        RECT 199.645 1707.475 200.495 1707.570 ;
        RECT 199.915 1703.845 200.235 1704.505 ;
        RECT 202.705 1704.465 203.555 1704.565 ;
        RECT 217.045 1704.465 217.365 1704.585 ;
        RECT 202.705 1704.325 220.540 1704.465 ;
        RECT 202.705 1704.245 203.555 1704.325 ;
        RECT 217.325 1703.845 217.645 1703.965 ;
        RECT 199.915 1703.705 220.540 1703.845 ;
        RECT 199.915 1703.415 200.235 1703.705 ;
        RECT 202.975 1702.700 203.295 1703.155 ;
        RECT 217.625 1702.700 217.945 1702.820 ;
        RECT 202.975 1702.560 220.540 1702.700 ;
        RECT 202.975 1702.065 203.295 1702.560 ;
        RECT 199.645 1701.730 200.495 1701.815 ;
        RECT 217.905 1701.730 218.225 1701.850 ;
        RECT 199.645 1701.590 220.540 1701.730 ;
        RECT 199.645 1701.495 200.495 1701.590 ;
        RECT 199.915 1697.865 200.235 1698.525 ;
        RECT 202.705 1698.485 203.555 1698.585 ;
        RECT 217.605 1698.485 217.925 1698.605 ;
        RECT 202.705 1698.345 220.540 1698.485 ;
        RECT 202.705 1698.265 203.555 1698.345 ;
        RECT 217.885 1697.865 218.205 1697.985 ;
        RECT 199.915 1697.725 220.540 1697.865 ;
        RECT 199.915 1697.435 200.235 1697.725 ;
        RECT 199.915 1691.885 200.235 1692.545 ;
        RECT 202.705 1692.505 203.555 1692.605 ;
        RECT 218.165 1692.505 218.485 1692.625 ;
        RECT 202.705 1692.365 220.540 1692.505 ;
        RECT 202.705 1692.285 203.555 1692.365 ;
        RECT 218.445 1691.885 218.765 1692.005 ;
        RECT 199.915 1691.745 220.540 1691.885 ;
        RECT 199.915 1691.455 200.235 1691.745 ;
        RECT 199.915 1685.905 200.235 1686.565 ;
        RECT 202.705 1686.525 203.555 1686.625 ;
        RECT 218.725 1686.525 219.045 1686.645 ;
        RECT 202.705 1686.385 220.540 1686.525 ;
        RECT 202.705 1686.305 203.555 1686.385 ;
        RECT 219.005 1685.905 219.325 1686.025 ;
        RECT 199.915 1685.765 220.540 1685.905 ;
        RECT 199.915 1685.475 200.235 1685.765 ;
        RECT 199.915 1679.925 200.235 1680.585 ;
        RECT 202.705 1680.545 203.555 1680.645 ;
        RECT 219.285 1680.545 219.605 1680.665 ;
        RECT 202.705 1680.405 220.540 1680.545 ;
        RECT 202.705 1680.325 203.555 1680.405 ;
        RECT 219.565 1679.925 219.885 1680.045 ;
        RECT 199.915 1679.785 220.540 1679.925 ;
        RECT 199.915 1679.495 200.235 1679.785 ;
        RECT 199.915 1673.945 200.235 1674.605 ;
        RECT 202.705 1674.565 203.555 1674.665 ;
        RECT 219.845 1674.565 220.165 1674.685 ;
        RECT 202.705 1674.425 220.540 1674.565 ;
        RECT 202.705 1674.345 203.555 1674.425 ;
        RECT 220.125 1673.945 220.445 1674.065 ;
        RECT 199.915 1673.805 220.540 1673.945 ;
        RECT 199.915 1673.515 200.235 1673.805 ;
        RECT 1970.520 1129.670 1970.660 1129.765 ;
        RECT 670.520 1129.530 670.660 1129.625 ;
        RECT 674.735 1129.550 674.875 1129.625 ;
        RECT 670.520 1129.210 670.780 1129.530 ;
        RECT 674.735 1129.230 674.995 1129.550 ;
        RECT 675.880 1129.250 676.020 1129.625 ;
        RECT 670.520 1116.360 670.660 1129.210 ;
        RECT 670.440 1115.510 670.760 1116.360 ;
        RECT 674.735 1116.100 674.875 1129.230 ;
        RECT 675.880 1128.930 676.140 1129.250 ;
        RECT 676.500 1128.970 676.640 1129.625 ;
        RECT 679.745 1129.270 679.885 1129.625 ;
        RECT 674.240 1115.780 675.330 1116.100 ;
        RECT 675.880 1113.040 676.020 1128.930 ;
        RECT 676.500 1128.650 676.760 1128.970 ;
        RECT 679.745 1128.950 680.005 1129.270 ;
        RECT 680.715 1128.990 680.855 1129.625 ;
        RECT 676.500 1116.360 676.640 1128.650 ;
        RECT 676.420 1115.510 676.740 1116.360 ;
        RECT 679.745 1113.300 679.885 1128.950 ;
        RECT 680.715 1128.670 680.975 1128.990 ;
        RECT 681.860 1128.690 682.000 1129.625 ;
        RECT 680.715 1116.100 680.855 1128.670 ;
        RECT 681.860 1128.370 682.120 1128.690 ;
        RECT 682.480 1128.410 682.620 1129.625 ;
        RECT 685.725 1128.710 685.865 1129.625 ;
        RECT 680.220 1115.780 681.310 1116.100 ;
        RECT 675.590 1112.720 676.680 1113.040 ;
        RECT 679.650 1112.450 679.970 1113.300 ;
        RECT 681.860 1113.040 682.000 1128.370 ;
        RECT 682.480 1128.090 682.740 1128.410 ;
        RECT 685.725 1128.390 685.985 1128.710 ;
        RECT 686.695 1128.430 686.835 1129.625 ;
        RECT 682.480 1116.360 682.620 1128.090 ;
        RECT 682.400 1115.510 682.720 1116.360 ;
        RECT 685.725 1113.300 685.865 1128.390 ;
        RECT 686.695 1128.110 686.955 1128.430 ;
        RECT 687.840 1128.130 687.980 1129.625 ;
        RECT 686.695 1116.100 686.835 1128.110 ;
        RECT 687.840 1127.810 688.100 1128.130 ;
        RECT 688.460 1127.850 688.600 1129.625 ;
        RECT 691.705 1128.150 691.845 1129.625 ;
        RECT 686.200 1115.780 687.290 1116.100 ;
        RECT 681.570 1112.720 682.660 1113.040 ;
        RECT 685.630 1112.450 685.950 1113.300 ;
        RECT 687.840 1113.040 687.980 1127.810 ;
        RECT 688.460 1127.530 688.720 1127.850 ;
        RECT 691.705 1127.830 691.965 1128.150 ;
        RECT 692.675 1127.870 692.815 1129.625 ;
        RECT 688.460 1116.360 688.600 1127.530 ;
        RECT 688.380 1115.510 688.700 1116.360 ;
        RECT 691.705 1113.300 691.845 1127.830 ;
        RECT 692.675 1127.550 692.935 1127.870 ;
        RECT 693.820 1127.570 693.960 1129.625 ;
        RECT 692.675 1116.100 692.815 1127.550 ;
        RECT 693.820 1127.250 694.080 1127.570 ;
        RECT 694.440 1127.290 694.580 1129.625 ;
        RECT 697.685 1127.590 697.825 1129.625 ;
        RECT 692.180 1115.780 693.270 1116.100 ;
        RECT 687.550 1112.720 688.640 1113.040 ;
        RECT 691.610 1112.450 691.930 1113.300 ;
        RECT 693.820 1113.040 693.960 1127.250 ;
        RECT 694.440 1126.970 694.700 1127.290 ;
        RECT 697.685 1127.270 697.945 1127.590 ;
        RECT 698.655 1127.310 698.795 1129.625 ;
        RECT 694.440 1116.360 694.580 1126.970 ;
        RECT 694.360 1115.510 694.680 1116.360 ;
        RECT 697.685 1113.300 697.825 1127.270 ;
        RECT 698.655 1126.990 698.915 1127.310 ;
        RECT 699.800 1127.010 699.940 1129.625 ;
        RECT 698.655 1116.100 698.795 1126.990 ;
        RECT 699.800 1126.690 700.060 1127.010 ;
        RECT 700.420 1126.730 700.560 1129.625 ;
        RECT 703.665 1127.030 703.805 1129.625 ;
        RECT 698.160 1115.780 699.250 1116.100 ;
        RECT 693.530 1112.720 694.620 1113.040 ;
        RECT 697.590 1112.450 697.910 1113.300 ;
        RECT 699.800 1113.040 699.940 1126.690 ;
        RECT 700.420 1126.410 700.680 1126.730 ;
        RECT 703.665 1126.710 703.925 1127.030 ;
        RECT 704.635 1126.750 704.775 1129.625 ;
        RECT 700.420 1116.360 700.560 1126.410 ;
        RECT 700.340 1115.510 700.660 1116.360 ;
        RECT 703.665 1113.300 703.805 1126.710 ;
        RECT 704.515 1126.430 704.775 1126.750 ;
        RECT 704.635 1116.100 704.775 1126.430 ;
        RECT 705.780 1126.450 705.920 1129.625 ;
        RECT 705.780 1126.130 706.040 1126.450 ;
        RECT 706.400 1126.170 706.540 1129.625 ;
        RECT 709.645 1126.470 709.785 1129.625 ;
        RECT 704.140 1115.780 705.230 1116.100 ;
        RECT 699.510 1112.720 700.600 1113.040 ;
        RECT 703.570 1112.450 703.890 1113.300 ;
        RECT 705.780 1113.040 705.920 1126.130 ;
        RECT 706.400 1125.850 706.660 1126.170 ;
        RECT 709.645 1126.150 709.905 1126.470 ;
        RECT 710.615 1126.190 710.755 1129.625 ;
        RECT 706.400 1116.360 706.540 1125.850 ;
        RECT 706.320 1115.510 706.640 1116.360 ;
        RECT 709.645 1113.300 709.785 1126.150 ;
        RECT 710.615 1125.870 710.875 1126.190 ;
        RECT 711.760 1125.890 711.900 1129.625 ;
        RECT 710.615 1116.100 710.755 1125.870 ;
        RECT 711.760 1125.570 712.020 1125.890 ;
        RECT 712.380 1125.610 712.520 1129.625 ;
        RECT 715.625 1125.910 715.765 1129.625 ;
        RECT 710.120 1115.780 711.210 1116.100 ;
        RECT 705.490 1112.720 706.580 1113.040 ;
        RECT 709.550 1112.450 709.870 1113.300 ;
        RECT 711.760 1113.040 711.900 1125.570 ;
        RECT 712.380 1125.290 712.640 1125.610 ;
        RECT 715.625 1125.590 715.885 1125.910 ;
        RECT 716.595 1125.630 716.735 1129.625 ;
        RECT 712.380 1116.360 712.520 1125.290 ;
        RECT 712.300 1115.510 712.620 1116.360 ;
        RECT 715.625 1113.300 715.765 1125.590 ;
        RECT 716.475 1125.310 716.735 1125.630 ;
        RECT 716.595 1116.100 716.735 1125.310 ;
        RECT 717.740 1125.330 717.880 1129.625 ;
        RECT 717.740 1125.010 718.000 1125.330 ;
        RECT 718.360 1125.050 718.500 1129.625 ;
        RECT 721.605 1125.350 721.745 1129.625 ;
        RECT 716.100 1115.780 717.190 1116.100 ;
        RECT 711.470 1112.720 712.560 1113.040 ;
        RECT 715.530 1112.450 715.850 1113.300 ;
        RECT 717.740 1113.040 717.880 1125.010 ;
        RECT 718.360 1124.730 718.620 1125.050 ;
        RECT 721.605 1125.030 721.865 1125.350 ;
        RECT 722.575 1125.070 722.715 1129.625 ;
        RECT 718.360 1116.360 718.500 1124.730 ;
        RECT 718.280 1115.510 718.600 1116.360 ;
        RECT 721.605 1113.300 721.745 1125.030 ;
        RECT 722.575 1124.750 722.835 1125.070 ;
        RECT 723.720 1124.770 723.860 1129.625 ;
        RECT 722.575 1116.100 722.715 1124.750 ;
        RECT 723.720 1124.450 723.980 1124.770 ;
        RECT 724.340 1124.490 724.480 1129.625 ;
        RECT 727.585 1124.790 727.725 1129.625 ;
        RECT 722.080 1115.780 723.170 1116.100 ;
        RECT 717.450 1112.720 718.540 1113.040 ;
        RECT 721.510 1112.450 721.830 1113.300 ;
        RECT 723.720 1113.040 723.860 1124.450 ;
        RECT 724.340 1124.170 724.600 1124.490 ;
        RECT 727.585 1124.470 727.845 1124.790 ;
        RECT 728.555 1124.510 728.695 1129.625 ;
        RECT 724.340 1116.360 724.480 1124.170 ;
        RECT 724.260 1115.510 724.580 1116.360 ;
        RECT 727.585 1113.300 727.725 1124.470 ;
        RECT 728.555 1124.190 728.815 1124.510 ;
        RECT 729.700 1124.210 729.840 1129.625 ;
        RECT 728.555 1116.100 728.695 1124.190 ;
        RECT 729.700 1123.890 729.960 1124.210 ;
        RECT 730.320 1123.930 730.460 1129.625 ;
        RECT 733.565 1124.230 733.705 1129.625 ;
        RECT 728.060 1115.780 729.150 1116.100 ;
        RECT 723.430 1112.720 724.520 1113.040 ;
        RECT 727.490 1112.450 727.810 1113.300 ;
        RECT 729.700 1113.040 729.840 1123.890 ;
        RECT 730.320 1123.610 730.580 1123.930 ;
        RECT 733.565 1123.910 733.825 1124.230 ;
        RECT 734.535 1123.950 734.675 1129.625 ;
        RECT 730.320 1116.360 730.460 1123.610 ;
        RECT 730.240 1115.510 730.560 1116.360 ;
        RECT 733.565 1113.300 733.705 1123.910 ;
        RECT 734.535 1123.630 734.795 1123.950 ;
        RECT 735.680 1123.650 735.820 1129.625 ;
        RECT 734.535 1116.100 734.675 1123.630 ;
        RECT 735.680 1123.330 735.940 1123.650 ;
        RECT 736.300 1123.370 736.440 1129.625 ;
        RECT 739.545 1123.670 739.685 1129.625 ;
        RECT 734.040 1115.780 735.130 1116.100 ;
        RECT 729.410 1112.720 730.500 1113.040 ;
        RECT 733.470 1112.450 733.790 1113.300 ;
        RECT 735.680 1113.040 735.820 1123.330 ;
        RECT 736.300 1123.050 736.560 1123.370 ;
        RECT 739.545 1123.350 739.805 1123.670 ;
        RECT 740.515 1123.390 740.655 1129.625 ;
        RECT 736.300 1116.360 736.440 1123.050 ;
        RECT 736.220 1115.510 736.540 1116.360 ;
        RECT 739.545 1113.300 739.685 1123.350 ;
        RECT 740.515 1123.070 740.775 1123.390 ;
        RECT 741.660 1123.090 741.800 1129.625 ;
        RECT 740.515 1116.100 740.655 1123.070 ;
        RECT 741.660 1122.770 741.920 1123.090 ;
        RECT 742.280 1122.810 742.420 1129.625 ;
        RECT 745.525 1123.110 745.665 1129.625 ;
        RECT 740.020 1115.780 741.110 1116.100 ;
        RECT 735.390 1112.720 736.480 1113.040 ;
        RECT 739.450 1112.450 739.770 1113.300 ;
        RECT 741.660 1113.040 741.800 1122.770 ;
        RECT 742.280 1122.490 742.540 1122.810 ;
        RECT 745.525 1122.790 745.785 1123.110 ;
        RECT 746.495 1122.830 746.635 1129.625 ;
        RECT 742.280 1116.360 742.420 1122.490 ;
        RECT 742.200 1115.510 742.520 1116.360 ;
        RECT 745.525 1113.300 745.665 1122.790 ;
        RECT 746.495 1122.510 746.755 1122.830 ;
        RECT 747.640 1122.530 747.780 1129.625 ;
        RECT 746.495 1116.100 746.635 1122.510 ;
        RECT 747.640 1122.210 747.900 1122.530 ;
        RECT 748.260 1122.250 748.400 1129.625 ;
        RECT 751.505 1122.550 751.645 1129.625 ;
        RECT 746.000 1115.780 747.090 1116.100 ;
        RECT 741.370 1112.720 742.460 1113.040 ;
        RECT 745.430 1112.450 745.750 1113.300 ;
        RECT 747.640 1113.040 747.780 1122.210 ;
        RECT 748.260 1121.930 748.520 1122.250 ;
        RECT 751.505 1122.230 751.765 1122.550 ;
        RECT 752.475 1122.270 752.615 1129.625 ;
        RECT 748.260 1116.360 748.400 1121.930 ;
        RECT 748.180 1115.510 748.500 1116.360 ;
        RECT 751.505 1113.300 751.645 1122.230 ;
        RECT 752.475 1121.950 752.735 1122.270 ;
        RECT 753.620 1121.970 753.760 1129.625 ;
        RECT 752.475 1116.100 752.615 1121.950 ;
        RECT 753.620 1121.650 753.880 1121.970 ;
        RECT 754.240 1121.690 754.380 1129.625 ;
        RECT 757.485 1121.990 757.625 1129.625 ;
        RECT 751.980 1115.780 753.070 1116.100 ;
        RECT 747.350 1112.720 748.440 1113.040 ;
        RECT 751.410 1112.450 751.730 1113.300 ;
        RECT 753.620 1113.040 753.760 1121.650 ;
        RECT 754.240 1121.370 754.500 1121.690 ;
        RECT 757.485 1121.670 757.745 1121.990 ;
        RECT 758.455 1121.710 758.595 1129.625 ;
        RECT 754.240 1116.360 754.380 1121.370 ;
        RECT 754.160 1115.510 754.480 1116.360 ;
        RECT 757.485 1113.300 757.625 1121.670 ;
        RECT 758.455 1121.390 758.715 1121.710 ;
        RECT 759.600 1121.410 759.740 1129.625 ;
        RECT 763.465 1121.430 763.605 1129.625 ;
        RECT 758.455 1116.100 758.595 1121.390 ;
        RECT 759.600 1121.090 759.860 1121.410 ;
        RECT 763.465 1121.110 763.725 1121.430 ;
        RECT 764.435 1121.150 764.575 1129.625 ;
        RECT 757.960 1115.780 759.050 1116.100 ;
        RECT 753.330 1112.720 754.420 1113.040 ;
        RECT 757.390 1112.450 757.710 1113.300 ;
        RECT 759.600 1113.040 759.740 1121.090 ;
        RECT 763.465 1113.300 763.605 1121.110 ;
        RECT 764.435 1120.830 764.695 1121.150 ;
        RECT 769.445 1120.870 769.585 1129.625 ;
        RECT 764.435 1116.100 764.575 1120.830 ;
        RECT 769.445 1120.550 769.705 1120.870 ;
        RECT 770.415 1120.590 770.555 1129.625 ;
        RECT 763.940 1115.780 765.030 1116.100 ;
        RECT 769.445 1113.300 769.585 1120.550 ;
        RECT 770.415 1120.270 770.675 1120.590 ;
        RECT 775.425 1120.310 775.565 1129.625 ;
        RECT 770.415 1116.100 770.555 1120.270 ;
        RECT 775.425 1119.990 775.685 1120.310 ;
        RECT 776.395 1120.030 776.535 1129.625 ;
        RECT 769.920 1115.780 771.010 1116.100 ;
        RECT 775.425 1113.300 775.565 1119.990 ;
        RECT 776.275 1119.710 776.535 1120.030 ;
        RECT 776.395 1116.100 776.535 1119.710 ;
        RECT 781.405 1119.750 781.545 1129.625 ;
        RECT 781.405 1119.430 781.665 1119.750 ;
        RECT 782.375 1119.470 782.515 1129.625 ;
        RECT 775.900 1115.780 776.990 1116.100 ;
        RECT 781.405 1113.300 781.545 1119.430 ;
        RECT 782.375 1119.150 782.635 1119.470 ;
        RECT 787.385 1119.190 787.525 1129.625 ;
        RECT 782.375 1116.100 782.515 1119.150 ;
        RECT 787.385 1118.870 787.645 1119.190 ;
        RECT 788.355 1118.910 788.495 1129.625 ;
        RECT 781.880 1115.780 782.970 1116.100 ;
        RECT 787.385 1113.300 787.525 1118.870 ;
        RECT 788.235 1118.590 788.495 1118.910 ;
        RECT 788.355 1116.100 788.495 1118.590 ;
        RECT 793.365 1118.630 793.505 1129.625 ;
        RECT 793.365 1118.310 793.625 1118.630 ;
        RECT 794.335 1118.350 794.475 1129.625 ;
        RECT 1970.520 1129.350 1970.780 1129.670 ;
        RECT 1975.880 1129.390 1976.020 1129.765 ;
        RECT 787.860 1115.780 788.950 1116.100 ;
        RECT 793.365 1114.240 793.505 1118.310 ;
        RECT 794.335 1118.030 794.595 1118.350 ;
        RECT 794.335 1116.100 794.475 1118.030 ;
        RECT 1970.520 1116.360 1970.660 1129.350 ;
        RECT 1975.880 1129.070 1976.140 1129.390 ;
        RECT 1976.500 1129.110 1976.640 1129.765 ;
        RECT 793.840 1115.780 794.930 1116.100 ;
        RECT 1970.440 1115.510 1970.760 1116.360 ;
        RECT 793.365 1114.100 794.140 1114.240 ;
        RECT 759.310 1112.720 760.400 1113.040 ;
        RECT 763.370 1112.450 763.690 1113.300 ;
        RECT 769.350 1112.450 769.670 1113.300 ;
        RECT 775.330 1112.450 775.650 1113.300 ;
        RECT 781.310 1112.450 781.630 1113.300 ;
        RECT 787.290 1112.450 787.610 1113.300 ;
        RECT 794.000 1113.040 794.140 1114.100 ;
        RECT 1975.880 1113.040 1976.020 1129.070 ;
        RECT 1976.500 1128.790 1976.760 1129.110 ;
        RECT 1981.860 1128.830 1982.000 1129.765 ;
        RECT 1976.500 1116.360 1976.640 1128.790 ;
        RECT 1981.860 1128.510 1982.120 1128.830 ;
        RECT 1982.480 1128.550 1982.620 1129.765 ;
        RECT 1976.420 1115.510 1976.740 1116.360 ;
        RECT 1981.860 1113.040 1982.000 1128.510 ;
        RECT 1982.480 1128.230 1982.740 1128.550 ;
        RECT 1987.840 1128.270 1987.980 1129.765 ;
        RECT 1982.480 1116.360 1982.620 1128.230 ;
        RECT 1987.840 1127.950 1988.100 1128.270 ;
        RECT 1988.460 1127.990 1988.600 1129.765 ;
        RECT 1982.400 1115.510 1982.720 1116.360 ;
        RECT 1987.840 1113.040 1987.980 1127.950 ;
        RECT 1988.460 1127.670 1988.720 1127.990 ;
        RECT 1993.820 1127.710 1993.960 1129.765 ;
        RECT 1988.460 1116.360 1988.600 1127.670 ;
        RECT 1993.820 1127.390 1994.080 1127.710 ;
        RECT 1994.440 1127.430 1994.580 1129.765 ;
        RECT 1988.380 1115.510 1988.700 1116.360 ;
        RECT 1993.820 1113.040 1993.960 1127.390 ;
        RECT 1994.440 1127.110 1994.700 1127.430 ;
        RECT 1999.800 1127.150 1999.940 1129.765 ;
        RECT 1994.440 1116.360 1994.580 1127.110 ;
        RECT 1999.800 1126.830 2000.060 1127.150 ;
        RECT 2000.420 1126.870 2000.560 1129.765 ;
        RECT 1994.360 1115.510 1994.680 1116.360 ;
        RECT 1999.800 1113.040 1999.940 1126.830 ;
        RECT 2000.420 1126.550 2000.680 1126.870 ;
        RECT 2005.780 1126.590 2005.920 1129.765 ;
        RECT 2000.420 1116.360 2000.560 1126.550 ;
        RECT 2005.780 1126.270 2006.040 1126.590 ;
        RECT 2006.400 1126.310 2006.540 1129.765 ;
        RECT 2000.340 1115.510 2000.660 1116.360 ;
        RECT 2005.780 1113.040 2005.920 1126.270 ;
        RECT 2006.400 1125.990 2006.660 1126.310 ;
        RECT 2011.760 1126.030 2011.900 1129.765 ;
        RECT 2006.400 1116.360 2006.540 1125.990 ;
        RECT 2011.760 1125.710 2012.020 1126.030 ;
        RECT 2012.380 1125.750 2012.520 1129.765 ;
        RECT 2006.320 1115.510 2006.640 1116.360 ;
        RECT 2011.760 1113.040 2011.900 1125.710 ;
        RECT 2012.380 1125.430 2012.640 1125.750 ;
        RECT 2017.740 1125.470 2017.880 1129.765 ;
        RECT 2012.380 1116.360 2012.520 1125.430 ;
        RECT 2017.740 1125.150 2018.000 1125.470 ;
        RECT 2018.360 1125.190 2018.500 1129.765 ;
        RECT 2012.300 1115.510 2012.620 1116.360 ;
        RECT 2017.740 1113.040 2017.880 1125.150 ;
        RECT 2018.360 1124.870 2018.620 1125.190 ;
        RECT 2023.720 1124.910 2023.860 1129.765 ;
        RECT 2018.360 1116.360 2018.500 1124.870 ;
        RECT 2023.720 1124.590 2023.980 1124.910 ;
        RECT 2024.340 1124.630 2024.480 1129.765 ;
        RECT 2018.280 1115.510 2018.600 1116.360 ;
        RECT 2023.720 1113.040 2023.860 1124.590 ;
        RECT 2024.340 1124.310 2024.600 1124.630 ;
        RECT 2029.700 1124.350 2029.840 1129.765 ;
        RECT 2024.340 1116.360 2024.480 1124.310 ;
        RECT 2029.700 1124.030 2029.960 1124.350 ;
        RECT 2030.320 1124.070 2030.460 1129.765 ;
        RECT 2024.260 1115.510 2024.580 1116.360 ;
        RECT 2029.700 1113.040 2029.840 1124.030 ;
        RECT 2030.320 1123.750 2030.580 1124.070 ;
        RECT 2035.680 1123.790 2035.820 1129.765 ;
        RECT 2030.320 1116.360 2030.460 1123.750 ;
        RECT 2035.680 1123.470 2035.940 1123.790 ;
        RECT 2036.300 1123.510 2036.440 1129.765 ;
        RECT 2030.240 1115.510 2030.560 1116.360 ;
        RECT 2035.680 1113.040 2035.820 1123.470 ;
        RECT 2036.300 1123.190 2036.560 1123.510 ;
        RECT 2041.660 1123.230 2041.800 1129.765 ;
        RECT 2036.300 1116.360 2036.440 1123.190 ;
        RECT 2041.660 1122.910 2041.920 1123.230 ;
        RECT 2042.280 1122.950 2042.420 1129.765 ;
        RECT 2036.220 1115.510 2036.540 1116.360 ;
        RECT 2041.660 1113.040 2041.800 1122.910 ;
        RECT 2042.280 1122.630 2042.540 1122.950 ;
        RECT 2047.640 1122.670 2047.780 1129.765 ;
        RECT 2042.280 1116.360 2042.420 1122.630 ;
        RECT 2047.640 1122.350 2047.900 1122.670 ;
        RECT 2048.260 1122.390 2048.400 1129.765 ;
        RECT 2042.200 1115.510 2042.520 1116.360 ;
        RECT 2047.640 1113.040 2047.780 1122.350 ;
        RECT 2048.260 1122.070 2048.520 1122.390 ;
        RECT 2053.620 1122.110 2053.760 1129.765 ;
        RECT 2048.260 1116.360 2048.400 1122.070 ;
        RECT 2053.620 1121.790 2053.880 1122.110 ;
        RECT 2054.240 1121.830 2054.380 1129.765 ;
        RECT 2048.180 1115.510 2048.500 1116.360 ;
        RECT 2053.620 1113.040 2053.760 1121.790 ;
        RECT 2054.240 1121.510 2054.500 1121.830 ;
        RECT 2059.600 1121.550 2059.740 1129.765 ;
        RECT 2054.240 1116.360 2054.380 1121.510 ;
        RECT 2059.600 1121.230 2059.860 1121.550 ;
        RECT 2060.220 1121.270 2060.360 1129.765 ;
        RECT 2054.160 1115.510 2054.480 1116.360 ;
        RECT 2059.600 1113.040 2059.740 1121.230 ;
        RECT 2060.220 1120.950 2060.480 1121.270 ;
        RECT 2065.580 1120.990 2065.720 1129.765 ;
        RECT 2060.220 1116.360 2060.360 1120.950 ;
        RECT 2065.580 1120.670 2065.840 1120.990 ;
        RECT 2066.200 1120.710 2066.340 1129.765 ;
        RECT 2060.140 1115.510 2060.460 1116.360 ;
        RECT 2065.580 1113.040 2065.720 1120.670 ;
        RECT 2066.200 1120.390 2066.460 1120.710 ;
        RECT 2071.560 1120.430 2071.700 1129.765 ;
        RECT 2066.200 1116.360 2066.340 1120.390 ;
        RECT 2071.560 1120.110 2071.820 1120.430 ;
        RECT 2072.180 1120.150 2072.320 1129.765 ;
        RECT 2066.120 1115.510 2066.440 1116.360 ;
        RECT 2071.560 1113.040 2071.700 1120.110 ;
        RECT 2072.180 1119.830 2072.440 1120.150 ;
        RECT 2077.540 1119.870 2077.680 1129.765 ;
        RECT 2072.180 1116.360 2072.320 1119.830 ;
        RECT 2077.540 1119.550 2077.800 1119.870 ;
        RECT 2078.160 1119.590 2078.300 1129.765 ;
        RECT 2072.100 1115.510 2072.420 1116.360 ;
        RECT 2077.540 1113.040 2077.680 1119.550 ;
        RECT 2078.160 1119.270 2078.420 1119.590 ;
        RECT 2083.520 1119.310 2083.660 1129.765 ;
        RECT 2078.160 1116.360 2078.300 1119.270 ;
        RECT 2083.520 1118.990 2083.780 1119.310 ;
        RECT 2084.140 1119.030 2084.280 1129.765 ;
        RECT 2078.080 1115.510 2078.400 1116.360 ;
        RECT 2083.520 1113.040 2083.660 1118.990 ;
        RECT 2084.140 1118.710 2084.400 1119.030 ;
        RECT 2089.500 1118.750 2089.640 1129.765 ;
        RECT 2084.140 1116.360 2084.280 1118.710 ;
        RECT 2089.500 1118.430 2089.760 1118.750 ;
        RECT 2090.120 1118.470 2090.260 1129.765 ;
        RECT 2084.060 1115.510 2084.380 1116.360 ;
        RECT 2089.500 1114.170 2089.640 1118.430 ;
        RECT 2090.120 1118.150 2090.380 1118.470 ;
        RECT 2090.120 1116.360 2090.260 1118.150 ;
        RECT 2090.040 1115.510 2090.360 1116.360 ;
        RECT 2089.500 1114.030 2090.275 1114.170 ;
        RECT 2090.135 1113.300 2090.275 1114.030 ;
        RECT 793.340 1112.720 794.430 1113.040 ;
        RECT 1975.590 1112.720 1976.680 1113.040 ;
        RECT 1981.570 1112.720 1982.660 1113.040 ;
        RECT 1987.550 1112.720 1988.640 1113.040 ;
        RECT 1993.530 1112.720 1994.620 1113.040 ;
        RECT 1999.510 1112.720 2000.600 1113.040 ;
        RECT 2005.490 1112.720 2006.580 1113.040 ;
        RECT 2011.470 1112.720 2012.560 1113.040 ;
        RECT 2017.450 1112.720 2018.540 1113.040 ;
        RECT 2023.430 1112.720 2024.520 1113.040 ;
        RECT 2029.410 1112.720 2030.500 1113.040 ;
        RECT 2035.390 1112.720 2036.480 1113.040 ;
        RECT 2041.370 1112.720 2042.460 1113.040 ;
        RECT 2047.350 1112.720 2048.440 1113.040 ;
        RECT 2053.330 1112.720 2054.420 1113.040 ;
        RECT 2059.310 1112.720 2060.400 1113.040 ;
        RECT 2065.290 1112.720 2066.380 1113.040 ;
        RECT 2071.270 1112.720 2072.360 1113.040 ;
        RECT 2077.250 1112.720 2078.340 1113.040 ;
        RECT 2083.230 1112.720 2084.320 1113.040 ;
        RECT 2090.050 1112.450 2090.370 1113.300 ;
  END
END gpio_signal_buffering
END LIBRARY

