VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO empty_macro
  CLASS BLOCK ;
  FOREIGN empty_macro ;
  ORIGIN 0.000 0.000 ;
  SIZE 3141.260 BY 572.000 ;
END empty_macro
END LIBRARY

