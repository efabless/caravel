VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_id_textblock
  CLASS BLOCK ;
  FOREIGN user_id_textblock ;
  ORIGIN 0.000 0.000 ;
  SIZE 40.000 BY 25.000 ;
END user_id_textblock
END LIBRARY

