* NGSPICE file created from gpio_control_block.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dfbbn_1 abstract view
.subckt sky130_fd_sc_hd__dfbbn_1 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_2 abstract view
.subckt sky130_fd_sc_hd__einvp_2 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_1 abstract view
.subckt sky130_fd_sc_hd__ebufn_1 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for gpio_logic_high abstract view
.subckt gpio_logic_high gpio_logic1 vccd1 vssd1
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

.subckt gpio_control_block gpio_defaults[0] gpio_defaults[10] gpio_defaults[11] gpio_defaults[12]
+ gpio_defaults[1] gpio_defaults[2] gpio_defaults[3] gpio_defaults[4] gpio_defaults[5]
+ gpio_defaults[6] gpio_defaults[7] gpio_defaults[8] gpio_defaults[9] mgmt_gpio_in
+ mgmt_gpio_oeb mgmt_gpio_out one pad_gpio_ana_en pad_gpio_ana_pol pad_gpio_ana_sel
+ pad_gpio_dm[0] pad_gpio_dm[1] pad_gpio_dm[2] pad_gpio_holdover pad_gpio_ib_mode_sel
+ pad_gpio_in pad_gpio_inenb pad_gpio_out pad_gpio_outenb pad_gpio_slow_sel pad_gpio_vtrip_sel
+ resetn resetn_out serial_clock serial_clock_out serial_data_in serial_data_out serial_load
+ serial_load_out user_gpio_in user_gpio_oeb user_gpio_out vccd vccd1 vssd vssd1 zero
X_200_ _162_/X _220_/D _166_/X _164_/X vssd vssd vccd vccd _200_/Q _200_/Q_N sky130_fd_sc_hd__dfbbn_1
X_131_ _131_/A vssd vssd vccd vccd _131_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_5 gpio_defaults[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_78 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_114_ _190_/A _116_/B vssd vssd vccd vccd _115_/A sky130_fd_sc_hd__or2b_1
Xoutput31 _202_/Q vssd vssd vccd vccd pad_gpio_inenb sky130_fd_sc_hd__buf_2
X_130_ _130_/A vssd vssd vccd vccd _131_/A sky130_fd_sc_hd__clkbuf_1
X_113_ _113_/A vssd vssd vccd vccd _113_/X sky130_fd_sc_hd__clkbuf_1
Xoutput32 _196_/X vssd vssd vccd vccd pad_gpio_out sky130_fd_sc_hd__buf_2
XFILLER_6_46 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_6 gpio_defaults[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_189_ _189_/A vssd vssd vccd vccd _189_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_112_ _130_/A vssd vssd vccd vccd _113_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_7 gpio_defaults[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput33 _193_/X vssd vssd vccd vccd pad_gpio_outenb sky130_fd_sc_hd__buf_2
XFILLER_3_26 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_188_ _188_/A vssd vssd vccd vccd _189_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_15_9 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_14 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_111_ _111_/A vssd vssd vccd vccd _111_/X sky130_fd_sc_hd__clkbuf_1
Xoutput34 _200_/Q vssd vssd vccd vccd pad_gpio_slow_sel sky130_fd_sc_hd__buf_2
Xoutput23 _208_/Q vssd vssd vccd vccd pad_gpio_ana_en sky130_fd_sc_hd__buf_2
XANTENNA_8 gpio_defaults[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_187_ _187_/A vssd vssd vccd vccd _187_/X sky130_fd_sc_hd__clkbuf_1
X_110_ _190_/A _110_/B vssd vssd vccd vccd _111_/A sky130_fd_sc_hd__or2_1
XFILLER_1_93 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput35 _201_/Q vssd vssd vccd vccd pad_gpio_vtrip_sel sky130_fd_sc_hd__buf_2
XANTENNA_9 gpio_defaults[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xoutput24 _210_/Q vssd vssd vccd vccd pad_gpio_ana_pol sky130_fd_sc_hd__buf_2
XFILLER_7_92 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_15 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_186_ one _223_/Q vssd vssd vccd vccd _187_/A sky130_fd_sc_hd__and2_1
X_169_ _190_/A _171_/B vssd vssd vccd vccd _170_/A sky130_fd_sc_hd__or2b_1
Xoutput36 _190_/X vssd vssd vccd vccd resetn_out sky130_fd_sc_hd__buf_2
Xoutput25 _209_/Q vssd vssd vccd vccd pad_gpio_ana_sel sky130_fd_sc_hd__buf_2
XPHY_0 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_92 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_185_ _197_/A vssd vssd vccd vccd _185_/Y sky130_fd_sc_hd__inv_2
XFILLER_4_61 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_168_ _168_/A vssd vssd vccd vccd _168_/X sky130_fd_sc_hd__clkbuf_1
Xoutput37 _191_/X vssd vssd vccd vccd serial_clock_out sky130_fd_sc_hd__clkbuf_1
Xoutput26 _205_/Q vssd vssd vccd vccd pad_gpio_dm[0] sky130_fd_sc_hd__buf_2
XPHY_1 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xconst_source vssd vssd vccd vccd one zero sky130_fd_sc_hd__conb_1
X_184_ _184_/A vssd vssd vccd vccd _194_/S sky130_fd_sc_hd__clkbuf_1
X_219_ _191_/A _219_/D _190_/A vssd vssd vccd vccd _220_/D sky130_fd_sc_hd__dfrtp_1
X_167_ _188_/A vssd vssd vccd vccd _168_/A sky130_fd_sc_hd__clkbuf_1
Xoutput38 _187_/X vssd vssd vccd vccd serial_data_out sky130_fd_sc_hd__buf_2
XFILLER_15_39 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xoutput27 _206_/Q vssd vssd vccd vccd pad_gpio_dm[1] sky130_fd_sc_hd__buf_2
XPHY_2 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_166_ _166_/A vssd vssd vccd vccd _166_/X sky130_fd_sc_hd__clkbuf_1
X_183_ _207_/Q _206_/Q vssd vssd vccd vccd _184_/A sky130_fd_sc_hd__or2b_1
XFILLER_1_86 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xoutput39 _192_/X vssd vssd vccd vccd serial_load_out sky130_fd_sc_hd__buf_2
Xoutput28 _207_/Q vssd vssd vccd vccd pad_gpio_dm[2] sky130_fd_sc_hd__buf_2
X_149_ _161_/A vssd vssd vccd vccd _150_/A sky130_fd_sc_hd__clkbuf_1
X_218_ _223_/CLK _218_/D _190_/A vssd vssd vccd vccd _219_/D sky130_fd_sc_hd__dfrtp_1
XPHY_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_182_ _182_/A vssd vssd vccd vccd _182_/X sky130_fd_sc_hd__clkbuf_1
X_165_ _190_/A _165_/B vssd vssd vccd vccd _166_/A sky130_fd_sc_hd__or2_1
X_217_ _223_/CLK _217_/D _190_/A vssd vssd vccd vccd _218_/D sky130_fd_sc_hd__dfrtp_1
X_148_ _148_/A vssd vssd vccd vccd _148_/X sky130_fd_sc_hd__clkbuf_1
Xoutput29 _199_/Q vssd vssd vccd vccd pad_gpio_holdover sky130_fd_sc_hd__buf_2
XPHY_4 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_181_ _204_/Q _195_/S vssd vssd vccd vccd _182_/A sky130_fd_sc_hd__and2_1
X_164_ _164_/A vssd vssd vccd vccd _164_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_77 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_20 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_216_ _223_/CLK _216_/D _190_/A vssd vssd vccd vccd _217_/D sky130_fd_sc_hd__dfrtp_1
X_147_ _190_/A _147_/B vssd vssd vccd vccd _148_/A sky130_fd_sc_hd__or2_1
XFILLER_16_85 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_5 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_180_ _180_/A vssd vssd vccd vccd _180_/X sky130_fd_sc_hd__clkbuf_1
X_163_ _190_/A _165_/B vssd vssd vccd vccd _164_/A sky130_fd_sc_hd__or2b_1
XFILLER_1_67 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_6 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_146_ _146_/A vssd vssd vccd vccd _146_/X sky130_fd_sc_hd__clkbuf_1
X_129_ _129_/A vssd vssd vccd vccd _129_/X sky130_fd_sc_hd__clkbuf_1
X_215_ _223_/CLK _215_/D _190_/A vssd vssd vccd vccd _216_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_13_65 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_162_ _162_/A vssd vssd vccd vccd _162_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_10 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xinput1 gpio_defaults[0] vssd vssd vccd vccd _177_/A sky130_fd_sc_hd__clkbuf_1
X_145_ _190_/A _147_/B vssd vssd vccd vccd _146_/A sky130_fd_sc_hd__or2b_1
X_214_ _191_/A _214_/D _190_/A vssd vssd vccd vccd _215_/D sky130_fd_sc_hd__dfrtp_1
X_128_ _190_/A _128_/B vssd vssd vccd vccd _129_/A sky130_fd_sc_hd__or2_1
XPHY_7 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xgpio_in_buf _185_/Y gpio_in_buf/TE vssd vssd vccd vccd output40/A sky130_fd_sc_hd__einvp_2
X_161_ _161_/A vssd vssd vccd vccd _162_/A sky130_fd_sc_hd__clkbuf_1
Xinput2 gpio_defaults[10] vssd vssd vccd vccd _134_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_16_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_213_ _191_/A _213_/D _190_/A vssd vssd vccd vccd _214_/D sky130_fd_sc_hd__dfrtp_1
X_127_ _127_/A vssd vssd vccd vccd _127_/X sky130_fd_sc_hd__clkbuf_1
X_144_ _144_/A vssd vssd vccd vccd _144_/X sky130_fd_sc_hd__clkbuf_1
XPHY_8 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_160_ _160_/A vssd vssd vccd vccd _160_/X sky130_fd_sc_hd__clkbuf_1
X_212_ _191_/A _212_/D _190_/A vssd vssd vccd vccd _213_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_10_68 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_13 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_26 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_143_ _161_/A vssd vssd vccd vccd _144_/A sky130_fd_sc_hd__clkbuf_1
Xinput3 gpio_defaults[11] vssd vssd vccd vccd _128_/B sky130_fd_sc_hd__clkbuf_1
X_126_ _190_/A _128_/B vssd vssd vccd vccd _127_/A sky130_fd_sc_hd__or2b_1
XPHY_9 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_57 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_109_ _109_/A vssd vssd vccd vccd _109_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_80 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput4 gpio_defaults[12] vssd vssd vccd vccd _122_/B sky130_fd_sc_hd__clkbuf_1
X_211_ _191_/A _211_/D _190_/A vssd vssd vccd vccd _212_/D sky130_fd_sc_hd__dfrtp_1
X_142_ _142_/A vssd vssd vccd vccd _142_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_20 gpio_defaults[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_125_ _125_/A vssd vssd vccd vccd _125_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_13 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_108_ _190_/A _110_/B vssd vssd vccd vccd _109_/A sky130_fd_sc_hd__or2b_1
XTAP_50 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_141_ _190_/A _141_/B vssd vssd vccd vccd _142_/A sky130_fd_sc_hd__or2_1
XFILLER_10_37 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xinput5 gpio_defaults[1] vssd vssd vccd vccd _141_/B sky130_fd_sc_hd__clkbuf_1
X_210_ _189_/X _219_/D _105_/X _103_/X vssd vssd vccd vccd _210_/Q _210_/Q_N sky130_fd_sc_hd__dfbbn_1
Xclkbuf_1_1_0_serial_clock clkbuf_0_serial_clock/X vssd vssd vccd vccd _191_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_21 serial_load vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_124_ _130_/A vssd vssd vccd vccd _125_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_10 gpio_defaults[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_93 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_107_ _188_/A vssd vssd vccd vccd _130_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_5_93 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_51 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_140_ _140_/A vssd vssd vccd vccd _140_/X sky130_fd_sc_hd__clkbuf_1
Xinput6 gpio_defaults[2] vssd vssd vccd vccd _171_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA_11 gpio_defaults[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XTAP_40 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_106_ _192_/A vssd vssd vccd vccd _188_/A sky130_fd_sc_hd__inv_2
Xinput20 user_gpio_oeb vssd vssd vccd vccd _193_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_16_7 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_92 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_123_ _123_/A vssd vssd vccd vccd _123_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_13_49 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_52 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 gpio_defaults[3] vssd vssd vccd vccd _153_/B sky130_fd_sc_hd__clkbuf_1
XTAP_41 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput21 user_gpio_out vssd vssd vccd vccd _196_/A0 sky130_fd_sc_hd__clkbuf_1
X_199_ _168_/X _214_/D _172_/X _170_/X vssd vssd vccd vccd _199_/Q _199_/Q_N sky130_fd_sc_hd__dfbbn_1
XANTENNA_12 mgmt_gpio_oeb vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_122_ _190_/A _122_/B vssd vssd vccd vccd _123_/A sky130_fd_sc_hd__or2_1
Xinput10 gpio_defaults[6] vssd vssd vccd vccd _110_/B sky130_fd_sc_hd__clkbuf_1
X_105_ _105_/A vssd vssd vccd vccd _105_/X sky130_fd_sc_hd__clkbuf_1
X_198_ _174_/X _212_/D _178_/X _176_/X vssd vssd vccd vccd _198_/Q _198_/Q_N sky130_fd_sc_hd__dfbbn_1
XTAP_53 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 gpio_defaults[4] vssd vssd vccd vccd _147_/B sky130_fd_sc_hd__clkbuf_1
XTAP_42 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_29 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_13 mgmt_gpio_out vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_104_ _190_/A _104_/B vssd vssd vccd vccd _105_/A sky130_fd_sc_hd__or2_1
X_121_ _121_/A vssd vssd vccd vccd _121_/X sky130_fd_sc_hd__clkbuf_1
Xinput11 gpio_defaults[7] vssd vssd vccd vccd _104_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_12_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_54 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 gpio_defaults[5] vssd vssd vccd vccd _116_/B sky130_fd_sc_hd__clkbuf_1
XTAP_43 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_197_ _197_/A _180_/X vssd vssd vccd vccd mgmt_gpio_in sky130_fd_sc_hd__ebufn_1
XANTENNA_14 one vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xinput12 gpio_defaults[8] vssd vssd vccd vccd _165_/B sky130_fd_sc_hd__clkbuf_1
X_120_ _190_/A _122_/B vssd vssd vccd vccd _121_/A sky130_fd_sc_hd__or2b_1
XFILLER_16_18 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_103_ _103_/A vssd vssd vccd vccd _103_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_53 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_196_ _196_/A0 _195_/X _198_/Q vssd vssd vccd vccd _196_/X sky130_fd_sc_hd__mux2_1
XTAP_55 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_44 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_15 one vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_179_ _202_/Q _204_/Q vssd vssd vccd vccd _180_/A sky130_fd_sc_hd__or2b_1
Xinput13 gpio_defaults[9] vssd vssd vccd vccd _159_/B sky130_fd_sc_hd__clkbuf_1
X_102_ _190_/A _104_/B vssd vssd vccd vccd _103_/A sky130_fd_sc_hd__or2b_1
XFILLER_8_20 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_56 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_45 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xgpio_logic_high gpio_in_buf/TE vccd1 vssd1 gpio_logic_high
XTAP_34 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_16 pad_gpio_in vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_195_ _195_/A0 _194_/X _195_/S vssd vssd vccd vccd _195_/X sky130_fd_sc_hd__mux2_1
Xinput14 mgmt_gpio_oeb vssd vssd vccd vccd _195_/S sky130_fd_sc_hd__clkbuf_1
X_178_ _178_/A vssd vssd vccd vccd _178_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_8_10 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XTAP_57 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_194_ _194_/A0 _195_/A0 _194_/S vssd vssd vccd vccd _194_/X sky130_fd_sc_hd__mux2_1
XTAP_46 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_35 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_17 serial_data_in vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_177_ _177_/A _190_/A vssd vssd vccd vccd _178_/A sky130_fd_sc_hd__or2_1
Xinput15 mgmt_gpio_out vssd vssd vccd vccd _195_/A0 sky130_fd_sc_hd__clkbuf_1
XFILLER_8_33 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XTAP_58 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_47 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_36 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_18 user_gpio_oeb vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_31 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_193_ _193_/A0 _182_/X _198_/Q vssd vssd vccd vccd _193_/X sky130_fd_sc_hd__mux2_1
XPHY_20 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_159_ _190_/A _159_/B vssd vssd vccd vccd _160_/A sky130_fd_sc_hd__or2_1
X_176_ _176_/A vssd vssd vccd vccd _176_/X sky130_fd_sc_hd__clkbuf_1
Xinput16 pad_gpio_in vssd vssd vccd vccd _197_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_8_45 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_192_ _192_/A vssd vssd vccd vccd _192_/X sky130_fd_sc_hd__clkbuf_1
XPHY_21 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_48 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XTAP_37 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput17 resetn vssd vssd vccd vccd _190_/A sky130_fd_sc_hd__buf_12
XANTENNA_19 user_gpio_out vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_175_ _190_/A _177_/A vssd vssd vccd vccd _176_/A sky130_fd_sc_hd__or2b_1
XFILLER_11_78 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_12 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_158_ _158_/A vssd vssd vccd vccd _158_/X sky130_fd_sc_hd__clkbuf_1
XTAP_49 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_38 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0_0_serial_clock clkbuf_0_serial_clock/X vssd vssd vccd vccd _223_/CLK sky130_fd_sc_hd__clkbuf_2
XPHY_33 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_191_ _191_/A vssd vssd vccd vccd _191_/X sky130_fd_sc_hd__buf_2
XFILLER_11_57 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_46 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_22 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xclkbuf_0_serial_clock serial_clock vssd vssd vccd vccd clkbuf_0_serial_clock/X sky130_fd_sc_hd__clkbuf_16
XPHY_11 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_174_ _174_/A vssd vssd vccd vccd _174_/X sky130_fd_sc_hd__clkbuf_1
Xinput18 serial_data_in vssd vssd vccd vccd _211_/D sky130_fd_sc_hd__clkbuf_1
X_157_ _190_/A _159_/B vssd vssd vccd vccd _158_/A sky130_fd_sc_hd__or2b_1
XFILLER_5_26 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_209_ _130_/A _218_/D _111_/X _109_/X vssd vssd vccd vccd _209_/Q _209_/Q_N sky130_fd_sc_hd__dfbbn_1
XTAP_39 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_23 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_173_ _188_/A vssd vssd vccd vccd _174_/A sky130_fd_sc_hd__clkbuf_1
X_190_ _190_/A vssd vssd vccd vccd _190_/X sky130_fd_sc_hd__clkbuf_1
Xinput19 serial_load vssd vssd vccd vccd _192_/A sky130_fd_sc_hd__clkbuf_1
X_156_ _156_/A vssd vssd vccd vccd _156_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_92 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_139_ _190_/A _141_/B vssd vssd vccd vccd _140_/A sky130_fd_sc_hd__or2b_1
X_208_ _113_/X _217_/D _117_/X _115_/X vssd vssd vccd vccd _208_/Q _208_/Q_N sky130_fd_sc_hd__dfbbn_1
XPHY_24 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_13 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_155_ _161_/A vssd vssd vccd vccd _156_/A sky130_fd_sc_hd__clkbuf_1
X_172_ _172_/A vssd vssd vccd vccd _172_/X sky130_fd_sc_hd__clkbuf_1
X_138_ _138_/A vssd vssd vccd vccd _138_/X sky130_fd_sc_hd__clkbuf_1
X_207_ _119_/X _223_/Q _123_/X _121_/X vssd vssd vccd vccd _207_/Q _207_/Q_N sky130_fd_sc_hd__dfbbn_1
XFILLER_14_15 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_25 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_171_ _190_/A _171_/B vssd vssd vccd vccd _172_/A sky130_fd_sc_hd__or2_1
XPHY_14 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_154_ _154_/A vssd vssd vccd vccd _154_/X sky130_fd_sc_hd__clkbuf_1
X_223_ _223_/CLK _223_/D _190_/A vssd vssd vccd vccd _223_/Q sky130_fd_sc_hd__dfrtp_1
X_137_ _161_/A vssd vssd vccd vccd _138_/A sky130_fd_sc_hd__clkbuf_1
X_206_ _125_/X _223_/D _129_/X _127_/X vssd vssd vccd vccd _206_/Q _206_/Q_N sky130_fd_sc_hd__dfbbn_1
XFILLER_15_81 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_26 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_170_ _170_/A vssd vssd vccd vccd _170_/X sky130_fd_sc_hd__clkbuf_1
X_205_ _131_/X _222_/D _135_/X _133_/X vssd vssd vccd vccd _205_/Q _194_/A0 sky130_fd_sc_hd__dfbbn_1
X_136_ _188_/A vssd vssd vccd vccd _161_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_222_ _223_/CLK _222_/D _190_/A vssd vssd vccd vccd _223_/D sky130_fd_sc_hd__dfrtp_1
X_153_ _190_/A _153_/B vssd vssd vccd vccd _154_/A sky130_fd_sc_hd__or2_1
XFILLER_0_85 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_119_ _119_/A vssd vssd vccd vccd _119_/X sky130_fd_sc_hd__clkbuf_1
XPHY_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_16 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_0 gpio_defaults[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_221_ _191_/A _221_/D _190_/A vssd vssd vccd vccd _222_/D sky130_fd_sc_hd__dfrtp_1
XFILLER_12_72 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_152_ _152_/A vssd vssd vccd vccd _152_/X sky130_fd_sc_hd__clkbuf_1
X_204_ _138_/X _213_/D _142_/X _140_/X vssd vssd vccd vccd _204_/Q _204_/Q_N sky130_fd_sc_hd__dfbbn_1
X_135_ _135_/A vssd vssd vccd vccd _135_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_118_ _130_/A vssd vssd vccd vccd _119_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_14_29 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_28 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_17 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_1 gpio_defaults[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_19 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_220_ _191_/A _220_/D _190_/A vssd vssd vccd vccd _221_/D sky130_fd_sc_hd__dfrtp_1
X_134_ _190_/A _134_/B vssd vssd vccd vccd _135_/A sky130_fd_sc_hd__or2_1
X_203_ _144_/X _216_/D _148_/X _146_/X vssd vssd vccd vccd _203_/Q _203_/Q_N sky130_fd_sc_hd__dfbbn_1
X_151_ _190_/A _153_/B vssd vssd vccd vccd _152_/A sky130_fd_sc_hd__or2b_1
XFILLER_15_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_63 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_117_ _117_/A vssd vssd vccd vccd _117_/X sky130_fd_sc_hd__clkbuf_1
XPHY_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_8 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_18 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_2 gpio_defaults[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_41 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_150_ _150_/A vssd vssd vccd vccd _150_/X sky130_fd_sc_hd__clkbuf_1
X_202_ _150_/X _215_/D _154_/X _152_/X vssd vssd vccd vccd _202_/Q _202_/Q_N sky130_fd_sc_hd__dfbbn_1
X_133_ _133_/A vssd vssd vccd vccd _133_/X sky130_fd_sc_hd__clkbuf_1
XPHY_19 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_3 gpio_defaults[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_116_ _190_/A _116_/B vssd vssd vccd vccd _117_/A sky130_fd_sc_hd__or2_1
Xoutput40 output40/A vssd vssd vccd vccd user_gpio_in sky130_fd_sc_hd__buf_2
X_201_ _156_/X _221_/D _160_/X _158_/X vssd vssd vccd vccd _201_/Q _201_/Q_N sky130_fd_sc_hd__dfbbn_1
X_132_ _190_/A _134_/B vssd vssd vccd vccd _133_/A sky130_fd_sc_hd__or2b_1
X_115_ _115_/A vssd vssd vccd vccd _115_/X sky130_fd_sc_hd__clkbuf_1
Xoutput30 _203_/Q vssd vssd vccd vccd pad_gpio_ib_mode_sel sky130_fd_sc_hd__buf_2
XANTENNA_4 gpio_defaults[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
.ends

