magic
tech sky130A
magscale 1 2
timestamp 1668092855
<< metal1 >>
rect 366174 1027828 366180 1027880
rect 366232 1027868 366238 1027880
rect 366542 1027868 366548 1027880
rect 366232 1027840 366548 1027868
rect 366232 1027828 366238 1027840
rect 366542 1027828 366548 1027840
rect 366600 1027828 366606 1027880
rect 366174 1024360 366180 1024412
rect 366232 1024400 366238 1024412
rect 366542 1024400 366548 1024412
rect 366232 1024372 366548 1024400
rect 366232 1024360 366238 1024372
rect 366542 1024360 366548 1024372
rect 366600 1024360 366606 1024412
rect 200022 1007360 200028 1007412
rect 200080 1007400 200086 1007412
rect 202690 1007400 202696 1007412
rect 200080 1007372 202696 1007400
rect 200080 1007360 200086 1007372
rect 202690 1007360 202696 1007372
rect 202748 1007360 202754 1007412
rect 505370 1007088 505376 1007140
rect 505428 1007128 505434 1007140
rect 513834 1007128 513840 1007140
rect 505428 1007100 513840 1007128
rect 505428 1007088 505434 1007100
rect 513834 1007088 513840 1007100
rect 513892 1007088 513898 1007140
rect 427998 1006884 428004 1006936
rect 428056 1006924 428062 1006936
rect 428056 1006896 441614 1006924
rect 428056 1006884 428062 1006896
rect 357710 1006816 357716 1006868
rect 357768 1006856 357774 1006868
rect 369854 1006856 369860 1006868
rect 357768 1006828 369860 1006856
rect 357768 1006816 357774 1006828
rect 369854 1006816 369860 1006828
rect 369912 1006816 369918 1006868
rect 430850 1006748 430856 1006800
rect 430908 1006788 430914 1006800
rect 434622 1006788 434628 1006800
rect 430908 1006760 434628 1006788
rect 430908 1006748 430914 1006760
rect 434622 1006748 434628 1006760
rect 434680 1006748 434686 1006800
rect 360194 1006680 360200 1006732
rect 360252 1006720 360258 1006732
rect 373258 1006720 373264 1006732
rect 360252 1006692 373264 1006720
rect 360252 1006680 360258 1006692
rect 373258 1006680 373264 1006692
rect 373316 1006680 373322 1006732
rect 145742 1006544 145748 1006596
rect 145800 1006584 145806 1006596
rect 153746 1006584 153752 1006596
rect 145800 1006556 153752 1006584
rect 145800 1006544 145806 1006556
rect 153746 1006544 153752 1006556
rect 153804 1006544 153810 1006596
rect 430022 1006476 430028 1006528
rect 430080 1006516 430086 1006528
rect 433978 1006516 433984 1006528
rect 430080 1006488 433984 1006516
rect 430080 1006476 430086 1006488
rect 433978 1006476 433984 1006488
rect 434036 1006476 434042 1006528
rect 93302 1006408 93308 1006460
rect 93360 1006448 93366 1006460
rect 102318 1006448 102324 1006460
rect 93360 1006420 102324 1006448
rect 93360 1006408 93366 1006420
rect 102318 1006408 102324 1006420
rect 102376 1006408 102382 1006460
rect 145558 1006408 145564 1006460
rect 145616 1006448 145622 1006460
rect 152090 1006448 152096 1006460
rect 145616 1006420 152096 1006448
rect 145616 1006408 145622 1006420
rect 152090 1006408 152096 1006420
rect 152148 1006408 152154 1006460
rect 157426 1006408 157432 1006460
rect 157484 1006448 157490 1006460
rect 166258 1006448 166264 1006460
rect 157484 1006420 166264 1006448
rect 157484 1006408 157490 1006420
rect 166258 1006408 166264 1006420
rect 166316 1006408 166322 1006460
rect 171778 1006448 171784 1006460
rect 171106 1006420 171784 1006448
rect 101950 1006312 101956 1006324
rect 94332 1006284 101956 1006312
rect 93118 1006000 93124 1006052
rect 93176 1006040 93182 1006052
rect 94332 1006040 94360 1006284
rect 101950 1006272 101956 1006284
rect 102008 1006272 102014 1006324
rect 144178 1006272 144184 1006324
rect 144236 1006312 144242 1006324
rect 151722 1006312 151728 1006324
rect 144236 1006284 151728 1006312
rect 144236 1006272 144242 1006284
rect 151722 1006272 151728 1006284
rect 151780 1006272 151786 1006324
rect 158254 1006272 158260 1006324
rect 158312 1006312 158318 1006324
rect 171106 1006312 171134 1006420
rect 171778 1006408 171784 1006420
rect 171836 1006408 171842 1006460
rect 206186 1006408 206192 1006460
rect 206244 1006448 206250 1006460
rect 210050 1006448 210056 1006460
rect 206244 1006420 210056 1006448
rect 206244 1006408 206250 1006420
rect 210050 1006408 210056 1006420
rect 210108 1006408 210114 1006460
rect 300302 1006408 300308 1006460
rect 300360 1006448 300366 1006460
rect 306926 1006448 306932 1006460
rect 300360 1006420 306932 1006448
rect 300360 1006408 300366 1006420
rect 306926 1006408 306932 1006420
rect 306984 1006408 306990 1006460
rect 441586 1006448 441614 1006896
rect 505370 1006884 505376 1006936
rect 505428 1006924 505434 1006936
rect 518158 1006924 518164 1006936
rect 505428 1006896 518164 1006924
rect 505428 1006884 505434 1006896
rect 518158 1006884 518164 1006896
rect 518216 1006884 518222 1006936
rect 554774 1006884 554780 1006936
rect 554832 1006924 554838 1006936
rect 569218 1006924 569224 1006936
rect 554832 1006896 569224 1006924
rect 554832 1006884 554838 1006896
rect 569218 1006884 569224 1006896
rect 569276 1006884 569282 1006936
rect 506198 1006748 506204 1006800
rect 506256 1006788 506262 1006800
rect 506256 1006760 509234 1006788
rect 506256 1006748 506262 1006760
rect 509206 1006720 509234 1006760
rect 555970 1006748 555976 1006800
rect 556028 1006788 556034 1006800
rect 565814 1006788 565820 1006800
rect 556028 1006760 565820 1006788
rect 556028 1006748 556034 1006760
rect 565814 1006748 565820 1006760
rect 565872 1006748 565878 1006800
rect 520918 1006720 520924 1006732
rect 509206 1006692 520924 1006720
rect 520918 1006680 520924 1006692
rect 520976 1006680 520982 1006732
rect 447778 1006448 447784 1006460
rect 441586 1006420 447784 1006448
rect 447778 1006408 447784 1006420
rect 447836 1006408 447842 1006460
rect 508222 1006408 508228 1006460
rect 508280 1006448 508286 1006460
rect 508280 1006420 518894 1006448
rect 508280 1006408 508286 1006420
rect 158312 1006284 171134 1006312
rect 158312 1006272 158318 1006284
rect 210418 1006272 210424 1006324
rect 210476 1006312 210482 1006324
rect 228358 1006312 228364 1006324
rect 210476 1006284 228364 1006312
rect 210476 1006272 210482 1006284
rect 228358 1006272 228364 1006284
rect 228416 1006272 228422 1006324
rect 249242 1006272 249248 1006324
rect 249300 1006312 249306 1006324
rect 256142 1006312 256148 1006324
rect 249300 1006284 256148 1006312
rect 249300 1006272 249306 1006284
rect 256142 1006272 256148 1006284
rect 256200 1006272 256206 1006324
rect 298922 1006272 298928 1006324
rect 298980 1006312 298986 1006324
rect 311802 1006312 311808 1006324
rect 298980 1006284 311808 1006312
rect 298980 1006272 298986 1006284
rect 311802 1006272 311808 1006284
rect 311860 1006272 311866 1006324
rect 361390 1006272 361396 1006324
rect 361448 1006312 361454 1006324
rect 375006 1006312 375012 1006324
rect 361448 1006284 375012 1006312
rect 361448 1006272 361454 1006284
rect 375006 1006272 375012 1006284
rect 375064 1006272 375070 1006324
rect 402238 1006272 402244 1006324
rect 402296 1006312 402302 1006324
rect 429194 1006312 429200 1006324
rect 402296 1006284 429200 1006312
rect 402296 1006272 402302 1006284
rect 429194 1006272 429200 1006284
rect 429252 1006272 429258 1006324
rect 434622 1006272 434628 1006324
rect 434680 1006312 434686 1006324
rect 469858 1006312 469864 1006324
rect 434680 1006284 469864 1006312
rect 434680 1006272 434686 1006284
rect 469858 1006272 469864 1006284
rect 469916 1006272 469922 1006324
rect 518866 1006312 518894 1006420
rect 556982 1006408 556988 1006460
rect 557040 1006448 557046 1006460
rect 559650 1006448 559656 1006460
rect 557040 1006420 559656 1006448
rect 557040 1006408 557046 1006420
rect 559650 1006408 559656 1006420
rect 559708 1006408 559714 1006460
rect 522298 1006312 522304 1006324
rect 518866 1006284 522304 1006312
rect 522298 1006272 522304 1006284
rect 522356 1006272 522362 1006324
rect 431678 1006204 431684 1006256
rect 431736 1006244 431742 1006256
rect 431736 1006216 434392 1006244
rect 431736 1006204 431742 1006216
rect 101398 1006136 101404 1006188
rect 101456 1006176 101462 1006188
rect 103974 1006176 103980 1006188
rect 101456 1006148 103980 1006176
rect 101456 1006136 101462 1006148
rect 103974 1006136 103980 1006148
rect 104032 1006136 104038 1006188
rect 107654 1006136 107660 1006188
rect 107712 1006176 107718 1006188
rect 124858 1006176 124864 1006188
rect 107712 1006148 124864 1006176
rect 107712 1006136 107718 1006148
rect 124858 1006136 124864 1006148
rect 124916 1006136 124922 1006188
rect 144730 1006136 144736 1006188
rect 144788 1006176 144794 1006188
rect 150894 1006176 150900 1006188
rect 144788 1006148 150900 1006176
rect 144788 1006136 144794 1006148
rect 150894 1006136 150900 1006148
rect 150952 1006136 150958 1006188
rect 160278 1006136 160284 1006188
rect 160336 1006176 160342 1006188
rect 164878 1006176 164884 1006188
rect 160336 1006148 164884 1006176
rect 160336 1006136 160342 1006148
rect 164878 1006136 164884 1006148
rect 164936 1006136 164942 1006188
rect 166258 1006136 166264 1006188
rect 166316 1006176 166322 1006188
rect 175918 1006176 175924 1006188
rect 166316 1006148 175924 1006176
rect 166316 1006136 166322 1006148
rect 175918 1006136 175924 1006148
rect 175976 1006136 175982 1006188
rect 208394 1006136 208400 1006188
rect 208452 1006176 208458 1006188
rect 208452 1006148 214604 1006176
rect 208452 1006136 208458 1006148
rect 93176 1006012 94360 1006040
rect 93176 1006000 93182 1006012
rect 94498 1006000 94504 1006052
rect 94556 1006040 94562 1006052
rect 98270 1006040 98276 1006052
rect 94556 1006012 98276 1006040
rect 94556 1006000 94562 1006012
rect 98270 1006000 98276 1006012
rect 98328 1006000 98334 1006052
rect 102778 1006000 102784 1006052
rect 102836 1006040 102842 1006052
rect 104802 1006040 104808 1006052
rect 102836 1006012 104808 1006040
rect 102836 1006000 102842 1006012
rect 104802 1006000 104808 1006012
rect 104860 1006000 104866 1006052
rect 108482 1006000 108488 1006052
rect 108540 1006040 108546 1006052
rect 126238 1006040 126244 1006052
rect 108540 1006012 126244 1006040
rect 108540 1006000 108546 1006012
rect 126238 1006000 126244 1006012
rect 126296 1006000 126302 1006052
rect 147582 1006000 147588 1006052
rect 147640 1006040 147646 1006052
rect 150066 1006040 150072 1006052
rect 147640 1006012 150072 1006040
rect 147640 1006000 147646 1006012
rect 150066 1006000 150072 1006012
rect 150124 1006000 150130 1006052
rect 159450 1006000 159456 1006052
rect 159508 1006040 159514 1006052
rect 177298 1006040 177304 1006052
rect 159508 1006012 177304 1006040
rect 159508 1006000 159514 1006012
rect 177298 1006000 177304 1006012
rect 177356 1006000 177362 1006052
rect 196802 1006000 196808 1006052
rect 196860 1006040 196866 1006052
rect 201034 1006040 201040 1006052
rect 196860 1006012 201040 1006040
rect 196860 1006000 196866 1006012
rect 201034 1006000 201040 1006012
rect 201092 1006000 201098 1006052
rect 209222 1006000 209228 1006052
rect 209280 1006040 209286 1006052
rect 211798 1006040 211804 1006052
rect 209280 1006012 211804 1006040
rect 209280 1006000 209286 1006012
rect 211798 1006000 211804 1006012
rect 211856 1006000 211862 1006052
rect 214576 1006040 214604 1006148
rect 249058 1006136 249064 1006188
rect 249116 1006176 249122 1006188
rect 255314 1006176 255320 1006188
rect 249116 1006148 255320 1006176
rect 249116 1006136 249122 1006148
rect 255314 1006136 255320 1006148
rect 255372 1006136 255378 1006188
rect 261846 1006136 261852 1006188
rect 261904 1006176 261910 1006188
rect 279418 1006176 279424 1006188
rect 261904 1006148 279424 1006176
rect 261904 1006136 261910 1006148
rect 279418 1006136 279424 1006148
rect 279476 1006136 279482 1006188
rect 300118 1006136 300124 1006188
rect 300176 1006176 300182 1006188
rect 306098 1006176 306104 1006188
rect 300176 1006148 306104 1006176
rect 300176 1006136 300182 1006148
rect 306098 1006136 306104 1006148
rect 306156 1006136 306162 1006188
rect 357342 1006136 357348 1006188
rect 357400 1006176 357406 1006188
rect 362218 1006176 362224 1006188
rect 357400 1006148 362224 1006176
rect 357400 1006136 357406 1006148
rect 362218 1006136 362224 1006148
rect 362276 1006136 362282 1006188
rect 431494 1006176 431500 1006188
rect 412606 1006148 431500 1006176
rect 229738 1006040 229744 1006052
rect 214576 1006012 229744 1006040
rect 229738 1006000 229744 1006012
rect 229796 1006000 229802 1006052
rect 247034 1006000 247040 1006052
rect 247092 1006040 247098 1006052
rect 252462 1006040 252468 1006052
rect 247092 1006012 252468 1006040
rect 247092 1006000 247098 1006012
rect 252462 1006000 252468 1006012
rect 252520 1006000 252526 1006052
rect 260190 1006000 260196 1006052
rect 260248 1006040 260254 1006052
rect 280798 1006040 280804 1006052
rect 260248 1006012 280804 1006040
rect 260248 1006000 260254 1006012
rect 280798 1006000 280804 1006012
rect 280856 1006000 280862 1006052
rect 298738 1006000 298744 1006052
rect 298796 1006040 298802 1006052
rect 298796 1006012 299474 1006040
rect 298796 1006000 298802 1006012
rect 299446 1005836 299474 1006012
rect 303246 1006000 303252 1006052
rect 303304 1006040 303310 1006052
rect 304074 1006040 304080 1006052
rect 303304 1006012 304080 1006040
rect 303304 1006000 303310 1006012
rect 304074 1006000 304080 1006012
rect 304132 1006000 304138 1006052
rect 314654 1006000 314660 1006052
rect 314712 1006040 314718 1006052
rect 319438 1006040 319444 1006052
rect 314712 1006012 319444 1006040
rect 314712 1006000 314718 1006012
rect 319438 1006000 319444 1006012
rect 319496 1006000 319502 1006052
rect 356882 1006000 356888 1006052
rect 356940 1006040 356946 1006052
rect 360838 1006040 360844 1006052
rect 356940 1006012 360844 1006040
rect 356940 1006000 356946 1006012
rect 360838 1006000 360844 1006012
rect 360896 1006000 360902 1006052
rect 363414 1006000 363420 1006052
rect 363472 1006040 363478 1006052
rect 382918 1006040 382924 1006052
rect 363472 1006012 382924 1006040
rect 363472 1006000 363478 1006012
rect 382918 1006000 382924 1006012
rect 382976 1006000 382982 1006052
rect 400858 1006000 400864 1006052
rect 400916 1006040 400922 1006052
rect 412606 1006040 412634 1006148
rect 431494 1006136 431500 1006148
rect 431552 1006136 431558 1006188
rect 434364 1006176 434392 1006216
rect 434364 1006148 441614 1006176
rect 400916 1006012 412634 1006040
rect 400916 1006000 400922 1006012
rect 428366 1006000 428372 1006052
rect 428424 1006040 428430 1006052
rect 438118 1006040 438124 1006052
rect 428424 1006012 438124 1006040
rect 428424 1006000 428430 1006012
rect 438118 1006000 438124 1006012
rect 438176 1006000 438182 1006052
rect 441586 1006040 441614 1006148
rect 507026 1006136 507032 1006188
rect 507084 1006176 507090 1006188
rect 507084 1006148 518894 1006176
rect 507084 1006136 507090 1006148
rect 471238 1006040 471244 1006052
rect 441586 1006012 471244 1006040
rect 471238 1006000 471244 1006012
rect 471296 1006000 471302 1006052
rect 496722 1006000 496728 1006052
rect 496780 1006040 496786 1006052
rect 498838 1006040 498844 1006052
rect 496780 1006012 498844 1006040
rect 496780 1006000 496786 1006012
rect 498838 1006000 498844 1006012
rect 498896 1006000 498902 1006052
rect 502518 1006000 502524 1006052
rect 502576 1006040 502582 1006052
rect 505738 1006040 505744 1006052
rect 502576 1006012 505744 1006040
rect 502576 1006000 502582 1006012
rect 505738 1006000 505744 1006012
rect 505796 1006000 505802 1006052
rect 509050 1006000 509056 1006052
rect 509108 1006040 509114 1006052
rect 518866 1006040 518894 1006148
rect 556798 1006136 556804 1006188
rect 556856 1006176 556862 1006188
rect 567838 1006176 567844 1006188
rect 556856 1006148 567844 1006176
rect 556856 1006136 556862 1006148
rect 567838 1006136 567844 1006148
rect 567896 1006136 567902 1006188
rect 523678 1006040 523684 1006052
rect 509108 1006012 509234 1006040
rect 518866 1006012 523684 1006040
rect 509108 1006000 509114 1006012
rect 509206 1005972 509234 1006012
rect 523678 1006000 523684 1006012
rect 523736 1006000 523742 1006052
rect 555142 1006000 555148 1006052
rect 555200 1006040 555206 1006052
rect 556430 1006040 556436 1006052
rect 555200 1006012 556436 1006040
rect 555200 1006000 555206 1006012
rect 556430 1006000 556436 1006012
rect 556488 1006000 556494 1006052
rect 557166 1006000 557172 1006052
rect 557224 1006040 557230 1006052
rect 571978 1006040 571984 1006052
rect 557224 1006012 571984 1006040
rect 557224 1006000 557230 1006012
rect 571978 1006000 571984 1006012
rect 572036 1006000 572042 1006052
rect 514018 1005972 514024 1005984
rect 509206 1005944 514024 1005972
rect 514018 1005932 514024 1005944
rect 514076 1005932 514082 1005984
rect 304074 1005836 304080 1005848
rect 299446 1005808 304080 1005836
rect 304074 1005796 304080 1005808
rect 304132 1005796 304138 1005848
rect 425514 1005660 425520 1005712
rect 425572 1005700 425578 1005712
rect 452562 1005700 452568 1005712
rect 425572 1005672 452568 1005700
rect 425572 1005660 425578 1005672
rect 452562 1005660 452568 1005672
rect 452620 1005660 452626 1005712
rect 505002 1005660 505008 1005712
rect 505060 1005700 505066 1005712
rect 515398 1005700 515404 1005712
rect 505060 1005672 515404 1005700
rect 505060 1005660 505066 1005672
rect 515398 1005660 515404 1005672
rect 515456 1005660 515462 1005712
rect 360562 1005524 360568 1005576
rect 360620 1005564 360626 1005576
rect 378778 1005564 378784 1005576
rect 360620 1005536 378784 1005564
rect 360620 1005524 360626 1005536
rect 378778 1005524 378784 1005536
rect 378836 1005524 378842 1005576
rect 427170 1005524 427176 1005576
rect 427228 1005564 427234 1005576
rect 458818 1005564 458824 1005576
rect 427228 1005536 458824 1005564
rect 427228 1005524 427234 1005536
rect 458818 1005524 458824 1005536
rect 458876 1005524 458882 1005576
rect 556430 1005524 556436 1005576
rect 556488 1005564 556494 1005576
rect 573358 1005564 573364 1005576
rect 556488 1005536 573364 1005564
rect 556488 1005524 556494 1005536
rect 573358 1005524 573364 1005536
rect 573416 1005524 573422 1005576
rect 358538 1005388 358544 1005440
rect 358596 1005428 358602 1005440
rect 371878 1005428 371884 1005440
rect 358596 1005400 371884 1005428
rect 358596 1005388 358602 1005400
rect 371878 1005388 371884 1005400
rect 371936 1005388 371942 1005440
rect 428366 1005388 428372 1005440
rect 428424 1005428 428430 1005440
rect 465718 1005428 465724 1005440
rect 428424 1005400 465724 1005428
rect 428424 1005388 428430 1005400
rect 465718 1005388 465724 1005400
rect 465776 1005388 465782 1005440
rect 502150 1005388 502156 1005440
rect 502208 1005428 502214 1005440
rect 519538 1005428 519544 1005440
rect 502208 1005400 519544 1005428
rect 502208 1005388 502214 1005400
rect 519538 1005388 519544 1005400
rect 519596 1005388 519602 1005440
rect 553118 1005388 553124 1005440
rect 553176 1005428 553182 1005440
rect 570598 1005428 570604 1005440
rect 553176 1005400 570604 1005428
rect 553176 1005388 553182 1005400
rect 570598 1005388 570604 1005400
rect 570656 1005388 570662 1005440
rect 149698 1005320 149704 1005372
rect 149756 1005360 149762 1005372
rect 152918 1005360 152924 1005372
rect 149756 1005332 152924 1005360
rect 149756 1005320 149762 1005332
rect 152918 1005320 152924 1005332
rect 152976 1005320 152982 1005372
rect 357710 1005252 357716 1005304
rect 357768 1005292 357774 1005304
rect 376754 1005292 376760 1005304
rect 357768 1005264 376760 1005292
rect 357768 1005252 357774 1005264
rect 376754 1005252 376760 1005264
rect 376812 1005252 376818 1005304
rect 423490 1005252 423496 1005304
rect 423548 1005292 423554 1005304
rect 467098 1005292 467104 1005304
rect 423548 1005264 467104 1005292
rect 423548 1005252 423554 1005264
rect 467098 1005252 467104 1005264
rect 467156 1005252 467162 1005304
rect 499666 1005252 499672 1005304
rect 499724 1005292 499730 1005304
rect 516778 1005292 516784 1005304
rect 499724 1005264 516784 1005292
rect 499724 1005252 499730 1005264
rect 516778 1005252 516784 1005264
rect 516836 1005252 516842 1005304
rect 551462 1005252 551468 1005304
rect 551520 1005292 551526 1005304
rect 574738 1005292 574744 1005304
rect 551520 1005264 574744 1005292
rect 551520 1005252 551526 1005264
rect 574738 1005252 574744 1005264
rect 574796 1005252 574802 1005304
rect 208394 1005116 208400 1005168
rect 208452 1005156 208458 1005168
rect 209866 1005156 209872 1005168
rect 208452 1005128 209872 1005156
rect 208452 1005116 208458 1005128
rect 209866 1005116 209872 1005128
rect 209924 1005116 209930 1005168
rect 149882 1005048 149888 1005100
rect 149940 1005088 149946 1005100
rect 152918 1005088 152924 1005100
rect 149940 1005060 152924 1005088
rect 149940 1005048 149946 1005060
rect 152918 1005048 152924 1005060
rect 152976 1005048 152982 1005100
rect 500494 1005048 500500 1005100
rect 500552 1005088 500558 1005100
rect 508498 1005088 508504 1005100
rect 500552 1005060 508504 1005088
rect 500552 1005048 500558 1005060
rect 508498 1005048 508504 1005060
rect 508556 1005048 508562 1005100
rect 207566 1004980 207572 1005032
rect 207624 1005020 207630 1005032
rect 210050 1005020 210056 1005032
rect 207624 1004992 210056 1005020
rect 207624 1004980 207630 1004992
rect 210050 1004980 210056 1004992
rect 210108 1004980 210114 1005032
rect 151078 1004912 151084 1004964
rect 151136 1004952 151142 1004964
rect 153746 1004952 153752 1004964
rect 151136 1004924 153752 1004952
rect 151136 1004912 151142 1004924
rect 153746 1004912 153752 1004924
rect 153804 1004912 153810 1004964
rect 158622 1004912 158628 1004964
rect 158680 1004952 158686 1004964
rect 162118 1004952 162124 1004964
rect 158680 1004924 162124 1004952
rect 158680 1004912 158686 1004924
rect 162118 1004912 162124 1004924
rect 162176 1004912 162182 1004964
rect 263042 1004912 263048 1004964
rect 263100 1004952 263106 1004964
rect 268378 1004952 268384 1004964
rect 263100 1004924 268384 1004952
rect 263100 1004912 263106 1004924
rect 268378 1004912 268384 1004924
rect 268436 1004912 268442 1004964
rect 313826 1004912 313832 1004964
rect 313884 1004952 313890 1004964
rect 316034 1004952 316040 1004964
rect 313884 1004924 316040 1004952
rect 313884 1004912 313890 1004924
rect 316034 1004912 316040 1004924
rect 316092 1004912 316098 1004964
rect 361390 1004912 361396 1004964
rect 361448 1004952 361454 1004964
rect 364886 1004952 364892 1004964
rect 361448 1004924 364892 1004952
rect 361448 1004912 361454 1004924
rect 364886 1004912 364892 1004924
rect 364944 1004912 364950 1004964
rect 431218 1004912 431224 1004964
rect 431276 1004952 431282 1004964
rect 433518 1004952 433524 1004964
rect 431276 1004924 433524 1004952
rect 431276 1004912 431282 1004924
rect 433518 1004912 433524 1004924
rect 433576 1004912 433582 1004964
rect 160646 1004776 160652 1004828
rect 160704 1004816 160710 1004828
rect 163130 1004816 163136 1004828
rect 160704 1004788 163136 1004816
rect 160704 1004776 160710 1004788
rect 163130 1004776 163136 1004788
rect 163188 1004776 163194 1004828
rect 209222 1004776 209228 1004828
rect 209280 1004816 209286 1004828
rect 211154 1004816 211160 1004828
rect 209280 1004788 211160 1004816
rect 209280 1004776 209286 1004788
rect 211154 1004776 211160 1004788
rect 211212 1004776 211218 1004828
rect 314654 1004776 314660 1004828
rect 314712 1004816 314718 1004828
rect 316678 1004816 316684 1004828
rect 314712 1004788 316684 1004816
rect 314712 1004776 314718 1004788
rect 316678 1004776 316684 1004788
rect 316736 1004776 316742 1004828
rect 353202 1004776 353208 1004828
rect 353260 1004816 353266 1004828
rect 355686 1004816 355692 1004828
rect 353260 1004788 355692 1004816
rect 353260 1004776 353266 1004788
rect 355686 1004776 355692 1004788
rect 355744 1004776 355750 1004828
rect 362586 1004776 362592 1004828
rect 362644 1004816 362650 1004828
rect 365254 1004816 365260 1004828
rect 362644 1004788 365260 1004816
rect 362644 1004776 362650 1004788
rect 365254 1004776 365260 1004788
rect 365312 1004776 365318 1004828
rect 420638 1004776 420644 1004828
rect 420696 1004816 420702 1004828
rect 422662 1004816 422668 1004828
rect 420696 1004788 422668 1004816
rect 420696 1004776 420702 1004788
rect 422662 1004776 422668 1004788
rect 422720 1004776 422726 1004828
rect 432046 1004776 432052 1004828
rect 432104 1004816 432110 1004828
rect 435542 1004816 435548 1004828
rect 432104 1004788 435548 1004816
rect 432104 1004776 432110 1004788
rect 435542 1004776 435548 1004788
rect 435600 1004776 435606 1004828
rect 498102 1004776 498108 1004828
rect 498160 1004816 498166 1004828
rect 500494 1004816 500500 1004828
rect 498160 1004788 500500 1004816
rect 498160 1004776 498166 1004788
rect 500494 1004776 500500 1004788
rect 500552 1004776 500558 1004828
rect 507854 1004776 507860 1004828
rect 507912 1004816 507918 1004828
rect 509694 1004816 509700 1004828
rect 507912 1004788 509700 1004816
rect 507912 1004776 507918 1004788
rect 509694 1004776 509700 1004788
rect 509752 1004776 509758 1004828
rect 555970 1004776 555976 1004828
rect 556028 1004816 556034 1004828
rect 558178 1004816 558184 1004828
rect 556028 1004788 558184 1004816
rect 556028 1004776 556034 1004788
rect 558178 1004776 558184 1004788
rect 558236 1004776 558242 1004828
rect 151262 1004640 151268 1004692
rect 151320 1004680 151326 1004692
rect 154114 1004680 154120 1004692
rect 151320 1004652 154120 1004680
rect 151320 1004640 151326 1004652
rect 154114 1004640 154120 1004652
rect 154172 1004640 154178 1004692
rect 161106 1004640 161112 1004692
rect 161164 1004680 161170 1004692
rect 162946 1004680 162952 1004692
rect 161164 1004652 162952 1004680
rect 161164 1004640 161170 1004652
rect 162946 1004640 162952 1004652
rect 163004 1004640 163010 1004692
rect 212534 1004640 212540 1004692
rect 212592 1004680 212598 1004692
rect 217318 1004680 217324 1004692
rect 212592 1004652 217324 1004680
rect 212592 1004640 212598 1004652
rect 217318 1004640 217324 1004652
rect 217376 1004640 217382 1004692
rect 315482 1004640 315488 1004692
rect 315540 1004680 315546 1004692
rect 318058 1004680 318064 1004692
rect 315540 1004652 318064 1004680
rect 315540 1004640 315546 1004652
rect 318058 1004640 318064 1004652
rect 318116 1004640 318122 1004692
rect 354398 1004640 354404 1004692
rect 354456 1004680 354462 1004692
rect 356514 1004680 356520 1004692
rect 354456 1004652 356520 1004680
rect 354456 1004640 354462 1004652
rect 356514 1004640 356520 1004652
rect 356572 1004640 356578 1004692
rect 364242 1004640 364248 1004692
rect 364300 1004680 364306 1004692
rect 366358 1004680 366364 1004692
rect 364300 1004652 366364 1004680
rect 364300 1004640 364306 1004652
rect 366358 1004640 366364 1004652
rect 366416 1004640 366422 1004692
rect 430022 1004640 430028 1004692
rect 430080 1004680 430086 1004692
rect 431954 1004680 431960 1004692
rect 430080 1004652 431960 1004680
rect 430080 1004640 430086 1004652
rect 431954 1004640 431960 1004652
rect 432012 1004640 432018 1004692
rect 499482 1004640 499488 1004692
rect 499540 1004680 499546 1004692
rect 501322 1004680 501328 1004692
rect 499540 1004652 501328 1004680
rect 499540 1004640 499546 1004652
rect 501322 1004640 501328 1004652
rect 501380 1004640 501386 1004692
rect 507394 1004640 507400 1004692
rect 507452 1004680 507458 1004692
rect 509234 1004680 509240 1004692
rect 507452 1004652 509240 1004680
rect 507452 1004640 507458 1004652
rect 509234 1004640 509240 1004652
rect 509292 1004640 509298 1004692
rect 557626 1004640 557632 1004692
rect 557684 1004680 557690 1004692
rect 559558 1004680 559564 1004692
rect 557684 1004652 559564 1004680
rect 557684 1004640 557690 1004652
rect 559558 1004640 559564 1004652
rect 559616 1004640 559622 1004692
rect 560846 1004640 560852 1004692
rect 560904 1004680 560910 1004692
rect 566458 1004680 566464 1004692
rect 560904 1004652 566464 1004680
rect 560904 1004640 560910 1004652
rect 566458 1004640 566464 1004652
rect 566516 1004640 566522 1004692
rect 424686 1004028 424692 1004080
rect 424744 1004068 424750 1004080
rect 446030 1004068 446036 1004080
rect 424744 1004040 446036 1004068
rect 424744 1004028 424750 1004040
rect 446030 1004028 446036 1004040
rect 446088 1004028 446094 1004080
rect 551094 1004028 551100 1004080
rect 551152 1004068 551158 1004080
rect 564434 1004068 564440 1004080
rect 551152 1004040 564440 1004068
rect 551152 1004028 551158 1004040
rect 564434 1004028 564440 1004040
rect 564492 1004028 564498 1004080
rect 360562 1003892 360568 1003944
rect 360620 1003932 360626 1003944
rect 375374 1003932 375380 1003944
rect 360620 1003904 375380 1003932
rect 360620 1003892 360626 1003904
rect 375374 1003892 375380 1003904
rect 375432 1003892 375438 1003944
rect 426342 1003892 426348 1003944
rect 426400 1003932 426406 1003944
rect 449894 1003932 449900 1003944
rect 426400 1003904 449900 1003932
rect 426400 1003892 426406 1003904
rect 449894 1003892 449900 1003904
rect 449952 1003892 449958 1003944
rect 452562 1003892 452568 1003944
rect 452620 1003932 452626 1003944
rect 460934 1003932 460940 1003944
rect 452620 1003904 460940 1003932
rect 452620 1003892 452626 1003904
rect 460934 1003892 460940 1003904
rect 460992 1003892 460998 1003944
rect 504542 1003892 504548 1003944
rect 504600 1003932 504606 1003944
rect 520274 1003932 520280 1003944
rect 504600 1003904 520280 1003932
rect 504600 1003892 504606 1003904
rect 520274 1003892 520280 1003904
rect 520332 1003892 520338 1003944
rect 552290 1003892 552296 1003944
rect 552348 1003932 552354 1003944
rect 567378 1003932 567384 1003944
rect 552348 1003904 567384 1003932
rect 552348 1003892 552354 1003904
rect 567378 1003892 567384 1003904
rect 567436 1003892 567442 1003944
rect 565814 1003620 565820 1003672
rect 565872 1003660 565878 1003672
rect 568574 1003660 568580 1003672
rect 565872 1003632 568580 1003660
rect 565872 1003620 565878 1003632
rect 568574 1003620 568580 1003632
rect 568632 1003620 568638 1003672
rect 513834 1003348 513840 1003400
rect 513892 1003388 513898 1003400
rect 518894 1003388 518900 1003400
rect 513892 1003360 518900 1003388
rect 513892 1003348 513898 1003360
rect 518894 1003348 518900 1003360
rect 518952 1003348 518958 1003400
rect 355686 1003280 355692 1003332
rect 355744 1003320 355750 1003332
rect 363598 1003320 363604 1003332
rect 355744 1003292 363604 1003320
rect 355744 1003280 355750 1003292
rect 363598 1003280 363604 1003292
rect 363656 1003280 363662 1003332
rect 375006 1003212 375012 1003264
rect 375064 1003252 375070 1003264
rect 379422 1003252 379428 1003264
rect 375064 1003224 379428 1003252
rect 375064 1003212 375070 1003224
rect 379422 1003212 379428 1003224
rect 379480 1003212 379486 1003264
rect 421834 1002668 421840 1002720
rect 421892 1002708 421898 1002720
rect 462958 1002708 462964 1002720
rect 421892 1002680 462964 1002708
rect 421892 1002668 421898 1002680
rect 462958 1002668 462964 1002680
rect 463016 1002668 463022 1002720
rect 97442 1002600 97448 1002652
rect 97500 1002640 97506 1002652
rect 100294 1002640 100300 1002652
rect 97500 1002612 100300 1002640
rect 97500 1002600 97506 1002612
rect 100294 1002600 100300 1002612
rect 100352 1002600 100358 1002652
rect 106826 1002600 106832 1002652
rect 106884 1002640 106890 1002652
rect 109494 1002640 109500 1002652
rect 106884 1002612 109500 1002640
rect 106884 1002600 106890 1002612
rect 109494 1002600 109500 1002612
rect 109552 1002600 109558 1002652
rect 253198 1002600 253204 1002652
rect 253256 1002640 253262 1002652
rect 256142 1002640 256148 1002652
rect 253256 1002612 256148 1002640
rect 253256 1002600 253262 1002612
rect 256142 1002600 256148 1002612
rect 256200 1002600 256206 1002652
rect 558822 1002600 558828 1002652
rect 558880 1002640 558886 1002652
rect 562502 1002640 562508 1002652
rect 558880 1002612 562508 1002640
rect 558880 1002600 558886 1002612
rect 562502 1002600 562508 1002612
rect 562560 1002600 562566 1002652
rect 358538 1002532 358544 1002584
rect 358596 1002572 358602 1002584
rect 371142 1002572 371148 1002584
rect 358596 1002544 371148 1002572
rect 358596 1002532 358602 1002544
rect 371142 1002532 371148 1002544
rect 371200 1002532 371206 1002584
rect 423490 1002532 423496 1002584
rect 423548 1002572 423554 1002584
rect 468478 1002572 468484 1002584
rect 423548 1002544 468484 1002572
rect 423548 1002532 423554 1002544
rect 468478 1002532 468484 1002544
rect 468536 1002532 468542 1002584
rect 92658 1002464 92664 1002516
rect 92716 1002504 92722 1002516
rect 99466 1002504 99472 1002516
rect 92716 1002476 99472 1002504
rect 92716 1002464 92722 1002476
rect 99466 1002464 99472 1002476
rect 99524 1002464 99530 1002516
rect 100018 1002464 100024 1002516
rect 100076 1002504 100082 1002516
rect 103146 1002504 103152 1002516
rect 100076 1002476 103152 1002504
rect 100076 1002464 100082 1002476
rect 103146 1002464 103152 1002476
rect 103204 1002464 103210 1002516
rect 108022 1002464 108028 1002516
rect 108080 1002504 108086 1002516
rect 110690 1002504 110696 1002516
rect 108080 1002476 110696 1002504
rect 108080 1002464 108086 1002476
rect 110690 1002464 110696 1002476
rect 110748 1002464 110754 1002516
rect 153838 1002464 153844 1002516
rect 153896 1002504 153902 1002516
rect 155770 1002504 155776 1002516
rect 153896 1002476 155776 1002504
rect 153896 1002464 153902 1002476
rect 155770 1002464 155776 1002476
rect 155828 1002464 155834 1002516
rect 211246 1002464 211252 1002516
rect 211304 1002504 211310 1002516
rect 215938 1002504 215944 1002516
rect 211304 1002476 215944 1002504
rect 211304 1002464 211310 1002476
rect 215938 1002464 215944 1002476
rect 215996 1002464 216002 1002516
rect 251818 1002464 251824 1002516
rect 251876 1002504 251882 1002516
rect 254486 1002504 254492 1002516
rect 251876 1002476 254492 1002504
rect 251876 1002464 251882 1002476
rect 254486 1002464 254492 1002476
rect 254544 1002464 254550 1002516
rect 560846 1002464 560852 1002516
rect 560904 1002504 560910 1002516
rect 565078 1002504 565084 1002516
rect 560904 1002476 565084 1002504
rect 560904 1002464 560910 1002476
rect 565078 1002464 565084 1002476
rect 565136 1002464 565142 1002516
rect 97258 1002328 97264 1002380
rect 97316 1002368 97322 1002380
rect 100294 1002368 100300 1002380
rect 97316 1002340 100300 1002368
rect 97316 1002328 97322 1002340
rect 100294 1002328 100300 1002340
rect 100352 1002328 100358 1002380
rect 105998 1002328 106004 1002380
rect 106056 1002368 106062 1002380
rect 108298 1002368 108304 1002380
rect 106056 1002340 108304 1002368
rect 106056 1002328 106062 1002340
rect 108298 1002328 108304 1002340
rect 108356 1002328 108362 1002380
rect 156598 1002328 156604 1002380
rect 156656 1002368 156662 1002380
rect 158714 1002368 158720 1002380
rect 156656 1002340 158720 1002368
rect 156656 1002328 156662 1002340
rect 158714 1002328 158720 1002340
rect 158772 1002328 158778 1002380
rect 261018 1002328 261024 1002380
rect 261076 1002368 261082 1002380
rect 264238 1002368 264244 1002380
rect 261076 1002340 264244 1002368
rect 261076 1002328 261082 1002340
rect 264238 1002328 264244 1002340
rect 264296 1002328 264302 1002380
rect 500862 1002328 500868 1002380
rect 500920 1002368 500926 1002380
rect 503346 1002368 503352 1002380
rect 500920 1002340 503352 1002368
rect 500920 1002328 500926 1002340
rect 503346 1002328 503352 1002340
rect 503404 1002328 503410 1002380
rect 557994 1002328 558000 1002380
rect 558052 1002368 558058 1002380
rect 560938 1002368 560944 1002380
rect 558052 1002340 560944 1002368
rect 558052 1002328 558058 1002340
rect 560938 1002328 560944 1002340
rect 560996 1002328 561002 1002380
rect 365070 1002260 365076 1002312
rect 365128 1002300 365134 1002312
rect 367922 1002300 367928 1002312
rect 365128 1002272 367928 1002300
rect 365128 1002260 365134 1002272
rect 367922 1002260 367928 1002272
rect 367980 1002260 367986 1002312
rect 98822 1002192 98828 1002244
rect 98880 1002232 98886 1002244
rect 101122 1002232 101128 1002244
rect 98880 1002204 101128 1002232
rect 98880 1002192 98886 1002204
rect 101122 1002192 101128 1002204
rect 101180 1002192 101186 1002244
rect 105630 1002192 105636 1002244
rect 105688 1002232 105694 1002244
rect 107930 1002232 107936 1002244
rect 105688 1002204 107936 1002232
rect 105688 1002192 105694 1002204
rect 107930 1002192 107936 1002204
rect 107988 1002192 107994 1002244
rect 108850 1002192 108856 1002244
rect 108908 1002232 108914 1002244
rect 112070 1002232 112076 1002244
rect 108908 1002204 112076 1002232
rect 108908 1002192 108914 1002204
rect 112070 1002192 112076 1002204
rect 112128 1002192 112134 1002244
rect 148502 1002192 148508 1002244
rect 148560 1002232 148566 1002244
rect 151722 1002232 151728 1002244
rect 148560 1002204 151728 1002232
rect 148560 1002192 148566 1002204
rect 151722 1002192 151728 1002204
rect 151780 1002192 151786 1002244
rect 155770 1002192 155776 1002244
rect 155828 1002232 155834 1002244
rect 157334 1002232 157340 1002244
rect 155828 1002204 157340 1002232
rect 155828 1002192 155834 1002204
rect 157334 1002192 157340 1002204
rect 157392 1002192 157398 1002244
rect 211246 1002192 211252 1002244
rect 211304 1002232 211310 1002244
rect 213178 1002232 213184 1002244
rect 211304 1002204 213184 1002232
rect 211304 1002192 211310 1002204
rect 213178 1002192 213184 1002204
rect 213236 1002192 213242 1002244
rect 262674 1002192 262680 1002244
rect 262732 1002232 262738 1002244
rect 265802 1002232 265808 1002244
rect 262732 1002204 265808 1002232
rect 262732 1002192 262738 1002204
rect 265802 1002192 265808 1002204
rect 265860 1002192 265866 1002244
rect 357342 1002192 357348 1002244
rect 357400 1002232 357406 1002244
rect 359366 1002232 359372 1002244
rect 357400 1002204 359372 1002232
rect 357400 1002192 357406 1002204
rect 359366 1002192 359372 1002204
rect 359424 1002192 359430 1002244
rect 502242 1002192 502248 1002244
rect 502300 1002232 502306 1002244
rect 504174 1002232 504180 1002244
rect 502300 1002204 504180 1002232
rect 502300 1002192 502306 1002204
rect 504174 1002192 504180 1002204
rect 504232 1002192 504238 1002244
rect 553302 1002192 553308 1002244
rect 553360 1002232 553366 1002244
rect 553946 1002232 553952 1002244
rect 553360 1002204 553952 1002232
rect 553360 1002192 553366 1002204
rect 553946 1002192 553952 1002204
rect 554004 1002192 554010 1002244
rect 560478 1002192 560484 1002244
rect 560536 1002232 560542 1002244
rect 563054 1002232 563060 1002244
rect 560536 1002204 563060 1002232
rect 560536 1002192 560542 1002204
rect 563054 1002192 563060 1002204
rect 563112 1002192 563118 1002244
rect 365898 1002124 365904 1002176
rect 365956 1002164 365962 1002176
rect 369118 1002164 369124 1002176
rect 365956 1002136 369124 1002164
rect 365956 1002124 365962 1002136
rect 369118 1002124 369124 1002136
rect 369176 1002124 369182 1002176
rect 95878 1002056 95884 1002108
rect 95936 1002096 95942 1002108
rect 99098 1002096 99104 1002108
rect 95936 1002068 99104 1002096
rect 95936 1002056 95942 1002068
rect 99098 1002056 99104 1002068
rect 99156 1002056 99162 1002108
rect 101950 1002096 101956 1002108
rect 99484 1002068 101956 1002096
rect 96062 1001920 96068 1001972
rect 96120 1001960 96126 1001972
rect 98270 1001960 98276 1001972
rect 96120 1001932 98276 1001960
rect 96120 1001920 96126 1001932
rect 98270 1001920 98276 1001932
rect 98328 1001920 98334 1001972
rect 98638 1001920 98644 1001972
rect 98696 1001960 98702 1001972
rect 99484 1001960 99512 1002068
rect 101950 1002056 101956 1002068
rect 102008 1002056 102014 1002108
rect 106826 1002056 106832 1002108
rect 106884 1002096 106890 1002108
rect 109034 1002096 109040 1002108
rect 106884 1002068 109040 1002096
rect 106884 1002056 106890 1002068
rect 109034 1002056 109040 1002068
rect 109092 1002056 109098 1002108
rect 109678 1002056 109684 1002108
rect 109736 1002096 109742 1002108
rect 111886 1002096 111892 1002108
rect 109736 1002068 111892 1002096
rect 109736 1002056 109742 1002068
rect 111886 1002056 111892 1002068
rect 111944 1002056 111950 1002108
rect 143994 1002056 144000 1002108
rect 144052 1002096 144058 1002108
rect 147582 1002096 147588 1002108
rect 144052 1002068 147588 1002096
rect 144052 1002056 144058 1002068
rect 147582 1002056 147588 1002068
rect 147640 1002056 147646 1002108
rect 148318 1002056 148324 1002108
rect 148376 1002096 148382 1002108
rect 150894 1002096 150900 1002108
rect 148376 1002068 150900 1002096
rect 148376 1002056 148382 1002068
rect 150894 1002056 150900 1002068
rect 150952 1002056 150958 1002108
rect 155218 1002056 155224 1002108
rect 155276 1002096 155282 1002108
rect 156598 1002096 156604 1002108
rect 155276 1002068 156604 1002096
rect 155276 1002056 155282 1002068
rect 156598 1002056 156604 1002068
rect 156656 1002056 156662 1002108
rect 203518 1002056 203524 1002108
rect 203576 1002096 203582 1002108
rect 206370 1002096 206376 1002108
rect 203576 1002068 206376 1002096
rect 203576 1002056 203582 1002068
rect 206370 1002056 206376 1002068
rect 206428 1002056 206434 1002108
rect 210878 1002056 210884 1002108
rect 210936 1002096 210942 1002108
rect 212534 1002096 212540 1002108
rect 210936 1002068 212540 1002096
rect 210936 1002056 210942 1002068
rect 212534 1002056 212540 1002068
rect 212592 1002056 212598 1002108
rect 252002 1002056 252008 1002108
rect 252060 1002096 252066 1002108
rect 254118 1002096 254124 1002108
rect 252060 1002068 254124 1002096
rect 252060 1002056 252066 1002068
rect 254118 1002056 254124 1002068
rect 254176 1002056 254182 1002108
rect 263870 1002056 263876 1002108
rect 263928 1002096 263934 1002108
rect 266998 1002096 267004 1002108
rect 263928 1002068 267004 1002096
rect 263928 1002056 263934 1002068
rect 266998 1002056 267004 1002068
rect 267056 1002056 267062 1002108
rect 301498 1002056 301504 1002108
rect 301556 1002096 301562 1002108
rect 304902 1002096 304908 1002108
rect 301556 1002068 304908 1002096
rect 301556 1002056 301562 1002068
rect 304902 1002056 304908 1002068
rect 304960 1002056 304966 1002108
rect 310146 1002056 310152 1002108
rect 310204 1002096 310210 1002108
rect 311894 1002096 311900 1002108
rect 310204 1002068 311900 1002096
rect 310204 1002056 310210 1002068
rect 311894 1002056 311900 1002068
rect 311952 1002056 311958 1002108
rect 424502 1002056 424508 1002108
rect 424560 1002096 424566 1002108
rect 425514 1002096 425520 1002108
rect 424560 1002068 425520 1002096
rect 424560 1002056 424566 1002068
rect 425514 1002056 425520 1002068
rect 425572 1002056 425578 1002108
rect 427538 1002056 427544 1002108
rect 427596 1002096 427602 1002108
rect 429838 1002096 429844 1002108
rect 427596 1002068 429844 1002096
rect 427596 1002056 427602 1002068
rect 429838 1002056 429844 1002068
rect 429896 1002056 429902 1002108
rect 433334 1002056 433340 1002108
rect 433392 1002096 433398 1002108
rect 435358 1002096 435364 1002108
rect 433392 1002068 435364 1002096
rect 433392 1002056 433398 1002068
rect 435358 1002056 435364 1002068
rect 435416 1002056 435422 1002108
rect 502518 1002056 502524 1002108
rect 502576 1002096 502582 1002108
rect 503714 1002096 503720 1002108
rect 502576 1002068 503720 1002096
rect 502576 1002056 502582 1002068
rect 503714 1002056 503720 1002068
rect 503772 1002056 503778 1002108
rect 509878 1002056 509884 1002108
rect 509936 1002096 509942 1002108
rect 512822 1002096 512828 1002108
rect 509936 1002068 512828 1002096
rect 509936 1002056 509942 1002068
rect 512822 1002056 512828 1002068
rect 512880 1002056 512886 1002108
rect 560018 1002056 560024 1002108
rect 560076 1002096 560082 1002108
rect 562318 1002096 562324 1002108
rect 560076 1002068 562324 1002096
rect 560076 1002056 560082 1002068
rect 562318 1002056 562324 1002068
rect 562376 1002056 562382 1002108
rect 365070 1001988 365076 1002040
rect 365128 1002028 365134 1002040
rect 367738 1002028 367744 1002040
rect 365128 1002000 367744 1002028
rect 365128 1001988 365134 1002000
rect 367738 1001988 367744 1002000
rect 367796 1001988 367802 1002040
rect 369854 1001988 369860 1002040
rect 369912 1002028 369918 1002040
rect 374638 1002028 374644 1002040
rect 369912 1002000 374644 1002028
rect 369912 1001988 369918 1002000
rect 374638 1001988 374644 1002000
rect 374696 1001988 374702 1002040
rect 423582 1001988 423588 1002040
rect 423640 1002028 423646 1002040
rect 424318 1002028 424324 1002040
rect 423640 1002000 424324 1002028
rect 423640 1001988 423646 1002000
rect 424318 1001988 424324 1002000
rect 424376 1001988 424382 1002040
rect 98696 1001932 99512 1001960
rect 98696 1001920 98702 1001932
rect 100202 1001920 100208 1001972
rect 100260 1001960 100266 1001972
rect 103146 1001960 103152 1001972
rect 100260 1001932 103152 1001960
rect 100260 1001920 100266 1001932
rect 103146 1001920 103152 1001932
rect 103204 1001920 103210 1001972
rect 105998 1001920 106004 1001972
rect 106056 1001960 106062 1001972
rect 107746 1001960 107752 1001972
rect 106056 1001932 107752 1001960
rect 106056 1001920 106062 1001932
rect 107746 1001920 107752 1001932
rect 107804 1001920 107810 1001972
rect 108850 1001920 108856 1001972
rect 108908 1001960 108914 1001972
rect 110506 1001960 110512 1001972
rect 108908 1001932 110512 1001960
rect 108908 1001920 108914 1001932
rect 110506 1001920 110512 1001932
rect 110564 1001920 110570 1001972
rect 146938 1001920 146944 1001972
rect 146996 1001960 147002 1001972
rect 149238 1001960 149244 1001972
rect 146996 1001932 149244 1001960
rect 146996 1001920 147002 1001932
rect 149238 1001920 149244 1001932
rect 149296 1001920 149302 1001972
rect 152458 1001920 152464 1001972
rect 152516 1001960 152522 1001972
rect 154574 1001960 154580 1001972
rect 152516 1001932 154580 1001960
rect 152516 1001920 152522 1001932
rect 154574 1001920 154580 1001932
rect 154632 1001920 154638 1001972
rect 154942 1001920 154948 1001972
rect 155000 1001960 155006 1001972
rect 155954 1001960 155960 1001972
rect 155000 1001932 155960 1001960
rect 155000 1001920 155006 1001932
rect 155954 1001920 155960 1001932
rect 156012 1001920 156018 1001972
rect 157794 1001920 157800 1001972
rect 157852 1001960 157858 1001972
rect 160094 1001960 160100 1001972
rect 157852 1001932 160100 1001960
rect 157852 1001920 157858 1001932
rect 160094 1001920 160100 1001932
rect 160152 1001920 160158 1001972
rect 204162 1001920 204168 1001972
rect 204220 1001960 204226 1001972
rect 205542 1001960 205548 1001972
rect 204220 1001932 205548 1001960
rect 204220 1001920 204226 1001932
rect 205542 1001920 205548 1001932
rect 205600 1001920 205606 1001972
rect 206738 1001920 206744 1001972
rect 206796 1001960 206802 1001972
rect 208394 1001960 208400 1001972
rect 206796 1001932 208400 1001960
rect 206796 1001920 206802 1001932
rect 208394 1001920 208400 1001932
rect 208452 1001920 208458 1001972
rect 212074 1001920 212080 1001972
rect 212132 1001960 212138 1001972
rect 213914 1001960 213920 1001972
rect 212132 1001932 213920 1001960
rect 212132 1001920 212138 1001932
rect 213914 1001920 213920 1001932
rect 213972 1001920 213978 1001972
rect 253382 1001920 253388 1001972
rect 253440 1001960 253446 1001972
rect 255314 1001960 255320 1001972
rect 253440 1001932 255320 1001960
rect 253440 1001920 253446 1001932
rect 255314 1001920 255320 1001932
rect 255372 1001920 255378 1001972
rect 263502 1001920 263508 1001972
rect 263560 1001960 263566 1001972
rect 265618 1001960 265624 1001972
rect 263560 1001932 265624 1001960
rect 263560 1001920 263566 1001932
rect 265618 1001920 265624 1001932
rect 265676 1001920 265682 1001972
rect 310974 1001920 310980 1001972
rect 311032 1001960 311038 1001972
rect 313274 1001960 313280 1001972
rect 311032 1001932 313280 1001960
rect 311032 1001920 311038 1001932
rect 313274 1001920 313280 1001932
rect 313332 1001920 313338 1001972
rect 351822 1001920 351828 1001972
rect 351880 1001960 351886 1001972
rect 354030 1001960 354036 1001972
rect 351880 1001932 354036 1001960
rect 351880 1001920 351886 1001932
rect 354030 1001920 354036 1001932
rect 354088 1001920 354094 1001972
rect 358722 1001920 358728 1001972
rect 358780 1001960 358786 1001972
rect 359366 1001960 359372 1001972
rect 358780 1001932 359372 1001960
rect 358780 1001920 358786 1001932
rect 359366 1001920 359372 1001932
rect 359424 1001920 359430 1001972
rect 419442 1001920 419448 1001972
rect 419500 1001960 419506 1001972
rect 421466 1001960 421472 1001972
rect 419500 1001932 421472 1001960
rect 419500 1001920 419506 1001932
rect 421466 1001920 421472 1001932
rect 421524 1001920 421530 1001972
rect 429194 1001920 429200 1001972
rect 429252 1001960 429258 1001972
rect 431218 1001960 431224 1001972
rect 429252 1001932 431224 1001960
rect 429252 1001920 429258 1001932
rect 431218 1001920 431224 1001932
rect 431276 1001920 431282 1001972
rect 432874 1001920 432880 1001972
rect 432932 1001960 432938 1001972
rect 436738 1001960 436744 1001972
rect 432932 1001932 436744 1001960
rect 432932 1001920 432938 1001932
rect 436738 1001920 436744 1001932
rect 436796 1001920 436802 1001972
rect 496538 1001920 496544 1001972
rect 496596 1001960 496602 1001972
rect 498470 1001960 498476 1001972
rect 496596 1001932 498476 1001960
rect 496596 1001920 496602 1001932
rect 498470 1001920 498476 1001932
rect 498528 1001920 498534 1001972
rect 501690 1001920 501696 1001972
rect 501748 1001960 501754 1001972
rect 502978 1001960 502984 1001972
rect 501748 1001932 502984 1001960
rect 501748 1001920 501754 1001932
rect 502978 1001920 502984 1001932
rect 503036 1001920 503042 1001972
rect 503346 1001920 503352 1001972
rect 503404 1001960 503410 1001972
rect 504358 1001960 504364 1001972
rect 503404 1001932 504364 1001960
rect 503404 1001920 503410 1001932
rect 504358 1001920 504364 1001932
rect 504416 1001920 504422 1001972
rect 510338 1001920 510344 1001972
rect 510396 1001960 510402 1001972
rect 512638 1001960 512644 1001972
rect 510396 1001932 512644 1001960
rect 510396 1001920 510402 1001932
rect 512638 1001920 512644 1001932
rect 512696 1001920 512702 1001972
rect 558822 1001920 558828 1001972
rect 558880 1001960 558886 1001972
rect 560294 1001960 560300 1001972
rect 558880 1001932 560300 1001960
rect 558880 1001920 558886 1001932
rect 560294 1001920 560300 1001932
rect 560352 1001920 560358 1001972
rect 561674 1001920 561680 1001972
rect 561732 1001960 561738 1001972
rect 563698 1001960 563704 1001972
rect 561732 1001932 563704 1001960
rect 561732 1001920 561738 1001932
rect 563698 1001920 563704 1001932
rect 563756 1001920 563762 1001972
rect 354858 1001308 354864 1001360
rect 354916 1001348 354922 1001360
rect 377950 1001348 377956 1001360
rect 354916 1001320 377956 1001348
rect 354916 1001308 354922 1001320
rect 377950 1001308 377956 1001320
rect 378008 1001308 378014 1001360
rect 499482 1001308 499488 1001360
rect 499540 1001348 499546 1001360
rect 516962 1001348 516968 1001360
rect 499540 1001320 516968 1001348
rect 499540 1001308 499546 1001320
rect 516962 1001308 516968 1001320
rect 517020 1001308 517026 1001360
rect 353202 1001172 353208 1001224
rect 353260 1001212 353266 1001224
rect 380894 1001212 380900 1001224
rect 353260 1001184 380900 1001212
rect 353260 1001172 353266 1001184
rect 380894 1001172 380900 1001184
rect 380952 1001172 380958 1001224
rect 429838 1001172 429844 1001224
rect 429896 1001212 429902 1001224
rect 447134 1001212 447140 1001224
rect 429896 1001184 447140 1001212
rect 429896 1001172 429902 1001184
rect 447134 1001172 447140 1001184
rect 447192 1001172 447198 1001224
rect 496538 1001172 496544 1001224
rect 496596 1001212 496602 1001224
rect 522758 1001212 522764 1001224
rect 496596 1001184 522764 1001212
rect 496596 1001172 496602 1001184
rect 522758 1001172 522764 1001184
rect 522816 1001172 522822 1001224
rect 550266 1001172 550272 1001224
rect 550324 1001212 550330 1001224
rect 574094 1001212 574100 1001224
rect 550324 1001184 574100 1001212
rect 550324 1001172 550330 1001184
rect 574094 1001172 574100 1001184
rect 574152 1001172 574158 1001224
rect 449894 1001104 449900 1001156
rect 449952 1001144 449958 1001156
rect 453758 1001144 453764 1001156
rect 449952 1001116 453764 1001144
rect 449952 1001104 449958 1001116
rect 453758 1001104 453764 1001116
rect 453816 1001104 453822 1001156
rect 447778 1000764 447784 1000816
rect 447836 1000804 447842 1000816
rect 449894 1000804 449900 1000816
rect 447836 1000776 449900 1000804
rect 447836 1000764 447842 1000776
rect 449894 1000764 449900 1000776
rect 449952 1000764 449958 1000816
rect 97994 1000492 98000 1000544
rect 98052 1000532 98058 1000544
rect 100202 1000532 100208 1000544
rect 98052 1000504 100208 1000532
rect 98052 1000492 98058 1000504
rect 100202 1000492 100208 1000504
rect 100260 1000492 100266 1000544
rect 447134 1000016 447140 1000068
rect 447192 1000056 447198 1000068
rect 450078 1000056 450084 1000068
rect 447192 1000028 450084 1000056
rect 447192 1000016 447198 1000028
rect 450078 1000016 450084 1000028
rect 450136 1000016 450142 1000068
rect 95142 999132 95148 999184
rect 95200 999172 95206 999184
rect 98822 999172 98828 999184
rect 95200 999144 98828 999172
rect 95200 999132 95206 999144
rect 98822 999132 98828 999144
rect 98880 999132 98886 999184
rect 376754 999132 376760 999184
rect 376812 999172 376818 999184
rect 383378 999172 383384 999184
rect 376812 999144 383384 999172
rect 376812 999132 376818 999144
rect 383378 999132 383384 999144
rect 383436 999132 383442 999184
rect 618162 999132 618168 999184
rect 618220 999172 618226 999184
rect 625522 999172 625528 999184
rect 618220 999144 625528 999172
rect 618220 999132 618226 999144
rect 625522 999132 625528 999144
rect 625580 999132 625586 999184
rect 564434 999064 564440 999116
rect 564492 999104 564498 999116
rect 567930 999104 567936 999116
rect 564492 999076 567936 999104
rect 564492 999064 564498 999076
rect 567930 999064 567936 999076
rect 567988 999064 567994 999116
rect 196618 998792 196624 998844
rect 196676 998832 196682 998844
rect 203886 998832 203892 998844
rect 196676 998804 203892 998832
rect 196676 998792 196682 998804
rect 203886 998792 203892 998804
rect 203944 998792 203950 998844
rect 449894 998792 449900 998844
rect 449952 998832 449958 998844
rect 472618 998832 472624 998844
rect 449952 998804 472624 998832
rect 449952 998792 449958 998804
rect 472618 998792 472624 998804
rect 472676 998792 472682 998844
rect 515398 998792 515404 998844
rect 515456 998832 515462 998844
rect 517146 998832 517152 998844
rect 515456 998804 517152 998832
rect 515456 998792 515462 998804
rect 517146 998792 517152 998804
rect 517204 998792 517210 998844
rect 197998 998656 198004 998708
rect 198056 998696 198062 998708
rect 202690 998696 202696 998708
rect 198056 998668 202696 998696
rect 198056 998656 198062 998668
rect 202690 998656 202696 998668
rect 202748 998656 202754 998708
rect 427078 998656 427084 998708
rect 427136 998696 427142 998708
rect 472434 998696 472440 998708
rect 427136 998668 472440 998696
rect 427136 998656 427142 998668
rect 472434 998656 472440 998668
rect 472492 998656 472498 998708
rect 201034 998520 201040 998572
rect 201092 998560 201098 998572
rect 203886 998560 203892 998572
rect 201092 998532 203892 998560
rect 201092 998520 201098 998532
rect 203886 998520 203892 998532
rect 203944 998520 203950 998572
rect 303246 998520 303252 998572
rect 303304 998560 303310 998572
rect 308950 998560 308956 998572
rect 303304 998532 308956 998560
rect 303304 998520 303310 998532
rect 308950 998520 308956 998532
rect 309008 998520 309014 998572
rect 371878 998520 371884 998572
rect 371936 998560 371942 998572
rect 382734 998560 382740 998572
rect 371936 998532 382740 998560
rect 371936 998520 371942 998532
rect 382734 998520 382740 998532
rect 382792 998520 382798 998572
rect 424502 998520 424508 998572
rect 424560 998560 424566 998572
rect 472250 998560 472256 998572
rect 424560 998532 472256 998560
rect 424560 998520 424566 998532
rect 472250 998520 472256 998532
rect 472308 998520 472314 998572
rect 502242 998520 502248 998572
rect 502300 998560 502306 998572
rect 516502 998560 516508 998572
rect 502300 998532 516508 998560
rect 502300 998520 502306 998532
rect 516502 998520 516508 998532
rect 516560 998520 516566 998572
rect 92290 998384 92296 998436
rect 92348 998424 92354 998436
rect 97994 998424 98000 998436
rect 92348 998396 98000 998424
rect 92348 998384 92354 998396
rect 97994 998384 98000 998396
rect 98052 998384 98058 998436
rect 143718 998384 143724 998436
rect 143776 998424 143782 998436
rect 153838 998424 153844 998436
rect 143776 998396 153844 998424
rect 143776 998384 143782 998396
rect 153838 998384 153844 998396
rect 153896 998384 153902 998436
rect 195238 998384 195244 998436
rect 195296 998424 195302 998436
rect 204162 998424 204168 998436
rect 195296 998396 204168 998424
rect 195296 998384 195302 998396
rect 204162 998384 204168 998396
rect 204220 998384 204226 998436
rect 304258 998384 304264 998436
rect 304316 998424 304322 998436
rect 307294 998424 307300 998436
rect 304316 998396 307300 998424
rect 304316 998384 304322 998396
rect 307294 998384 307300 998396
rect 307352 998384 307358 998436
rect 351822 998384 351828 998436
rect 351880 998424 351886 998436
rect 382274 998424 382280 998436
rect 351880 998396 382280 998424
rect 351880 998384 351886 998396
rect 382274 998384 382280 998396
rect 382332 998384 382338 998436
rect 423582 998384 423588 998436
rect 423640 998424 423646 998436
rect 472066 998424 472072 998436
rect 423640 998396 472072 998424
rect 423640 998384 423646 998396
rect 472066 998384 472072 998396
rect 472124 998384 472130 998436
rect 503714 998384 503720 998436
rect 503772 998424 503778 998436
rect 524046 998424 524052 998436
rect 503772 998396 524052 998424
rect 503772 998384 503778 998396
rect 524046 998384 524052 998396
rect 524104 998384 524110 998436
rect 552290 998384 552296 998436
rect 552348 998424 552354 998436
rect 570782 998424 570788 998436
rect 552348 998396 570788 998424
rect 552348 998384 552354 998396
rect 570782 998384 570788 998396
rect 570840 998384 570846 998436
rect 247218 998248 247224 998300
rect 247276 998288 247282 998300
rect 247276 998260 253934 998288
rect 247276 998248 247282 998260
rect 199378 998112 199384 998164
rect 199436 998152 199442 998164
rect 201862 998152 201868 998164
rect 199436 998124 201868 998152
rect 199436 998112 199442 998124
rect 201862 998112 201868 998124
rect 201920 998112 201926 998164
rect 250438 998112 250444 998164
rect 250496 998152 250502 998164
rect 253658 998152 253664 998164
rect 250496 998124 253664 998152
rect 250496 998112 250502 998124
rect 253658 998112 253664 998124
rect 253716 998112 253722 998164
rect 195790 997976 195796 998028
rect 195848 998016 195854 998028
rect 200666 998016 200672 998028
rect 195848 997988 200672 998016
rect 195848 997976 195854 997988
rect 200666 997976 200672 997988
rect 200724 997976 200730 998028
rect 202322 997976 202328 998028
rect 202380 998016 202386 998028
rect 205542 998016 205548 998028
rect 202380 997988 205548 998016
rect 202380 997976 202386 997988
rect 205542 997976 205548 997988
rect 205600 997976 205606 998028
rect 250622 997908 250628 997960
rect 250680 997948 250686 997960
rect 253658 997948 253664 997960
rect 250680 997920 253664 997948
rect 250680 997908 250686 997920
rect 253658 997908 253664 997920
rect 253716 997908 253722 997960
rect 144178 997840 144184 997892
rect 144236 997880 144242 997892
rect 151262 997880 151268 997892
rect 144236 997852 151268 997880
rect 144236 997840 144242 997852
rect 151262 997840 151268 997852
rect 151320 997840 151326 997892
rect 195422 997840 195428 997892
rect 195480 997880 195486 997892
rect 200022 997880 200028 997892
rect 195480 997852 200028 997880
rect 195480 997840 195486 997852
rect 200022 997840 200028 997852
rect 200080 997840 200086 997892
rect 202138 997840 202144 997892
rect 202196 997880 202202 997892
rect 204714 997880 204720 997892
rect 202196 997852 204720 997880
rect 202196 997840 202202 997852
rect 204714 997840 204720 997852
rect 204772 997840 204778 997892
rect 246574 997840 246580 997892
rect 246632 997880 246638 997892
rect 247034 997880 247040 997892
rect 246632 997852 247040 997880
rect 246632 997840 246638 997852
rect 247034 997840 247040 997852
rect 247092 997840 247098 997892
rect 247678 997772 247684 997824
rect 247736 997812 247742 997824
rect 252462 997812 252468 997824
rect 247736 997784 252468 997812
rect 247736 997772 247742 997784
rect 252462 997772 252468 997784
rect 252520 997772 252526 997824
rect 253906 997812 253934 998260
rect 259362 998248 259368 998300
rect 259420 998288 259426 998300
rect 260926 998288 260932 998300
rect 259420 998260 260932 998288
rect 259420 998248 259426 998260
rect 260926 998248 260932 998260
rect 260984 998248 260990 998300
rect 302878 998248 302884 998300
rect 302936 998288 302942 998300
rect 306098 998288 306104 998300
rect 302936 998260 306104 998288
rect 302936 998248 302942 998260
rect 306098 998248 306104 998260
rect 306156 998248 306162 998300
rect 258166 998112 258172 998164
rect 258224 998152 258230 998164
rect 259454 998152 259460 998164
rect 258224 998124 259460 998152
rect 258224 998112 258230 998124
rect 259454 998112 259460 998124
rect 259512 998112 259518 998164
rect 305638 998112 305644 998164
rect 305696 998152 305702 998164
rect 308122 998152 308128 998164
rect 305696 998124 308128 998152
rect 305696 998112 305702 998124
rect 308122 998112 308128 998124
rect 308180 998112 308186 998164
rect 254762 998044 254768 998096
rect 254820 998084 254826 998096
rect 257338 998084 257344 998096
rect 254820 998056 257344 998084
rect 254820 998044 254826 998056
rect 257338 998044 257344 998056
rect 257396 998044 257402 998096
rect 259822 998044 259828 998096
rect 259880 998084 259886 998096
rect 262306 998084 262312 998096
rect 259880 998056 262312 998084
rect 259880 998044 259886 998056
rect 262306 998044 262312 998056
rect 262364 998044 262370 998096
rect 304442 997976 304448 998028
rect 304500 998016 304506 998028
rect 306926 998016 306932 998028
rect 304500 997988 306932 998016
rect 304500 997976 304506 997988
rect 306926 997976 306932 997988
rect 306984 997976 306990 998028
rect 308398 997976 308404 998028
rect 308456 998016 308462 998028
rect 310606 998016 310612 998028
rect 308456 997988 310612 998016
rect 308456 997976 308462 997988
rect 310606 997976 310612 997988
rect 310664 997976 310670 998028
rect 549162 997976 549168 998028
rect 549220 998016 549226 998028
rect 551462 998016 551468 998028
rect 549220 997988 551468 998016
rect 549220 997976 549226 997988
rect 551462 997976 551468 997988
rect 551520 997976 551526 998028
rect 254578 997908 254584 997960
rect 254636 997948 254642 997960
rect 256510 997948 256516 997960
rect 254636 997920 256516 997948
rect 254636 997908 254642 997920
rect 256510 997908 256516 997920
rect 256568 997908 256574 997960
rect 260190 997908 260196 997960
rect 260248 997948 260254 997960
rect 262490 997948 262496 997960
rect 260248 997920 262496 997948
rect 260248 997908 260254 997920
rect 262490 997908 262496 997920
rect 262548 997908 262554 997960
rect 379422 997908 379428 997960
rect 379480 997948 379486 997960
rect 383194 997948 383200 997960
rect 379480 997920 383200 997948
rect 379480 997908 379486 997920
rect 383194 997908 383200 997920
rect 383252 997908 383258 997960
rect 303062 997840 303068 997892
rect 303120 997880 303126 997892
rect 305270 997880 305276 997892
rect 303120 997852 305276 997880
rect 303120 997840 303126 997852
rect 305270 997840 305276 997852
rect 305328 997840 305334 997892
rect 307018 997840 307024 997892
rect 307076 997880 307082 997892
rect 308950 997880 308956 997892
rect 307076 997852 308956 997880
rect 307076 997840 307082 997852
rect 308950 997840 308956 997852
rect 309008 997840 309014 997892
rect 551554 997840 551560 997892
rect 551612 997880 551618 997892
rect 553118 997880 553124 997892
rect 551612 997852 553124 997880
rect 551612 997840 551618 997852
rect 553118 997840 553124 997852
rect 553176 997840 553182 997892
rect 278130 997812 278136 997824
rect 253906 997784 278136 997812
rect 278130 997772 278136 997784
rect 278188 997772 278194 997824
rect 378778 997772 378784 997824
rect 378836 997812 378842 997824
rect 383562 997812 383568 997824
rect 378836 997784 383568 997812
rect 378836 997772 378842 997784
rect 383562 997772 383568 997784
rect 383620 997772 383626 997824
rect 520274 997772 520280 997824
rect 520332 997812 520338 997824
rect 523862 997812 523868 997824
rect 520332 997784 523868 997812
rect 520332 997772 520338 997784
rect 523862 997772 523868 997784
rect 523920 997772 523926 997824
rect 625706 997812 625712 997824
rect 591316 997784 625712 997812
rect 108298 997704 108304 997756
rect 108356 997744 108362 997756
rect 116302 997744 116308 997756
rect 108356 997716 116308 997744
rect 108356 997704 108362 997716
rect 116302 997704 116308 997716
rect 116360 997704 116366 997756
rect 143810 997704 143816 997756
rect 143868 997744 143874 997756
rect 160094 997744 160100 997756
rect 143868 997716 160100 997744
rect 143868 997704 143874 997716
rect 160094 997704 160100 997716
rect 160152 997704 160158 997756
rect 162118 997704 162124 997756
rect 162176 997744 162182 997756
rect 170306 997744 170312 997756
rect 162176 997716 170312 997744
rect 162176 997704 162182 997716
rect 170306 997704 170312 997716
rect 170364 997704 170370 997756
rect 195606 997704 195612 997756
rect 195664 997744 195670 997756
rect 207014 997744 207020 997756
rect 195664 997716 207020 997744
rect 195664 997704 195670 997716
rect 207014 997704 207020 997716
rect 207072 997704 207078 997756
rect 298738 997704 298744 997756
rect 298796 997744 298802 997756
rect 311894 997744 311900 997756
rect 298796 997716 311900 997744
rect 298796 997704 298802 997716
rect 311894 997704 311900 997716
rect 311952 997704 311958 997756
rect 371142 997704 371148 997756
rect 371200 997744 371206 997756
rect 372522 997744 372528 997756
rect 371200 997716 372528 997744
rect 371200 997704 371206 997716
rect 372522 997704 372528 997716
rect 372580 997704 372586 997756
rect 375374 997704 375380 997756
rect 375432 997744 375438 997756
rect 378594 997744 378600 997756
rect 375432 997716 378600 997744
rect 375432 997704 375438 997716
rect 378594 997704 378600 997716
rect 378652 997704 378658 997756
rect 399938 997704 399944 997756
rect 399996 997744 400002 997756
rect 431954 997744 431960 997756
rect 399996 997716 431960 997744
rect 399996 997704 400002 997716
rect 431954 997704 431960 997716
rect 432012 997704 432018 997756
rect 438118 997704 438124 997756
rect 438176 997744 438182 997756
rect 439866 997744 439872 997756
rect 438176 997716 439872 997744
rect 438176 997704 438182 997716
rect 439866 997704 439872 997716
rect 439924 997704 439930 997756
rect 488994 997704 489000 997756
rect 489052 997744 489058 997756
rect 506474 997744 506480 997756
rect 489052 997716 506480 997744
rect 489052 997704 489058 997716
rect 506474 997704 506480 997716
rect 506532 997704 506538 997756
rect 509694 997704 509700 997756
rect 509752 997744 509758 997756
rect 517330 997744 517336 997756
rect 509752 997716 517336 997744
rect 509752 997704 509758 997716
rect 517330 997704 517336 997716
rect 517388 997704 517394 997756
rect 540882 997704 540888 997756
rect 540940 997744 540946 997756
rect 556982 997744 556988 997756
rect 540940 997716 556988 997744
rect 540940 997704 540946 997716
rect 556982 997704 556988 997716
rect 557040 997704 557046 997756
rect 246942 997636 246948 997688
rect 247000 997676 247006 997688
rect 258074 997676 258080 997688
rect 247000 997648 258080 997676
rect 247000 997636 247006 997648
rect 258074 997636 258080 997648
rect 258132 997636 258138 997688
rect 571978 997636 571984 997688
rect 572036 997676 572042 997688
rect 590562 997676 590568 997688
rect 572036 997648 590568 997676
rect 572036 997636 572042 997648
rect 590562 997636 590568 997648
rect 590620 997636 590626 997688
rect 92474 997568 92480 997620
rect 92532 997608 92538 997620
rect 100018 997608 100024 997620
rect 92532 997580 100024 997608
rect 92532 997568 92538 997580
rect 100018 997568 100024 997580
rect 100076 997568 100082 997620
rect 109494 997568 109500 997620
rect 109552 997608 109558 997620
rect 117222 997608 117228 997620
rect 109552 997580 117228 997608
rect 109552 997568 109558 997580
rect 117222 997568 117228 997580
rect 117280 997568 117286 997620
rect 144822 997568 144828 997620
rect 144880 997608 144886 997620
rect 158714 997608 158720 997620
rect 144880 997580 158720 997608
rect 144880 997568 144886 997580
rect 158714 997568 158720 997580
rect 158772 997568 158778 997620
rect 299382 997568 299388 997620
rect 299440 997608 299446 997620
rect 310514 997608 310520 997620
rect 299440 997580 310520 997608
rect 299440 997568 299446 997580
rect 310514 997568 310520 997580
rect 310572 997568 310578 997620
rect 365254 997568 365260 997620
rect 365312 997608 365318 997620
rect 372338 997608 372344 997620
rect 365312 997580 372344 997608
rect 365312 997568 365318 997580
rect 372338 997568 372344 997580
rect 372396 997568 372402 997620
rect 431218 997568 431224 997620
rect 431276 997608 431282 997620
rect 439682 997608 439688 997620
rect 431276 997580 439688 997608
rect 431276 997568 431282 997580
rect 439682 997568 439688 997580
rect 439740 997568 439746 997620
rect 498102 997568 498108 997620
rect 498160 997608 498166 997620
rect 516870 997608 516876 997620
rect 498160 997580 516876 997608
rect 498160 997568 498166 997580
rect 516870 997568 516876 997580
rect 516928 997568 516934 997620
rect 246758 997500 246764 997552
rect 246816 997540 246822 997552
rect 255958 997540 255964 997552
rect 246816 997512 255964 997540
rect 246816 997500 246822 997512
rect 255958 997500 255964 997512
rect 256016 997500 256022 997552
rect 553302 997500 553308 997552
rect 553360 997540 553366 997552
rect 591316 997540 591344 997784
rect 625706 997772 625712 997784
rect 625764 997772 625770 997824
rect 553360 997512 591344 997540
rect 553360 997500 553366 997512
rect 504358 997432 504364 997484
rect 504416 997472 504422 997484
rect 516686 997472 516692 997484
rect 504416 997444 516692 997472
rect 504416 997432 504422 997444
rect 516686 997432 516692 997444
rect 516744 997432 516750 997484
rect 568574 997364 568580 997416
rect 568632 997404 568638 997416
rect 590378 997404 590384 997416
rect 568632 997376 590384 997404
rect 568632 997364 568638 997376
rect 590378 997364 590384 997376
rect 590436 997364 590442 997416
rect 551554 997296 551560 997348
rect 551612 997336 551618 997348
rect 567562 997336 567568 997348
rect 551612 997308 567568 997336
rect 551612 997296 551618 997308
rect 567562 997296 567568 997308
rect 567620 997296 567626 997348
rect 591298 997296 591304 997348
rect 591356 997336 591362 997348
rect 618162 997336 618168 997348
rect 591356 997308 618168 997336
rect 591356 997296 591362 997308
rect 618162 997296 618168 997308
rect 618220 997296 618226 997348
rect 200206 997228 200212 997280
rect 200264 997268 200270 997280
rect 206186 997268 206192 997280
rect 200264 997240 206192 997268
rect 200264 997228 200270 997240
rect 206186 997228 206192 997240
rect 206244 997228 206250 997280
rect 303246 997228 303252 997280
rect 303304 997268 303310 997280
rect 304442 997268 304448 997280
rect 303304 997240 304448 997268
rect 303304 997228 303310 997240
rect 304442 997228 304448 997240
rect 304500 997228 304506 997280
rect 446030 997228 446036 997280
rect 446088 997268 446094 997280
rect 446088 997240 448744 997268
rect 446088 997228 446094 997240
rect 160738 997160 160744 997212
rect 160796 997200 160802 997212
rect 162946 997200 162952 997212
rect 160796 997172 162952 997200
rect 160796 997160 160802 997172
rect 162946 997160 162952 997172
rect 163004 997160 163010 997212
rect 362218 997160 362224 997212
rect 362276 997200 362282 997212
rect 372706 997200 372712 997212
rect 362276 997172 372712 997200
rect 362276 997160 362282 997172
rect 372706 997160 372712 997172
rect 372764 997160 372770 997212
rect 400122 997092 400128 997144
rect 400180 997132 400186 997144
rect 446122 997132 446128 997144
rect 400180 997104 446128 997132
rect 400180 997092 400186 997104
rect 446122 997092 446128 997104
rect 446180 997092 446186 997144
rect 106918 997024 106924 997076
rect 106976 997064 106982 997076
rect 111886 997064 111892 997076
rect 106976 997036 111892 997064
rect 106976 997024 106982 997036
rect 111886 997024 111892 997036
rect 111944 997024 111950 997076
rect 298370 997024 298376 997076
rect 298428 997064 298434 997076
rect 307202 997064 307208 997076
rect 298428 997036 307208 997064
rect 298428 997024 298434 997036
rect 307202 997024 307208 997036
rect 307260 997024 307266 997076
rect 357342 997024 357348 997076
rect 357400 997064 357406 997076
rect 372338 997064 372344 997076
rect 357400 997036 372344 997064
rect 357400 997024 357406 997036
rect 372338 997024 372344 997036
rect 372396 997024 372402 997076
rect 448716 997064 448744 997240
rect 450078 997160 450084 997212
rect 450136 997200 450142 997212
rect 471882 997200 471888 997212
rect 450136 997172 471888 997200
rect 450136 997160 450142 997172
rect 471882 997160 471888 997172
rect 471940 997160 471946 997212
rect 553486 997160 553492 997212
rect 553544 997200 553550 997212
rect 570138 997200 570144 997212
rect 553544 997172 570144 997200
rect 553544 997160 553550 997172
rect 570138 997160 570144 997172
rect 570196 997160 570202 997212
rect 573358 997160 573364 997212
rect 573416 997200 573422 997212
rect 622394 997200 622400 997212
rect 573416 997172 622400 997200
rect 573416 997160 573422 997172
rect 622394 997160 622400 997172
rect 622452 997160 622458 997212
rect 469214 997064 469220 997076
rect 448716 997036 469220 997064
rect 469214 997024 469220 997036
rect 469272 997024 469278 997076
rect 500862 997024 500868 997076
rect 500920 997064 500926 997076
rect 522942 997064 522948 997076
rect 500920 997036 522948 997064
rect 500920 997024 500926 997036
rect 522942 997024 522948 997036
rect 523000 997024 523006 997076
rect 567378 997024 567384 997076
rect 567436 997064 567442 997076
rect 620278 997064 620284 997076
rect 567436 997036 620284 997064
rect 567436 997024 567442 997036
rect 620278 997024 620284 997036
rect 620336 997024 620342 997076
rect 92474 996956 92480 997008
rect 92532 996996 92538 997008
rect 100754 996996 100760 997008
rect 92532 996968 100760 996996
rect 92532 996956 92538 996968
rect 100754 996956 100760 996968
rect 100812 996956 100818 997008
rect 569218 996888 569224 996940
rect 569276 996928 569282 996940
rect 590562 996928 590568 996940
rect 569276 996900 590568 996928
rect 569276 996888 569282 996900
rect 590562 996888 590568 996900
rect 590620 996888 590626 996940
rect 143810 996684 143816 996736
rect 143868 996724 143874 996736
rect 148502 996724 148508 996736
rect 143868 996696 148508 996724
rect 143868 996684 143874 996696
rect 148502 996684 148508 996696
rect 148560 996684 148566 996736
rect 200758 996684 200764 996736
rect 200816 996724 200822 996736
rect 202506 996724 202512 996736
rect 200816 996696 202512 996724
rect 200816 996684 200822 996696
rect 202506 996684 202512 996696
rect 202564 996684 202570 996736
rect 251634 996684 251640 996736
rect 251692 996724 251698 996736
rect 253382 996724 253388 996736
rect 251692 996696 253388 996724
rect 251692 996684 251698 996696
rect 253382 996684 253388 996696
rect 253440 996684 253446 996736
rect 199378 996384 199384 996396
rect 195624 996356 199384 996384
rect 195624 996260 195652 996356
rect 199378 996344 199384 996356
rect 199436 996344 199442 996396
rect 195606 996208 195612 996260
rect 195664 996208 195670 996260
rect 246942 996208 246948 996260
rect 247000 996248 247006 996260
rect 252002 996248 252008 996260
rect 247000 996220 252008 996248
rect 247000 996208 247006 996220
rect 252002 996208 252008 996220
rect 252060 996208 252066 996260
rect 143994 996072 144000 996124
rect 144052 996112 144058 996124
rect 144052 996084 151814 996112
rect 144052 996072 144058 996084
rect 143810 995976 143816 995988
rect 136468 995948 143816 995976
rect 136468 995852 136496 995948
rect 143810 995936 143816 995948
rect 143868 995936 143874 995988
rect 136450 995800 136456 995852
rect 136508 995800 136514 995852
rect 137738 995800 137744 995852
rect 137796 995840 137802 995852
rect 144638 995840 144644 995852
rect 137796 995812 144644 995840
rect 137796 995800 137802 995812
rect 144638 995800 144644 995812
rect 144696 995800 144702 995852
rect 151786 995840 151814 996084
rect 171778 996072 171784 996124
rect 171836 996112 171842 996124
rect 211154 996112 211160 996124
rect 171836 996084 211160 996112
rect 171836 996072 171842 996084
rect 211154 996072 211160 996084
rect 211212 996072 211218 996124
rect 211798 996072 211804 996124
rect 211856 996112 211862 996124
rect 262490 996112 262496 996124
rect 211856 996084 262496 996112
rect 211856 996072 211862 996084
rect 262490 996072 262496 996084
rect 262548 996072 262554 996124
rect 265802 996072 265808 996124
rect 265860 996112 265866 996124
rect 316034 996112 316040 996124
rect 265860 996084 316040 996112
rect 265860 996072 265866 996084
rect 316034 996072 316040 996084
rect 316092 996072 316098 996124
rect 382918 996072 382924 996124
rect 382976 996112 382982 996124
rect 433518 996112 433524 996124
rect 382976 996084 433524 996112
rect 382976 996072 382982 996084
rect 433518 996072 433524 996084
rect 433576 996072 433582 996124
rect 522298 996072 522304 996124
rect 522356 996112 522362 996124
rect 563054 996112 563060 996124
rect 522356 996084 563060 996112
rect 522356 996072 522362 996084
rect 563054 996072 563060 996084
rect 563112 996072 563118 996124
rect 570598 996072 570604 996124
rect 570656 996112 570662 996124
rect 570656 996084 626534 996112
rect 570656 996072 570662 996084
rect 169386 995936 169392 995988
rect 169444 995976 169450 995988
rect 171502 995976 171508 995988
rect 169444 995948 171508 995976
rect 169444 995936 169450 995948
rect 171502 995936 171508 995948
rect 171560 995936 171566 995988
rect 175918 995936 175924 995988
rect 175976 995976 175982 995988
rect 209866 995976 209872 995988
rect 175976 995948 209872 995976
rect 175976 995936 175982 995948
rect 209866 995936 209872 995948
rect 209924 995936 209930 995988
rect 213178 995936 213184 995988
rect 213236 995976 213242 995988
rect 261110 995976 261116 995988
rect 213236 995948 261116 995976
rect 213236 995936 213242 995948
rect 261110 995936 261116 995948
rect 261168 995936 261174 995988
rect 280798 995936 280804 995988
rect 280856 995976 280862 995988
rect 313274 995976 313280 995988
rect 280856 995948 313280 995976
rect 280856 995936 280862 995948
rect 313274 995936 313280 995948
rect 313332 995936 313338 995988
rect 366358 995936 366364 995988
rect 366416 995976 366422 995988
rect 400858 995976 400864 995988
rect 366416 995948 400864 995976
rect 366416 995936 366422 995948
rect 400858 995936 400864 995948
rect 400916 995936 400922 995988
rect 470566 995948 480254 995976
rect 152458 995840 152464 995852
rect 151786 995812 152464 995840
rect 152458 995800 152464 995812
rect 152516 995800 152522 995852
rect 170674 995800 170680 995852
rect 170732 995840 170738 995852
rect 171686 995840 171692 995852
rect 170732 995812 171692 995840
rect 170732 995800 170738 995812
rect 171686 995800 171692 995812
rect 171744 995800 171750 995852
rect 177298 995800 177304 995852
rect 177356 995840 177362 995852
rect 212534 995840 212540 995852
rect 177356 995812 212540 995840
rect 177356 995800 177362 995812
rect 212534 995800 212540 995812
rect 212592 995800 212598 995852
rect 229738 995800 229744 995852
rect 229796 995840 229802 995852
rect 262306 995840 262312 995852
rect 229796 995812 262312 995840
rect 229796 995800 229802 995812
rect 262306 995800 262312 995812
rect 262364 995800 262370 995852
rect 264238 995800 264244 995852
rect 264296 995840 264302 995852
rect 298922 995840 298928 995852
rect 264296 995812 298928 995840
rect 264296 995800 264302 995812
rect 298922 995800 298928 995812
rect 298980 995800 298986 995852
rect 364886 995800 364892 995852
rect 364944 995840 364950 995852
rect 402238 995840 402244 995852
rect 364944 995812 402244 995840
rect 364944 995800 364950 995812
rect 402238 995800 402244 995812
rect 402296 995800 402302 995852
rect 453758 995800 453764 995852
rect 453816 995840 453822 995852
rect 470566 995840 470594 995948
rect 480226 995908 480254 995948
rect 558178 995936 558184 995988
rect 558236 995976 558242 995988
rect 625890 995976 625896 995988
rect 558236 995948 625896 995976
rect 558236 995936 558242 995948
rect 625890 995936 625896 995948
rect 625948 995936 625954 995988
rect 488902 995908 488908 995920
rect 480226 995880 488908 995908
rect 488902 995868 488908 995880
rect 488960 995868 488966 995920
rect 453816 995812 470594 995840
rect 453816 995800 453822 995812
rect 523678 995800 523684 995852
rect 523736 995840 523742 995852
rect 560294 995840 560300 995852
rect 523736 995812 560300 995840
rect 523736 995800 523742 995812
rect 560294 995800 560300 995812
rect 560352 995800 560358 995852
rect 626506 995840 626534 996084
rect 642082 995908 642088 995920
rect 634786 995880 642088 995908
rect 634786 995840 634814 995880
rect 642082 995868 642088 995880
rect 642140 995868 642146 995920
rect 626506 995812 634814 995840
rect 143442 995528 143448 995580
rect 143500 995568 143506 995580
rect 144178 995568 144184 995580
rect 143500 995540 144184 995568
rect 143500 995528 143506 995540
rect 144178 995528 144184 995540
rect 144236 995528 144242 995580
rect 171042 995528 171048 995580
rect 171100 995568 171106 995580
rect 171100 995540 171916 995568
rect 171100 995528 171106 995540
rect 171888 995415 171916 995540
rect 246206 995528 246212 995580
rect 246264 995568 246270 995580
rect 257338 995568 257344 995580
rect 246264 995540 257344 995568
rect 246264 995528 246270 995540
rect 257338 995528 257344 995540
rect 257396 995528 257402 995580
rect 382734 995528 382740 995580
rect 382792 995568 382798 995580
rect 384942 995568 384948 995580
rect 382792 995540 384948 995568
rect 382792 995528 382798 995540
rect 384942 995528 384948 995540
rect 385000 995528 385006 995580
rect 472618 995528 472624 995580
rect 472676 995568 472682 995580
rect 473354 995568 473360 995580
rect 472676 995540 473360 995568
rect 472676 995528 472682 995540
rect 473354 995528 473360 995540
rect 473412 995528 473418 995580
rect 496814 995528 496820 995580
rect 496872 995568 496878 995580
rect 520182 995568 520188 995580
rect 496872 995540 520188 995568
rect 496872 995528 496878 995540
rect 520182 995528 520188 995540
rect 520240 995528 520246 995580
rect 524046 995528 524052 995580
rect 524104 995568 524110 995580
rect 525334 995568 525340 995580
rect 524104 995540 525340 995568
rect 524104 995528 524110 995540
rect 525334 995528 525340 995540
rect 525392 995528 525398 995580
rect 386690 995460 386696 995512
rect 386748 995500 386754 995512
rect 388622 995500 388628 995512
rect 386748 995472 388628 995500
rect 386748 995460 386754 995472
rect 388622 995460 388628 995472
rect 388680 995460 388686 995512
rect 473814 995460 473820 995512
rect 473872 995500 473878 995512
rect 478230 995500 478236 995512
rect 473872 995472 478236 995500
rect 473872 995460 473878 995472
rect 478230 995460 478236 995472
rect 478288 995460 478294 995512
rect 529566 995460 529572 995512
rect 529624 995500 529630 995512
rect 530210 995500 530216 995512
rect 529624 995472 530216 995500
rect 529624 995460 529630 995472
rect 530210 995460 530216 995472
rect 530268 995460 530274 995512
rect 625890 995460 625896 995512
rect 625948 995500 625954 995512
rect 629662 995500 629668 995512
rect 625948 995472 629668 995500
rect 625948 995460 625954 995472
rect 629662 995460 629668 995472
rect 629720 995460 629726 995512
rect 415394 995392 415400 995444
rect 415452 995432 415458 995444
rect 415452 995404 415716 995432
rect 415452 995392 415458 995404
rect 415688 995387 415716 995404
rect 171686 995277 171692 995329
rect 171744 995277 171750 995329
rect 180702 995324 180708 995376
rect 180760 995364 180766 995376
rect 182634 995364 182640 995376
rect 180760 995336 182640 995364
rect 180760 995324 180766 995336
rect 182634 995324 182640 995336
rect 182692 995324 182698 995376
rect 193122 995324 193128 995376
rect 193180 995364 193186 995376
rect 195054 995364 195060 995376
rect 193180 995336 195060 995364
rect 193180 995324 193186 995336
rect 195054 995324 195060 995336
rect 195112 995324 195118 995376
rect 245562 995324 245568 995376
rect 245620 995364 245626 995376
rect 246758 995364 246764 995376
rect 245620 995336 246764 995364
rect 245620 995324 245626 995336
rect 246758 995324 246764 995336
rect 246816 995324 246822 995376
rect 415688 995359 415978 995387
rect 378134 995256 378140 995308
rect 378192 995296 378198 995308
rect 397638 995296 397644 995308
rect 378192 995268 397644 995296
rect 378192 995256 378198 995268
rect 397638 995256 397644 995268
rect 397696 995256 397702 995308
rect 171502 995165 171508 995217
rect 171560 995165 171566 995217
rect 180472 995188 180478 995240
rect 180530 995228 180536 995240
rect 184658 995228 184664 995240
rect 180530 995200 184664 995228
rect 180530 995188 180536 995200
rect 184658 995188 184664 995200
rect 184716 995188 184722 995240
rect 190362 995188 190368 995240
rect 190420 995228 190426 995240
rect 190546 995228 190552 995240
rect 190420 995200 190552 995228
rect 190420 995188 190426 995200
rect 190546 995188 190552 995200
rect 190604 995188 190610 995240
rect 192478 995188 192484 995240
rect 192536 995228 192542 995240
rect 194134 995228 194140 995240
rect 192536 995200 194140 995228
rect 192536 995188 192542 995200
rect 194134 995188 194140 995200
rect 194192 995188 194198 995240
rect 194318 995188 194324 995240
rect 194376 995228 194382 995240
rect 195238 995228 195244 995240
rect 194376 995200 195244 995228
rect 194376 995188 194382 995200
rect 195238 995188 195244 995200
rect 195296 995188 195302 995240
rect 234936 995188 234942 995240
rect 234994 995228 235000 995240
rect 253198 995228 253204 995240
rect 234994 995200 253204 995228
rect 234994 995188 235000 995200
rect 253198 995188 253204 995200
rect 253256 995188 253262 995240
rect 292482 995188 292488 995240
rect 292540 995228 292546 995240
rect 303062 995228 303068 995240
rect 292540 995200 303068 995228
rect 292540 995188 292546 995200
rect 303062 995188 303068 995200
rect 303120 995188 303126 995240
rect 416130 995235 416136 995287
rect 416188 995235 416194 995287
rect 360838 995120 360844 995172
rect 360896 995160 360902 995172
rect 389634 995160 389640 995172
rect 360896 995132 389640 995160
rect 360896 995120 360902 995132
rect 389634 995120 389640 995132
rect 389692 995120 389698 995172
rect 537754 995120 537760 995172
rect 537812 995160 537818 995172
rect 538398 995160 538404 995172
rect 537812 995132 538404 995160
rect 537812 995120 537818 995132
rect 538398 995120 538404 995132
rect 538456 995120 538462 995172
rect 172422 995092 172428 995104
rect 171428 995064 172428 995092
rect 172422 995052 172428 995064
rect 172480 995052 172486 995104
rect 181438 995052 181444 995104
rect 181496 995092 181502 995104
rect 210050 995092 210056 995104
rect 181496 995064 210056 995092
rect 181496 995052 181502 995064
rect 210050 995052 210056 995064
rect 210108 995052 210114 995104
rect 234522 995052 234528 995104
rect 234580 995092 234586 995104
rect 259454 995092 259460 995104
rect 234580 995064 259460 995092
rect 234580 995052 234586 995064
rect 259454 995052 259460 995064
rect 259512 995052 259518 995104
rect 283466 995052 283472 995104
rect 283524 995092 283530 995104
rect 305638 995092 305644 995104
rect 283524 995064 305644 995092
rect 283524 995052 283530 995064
rect 305638 995052 305644 995064
rect 305696 995052 305702 995104
rect 425698 995052 425704 995104
rect 425756 995092 425762 995104
rect 484118 995092 484124 995104
rect 425756 995064 484124 995092
rect 425756 995052 425762 995064
rect 484118 995052 484124 995064
rect 484176 995052 484182 995104
rect 505738 995052 505744 995104
rect 505796 995092 505802 995104
rect 528738 995092 528744 995104
rect 505796 995064 528744 995092
rect 505796 995052 505802 995064
rect 528738 995052 528744 995064
rect 528796 995052 528802 995104
rect 567562 995052 567568 995104
rect 567620 995092 567626 995104
rect 637022 995092 637028 995104
rect 567620 995064 637028 995092
rect 567620 995052 567626 995064
rect 637022 995052 637028 995064
rect 637080 995052 637086 995104
rect 358722 994984 358728 995036
rect 358780 995024 358786 995036
rect 398834 995024 398840 995036
rect 358780 994996 398840 995024
rect 358780 994984 358786 994996
rect 398834 994984 398840 994996
rect 398892 994984 398898 995036
rect 660408 995024 660436 995121
rect 643066 994996 660436 995024
rect 171244 994881 171272 994967
rect 180702 994916 180708 994968
rect 180760 994956 180766 994968
rect 208394 994956 208400 994968
rect 180760 994928 208400 994956
rect 180760 994916 180766 994928
rect 208394 994916 208400 994928
rect 208452 994916 208458 994968
rect 232866 994916 232872 994968
rect 232924 994956 232930 994968
rect 260926 994956 260932 994968
rect 232924 994928 260932 994956
rect 232924 994916 232930 994928
rect 260926 994916 260932 994928
rect 260984 994916 260990 994968
rect 284110 994916 284116 994968
rect 284168 994956 284174 994968
rect 308398 994956 308404 994968
rect 284168 994928 308404 994956
rect 284168 994916 284174 994928
rect 308398 994916 308404 994928
rect 308456 994916 308462 994968
rect 419442 994916 419448 994968
rect 419500 994956 419506 994968
rect 643066 994956 643094 994996
rect 660574 994983 660580 995035
rect 660632 994983 660638 995035
rect 419500 994928 643094 994956
rect 419500 994916 419506 994928
rect 80146 994780 80152 994832
rect 80204 994820 80210 994832
rect 103514 994820 103520 994832
rect 80204 994792 103520 994820
rect 80204 994780 80210 994792
rect 103514 994780 103520 994792
rect 103572 994780 103578 994832
rect 128446 994780 128452 994832
rect 128504 994820 128510 994832
rect 157334 994820 157340 994832
rect 128504 994792 157340 994820
rect 128504 994780 128510 994792
rect 157334 994780 157340 994792
rect 157392 994780 157398 994832
rect 170858 994829 170864 994881
rect 170916 994829 170922 994881
rect 171226 994829 171232 994881
rect 171284 994829 171290 994881
rect 372706 994848 372712 994900
rect 372764 994888 372770 994900
rect 393314 994888 393320 994900
rect 372764 994860 393320 994888
rect 372764 994848 372770 994860
rect 393314 994848 393320 994860
rect 393372 994848 393378 994900
rect 287146 994780 287152 994832
rect 287204 994820 287210 994832
rect 304258 994820 304264 994832
rect 287204 994792 304264 994820
rect 287204 994780 287210 994792
rect 304258 994780 304264 994792
rect 304316 994780 304322 994832
rect 433978 994780 433984 994832
rect 434036 994820 434042 994832
rect 509234 994820 509240 994832
rect 434036 994792 509240 994820
rect 434036 994780 434042 994792
rect 509234 994780 509240 994792
rect 509292 994780 509298 994832
rect 523862 994780 523868 994832
rect 523920 994820 523926 994832
rect 527910 994820 527916 994832
rect 523920 994792 527916 994820
rect 523920 994780 523926 994792
rect 527910 994780 527916 994792
rect 527968 994780 527974 994832
rect 529014 994780 529020 994832
rect 529072 994820 529078 994832
rect 538214 994820 538220 994832
rect 529072 994792 538220 994820
rect 529072 994780 529078 994792
rect 538214 994780 538220 994792
rect 538272 994780 538278 994832
rect 567930 994780 567936 994832
rect 567988 994820 567994 994832
rect 567988 994792 625154 994820
rect 567988 994780 567994 994792
rect 169386 994712 169392 994764
rect 169444 994752 169450 994764
rect 247678 994752 247684 994764
rect 169444 994724 247684 994752
rect 169444 994712 169450 994724
rect 247678 994712 247684 994724
rect 247736 994712 247742 994764
rect 378594 994712 378600 994764
rect 378652 994752 378658 994764
rect 396994 994752 397000 994764
rect 378652 994724 397000 994752
rect 378652 994712 378658 994724
rect 396994 994712 397000 994724
rect 397052 994712 397058 994764
rect 77662 994644 77668 994696
rect 77720 994684 77726 994696
rect 93302 994684 93308 994696
rect 77720 994656 93308 994684
rect 77720 994644 77726 994656
rect 93302 994644 93308 994656
rect 93360 994644 93366 994696
rect 104894 994644 104900 994696
rect 104952 994684 104958 994696
rect 110506 994684 110512 994696
rect 104952 994656 110512 994684
rect 104952 994644 104958 994656
rect 110506 994644 110512 994656
rect 110564 994644 110570 994696
rect 131574 994644 131580 994696
rect 131632 994684 131638 994696
rect 155954 994684 155960 994696
rect 131632 994656 155960 994684
rect 131632 994644 131638 994656
rect 155954 994644 155960 994656
rect 156012 994644 156018 994696
rect 420638 994644 420644 994696
rect 420696 994684 420702 994696
rect 590562 994684 590568 994696
rect 420696 994656 590568 994684
rect 420696 994644 420702 994656
rect 590562 994644 590568 994656
rect 590620 994644 590626 994696
rect 625126 994684 625154 994792
rect 625706 994780 625712 994832
rect 625764 994820 625770 994832
rect 630858 994820 630864 994832
rect 625764 994792 630864 994820
rect 625764 994780 625770 994792
rect 630858 994780 630864 994792
rect 630916 994780 630922 994832
rect 639506 994684 639512 994696
rect 625126 994656 639512 994684
rect 639506 994644 639512 994656
rect 639564 994644 639570 994696
rect 660776 994628 660804 994897
rect 171042 994576 171048 994628
rect 171100 994616 171106 994628
rect 298554 994616 298560 994628
rect 171100 994588 298560 994616
rect 171100 994576 171106 994588
rect 298554 994576 298560 994588
rect 298612 994576 298618 994628
rect 363598 994576 363604 994628
rect 363656 994616 363662 994628
rect 393958 994616 393964 994628
rect 363656 994588 393964 994616
rect 363656 994576 363662 994588
rect 393958 994576 393964 994588
rect 394016 994576 394022 994628
rect 660758 994576 660764 994628
rect 660816 994576 660822 994628
rect 660960 994560 660988 994785
rect 78306 994508 78312 994560
rect 78364 994548 78370 994560
rect 102778 994548 102784 994560
rect 78364 994520 102784 994548
rect 78364 994508 78370 994520
rect 102778 994508 102784 994520
rect 102836 994508 102842 994560
rect 129734 994508 129740 994560
rect 129792 994548 129798 994560
rect 155310 994548 155316 994560
rect 129792 994520 155316 994548
rect 129792 994508 129798 994520
rect 155310 994508 155316 994520
rect 155368 994508 155374 994560
rect 462958 994508 462964 994560
rect 463016 994548 463022 994560
rect 474642 994548 474648 994560
rect 463016 994520 474648 994548
rect 463016 994508 463022 994520
rect 474642 994508 474648 994520
rect 474700 994508 474706 994560
rect 485958 994548 485964 994560
rect 474844 994520 485964 994548
rect 180150 994440 180156 994492
rect 180208 994480 180214 994492
rect 207382 994480 207388 994492
rect 180208 994452 207388 994480
rect 180208 994440 180214 994452
rect 207382 994440 207388 994452
rect 207440 994440 207446 994492
rect 235902 994440 235908 994492
rect 235960 994480 235966 994492
rect 243722 994480 243728 994492
rect 235960 994452 243728 994480
rect 235960 994440 235966 994452
rect 243722 994440 243728 994452
rect 243780 994440 243786 994492
rect 354398 994440 354404 994492
rect 354456 994480 354462 994492
rect 392670 994480 392676 994492
rect 354456 994452 392676 994480
rect 354456 994440 354462 994452
rect 392670 994440 392676 994452
rect 392728 994440 392734 994492
rect 80698 994372 80704 994424
rect 80756 994412 80762 994424
rect 93118 994412 93124 994424
rect 80756 994384 93124 994412
rect 80756 994372 80762 994384
rect 93118 994372 93124 994384
rect 93176 994372 93182 994424
rect 132126 994372 132132 994424
rect 132184 994412 132190 994424
rect 145742 994412 145748 994424
rect 132184 994384 145748 994412
rect 132184 994372 132190 994384
rect 145742 994372 145748 994384
rect 145800 994372 145806 994424
rect 278130 994372 278136 994424
rect 278188 994412 278194 994424
rect 316402 994412 316408 994424
rect 278188 994384 316408 994412
rect 278188 994372 278194 994384
rect 316402 994372 316408 994384
rect 316460 994372 316466 994424
rect 465718 994372 465724 994424
rect 465776 994412 465782 994424
rect 474844 994412 474872 994520
rect 485958 994508 485964 994520
rect 486016 994508 486022 994560
rect 508498 994508 508504 994560
rect 508556 994548 508562 994560
rect 534350 994548 534356 994560
rect 508556 994520 534356 994548
rect 508556 994508 508562 994520
rect 534350 994508 534356 994520
rect 534408 994508 534414 994560
rect 567746 994508 567752 994560
rect 567804 994548 567810 994560
rect 639046 994548 639052 994560
rect 567804 994520 639052 994548
rect 567804 994508 567810 994520
rect 639046 994508 639052 994520
rect 639104 994508 639110 994560
rect 660942 994508 660948 994560
rect 661000 994508 661006 994560
rect 486602 994412 486608 994424
rect 465776 994384 474872 994412
rect 480226 994384 486608 994412
rect 465776 994372 465782 994384
rect 184658 994304 184664 994356
rect 184716 994344 184722 994356
rect 202322 994344 202328 994356
rect 184716 994316 202328 994344
rect 184716 994304 184722 994316
rect 202322 994304 202328 994316
rect 202380 994304 202386 994356
rect 231578 994304 231584 994356
rect 231636 994344 231642 994356
rect 243354 994344 243360 994356
rect 231636 994316 243360 994344
rect 231636 994304 231642 994316
rect 243354 994304 243360 994316
rect 243412 994304 243418 994356
rect 243538 994304 243544 994356
rect 243596 994344 243602 994356
rect 254578 994344 254584 994356
rect 243596 994316 254584 994344
rect 243596 994304 243602 994316
rect 254578 994304 254584 994316
rect 254636 994304 254642 994356
rect 88978 994236 88984 994288
rect 89036 994276 89042 994288
rect 121730 994276 121736 994288
rect 89036 994248 121736 994276
rect 89036 994236 89042 994248
rect 121730 994236 121736 994248
rect 121788 994236 121794 994288
rect 294138 994236 294144 994288
rect 294196 994276 294202 994288
rect 381170 994276 381176 994288
rect 294196 994248 381176 994276
rect 294196 994236 294202 994248
rect 381170 994236 381176 994248
rect 381228 994236 381234 994288
rect 474642 994236 474648 994288
rect 474700 994276 474706 994288
rect 480226 994276 480254 994384
rect 486602 994372 486608 994384
rect 486660 994372 486666 994424
rect 502978 994372 502984 994424
rect 503036 994412 503042 994424
rect 533706 994412 533712 994424
rect 503036 994384 533712 994412
rect 503036 994372 503042 994384
rect 533706 994372 533712 994384
rect 533764 994372 533770 994424
rect 570138 994372 570144 994424
rect 570196 994412 570202 994424
rect 591298 994412 591304 994424
rect 570196 994384 591304 994412
rect 570196 994372 570202 994384
rect 591298 994372 591304 994384
rect 591356 994372 591362 994424
rect 625522 994372 625528 994424
rect 625580 994412 625586 994424
rect 630214 994412 630220 994424
rect 625580 994384 630220 994412
rect 625580 994372 625586 994384
rect 630214 994372 630220 994384
rect 630272 994372 630278 994424
rect 474700 994248 480254 994276
rect 474700 994236 474706 994248
rect 494054 994236 494060 994288
rect 494112 994276 494118 994288
rect 511074 994276 511080 994288
rect 494112 994248 511080 994276
rect 494112 994236 494118 994248
rect 511074 994236 511080 994248
rect 511132 994236 511138 994288
rect 518158 994236 518164 994288
rect 518216 994276 518222 994288
rect 518216 994248 529244 994276
rect 518216 994236 518222 994248
rect 170674 994100 170680 994152
rect 170732 994140 170738 994152
rect 301498 994140 301504 994152
rect 170732 994112 301504 994140
rect 170732 994100 170738 994112
rect 301498 994100 301504 994112
rect 301556 994100 301562 994152
rect 519538 994100 519544 994152
rect 519596 994140 519602 994152
rect 529014 994140 529020 994152
rect 519596 994112 529020 994140
rect 519596 994100 519602 994112
rect 529014 994100 529020 994112
rect 529072 994100 529078 994152
rect 529216 994140 529244 994248
rect 529382 994236 529388 994288
rect 529440 994276 529446 994288
rect 539226 994276 539232 994288
rect 529440 994248 539232 994276
rect 529440 994236 529446 994248
rect 539226 994236 539232 994248
rect 539284 994236 539290 994288
rect 538398 994140 538404 994152
rect 529216 994112 538404 994140
rect 538398 994100 538404 994112
rect 538456 994100 538462 994152
rect 574094 994032 574100 994084
rect 574152 994072 574158 994084
rect 661144 994072 661172 994673
rect 574152 994044 661172 994072
rect 574152 994032 574158 994044
rect 232222 993964 232228 994016
rect 232280 994004 232286 994016
rect 243538 994004 243544 994016
rect 232280 993976 243544 994004
rect 232280 993964 232286 993976
rect 243538 993964 243544 993976
rect 243596 993964 243602 994016
rect 243722 993964 243728 994016
rect 243780 994004 243786 994016
rect 249242 994004 249248 994016
rect 243780 993976 249248 994004
rect 243780 993964 243786 993976
rect 249242 993964 249248 993976
rect 249300 993964 249306 994016
rect 286502 993964 286508 994016
rect 286560 994004 286566 994016
rect 298370 994004 298376 994016
rect 286560 993976 298376 994004
rect 286560 993964 286566 993976
rect 298370 993964 298376 993976
rect 298428 993964 298434 994016
rect 522942 993964 522948 994016
rect 523000 994004 523006 994016
rect 529382 994004 529388 994016
rect 523000 993976 529388 994004
rect 523000 993964 523006 993976
rect 529382 993964 529388 993976
rect 529440 993964 529446 994016
rect 142062 993896 142068 993948
rect 142120 993936 142126 993948
rect 142338 993936 142344 993948
rect 142120 993908 142344 993936
rect 142120 993896 142126 993908
rect 142338 993896 142344 993908
rect 142396 993896 142402 993948
rect 574738 993896 574744 993948
rect 574796 993936 574802 993948
rect 661328 993936 661356 994561
rect 574796 993908 661356 993936
rect 574796 993896 574802 993908
rect 243354 993828 243360 993880
rect 243412 993868 243418 993880
rect 246206 993868 246212 993880
rect 243412 993840 246212 993868
rect 243412 993828 243418 993840
rect 246206 993828 246212 993840
rect 246264 993828 246270 993880
rect 171226 993760 171232 993812
rect 171284 993800 171290 993812
rect 195790 993800 195796 993812
rect 171284 993772 195796 993800
rect 171284 993760 171290 993772
rect 195790 993760 195796 993772
rect 195848 993760 195854 993812
rect 522758 993760 522764 993812
rect 522816 993800 522822 993812
rect 660758 993800 660764 993812
rect 522816 993772 660764 993800
rect 522816 993760 522822 993772
rect 660758 993760 660764 993772
rect 660816 993760 660822 993812
rect 142062 993692 142068 993744
rect 142120 993732 142126 993744
rect 142120 993692 142154 993732
rect 142126 993664 142154 993692
rect 142246 993664 142252 993676
rect 142126 993636 142252 993664
rect 142246 993624 142252 993636
rect 142304 993624 142310 993676
rect 170858 993624 170864 993676
rect 170916 993664 170922 993676
rect 195606 993664 195612 993676
rect 170916 993636 195612 993664
rect 170916 993624 170922 993636
rect 195606 993624 195612 993636
rect 195664 993624 195670 993676
rect 516318 993624 516324 993676
rect 516376 993664 516382 993676
rect 660942 993664 660948 993676
rect 516376 993636 660948 993664
rect 516376 993624 516382 993636
rect 660942 993624 660948 993636
rect 661000 993624 661006 993676
rect 549162 993488 549168 993540
rect 549220 993528 549226 993540
rect 635826 993528 635832 993540
rect 549220 993500 635832 993528
rect 549220 993488 549226 993500
rect 635826 993488 635832 993500
rect 635884 993488 635890 993540
rect 554774 993352 554780 993404
rect 554832 993392 554838 993404
rect 640702 993392 640708 993404
rect 554832 993364 640708 993392
rect 554832 993352 554838 993364
rect 640702 993352 640708 993364
rect 640760 993352 640766 993404
rect 51718 993148 51724 993200
rect 51776 993188 51782 993200
rect 107930 993188 107936 993200
rect 51776 993160 107936 993188
rect 51776 993148 51782 993160
rect 107930 993148 107936 993160
rect 107988 993148 107994 993200
rect 50338 993012 50344 993064
rect 50396 993052 50402 993064
rect 107746 993052 107752 993064
rect 50396 993024 107752 993052
rect 50396 993012 50402 993024
rect 107746 993012 107752 993024
rect 107804 993012 107810 993064
rect 563698 993012 563704 993064
rect 563756 993052 563762 993064
rect 608594 993052 608600 993064
rect 563756 993024 608600 993052
rect 563756 993012 563762 993024
rect 608594 993012 608600 993024
rect 608652 993012 608658 993064
rect 55858 992876 55864 992928
rect 55916 992916 55922 992928
rect 146938 992916 146944 992928
rect 55916 992888 146944 992916
rect 55916 992876 55922 992888
rect 146938 992876 146944 992888
rect 146996 992876 147002 992928
rect 147674 992876 147680 992928
rect 147732 992916 147738 992928
rect 186498 992916 186504 992928
rect 147732 992888 186504 992916
rect 147732 992876 147738 992888
rect 186498 992876 186504 992888
rect 186556 992876 186562 992928
rect 202874 992876 202880 992928
rect 202932 992916 202938 992928
rect 213914 992916 213920 992928
rect 202932 992888 213920 992916
rect 202932 992876 202938 992888
rect 213914 992876 213920 992888
rect 213972 992876 213978 992928
rect 316678 992876 316684 992928
rect 316736 992916 316742 992928
rect 364978 992916 364984 992928
rect 316736 992888 364984 992916
rect 316736 992876 316742 992888
rect 364978 992876 364984 992888
rect 365036 992876 365042 992928
rect 367922 992876 367928 992928
rect 367980 992916 367986 992928
rect 429930 992916 429936 992928
rect 367980 992888 429936 992916
rect 367980 992876 367986 992888
rect 429930 992876 429936 992888
rect 429988 992876 429994 992928
rect 435542 992876 435548 992928
rect 435600 992916 435606 992928
rect 494698 992916 494704 992928
rect 435600 992888 494704 992916
rect 435600 992876 435606 992888
rect 494698 992876 494704 992888
rect 494756 992876 494762 992928
rect 512822 992876 512828 992928
rect 512880 992916 512886 992928
rect 527266 992916 527272 992928
rect 512880 992888 527272 992916
rect 512880 992876 512886 992888
rect 527266 992876 527272 992888
rect 527324 992876 527330 992928
rect 562502 992876 562508 992928
rect 562560 992916 562566 992928
rect 667198 992916 667204 992928
rect 562560 992888 667204 992916
rect 562560 992876 562566 992888
rect 667198 992876 667204 992888
rect 667256 992876 667262 992928
rect 638862 992264 638868 992316
rect 638920 992304 638926 992316
rect 640794 992304 640800 992316
rect 638920 992276 640800 992304
rect 638920 992264 638926 992276
rect 640794 992264 640800 992276
rect 640852 992264 640858 992316
rect 47578 991720 47584 991772
rect 47636 991760 47642 991772
rect 96062 991760 96068 991772
rect 47636 991732 96068 991760
rect 47636 991720 47642 991732
rect 96062 991720 96068 991732
rect 96120 991720 96126 991772
rect 48958 991584 48964 991636
rect 49016 991624 49022 991636
rect 110690 991624 110696 991636
rect 49016 991596 110696 991624
rect 49016 991584 49022 991596
rect 110690 991584 110696 991596
rect 110748 991584 110754 991636
rect 138290 991584 138296 991636
rect 138348 991624 138354 991636
rect 163130 991624 163136 991636
rect 138348 991596 163136 991624
rect 138348 991584 138354 991596
rect 163130 991584 163136 991596
rect 163188 991584 163194 991636
rect 54478 991448 54484 991500
rect 54536 991488 54542 991500
rect 148318 991488 148324 991500
rect 54536 991460 148324 991488
rect 54536 991448 54542 991460
rect 148318 991448 148324 991460
rect 148376 991448 148382 991500
rect 266998 991448 267004 991500
rect 267056 991488 267062 991500
rect 284294 991488 284300 991500
rect 267056 991460 284300 991488
rect 267056 991448 267062 991460
rect 284294 991448 284300 991460
rect 284352 991448 284358 991500
rect 318058 991448 318064 991500
rect 318116 991488 318122 991500
rect 349154 991488 349160 991500
rect 318116 991460 349160 991488
rect 318116 991448 318122 991460
rect 349154 991448 349160 991460
rect 349212 991448 349218 991500
rect 367738 991448 367744 991500
rect 367796 991488 367802 991500
rect 397822 991488 397828 991500
rect 367796 991460 397828 991488
rect 367796 991448 367802 991460
rect 397822 991448 397828 991460
rect 397880 991448 397886 991500
rect 435358 991448 435364 991500
rect 435416 991488 435422 991500
rect 478966 991488 478972 991500
rect 435416 991460 478972 991488
rect 435416 991448 435422 991460
rect 478966 991448 478972 991460
rect 479024 991448 479030 991500
rect 512638 991448 512644 991500
rect 512696 991488 512702 991500
rect 543826 991488 543832 991500
rect 512696 991460 543832 991488
rect 512696 991448 512702 991460
rect 543826 991448 543832 991460
rect 543884 991448 543890 991500
rect 559558 991448 559564 991500
rect 559616 991488 559622 991500
rect 658918 991488 658924 991500
rect 559616 991460 658924 991488
rect 559616 991448 559622 991460
rect 658918 991448 658924 991460
rect 658976 991448 658982 991500
rect 164878 990836 164884 990888
rect 164936 990876 164942 990888
rect 170766 990876 170772 990888
rect 164936 990848 170772 990876
rect 164936 990836 164942 990848
rect 170766 990836 170772 990848
rect 170824 990836 170830 990888
rect 265618 990836 265624 990888
rect 265676 990876 265682 990888
rect 267642 990876 267648 990888
rect 265676 990848 267648 990876
rect 265676 990836 265682 990848
rect 267642 990836 267648 990848
rect 267700 990836 267706 990888
rect 73430 990224 73436 990276
rect 73488 990264 73494 990276
rect 112070 990264 112076 990276
rect 73488 990236 112076 990264
rect 73488 990224 73494 990236
rect 112070 990224 112076 990236
rect 112128 990224 112134 990276
rect 562318 990224 562324 990276
rect 562376 990264 562382 990276
rect 669958 990264 669964 990276
rect 562376 990236 669964 990264
rect 562376 990224 562382 990236
rect 669958 990224 669964 990236
rect 670016 990224 670022 990276
rect 44818 990088 44824 990140
rect 44876 990128 44882 990140
rect 109034 990128 109040 990140
rect 44876 990100 109040 990128
rect 44876 990088 44882 990100
rect 109034 990088 109040 990100
rect 109092 990088 109098 990140
rect 319438 990088 319444 990140
rect 319496 990128 319502 990140
rect 332962 990128 332968 990140
rect 319496 990100 332968 990128
rect 319496 990088 319502 990100
rect 332962 990088 332968 990100
rect 333020 990088 333026 990140
rect 369118 990088 369124 990140
rect 369176 990128 369182 990140
rect 414106 990128 414112 990140
rect 369176 990100 414112 990128
rect 369176 990088 369182 990100
rect 414106 990088 414112 990100
rect 414164 990088 414170 990140
rect 560938 990088 560944 990140
rect 560996 990128 561002 990140
rect 668578 990128 668584 990140
rect 560996 990100 668584 990128
rect 560996 990088 561002 990100
rect 668578 990088 668584 990100
rect 668636 990088 668642 990140
rect 53282 988728 53288 988780
rect 53340 988768 53346 988780
rect 95878 988768 95884 988780
rect 53340 988740 95884 988768
rect 53340 988728 53346 988740
rect 95878 988728 95884 988740
rect 95936 988728 95942 988780
rect 104894 986620 104900 986672
rect 104952 986660 104958 986672
rect 105814 986660 105820 986672
rect 104952 986632 105820 986660
rect 104952 986620 104958 986632
rect 105814 986620 105820 986632
rect 105872 986620 105878 986672
rect 217318 986620 217324 986672
rect 217376 986660 217382 986672
rect 219434 986660 219440 986672
rect 217376 986632 219440 986660
rect 217376 986620 217382 986632
rect 219434 986620 219440 986632
rect 219492 986620 219498 986672
rect 566458 986076 566464 986128
rect 566516 986116 566522 986128
rect 592494 986116 592500 986128
rect 566516 986088 592500 986116
rect 566516 986076 566522 986088
rect 592494 986076 592500 986088
rect 592552 986076 592558 986128
rect 89622 985940 89628 985992
rect 89680 985980 89686 985992
rect 106918 985980 106924 985992
rect 89680 985952 106924 985980
rect 89680 985940 89686 985952
rect 106918 985940 106924 985952
rect 106976 985940 106982 985992
rect 215938 985940 215944 985992
rect 215996 985980 216002 985992
rect 235626 985980 235632 985992
rect 215996 985952 235632 985980
rect 215996 985940 216002 985952
rect 235626 985940 235632 985952
rect 235684 985940 235690 985992
rect 268378 985940 268384 985992
rect 268436 985980 268442 985992
rect 300486 985980 300492 985992
rect 268436 985952 300492 985980
rect 268436 985940 268442 985952
rect 300486 985940 300492 985952
rect 300544 985940 300550 985992
rect 436738 985940 436744 985992
rect 436796 985980 436802 985992
rect 462774 985980 462780 985992
rect 436796 985952 462780 985980
rect 436796 985940 436802 985952
rect 462774 985940 462780 985952
rect 462832 985940 462838 985992
rect 514018 985940 514024 985992
rect 514076 985980 514082 985992
rect 560110 985980 560116 985992
rect 514076 985952 560116 985980
rect 514076 985940 514082 985952
rect 560110 985940 560116 985952
rect 560168 985940 560174 985992
rect 565078 985940 565084 985992
rect 565136 985980 565142 985992
rect 624970 985980 624976 985992
rect 565136 985952 624976 985980
rect 565136 985940 565142 985952
rect 624970 985940 624976 985952
rect 625028 985940 625034 985992
rect 154482 985668 154488 985720
rect 154540 985708 154546 985720
rect 160738 985708 160744 985720
rect 154540 985680 160744 985708
rect 154540 985668 154546 985680
rect 160738 985668 160744 985680
rect 160796 985668 160802 985720
rect 43438 975672 43444 975724
rect 43496 975712 43502 975724
rect 62114 975712 62120 975724
rect 43496 975684 62120 975712
rect 43496 975672 43502 975684
rect 62114 975672 62120 975684
rect 62172 975672 62178 975724
rect 651650 975672 651656 975724
rect 651708 975712 651714 975724
rect 672718 975712 672724 975724
rect 651708 975684 672724 975712
rect 651708 975672 651714 975684
rect 672718 975672 672724 975684
rect 672776 975672 672782 975724
rect 43438 961868 43444 961920
rect 43496 961908 43502 961920
rect 62114 961908 62120 961920
rect 43496 961880 62120 961908
rect 43496 961868 43502 961880
rect 62114 961868 62120 961880
rect 62172 961868 62178 961920
rect 651466 961868 651472 961920
rect 651524 961908 651530 961920
rect 665818 961908 665824 961920
rect 651524 961880 665824 961908
rect 651524 961868 651530 961880
rect 665818 961868 665824 961880
rect 665876 961868 665882 961920
rect 36538 952416 36544 952468
rect 36596 952456 36602 952468
rect 41690 952456 41696 952468
rect 36596 952428 41696 952456
rect 36596 952416 36602 952428
rect 41690 952416 41696 952428
rect 41748 952416 41754 952468
rect 37918 952212 37924 952264
rect 37976 952252 37982 952264
rect 41690 952252 41696 952264
rect 37976 952224 41696 952252
rect 37976 952212 37982 952224
rect 41690 952212 41696 952224
rect 41748 952212 41754 952264
rect 675846 949424 675852 949476
rect 675904 949464 675910 949476
rect 682378 949464 682384 949476
rect 675904 949436 682384 949464
rect 675904 949424 675910 949436
rect 682378 949424 682384 949436
rect 682436 949424 682442 949476
rect 652202 948064 652208 948116
rect 652260 948104 652266 948116
rect 660298 948104 660304 948116
rect 652260 948076 660304 948104
rect 652260 948064 652266 948076
rect 660298 948064 660304 948076
rect 660356 948064 660362 948116
rect 45554 945956 45560 946008
rect 45612 945996 45618 946008
rect 62114 945996 62120 946008
rect 45612 945968 62120 945996
rect 45612 945956 45618 945968
rect 62114 945956 62120 945968
rect 62172 945956 62178 946008
rect 41230 942556 41236 942608
rect 41288 942596 41294 942608
rect 41690 942596 41696 942608
rect 41288 942568 41696 942596
rect 41288 942556 41294 942568
rect 41690 942556 41696 942568
rect 41748 942556 41754 942608
rect 41230 941196 41236 941248
rect 41288 941236 41294 941248
rect 41690 941236 41696 941248
rect 41288 941208 41696 941236
rect 41288 941196 41294 941208
rect 41690 941196 41696 941208
rect 41748 941196 41754 941248
rect 40954 938612 40960 938664
rect 41012 938652 41018 938664
rect 41414 938652 41420 938664
rect 41012 938624 41420 938652
rect 41012 938612 41018 938624
rect 41414 938612 41420 938624
rect 41472 938612 41478 938664
rect 41138 938408 41144 938460
rect 41196 938448 41202 938460
rect 41506 938448 41512 938460
rect 41196 938420 41512 938448
rect 41196 938408 41202 938420
rect 41506 938408 41512 938420
rect 41564 938408 41570 938460
rect 651466 936980 651472 937032
rect 651524 937020 651530 937032
rect 661678 937020 661684 937032
rect 651524 936992 661684 937020
rect 651524 936980 651530 936992
rect 661678 936980 661684 936992
rect 661736 936980 661742 937032
rect 675846 928752 675852 928804
rect 675904 928792 675910 928804
rect 683114 928792 683120 928804
rect 675904 928764 683120 928792
rect 675904 928752 675910 928764
rect 683114 928752 683120 928764
rect 683172 928752 683178 928804
rect 53098 923244 53104 923296
rect 53156 923284 53162 923296
rect 62114 923284 62120 923296
rect 53156 923256 62120 923284
rect 53156 923244 53162 923256
rect 62114 923244 62120 923256
rect 62172 923244 62178 923296
rect 651466 921816 651472 921868
rect 651524 921856 651530 921868
rect 663058 921856 663064 921868
rect 651524 921828 663064 921856
rect 651524 921816 651530 921828
rect 663058 921816 663064 921828
rect 663116 921816 663122 921868
rect 50338 909440 50344 909492
rect 50396 909480 50402 909492
rect 62114 909480 62120 909492
rect 50396 909452 62120 909480
rect 50396 909440 50402 909452
rect 62114 909440 62120 909452
rect 62172 909440 62178 909492
rect 652386 909440 652392 909492
rect 652444 909480 652450 909492
rect 665818 909480 665824 909492
rect 652444 909452 665824 909480
rect 652444 909440 652450 909452
rect 665818 909440 665824 909452
rect 665876 909440 665882 909492
rect 47762 896996 47768 897048
rect 47820 897036 47826 897048
rect 62114 897036 62120 897048
rect 47820 897008 62120 897036
rect 47820 896996 47826 897008
rect 62114 896996 62120 897008
rect 62172 896996 62178 897048
rect 651466 895636 651472 895688
rect 651524 895676 651530 895688
rect 671338 895676 671344 895688
rect 651524 895648 671344 895676
rect 651524 895636 651530 895648
rect 671338 895636 671344 895648
rect 671396 895636 671402 895688
rect 44082 892752 44088 892764
rect 42858 892724 44088 892752
rect 42858 892466 42886 892724
rect 44082 892712 44088 892724
rect 44140 892712 44146 892764
rect 42938 892322 42990 892328
rect 42938 892264 42990 892270
rect 43076 891948 43128 891954
rect 43076 891890 43128 891896
rect 44082 891868 44088 891880
rect 43194 891840 44088 891868
rect 44082 891828 44088 891840
rect 44140 891828 44146 891880
rect 651650 881832 651656 881884
rect 651708 881872 651714 881884
rect 664438 881872 664444 881884
rect 651708 881844 664444 881872
rect 651708 881832 651714 881844
rect 664438 881832 664444 881844
rect 664496 881832 664502 881884
rect 46198 870816 46204 870868
rect 46256 870856 46262 870868
rect 62114 870856 62120 870868
rect 46256 870828 62120 870856
rect 46256 870816 46262 870828
rect 62114 870816 62120 870828
rect 62172 870816 62178 870868
rect 651466 869388 651472 869440
rect 651524 869428 651530 869440
rect 658918 869428 658924 869440
rect 651524 869400 658924 869428
rect 651524 869388 651530 869400
rect 658918 869388 658924 869400
rect 658976 869388 658982 869440
rect 51718 858372 51724 858424
rect 51776 858412 51782 858424
rect 62114 858412 62120 858424
rect 51776 858384 62120 858412
rect 51776 858372 51782 858384
rect 62114 858372 62120 858384
rect 62172 858372 62178 858424
rect 651466 852116 651472 852168
rect 651524 852156 651530 852168
rect 664438 852156 664444 852168
rect 651524 852128 664444 852156
rect 651524 852116 651530 852128
rect 664438 852116 664444 852128
rect 664496 852116 664502 852168
rect 54478 844568 54484 844620
rect 54536 844608 54542 844620
rect 62114 844608 62120 844620
rect 54536 844580 62120 844608
rect 54536 844568 54542 844580
rect 62114 844568 62120 844580
rect 62172 844568 62178 844620
rect 651834 841780 651840 841832
rect 651892 841820 651898 841832
rect 669958 841820 669964 841832
rect 651892 841792 669964 841820
rect 651892 841780 651898 841792
rect 669958 841780 669964 841792
rect 670016 841780 670022 841832
rect 651466 829404 651472 829456
rect 651524 829444 651530 829456
rect 660298 829444 660304 829456
rect 651524 829416 660304 829444
rect 651524 829404 651530 829416
rect 660298 829404 660304 829416
rect 660356 829404 660362 829456
rect 47578 818320 47584 818372
rect 47636 818360 47642 818372
rect 62114 818360 62120 818372
rect 47636 818332 62120 818360
rect 47636 818320 47642 818332
rect 62114 818320 62120 818332
rect 62172 818320 62178 818372
rect 41230 817028 41236 817080
rect 41288 817068 41294 817080
rect 41690 817068 41696 817080
rect 41288 817040 41696 817068
rect 41288 817028 41294 817040
rect 41690 817028 41696 817040
rect 41748 817028 41754 817080
rect 41230 815600 41236 815652
rect 41288 815640 41294 815652
rect 41598 815640 41604 815652
rect 41288 815612 41604 815640
rect 41288 815600 41294 815612
rect 41598 815600 41604 815612
rect 41656 815600 41662 815652
rect 651466 815600 651472 815652
rect 651524 815640 651530 815652
rect 661678 815640 661684 815652
rect 651524 815612 661684 815640
rect 651524 815600 651530 815612
rect 661678 815600 661684 815612
rect 661736 815600 661742 815652
rect 40770 810704 40776 810756
rect 40828 810744 40834 810756
rect 41690 810744 41696 810756
rect 40828 810716 41696 810744
rect 40828 810704 40834 810716
rect 41690 810704 41696 810716
rect 41748 810704 41754 810756
rect 41138 807372 41144 807424
rect 41196 807412 41202 807424
rect 41598 807412 41604 807424
rect 41196 807384 41604 807412
rect 41196 807372 41202 807384
rect 41598 807372 41604 807384
rect 41656 807372 41662 807424
rect 50338 805944 50344 805996
rect 50396 805984 50402 805996
rect 62114 805984 62120 805996
rect 50396 805956 62120 805984
rect 50396 805944 50402 805956
rect 62114 805944 62120 805956
rect 62172 805944 62178 805996
rect 651466 803224 651472 803276
rect 651524 803264 651530 803276
rect 651524 803236 654134 803264
rect 651524 803224 651530 803236
rect 654106 803196 654134 803236
rect 667198 803196 667204 803208
rect 654106 803168 667204 803196
rect 667198 803156 667204 803168
rect 667256 803156 667262 803208
rect 33042 802408 33048 802460
rect 33100 802448 33106 802460
rect 41690 802448 41696 802460
rect 33100 802420 41696 802448
rect 33100 802408 33106 802420
rect 41690 802408 41696 802420
rect 41748 802408 41754 802460
rect 39298 801728 39304 801780
rect 39356 801768 39362 801780
rect 39356 801740 41414 801768
rect 39356 801728 39362 801740
rect 41386 801700 41414 801740
rect 41598 801700 41604 801712
rect 41386 801672 41604 801700
rect 41598 801660 41604 801672
rect 41656 801660 41662 801712
rect 55858 793568 55864 793620
rect 55916 793608 55922 793620
rect 62114 793608 62120 793620
rect 55916 793580 62120 793608
rect 55916 793568 55922 793580
rect 62114 793568 62120 793580
rect 62172 793568 62178 793620
rect 651466 789352 651472 789404
rect 651524 789392 651530 789404
rect 668578 789392 668584 789404
rect 651524 789364 668584 789392
rect 651524 789352 651530 789364
rect 668578 789352 668584 789364
rect 668636 789352 668642 789404
rect 652386 775548 652392 775600
rect 652444 775588 652450 775600
rect 668762 775588 668768 775600
rect 652444 775560 668768 775588
rect 652444 775548 652450 775560
rect 668762 775548 668768 775560
rect 668820 775548 668826 775600
rect 35802 772828 35808 772880
rect 35860 772868 35866 772880
rect 41690 772868 41696 772880
rect 35860 772840 41696 772868
rect 35860 772828 35866 772840
rect 41690 772828 41696 772840
rect 41748 772828 41754 772880
rect 35802 768952 35808 769004
rect 35860 768992 35866 769004
rect 40034 768992 40040 769004
rect 35860 768964 40040 768992
rect 35860 768952 35866 768964
rect 40034 768952 40040 768964
rect 40092 768952 40098 769004
rect 35526 768816 35532 768868
rect 35584 768856 35590 768868
rect 39298 768856 39304 768868
rect 35584 768828 39304 768856
rect 35584 768816 35590 768828
rect 39298 768816 39304 768828
rect 39356 768816 39362 768868
rect 35342 768680 35348 768732
rect 35400 768720 35406 768732
rect 41690 768720 41696 768732
rect 35400 768692 41696 768720
rect 35400 768680 35406 768692
rect 41690 768680 41696 768692
rect 41748 768680 41754 768732
rect 35802 767456 35808 767508
rect 35860 767496 35866 767508
rect 36538 767496 36544 767508
rect 35860 767468 36544 767496
rect 35860 767456 35866 767468
rect 36538 767456 36544 767468
rect 36596 767456 36602 767508
rect 35618 767320 35624 767372
rect 35676 767360 35682 767372
rect 41322 767360 41328 767372
rect 35676 767332 41328 767360
rect 35676 767320 35682 767332
rect 41322 767320 41328 767332
rect 41380 767320 41386 767372
rect 48958 767320 48964 767372
rect 49016 767360 49022 767372
rect 62114 767360 62120 767372
rect 49016 767332 62120 767360
rect 49016 767320 49022 767332
rect 62114 767320 62120 767332
rect 62172 767320 62178 767372
rect 40034 764736 40040 764788
rect 40092 764776 40098 764788
rect 41690 764776 41696 764788
rect 40092 764748 41696 764776
rect 40092 764736 40098 764748
rect 41690 764736 41696 764748
rect 41748 764736 41754 764788
rect 35802 763240 35808 763292
rect 35860 763280 35866 763292
rect 37918 763280 37924 763292
rect 35860 763252 37924 763280
rect 35860 763240 35866 763252
rect 37918 763240 37924 763252
rect 37976 763240 37982 763292
rect 651466 763240 651472 763292
rect 651524 763280 651530 763292
rect 651524 763252 654134 763280
rect 651524 763240 651530 763252
rect 654106 763212 654134 763252
rect 660298 763212 660304 763224
rect 654106 763184 660304 763212
rect 660298 763172 660304 763184
rect 660356 763172 660362 763224
rect 31018 759636 31024 759688
rect 31076 759676 31082 759688
rect 41690 759676 41696 759688
rect 31076 759648 41696 759676
rect 31076 759636 31082 759648
rect 41690 759636 41696 759648
rect 41748 759636 41754 759688
rect 35158 758276 35164 758328
rect 35216 758316 35222 758328
rect 40310 758316 40316 758328
rect 35216 758288 40316 758316
rect 35216 758276 35222 758288
rect 40310 758276 40316 758288
rect 40368 758276 40374 758328
rect 37918 757732 37924 757784
rect 37976 757772 37982 757784
rect 40310 757772 40316 757784
rect 37976 757744 40316 757772
rect 37976 757732 37982 757744
rect 40310 757732 40316 757744
rect 40368 757732 40374 757784
rect 676030 757120 676036 757172
rect 676088 757160 676094 757172
rect 683390 757160 683396 757172
rect 676088 757132 683396 757160
rect 676088 757120 676094 757132
rect 683390 757120 683396 757132
rect 683448 757120 683454 757172
rect 51718 753516 51724 753568
rect 51776 753556 51782 753568
rect 62114 753556 62120 753568
rect 51776 753528 62120 753556
rect 51776 753516 51782 753528
rect 62114 753516 62120 753528
rect 62172 753516 62178 753568
rect 651466 749368 651472 749420
rect 651524 749408 651530 749420
rect 665818 749408 665824 749420
rect 651524 749380 665824 749408
rect 651524 749368 651530 749380
rect 665818 749368 665824 749380
rect 665876 749368 665882 749420
rect 668394 742704 668400 742756
rect 668452 742744 668458 742756
rect 668762 742744 668768 742756
rect 668452 742716 668768 742744
rect 668452 742704 668458 742716
rect 668762 742704 668768 742716
rect 668820 742704 668826 742756
rect 54478 741072 54484 741124
rect 54536 741112 54542 741124
rect 62114 741112 62120 741124
rect 54536 741084 62120 741112
rect 54536 741072 54542 741084
rect 62114 741072 62120 741084
rect 62172 741072 62178 741124
rect 651834 735564 651840 735616
rect 651892 735604 651898 735616
rect 661862 735604 661868 735616
rect 651892 735576 661868 735604
rect 651892 735564 651898 735576
rect 661862 735564 661868 735576
rect 661920 735564 661926 735616
rect 35802 730056 35808 730108
rect 35860 730096 35866 730108
rect 41690 730096 41696 730108
rect 35860 730068 41696 730096
rect 35860 730056 35866 730068
rect 41690 730056 41696 730068
rect 41748 730056 41754 730108
rect 674380 728612 674432 728618
rect 674380 728554 674432 728560
rect 672166 728424 672172 728476
rect 672224 728464 672230 728476
rect 672224 728436 674268 728464
rect 672224 728424 672230 728436
rect 672350 728288 672356 728340
rect 672408 728328 672414 728340
rect 672408 728300 674176 728328
rect 672408 728288 672414 728300
rect 673178 728084 673184 728136
rect 673236 728124 673242 728136
rect 673236 728096 674058 728124
rect 673236 728084 673242 728096
rect 41322 725908 41328 725960
rect 41380 725948 41386 725960
rect 41690 725948 41696 725960
rect 41380 725920 41696 725948
rect 41380 725908 41386 725920
rect 41690 725908 41696 725920
rect 41748 725908 41754 725960
rect 41322 724752 41328 724804
rect 41380 724792 41386 724804
rect 41690 724792 41696 724804
rect 41380 724764 41696 724792
rect 41380 724752 41386 724764
rect 41690 724752 41696 724764
rect 41748 724752 41754 724804
rect 677318 724208 677324 724260
rect 677376 724248 677382 724260
rect 683206 724248 683212 724260
rect 677376 724220 683212 724248
rect 677376 724208 677382 724220
rect 683206 724208 683212 724220
rect 683264 724208 683270 724260
rect 651466 723120 651472 723172
rect 651524 723160 651530 723172
rect 663058 723160 663064 723172
rect 651524 723132 663064 723160
rect 651524 723120 651530 723132
rect 663058 723120 663064 723132
rect 663116 723120 663122 723172
rect 34146 720264 34152 720316
rect 34204 720304 34210 720316
rect 38654 720304 38660 720316
rect 34204 720276 38660 720304
rect 34204 720264 34210 720276
rect 38654 720264 38660 720276
rect 38712 720264 38718 720316
rect 36538 717340 36544 717392
rect 36596 717380 36602 717392
rect 41690 717380 41696 717392
rect 36596 717352 41696 717380
rect 36596 717340 36602 717352
rect 41690 717340 41696 717352
rect 41748 717340 41754 717392
rect 39298 716184 39304 716236
rect 39356 716224 39362 716236
rect 41506 716224 41512 716236
rect 39356 716196 41512 716224
rect 39356 716184 39362 716196
rect 41506 716184 41512 716196
rect 41564 716184 41570 716236
rect 34514 715504 34520 715556
rect 34572 715544 34578 715556
rect 40310 715544 40316 715556
rect 34572 715516 40316 715544
rect 34572 715504 34578 715516
rect 40310 715504 40316 715516
rect 40368 715504 40374 715556
rect 50338 714824 50344 714876
rect 50396 714864 50402 714876
rect 62114 714864 62120 714876
rect 50396 714836 62120 714864
rect 50396 714824 50402 714836
rect 62114 714824 62120 714836
rect 62172 714824 62178 714876
rect 652570 709316 652576 709368
rect 652628 709356 652634 709368
rect 664438 709356 664444 709368
rect 652628 709328 664444 709356
rect 652628 709316 652634 709328
rect 664438 709316 664444 709328
rect 664496 709316 664502 709368
rect 55858 701020 55864 701072
rect 55916 701060 55922 701072
rect 62114 701060 62120 701072
rect 55916 701032 62120 701060
rect 55916 701020 55922 701032
rect 62114 701020 62120 701032
rect 62172 701020 62178 701072
rect 652386 696940 652392 696992
rect 652444 696980 652450 696992
rect 669958 696980 669964 696992
rect 652444 696952 669964 696980
rect 652444 696940 652450 696952
rect 669958 696940 669964 696952
rect 670016 696940 670022 696992
rect 53098 688644 53104 688696
rect 53156 688684 53162 688696
rect 62114 688684 62120 688696
rect 53156 688656 62120 688684
rect 53156 688644 53162 688656
rect 62114 688644 62120 688656
rect 62172 688644 62178 688696
rect 35802 687216 35808 687268
rect 35860 687256 35866 687268
rect 41414 687256 41420 687268
rect 35860 687228 41420 687256
rect 35860 687216 35866 687228
rect 41414 687216 41420 687228
rect 41472 687216 41478 687268
rect 35802 683136 35808 683188
rect 35860 683176 35866 683188
rect 41690 683176 41696 683188
rect 35860 683148 41696 683176
rect 35860 683136 35866 683148
rect 41690 683136 41696 683148
rect 41748 683136 41754 683188
rect 651834 683136 651840 683188
rect 651892 683176 651898 683188
rect 658918 683176 658924 683188
rect 651892 683148 658924 683176
rect 651892 683136 651898 683148
rect 658918 683136 658924 683148
rect 658976 683136 658982 683188
rect 35802 681980 35808 682032
rect 35860 682020 35866 682032
rect 36538 682020 36544 682032
rect 35860 681992 36544 682020
rect 35860 681980 35866 681992
rect 36538 681980 36544 681992
rect 36596 681980 36602 682032
rect 35618 681844 35624 681896
rect 35676 681884 35682 681896
rect 41690 681884 41696 681896
rect 35676 681856 41696 681884
rect 35676 681844 35682 681856
rect 41690 681844 41696 681856
rect 41748 681844 41754 681896
rect 35434 681708 35440 681760
rect 35492 681748 35498 681760
rect 35492 681720 38654 681748
rect 35492 681708 35498 681720
rect 38626 681680 38654 681720
rect 41598 681680 41604 681692
rect 38626 681652 41604 681680
rect 41598 681640 41604 681652
rect 41656 681640 41662 681692
rect 51718 674840 51724 674892
rect 51776 674880 51782 674892
rect 62114 674880 62120 674892
rect 51776 674852 62120 674880
rect 51776 674840 51782 674852
rect 62114 674840 62120 674852
rect 62172 674840 62178 674892
rect 32398 672732 32404 672784
rect 32456 672772 32462 672784
rect 41598 672772 41604 672784
rect 32456 672744 41604 672772
rect 32456 672732 32462 672744
rect 41598 672732 41604 672744
rect 41656 672732 41662 672784
rect 36538 671644 36544 671696
rect 36596 671684 36602 671696
rect 39666 671684 39672 671696
rect 36596 671656 39672 671684
rect 36596 671644 36602 671656
rect 39666 671644 39672 671656
rect 39724 671644 39730 671696
rect 35158 671304 35164 671356
rect 35216 671344 35222 671356
rect 41322 671344 41328 671356
rect 35216 671316 41328 671344
rect 35216 671304 35222 671316
rect 41322 671304 41328 671316
rect 41380 671304 41386 671356
rect 652386 669332 652392 669384
rect 652444 669372 652450 669384
rect 668394 669372 668400 669384
rect 652444 669344 668400 669372
rect 652444 669332 652450 669344
rect 668394 669332 668400 669344
rect 668452 669332 668458 669384
rect 671982 665660 671988 665712
rect 672040 665700 672046 665712
rect 672994 665700 673000 665712
rect 672040 665672 673000 665700
rect 672040 665660 672046 665672
rect 672994 665660 673000 665672
rect 673052 665660 673058 665712
rect 47578 662396 47584 662448
rect 47636 662436 47642 662448
rect 62114 662436 62120 662448
rect 47636 662408 62120 662436
rect 47636 662396 47642 662408
rect 62114 662396 62120 662408
rect 62172 662396 62178 662448
rect 651650 656888 651656 656940
rect 651708 656928 651714 656940
rect 663058 656928 663064 656940
rect 651708 656900 663064 656928
rect 651708 656888 651714 656900
rect 663058 656888 663064 656900
rect 663116 656888 663122 656940
rect 54478 647844 54484 647896
rect 54536 647884 54542 647896
rect 62114 647884 62120 647896
rect 54536 647856 62120 647884
rect 54536 647844 54542 647856
rect 62114 647844 62120 647856
rect 62172 647844 62178 647896
rect 651466 643084 651472 643136
rect 651524 643124 651530 643136
rect 668578 643124 668584 643136
rect 651524 643096 668584 643124
rect 651524 643084 651530 643096
rect 668578 643084 668584 643096
rect 668636 643084 668642 643136
rect 35802 639072 35808 639124
rect 35860 639112 35866 639124
rect 36538 639112 36544 639124
rect 35860 639084 36544 639112
rect 35860 639072 35866 639084
rect 36538 639072 36544 639084
rect 36596 639072 36602 639124
rect 35618 638936 35624 638988
rect 35676 638976 35682 638988
rect 41506 638976 41512 638988
rect 35676 638948 41512 638976
rect 35676 638936 35682 638948
rect 41506 638936 41512 638948
rect 41564 638936 41570 638988
rect 35802 636828 35808 636880
rect 35860 636868 35866 636880
rect 41690 636868 41696 636880
rect 35860 636840 41696 636868
rect 35860 636828 35866 636840
rect 41690 636828 41696 636840
rect 41748 636828 41754 636880
rect 51718 636216 51724 636268
rect 51776 636256 51782 636268
rect 62114 636256 62120 636268
rect 51776 636228 62120 636256
rect 51776 636216 51782 636228
rect 62114 636216 62120 636228
rect 62172 636216 62178 636268
rect 675846 634176 675852 634228
rect 675904 634216 675910 634228
rect 682378 634216 682384 634228
rect 675904 634188 682384 634216
rect 675904 634176 675910 634188
rect 682378 634176 682384 634188
rect 682436 634176 682442 634228
rect 32398 629892 32404 629944
rect 32456 629932 32462 629944
rect 41690 629932 41696 629944
rect 32456 629904 41696 629932
rect 32456 629892 32462 629904
rect 41690 629892 41696 629904
rect 41748 629892 41754 629944
rect 651558 628532 651564 628584
rect 651616 628572 651622 628584
rect 667198 628572 667204 628584
rect 651616 628544 667204 628572
rect 651616 628532 651622 628544
rect 667198 628532 667204 628544
rect 667256 628532 667262 628584
rect 48958 623772 48964 623824
rect 49016 623812 49022 623824
rect 62114 623812 62120 623824
rect 49016 623784 62120 623812
rect 49016 623772 49022 623784
rect 62114 623772 62120 623784
rect 62172 623772 62178 623824
rect 675846 622820 675852 622872
rect 675904 622860 675910 622872
rect 676674 622860 676680 622872
rect 675904 622832 676680 622860
rect 675904 622820 675910 622832
rect 676674 622820 676680 622832
rect 676732 622820 676738 622872
rect 651466 616836 651472 616888
rect 651524 616876 651530 616888
rect 660298 616876 660304 616888
rect 651524 616848 660304 616876
rect 651524 616836 651530 616848
rect 660298 616836 660304 616848
rect 660356 616836 660362 616888
rect 43260 612944 43312 612950
rect 43260 612886 43312 612892
rect 43383 612768 43760 612796
rect 43383 612714 43411 612768
rect 43732 612728 43760 612768
rect 46934 612728 46940 612740
rect 43732 612700 46940 612728
rect 46934 612688 46940 612700
rect 46992 612688 46998 612740
rect 43714 612524 43720 612536
rect 43516 612496 43720 612524
rect 43714 612484 43720 612496
rect 43772 612484 43778 612536
rect 43582 612332 43634 612338
rect 43582 612274 43634 612280
rect 43898 612116 43904 612128
rect 43746 612088 43904 612116
rect 43898 612076 43904 612088
rect 43956 612076 43962 612128
rect 45554 611912 45560 611924
rect 43838 611884 45560 611912
rect 45554 611872 45560 611884
rect 45612 611872 45618 611924
rect 43931 611720 43983 611726
rect 43931 611662 43983 611668
rect 44910 611504 44916 611516
rect 44068 611476 44916 611504
rect 44910 611464 44916 611476
rect 44968 611464 44974 611516
rect 44149 611328 44155 611380
rect 44207 611328 44213 611380
rect 44726 611096 44732 611108
rect 44298 611068 44732 611096
rect 44726 611056 44732 611068
rect 44784 611056 44790 611108
rect 45738 610892 45744 610904
rect 44405 610864 45744 610892
rect 45738 610852 45744 610864
rect 45796 610852 45802 610904
rect 44502 610768 44554 610774
rect 44502 610710 44554 610716
rect 56042 608608 56048 608660
rect 56100 608648 56106 608660
rect 62114 608648 62120 608660
rect 56100 608620 62120 608648
rect 56100 608608 56106 608620
rect 62114 608608 62120 608620
rect 62172 608608 62178 608660
rect 651466 603100 651472 603152
rect 651524 603140 651530 603152
rect 661678 603140 661684 603152
rect 651524 603112 661684 603140
rect 651524 603100 651530 603112
rect 661678 603100 661684 603112
rect 661736 603100 661742 603152
rect 673454 598612 673460 598664
rect 673512 598652 673518 598664
rect 673822 598652 673828 598664
rect 673512 598624 673828 598652
rect 673512 598612 673518 598624
rect 673822 598612 673828 598624
rect 673880 598612 673886 598664
rect 48958 597524 48964 597576
rect 49016 597564 49022 597576
rect 62114 597564 62120 597576
rect 49016 597536 62120 597564
rect 49016 597524 49022 597536
rect 62114 597524 62120 597536
rect 62172 597524 62178 597576
rect 40862 592832 40868 592884
rect 40920 592872 40926 592884
rect 41598 592872 41604 592884
rect 40920 592844 41604 592872
rect 40920 592832 40926 592844
rect 41598 592832 41604 592844
rect 41656 592832 41662 592884
rect 673822 592424 673828 592476
rect 673880 592424 673886 592476
rect 40310 592288 40316 592340
rect 40368 592328 40374 592340
rect 41414 592328 41420 592340
rect 40368 592300 41420 592328
rect 40368 592288 40374 592300
rect 41414 592288 41420 592300
rect 41472 592288 41478 592340
rect 673546 592152 673552 592204
rect 673604 592192 673610 592204
rect 673840 592192 673868 592424
rect 673604 592164 673868 592192
rect 673604 592152 673610 592164
rect 675846 591336 675852 591388
rect 675904 591376 675910 591388
rect 682378 591376 682384 591388
rect 675904 591348 682384 591376
rect 675904 591336 675910 591348
rect 682378 591336 682384 591348
rect 682436 591336 682442 591388
rect 652386 590656 652392 590708
rect 652444 590696 652450 590708
rect 665818 590696 665824 590708
rect 652444 590668 665824 590696
rect 652444 590656 652450 590668
rect 665818 590656 665824 590668
rect 665876 590656 665882 590708
rect 33042 587120 33048 587172
rect 33100 587160 33106 587172
rect 40402 587160 40408 587172
rect 33100 587132 40408 587160
rect 33100 587120 33106 587132
rect 40402 587120 40408 587132
rect 40460 587120 40466 587172
rect 39942 586100 39948 586152
rect 40000 586140 40006 586152
rect 41690 586140 41696 586152
rect 40000 586112 41696 586140
rect 40000 586100 40006 586112
rect 41690 586100 41696 586112
rect 41748 586100 41754 586152
rect 35158 585896 35164 585948
rect 35216 585936 35222 585948
rect 41690 585936 41696 585948
rect 35216 585908 41696 585936
rect 35216 585896 35222 585908
rect 41690 585896 41696 585908
rect 41748 585896 41754 585948
rect 31018 585760 31024 585812
rect 31076 585800 31082 585812
rect 31076 585772 41414 585800
rect 31076 585760 31082 585772
rect 41386 585732 41414 585772
rect 41690 585732 41696 585744
rect 41386 585704 41696 585732
rect 41690 585692 41696 585704
rect 41748 585692 41754 585744
rect 40862 584536 40868 584588
rect 40920 584576 40926 584588
rect 41598 584576 41604 584588
rect 40920 584548 41604 584576
rect 40920 584536 40926 584548
rect 41598 584536 41604 584548
rect 41656 584536 41662 584588
rect 50338 583720 50344 583772
rect 50396 583760 50402 583772
rect 62114 583760 62120 583772
rect 50396 583732 62120 583760
rect 50396 583720 50402 583732
rect 62114 583720 62120 583732
rect 62172 583720 62178 583772
rect 672166 579028 672172 579080
rect 672224 579068 672230 579080
rect 673178 579068 673184 579080
rect 672224 579040 673184 579068
rect 672224 579028 672230 579040
rect 673178 579028 673184 579040
rect 673236 579028 673242 579080
rect 651466 576852 651472 576904
rect 651524 576892 651530 576904
rect 664438 576892 664444 576904
rect 651524 576864 664444 576892
rect 651524 576852 651530 576864
rect 664438 576852 664444 576864
rect 664496 576852 664502 576904
rect 651650 563048 651656 563100
rect 651708 563088 651714 563100
rect 658918 563088 658924 563100
rect 651708 563060 658924 563088
rect 651708 563048 651714 563060
rect 658918 563048 658924 563060
rect 658976 563048 658982 563100
rect 673638 558328 673644 558340
rect 673472 558300 673644 558328
rect 55858 558084 55864 558136
rect 55916 558124 55922 558136
rect 62114 558124 62120 558136
rect 55916 558096 62120 558124
rect 55916 558084 55922 558096
rect 62114 558084 62120 558096
rect 62172 558084 62178 558136
rect 35802 557540 35808 557592
rect 35860 557580 35866 557592
rect 41506 557580 41512 557592
rect 35860 557552 41512 557580
rect 35860 557540 35866 557552
rect 41506 557540 41512 557552
rect 41564 557540 41570 557592
rect 673472 557580 673500 558300
rect 673638 558288 673644 558300
rect 673696 558288 673702 558340
rect 673638 557812 673644 557864
rect 673696 557812 673702 557864
rect 673656 557728 673684 557812
rect 673638 557676 673644 557728
rect 673696 557676 673702 557728
rect 673472 557552 673592 557580
rect 673564 557456 673592 557552
rect 673546 557404 673552 557456
rect 673604 557404 673610 557456
rect 35802 554752 35808 554804
rect 35860 554792 35866 554804
rect 41690 554792 41696 554804
rect 35860 554764 41696 554792
rect 35860 554752 35866 554764
rect 41690 554752 41696 554764
rect 41748 554752 41754 554804
rect 35802 553392 35808 553444
rect 35860 553432 35866 553444
rect 41322 553432 41328 553444
rect 35860 553404 41328 553432
rect 35860 553392 35866 553404
rect 41322 553392 41328 553404
rect 41380 553392 41386 553444
rect 41322 552032 41328 552084
rect 41380 552072 41386 552084
rect 41690 552072 41696 552084
rect 41380 552044 41696 552072
rect 41380 552032 41386 552044
rect 41690 552032 41696 552044
rect 41748 552032 41754 552084
rect 651466 550604 651472 550656
rect 651524 550644 651530 550656
rect 660298 550644 660304 550656
rect 651524 550616 660304 550644
rect 651524 550604 651530 550616
rect 660298 550604 660304 550616
rect 660356 550604 660362 550656
rect 41230 548088 41236 548140
rect 41288 548128 41294 548140
rect 41690 548128 41696 548140
rect 41288 548100 41696 548128
rect 41288 548088 41294 548100
rect 41690 548088 41696 548100
rect 41748 548088 41754 548140
rect 31754 547816 31760 547868
rect 31812 547856 31818 547868
rect 38470 547856 38476 547868
rect 31812 547828 38476 547856
rect 31812 547816 31818 547828
rect 38470 547816 38476 547828
rect 38528 547816 38534 547868
rect 675846 546456 675852 546508
rect 675904 546496 675910 546508
rect 680998 546496 681004 546508
rect 675904 546468 681004 546496
rect 675904 546456 675910 546468
rect 680998 546456 681004 546468
rect 681056 546456 681062 546508
rect 47578 545096 47584 545148
rect 47636 545136 47642 545148
rect 62114 545136 62120 545148
rect 47636 545108 62120 545136
rect 47636 545096 47642 545108
rect 62114 545096 62120 545108
rect 62172 545096 62178 545148
rect 33778 542988 33784 543040
rect 33836 543028 33842 543040
rect 41506 543028 41512 543040
rect 33836 543000 41512 543028
rect 33836 542988 33842 543000
rect 41506 542988 41512 543000
rect 41564 542988 41570 543040
rect 38470 542308 38476 542360
rect 38528 542348 38534 542360
rect 41690 542348 41696 542360
rect 38528 542320 41696 542348
rect 38528 542308 38534 542320
rect 41690 542308 41696 542320
rect 41748 542308 41754 542360
rect 651466 536800 651472 536852
rect 651524 536840 651530 536852
rect 669406 536840 669412 536852
rect 651524 536812 669412 536840
rect 651524 536800 651530 536812
rect 669406 536800 669412 536812
rect 669464 536800 669470 536852
rect 50338 532720 50344 532772
rect 50396 532760 50402 532772
rect 62114 532760 62120 532772
rect 50396 532732 62120 532760
rect 50396 532720 50402 532732
rect 62114 532720 62120 532732
rect 62172 532720 62178 532772
rect 651834 522996 651840 523048
rect 651892 523036 651898 523048
rect 661862 523036 661868 523048
rect 651892 523008 661868 523036
rect 651892 522996 651898 523008
rect 661862 522996 661868 523008
rect 661920 522996 661926 523048
rect 676858 520276 676864 520328
rect 676916 520316 676922 520328
rect 683114 520316 683120 520328
rect 676916 520288 683120 520316
rect 676916 520276 676922 520288
rect 683114 520276 683120 520288
rect 683172 520276 683178 520328
rect 54478 518916 54484 518968
rect 54536 518956 54542 518968
rect 62114 518956 62120 518968
rect 54536 518928 62120 518956
rect 54536 518916 54542 518928
rect 62114 518916 62120 518928
rect 62172 518916 62178 518968
rect 675846 518780 675852 518832
rect 675904 518820 675910 518832
rect 677870 518820 677876 518832
rect 675904 518792 677876 518820
rect 675904 518780 675910 518792
rect 677870 518780 677876 518792
rect 677928 518780 677934 518832
rect 651466 510620 651472 510672
rect 651524 510660 651530 510672
rect 659102 510660 659108 510672
rect 651524 510632 659108 510660
rect 651524 510620 651530 510632
rect 659102 510620 659108 510632
rect 659160 510620 659166 510672
rect 46198 506472 46204 506524
rect 46256 506512 46262 506524
rect 62114 506512 62120 506524
rect 46256 506484 62120 506512
rect 46256 506472 46262 506484
rect 62114 506472 62120 506484
rect 62172 506472 62178 506524
rect 676030 502324 676036 502376
rect 676088 502364 676094 502376
rect 678238 502364 678244 502376
rect 676088 502336 678244 502364
rect 676088 502324 676094 502336
rect 678238 502324 678244 502336
rect 678296 502324 678302 502376
rect 675846 500896 675852 500948
rect 675904 500936 675910 500948
rect 680998 500936 681004 500948
rect 675904 500908 681004 500936
rect 675904 500896 675910 500908
rect 680998 500896 681004 500908
rect 681056 500896 681062 500948
rect 652570 494708 652576 494760
rect 652628 494748 652634 494760
rect 663242 494748 663248 494760
rect 652628 494720 663248 494748
rect 652628 494708 652634 494720
rect 663242 494708 663248 494720
rect 663300 494708 663306 494760
rect 48958 491920 48964 491972
rect 49016 491960 49022 491972
rect 62114 491960 62120 491972
rect 49016 491932 62120 491960
rect 49016 491920 49022 491932
rect 62114 491920 62120 491932
rect 62172 491920 62178 491972
rect 677502 491104 677508 491156
rect 677560 491144 677566 491156
rect 683298 491144 683304 491156
rect 677560 491116 683304 491144
rect 677560 491104 677566 491116
rect 683298 491104 683304 491116
rect 683356 491104 683362 491156
rect 651466 484440 651472 484492
rect 651524 484480 651530 484492
rect 651524 484452 654134 484480
rect 651524 484440 651530 484452
rect 654106 484412 654134 484452
rect 667198 484412 667204 484424
rect 654106 484384 667204 484412
rect 667198 484372 667204 484384
rect 667256 484372 667262 484424
rect 680998 481516 681004 481568
rect 681056 481556 681062 481568
rect 683114 481556 683120 481568
rect 681056 481528 683120 481556
rect 681056 481516 681062 481528
rect 683114 481516 683120 481528
rect 683172 481516 683178 481568
rect 51718 480224 51724 480276
rect 51776 480264 51782 480276
rect 62114 480264 62120 480276
rect 51776 480236 62120 480264
rect 51776 480224 51782 480236
rect 62114 480224 62120 480236
rect 62172 480224 62178 480276
rect 651466 470568 651472 470620
rect 651524 470608 651530 470620
rect 665818 470608 665824 470620
rect 651524 470580 665824 470608
rect 651524 470568 651530 470580
rect 665818 470568 665824 470580
rect 665876 470568 665882 470620
rect 51902 466420 51908 466472
rect 51960 466460 51966 466472
rect 62114 466460 62120 466472
rect 51960 466432 62120 466460
rect 51960 466420 51966 466432
rect 62114 466420 62120 466432
rect 62172 466420 62178 466472
rect 652386 456764 652392 456816
rect 652444 456804 652450 456816
rect 661678 456804 661684 456816
rect 652444 456776 661684 456804
rect 652444 456764 652450 456776
rect 661678 456764 661684 456776
rect 661736 456764 661742 456816
rect 673948 456204 674000 456210
rect 673948 456146 674000 456152
rect 673828 456000 673880 456006
rect 673828 455942 673880 455948
rect 673454 455812 673460 455864
rect 673512 455852 673518 455864
rect 673512 455824 673762 455852
rect 673512 455812 673518 455824
rect 673598 455660 673650 455666
rect 673598 455602 673650 455608
rect 673270 455336 673276 455388
rect 673328 455376 673334 455388
rect 673328 455348 673532 455376
rect 673328 455336 673334 455348
rect 673388 455252 673440 455258
rect 673388 455194 673440 455200
rect 672074 455064 672080 455116
rect 672132 455104 672138 455116
rect 672132 455076 673316 455104
rect 672132 455064 672138 455076
rect 673288 455022 673316 455076
rect 673040 454792 673046 454844
rect 673098 454792 673104 454844
rect 672902 454656 672908 454708
rect 672960 454696 672966 454708
rect 672960 454656 672994 454696
rect 672966 454410 672994 454656
rect 673058 454614 673086 454792
rect 673164 454640 673216 454646
rect 673164 454582 673216 454588
rect 672816 454232 672868 454238
rect 672816 454174 672868 454180
rect 53098 454044 53104 454096
rect 53156 454084 53162 454096
rect 62114 454084 62120 454096
rect 53156 454056 62120 454084
rect 53156 454044 53162 454056
rect 62114 454044 62120 454056
rect 62172 454044 62178 454096
rect 672724 453960 672776 453966
rect 672724 453902 672776 453908
rect 651466 444456 651472 444508
rect 651524 444496 651530 444508
rect 651524 444468 654134 444496
rect 651524 444456 651530 444468
rect 654106 444428 654134 444468
rect 668578 444428 668584 444440
rect 654106 444400 668584 444428
rect 668578 444388 668584 444400
rect 668636 444388 668642 444440
rect 50522 440240 50528 440292
rect 50580 440280 50586 440292
rect 62114 440280 62120 440292
rect 50580 440252 62120 440280
rect 50580 440240 50586 440252
rect 62114 440240 62120 440252
rect 62172 440240 62178 440292
rect 651466 430584 651472 430636
rect 651524 430624 651530 430636
rect 669958 430624 669964 430636
rect 651524 430596 669964 430624
rect 651524 430584 651530 430596
rect 669958 430584 669964 430596
rect 670016 430584 670022 430636
rect 54478 427796 54484 427848
rect 54536 427836 54542 427848
rect 62114 427836 62120 427848
rect 54536 427808 62120 427836
rect 54536 427796 54542 427808
rect 62114 427796 62120 427808
rect 62172 427796 62178 427848
rect 651834 416780 651840 416832
rect 651892 416820 651898 416832
rect 663058 416820 663064 416832
rect 651892 416792 663064 416820
rect 651892 416780 651898 416792
rect 663058 416780 663064 416792
rect 663116 416780 663122 416832
rect 33778 416032 33784 416084
rect 33836 416072 33842 416084
rect 41690 416072 41696 416084
rect 33836 416044 41696 416072
rect 33836 416032 33842 416044
rect 41690 416032 41696 416044
rect 41748 416032 41754 416084
rect 651466 404336 651472 404388
rect 651524 404376 651530 404388
rect 664438 404376 664444 404388
rect 651524 404348 664444 404376
rect 651524 404336 651530 404348
rect 664438 404336 664444 404348
rect 664496 404336 664502 404388
rect 55858 401616 55864 401668
rect 55916 401656 55922 401668
rect 62114 401656 62120 401668
rect 55916 401628 62120 401656
rect 55916 401616 55922 401628
rect 62114 401616 62120 401628
rect 62172 401616 62178 401668
rect 675846 395700 675852 395752
rect 675904 395740 675910 395752
rect 676398 395740 676404 395752
rect 675904 395712 676404 395740
rect 675904 395700 675910 395712
rect 676398 395700 676404 395712
rect 676456 395700 676462 395752
rect 652570 390532 652576 390584
rect 652628 390572 652634 390584
rect 658918 390572 658924 390584
rect 652628 390544 658924 390572
rect 652628 390532 652634 390544
rect 658918 390532 658924 390544
rect 658976 390532 658982 390584
rect 47762 389240 47768 389292
rect 47820 389280 47826 389292
rect 62114 389280 62120 389292
rect 47820 389252 62120 389280
rect 47820 389240 47826 389252
rect 62114 389240 62120 389252
rect 62172 389240 62178 389292
rect 35802 382508 35808 382560
rect 35860 382548 35866 382560
rect 40034 382548 40040 382560
rect 35860 382520 40040 382548
rect 35860 382508 35866 382520
rect 40034 382508 40040 382520
rect 40092 382508 40098 382560
rect 35618 382372 35624 382424
rect 35676 382412 35682 382424
rect 41690 382412 41696 382424
rect 35676 382384 41696 382412
rect 35676 382372 35682 382384
rect 41690 382372 41696 382384
rect 41748 382372 41754 382424
rect 35434 382236 35440 382288
rect 35492 382276 35498 382288
rect 41506 382276 41512 382288
rect 35492 382248 41512 382276
rect 35492 382236 35498 382248
rect 41506 382236 41512 382248
rect 41564 382236 41570 382288
rect 35526 381012 35532 381064
rect 35584 381052 35590 381064
rect 37918 381052 37924 381064
rect 35584 381024 37924 381052
rect 35584 381012 35590 381024
rect 37918 381012 37924 381024
rect 37976 381012 37982 381064
rect 35802 380876 35808 380928
rect 35860 380916 35866 380928
rect 41322 380916 41328 380928
rect 35860 380888 41328 380916
rect 35860 380876 35866 380888
rect 41322 380876 41328 380888
rect 41380 380876 41386 380928
rect 652386 378156 652392 378208
rect 652444 378196 652450 378208
rect 660298 378196 660304 378208
rect 652444 378168 660304 378196
rect 652444 378156 652450 378168
rect 660298 378156 660304 378168
rect 660356 378156 660362 378208
rect 35802 375980 35808 376032
rect 35860 376020 35866 376032
rect 39574 376020 39580 376032
rect 35860 375992 39580 376020
rect 35860 375980 35866 375992
rect 39574 375980 39580 375992
rect 39632 375980 39638 376032
rect 51902 375368 51908 375420
rect 51960 375408 51966 375420
rect 62114 375408 62120 375420
rect 51960 375380 62120 375408
rect 51960 375368 51966 375380
rect 62114 375368 62120 375380
rect 62172 375368 62178 375420
rect 651834 364352 651840 364404
rect 651892 364392 651898 364404
rect 661862 364392 661868 364404
rect 651892 364364 661868 364392
rect 651892 364352 651898 364364
rect 661862 364352 661868 364364
rect 661920 364352 661926 364404
rect 50338 362924 50344 362976
rect 50396 362964 50402 362976
rect 62114 362964 62120 362976
rect 50396 362936 62120 362964
rect 50396 362924 50402 362936
rect 62114 362924 62120 362936
rect 62172 362924 62178 362976
rect 44634 354968 44640 355020
rect 44692 355008 44698 355020
rect 44692 354980 45399 355008
rect 44692 354968 44698 354980
rect 44818 354560 44824 354612
rect 44876 354600 44882 354612
rect 44876 354572 45048 354600
rect 44876 354560 44882 354572
rect 44575 354544 44627 354550
rect 44575 354486 44627 354492
rect 44793 354464 44799 354476
rect 44712 354436 44799 354464
rect 44793 354424 44799 354436
rect 44851 354424 44857 354476
rect 45020 354396 45048 354572
rect 44928 354368 45048 354396
rect 44799 354340 44851 354346
rect 44799 354282 44851 354288
rect 44928 354110 44956 354368
rect 45371 354192 45399 354980
rect 45035 354164 45399 354192
rect 45035 353906 45063 354164
rect 45186 353812 45192 353864
rect 45244 353852 45250 353864
rect 45244 353824 45399 353852
rect 45244 353812 45250 353824
rect 45146 353728 45198 353734
rect 45146 353670 45198 353676
rect 45371 353648 45399 353824
rect 45250 353620 45399 353648
rect 45250 353498 45278 353620
rect 45359 353320 45411 353326
rect 45359 353262 45411 353268
rect 652386 350548 652392 350600
rect 652444 350588 652450 350600
rect 667198 350588 667204 350600
rect 652444 350560 667204 350588
rect 652444 350548 652450 350560
rect 667198 350548 667204 350560
rect 667256 350548 667262 350600
rect 46198 347012 46204 347064
rect 46256 347052 46262 347064
rect 62114 347052 62120 347064
rect 46256 347024 62120 347052
rect 46256 347012 46262 347024
rect 62114 347012 62120 347024
rect 62172 347012 62178 347064
rect 35802 343612 35808 343664
rect 35860 343652 35866 343664
rect 40218 343652 40224 343664
rect 35860 343624 40224 343652
rect 35860 343612 35866 343624
rect 40218 343612 40224 343624
rect 40276 343612 40282 343664
rect 35802 339464 35808 339516
rect 35860 339504 35866 339516
rect 37550 339504 37556 339516
rect 35860 339476 37556 339504
rect 35860 339464 35866 339476
rect 37550 339464 37556 339476
rect 37608 339464 37614 339516
rect 54478 336744 54484 336796
rect 54536 336784 54542 336796
rect 62114 336784 62120 336796
rect 54536 336756 62120 336784
rect 54536 336744 54542 336756
rect 62114 336744 62120 336756
rect 62172 336744 62178 336796
rect 651466 324300 651472 324352
rect 651524 324340 651530 324352
rect 666646 324340 666652 324352
rect 651524 324312 666652 324340
rect 651524 324300 651530 324312
rect 666646 324300 666652 324312
rect 666704 324300 666710 324352
rect 51718 310496 51724 310548
rect 51776 310536 51782 310548
rect 62114 310536 62120 310548
rect 51776 310508 62120 310536
rect 51776 310496 51782 310508
rect 62114 310496 62120 310508
rect 62172 310496 62178 310548
rect 651466 310496 651472 310548
rect 651524 310536 651530 310548
rect 667382 310536 667388 310548
rect 651524 310508 667388 310536
rect 651524 310496 651530 310508
rect 667382 310496 667388 310508
rect 667440 310496 667446 310548
rect 45462 298120 45468 298172
rect 45520 298160 45526 298172
rect 62114 298160 62120 298172
rect 45520 298132 62120 298160
rect 45520 298120 45526 298132
rect 62114 298120 62120 298132
rect 62172 298120 62178 298172
rect 675938 298052 675944 298104
rect 675996 298092 676002 298104
rect 678974 298092 678980 298104
rect 675996 298064 678980 298092
rect 675996 298052 676002 298064
rect 678974 298052 678980 298064
rect 679032 298052 679038 298104
rect 676214 297032 676220 297084
rect 676272 297072 676278 297084
rect 680998 297072 681004 297084
rect 676272 297044 681004 297072
rect 676272 297032 676278 297044
rect 680998 297032 681004 297044
rect 681056 297032 681062 297084
rect 41322 284928 41328 284980
rect 41380 284968 41386 284980
rect 41690 284968 41696 284980
rect 41380 284940 41696 284968
rect 41380 284928 41386 284940
rect 41690 284928 41696 284940
rect 41748 284928 41754 284980
rect 39298 284724 39304 284776
rect 39356 284764 39362 284776
rect 41690 284764 41696 284776
rect 39356 284736 41696 284764
rect 39356 284724 39362 284736
rect 41690 284724 41696 284736
rect 41748 284724 41754 284776
rect 651466 284316 651472 284368
rect 651524 284356 651530 284368
rect 667566 284356 667572 284368
rect 651524 284328 667572 284356
rect 651524 284316 651530 284328
rect 667566 284316 667572 284328
rect 667624 284316 667630 284368
rect 482830 276632 482836 276684
rect 482888 276672 482894 276684
rect 558822 276672 558828 276684
rect 482888 276644 558828 276672
rect 482888 276632 482894 276644
rect 558822 276632 558828 276644
rect 558880 276632 558886 276684
rect 103698 275952 103704 276004
rect 103756 275992 103762 276004
rect 160738 275992 160744 276004
rect 103756 275964 160744 275992
rect 103756 275952 103762 275964
rect 160738 275952 160744 275964
rect 160796 275952 160802 276004
rect 166350 275952 166356 276004
rect 166408 275992 166414 276004
rect 182082 275992 182088 276004
rect 166408 275964 182088 275992
rect 166408 275952 166414 275964
rect 182082 275952 182088 275964
rect 182140 275952 182146 276004
rect 188798 275952 188804 276004
rect 188856 275992 188862 276004
rect 221458 275992 221464 276004
rect 188856 275964 221464 275992
rect 188856 275952 188862 275964
rect 221458 275952 221464 275964
rect 221516 275952 221522 276004
rect 410058 275952 410064 276004
rect 410116 275992 410122 276004
rect 410116 275964 412634 275992
rect 410116 275952 410122 275964
rect 88334 275816 88340 275868
rect 88392 275856 88398 275868
rect 146938 275856 146944 275868
rect 88392 275828 146944 275856
rect 88392 275816 88398 275828
rect 146938 275816 146944 275828
rect 146996 275816 147002 275868
rect 149790 275816 149796 275868
rect 149848 275856 149854 275868
rect 187878 275856 187884 275868
rect 149848 275828 187884 275856
rect 149848 275816 149854 275828
rect 187878 275816 187884 275828
rect 187936 275816 187942 275868
rect 368842 275816 368848 275868
rect 368900 275856 368906 275868
rect 373258 275856 373264 275868
rect 368900 275828 373264 275856
rect 368900 275816 368906 275828
rect 373258 275816 373264 275828
rect 373316 275816 373322 275868
rect 393774 275816 393780 275868
rect 393832 275856 393838 275868
rect 411070 275856 411076 275868
rect 393832 275828 411076 275856
rect 393832 275816 393838 275828
rect 411070 275816 411076 275828
rect 411128 275816 411134 275868
rect 412606 275856 412634 275964
rect 419534 275952 419540 276004
rect 419592 275992 419598 276004
rect 439406 275992 439412 276004
rect 419592 275964 439412 275992
rect 419592 275952 419598 275964
rect 439406 275952 439412 275964
rect 439464 275952 439470 276004
rect 456058 275952 456064 276004
rect 456116 275992 456122 276004
rect 466638 275992 466644 276004
rect 456116 275964 466644 275992
rect 456116 275952 456122 275964
rect 466638 275952 466644 275964
rect 466696 275952 466702 276004
rect 466822 275952 466828 276004
rect 466880 275992 466886 276004
rect 523402 275992 523408 276004
rect 466880 275964 523408 275992
rect 466880 275952 466886 275964
rect 523402 275952 523408 275964
rect 523460 275952 523466 276004
rect 525794 275952 525800 276004
rect 525852 275992 525858 276004
rect 607306 275992 607312 276004
rect 525852 275964 607312 275992
rect 525852 275952 525858 275964
rect 607306 275952 607312 275964
rect 607364 275952 607370 276004
rect 424042 275856 424048 275868
rect 412606 275828 424048 275856
rect 424042 275816 424048 275828
rect 424100 275816 424106 275868
rect 432782 275816 432788 275868
rect 432840 275856 432846 275868
rect 487890 275856 487896 275868
rect 432840 275828 487896 275856
rect 432840 275816 432846 275828
rect 487890 275816 487896 275828
rect 487948 275816 487954 275868
rect 504726 275816 504732 275868
rect 504784 275856 504790 275868
rect 590746 275856 590752 275868
rect 504784 275828 590752 275856
rect 504784 275816 504790 275828
rect 590746 275816 590752 275828
rect 590804 275816 590810 275868
rect 220722 275748 220728 275800
rect 220780 275788 220786 275800
rect 224954 275788 224960 275800
rect 220780 275760 224960 275788
rect 220780 275748 220786 275760
rect 224954 275748 224960 275760
rect 225012 275748 225018 275800
rect 249058 275748 249064 275800
rect 249116 275788 249122 275800
rect 253474 275788 253480 275800
rect 249116 275760 253480 275788
rect 249116 275748 249122 275760
rect 253474 275748 253480 275760
rect 253532 275748 253538 275800
rect 277486 275748 277492 275800
rect 277544 275788 277550 275800
rect 285122 275788 285128 275800
rect 277544 275760 285128 275788
rect 277544 275748 277550 275760
rect 285122 275748 285128 275760
rect 285180 275748 285186 275800
rect 96614 275680 96620 275732
rect 96672 275720 96678 275732
rect 156598 275720 156604 275732
rect 96672 275692 156604 275720
rect 96672 275680 96678 275692
rect 156598 275680 156604 275692
rect 156656 275680 156662 275732
rect 174630 275680 174636 275732
rect 174688 275720 174694 275732
rect 208394 275720 208400 275732
rect 174688 275692 208400 275720
rect 174688 275680 174694 275692
rect 208394 275680 208400 275692
rect 208452 275680 208458 275732
rect 212442 275680 212448 275732
rect 212500 275720 212506 275732
rect 219894 275720 219900 275732
rect 212500 275692 219900 275720
rect 212500 275680 212506 275692
rect 219894 275680 219900 275692
rect 219952 275680 219958 275732
rect 232498 275680 232504 275732
rect 232556 275720 232562 275732
rect 245654 275720 245660 275732
rect 232556 275692 245660 275720
rect 232556 275680 232562 275692
rect 245654 275680 245660 275692
rect 245712 275680 245718 275732
rect 373258 275680 373264 275732
rect 373316 275720 373322 275732
rect 385034 275720 385040 275732
rect 373316 275692 385040 275720
rect 373316 275680 373322 275692
rect 385034 275680 385040 275692
rect 385092 275680 385098 275732
rect 400214 275680 400220 275732
rect 400272 275720 400278 275732
rect 418154 275720 418160 275732
rect 400272 275692 418160 275720
rect 400272 275680 400278 275692
rect 418154 275680 418160 275692
rect 418212 275680 418218 275732
rect 418338 275680 418344 275732
rect 418396 275720 418402 275732
rect 435910 275720 435916 275732
rect 418396 275692 435916 275720
rect 418396 275680 418402 275692
rect 435910 275680 435916 275692
rect 435968 275680 435974 275732
rect 491478 275720 491484 275732
rect 436112 275692 491484 275720
rect 259730 275612 259736 275664
rect 259788 275652 259794 275664
rect 266998 275652 267004 275664
rect 259788 275624 267004 275652
rect 259788 275612 259794 275624
rect 266998 275612 267004 275624
rect 267056 275612 267062 275664
rect 85942 275544 85948 275596
rect 86000 275584 86006 275596
rect 150802 275584 150808 275596
rect 86000 275556 150808 275584
rect 86000 275544 86006 275556
rect 150802 275544 150808 275556
rect 150860 275544 150866 275596
rect 160462 275544 160468 275596
rect 160520 275584 160526 275596
rect 172422 275584 172428 275596
rect 160520 275556 172428 275584
rect 160520 275544 160526 275556
rect 172422 275544 172428 275556
rect 172480 275544 172486 275596
rect 181714 275544 181720 275596
rect 181772 275584 181778 275596
rect 218606 275584 218612 275596
rect 181772 275556 218612 275584
rect 181772 275544 181778 275556
rect 218606 275544 218612 275556
rect 218664 275544 218670 275596
rect 225414 275544 225420 275596
rect 225472 275584 225478 275596
rect 243538 275584 243544 275596
rect 225472 275556 243544 275584
rect 225472 275544 225478 275556
rect 243538 275544 243544 275556
rect 243596 275544 243602 275596
rect 244366 275544 244372 275596
rect 244424 275584 244430 275596
rect 247034 275584 247040 275596
rect 244424 275556 247040 275584
rect 244424 275544 244430 275556
rect 247034 275544 247040 275556
rect 247092 275544 247098 275596
rect 283374 275544 283380 275596
rect 283432 275584 283438 275596
rect 289078 275584 289084 275596
rect 283432 275556 289084 275584
rect 283432 275544 283438 275556
rect 289078 275544 289084 275556
rect 289136 275544 289142 275596
rect 367830 275544 367836 275596
rect 367888 275584 367894 275596
rect 377950 275584 377956 275596
rect 367888 275556 377956 275584
rect 367888 275544 367894 275556
rect 377950 275544 377956 275556
rect 378008 275544 378014 275596
rect 382458 275544 382464 275596
rect 382516 275584 382522 275596
rect 400398 275584 400404 275596
rect 382516 275556 400404 275584
rect 382516 275544 382522 275556
rect 400398 275544 400404 275556
rect 400456 275544 400462 275596
rect 403434 275544 403440 275596
rect 403492 275584 403498 275596
rect 428826 275584 428832 275596
rect 403492 275556 428832 275584
rect 403492 275544 403498 275556
rect 428826 275544 428832 275556
rect 428884 275544 428890 275596
rect 435726 275544 435732 275596
rect 435784 275584 435790 275596
rect 436112 275584 436140 275692
rect 491478 275680 491484 275692
rect 491536 275680 491542 275732
rect 493870 275680 493876 275732
rect 493928 275720 493934 275732
rect 502058 275720 502064 275732
rect 493928 275692 502064 275720
rect 493928 275680 493934 275692
rect 502058 275680 502064 275692
rect 502116 275680 502122 275732
rect 505830 275680 505836 275732
rect 505888 275720 505894 275732
rect 512730 275720 512736 275732
rect 505888 275692 512736 275720
rect 505888 275680 505894 275692
rect 512730 275680 512736 275692
rect 512788 275680 512794 275732
rect 516410 275680 516416 275732
rect 516468 275720 516474 275732
rect 604914 275720 604920 275732
rect 516468 275692 604920 275720
rect 516468 275680 516474 275692
rect 604914 275680 604920 275692
rect 604972 275680 604978 275732
rect 605098 275680 605104 275732
rect 605156 275720 605162 275732
rect 616782 275720 616788 275732
rect 605156 275692 616788 275720
rect 605156 275680 605162 275692
rect 616782 275680 616788 275692
rect 616840 275680 616846 275732
rect 435784 275556 436140 275584
rect 435784 275544 435790 275556
rect 441338 275544 441344 275596
rect 441396 275584 441402 275596
rect 498562 275584 498568 275596
rect 441396 275556 498568 275584
rect 441396 275544 441402 275556
rect 498562 275544 498568 275556
rect 498620 275544 498626 275596
rect 510062 275544 510068 275596
rect 510120 275584 510126 275596
rect 519814 275584 519820 275596
rect 510120 275556 519820 275584
rect 510120 275544 510126 275556
rect 519814 275544 519820 275556
rect 519872 275544 519878 275596
rect 523034 275544 523040 275596
rect 523092 275584 523098 275596
rect 525610 275584 525616 275596
rect 523092 275556 525616 275584
rect 523092 275544 523098 275556
rect 525610 275544 525616 275556
rect 525668 275544 525674 275596
rect 525978 275544 525984 275596
rect 526036 275584 526042 275596
rect 619082 275584 619088 275596
rect 526036 275556 619088 275584
rect 526036 275544 526042 275556
rect 619082 275544 619088 275556
rect 619140 275544 619146 275596
rect 625798 275544 625804 275596
rect 625856 275584 625862 275596
rect 640426 275584 640432 275596
rect 625856 275556 640432 275584
rect 625856 275544 625862 275556
rect 640426 275544 640432 275556
rect 640484 275544 640490 275596
rect 76466 275408 76472 275460
rect 76524 275448 76530 275460
rect 143258 275448 143264 275460
rect 76524 275420 143264 275448
rect 76524 275408 76530 275420
rect 143258 275408 143264 275420
rect 143316 275408 143322 275460
rect 148594 275408 148600 275460
rect 148652 275448 148658 275460
rect 164142 275448 164148 275460
rect 148652 275420 164148 275448
rect 148652 275408 148658 275420
rect 164142 275408 164148 275420
rect 164200 275408 164206 275460
rect 167546 275408 167552 275460
rect 167604 275448 167610 275460
rect 209038 275448 209044 275460
rect 167604 275420 209044 275448
rect 167604 275408 167610 275420
rect 209038 275408 209044 275420
rect 209096 275408 209102 275460
rect 218330 275408 218336 275460
rect 218388 275448 218394 275460
rect 239398 275448 239404 275460
rect 218388 275420 239404 275448
rect 218388 275408 218394 275420
rect 239398 275408 239404 275420
rect 239456 275408 239462 275460
rect 253658 275408 253664 275460
rect 253716 275448 253722 275460
rect 261478 275448 261484 275460
rect 253716 275420 261484 275448
rect 253716 275408 253722 275420
rect 261478 275408 261484 275420
rect 261536 275408 261542 275460
rect 284570 275408 284576 275460
rect 284628 275448 284634 275460
rect 290090 275448 290096 275460
rect 284628 275420 290096 275448
rect 284628 275408 284634 275420
rect 290090 275408 290096 275420
rect 290148 275408 290154 275460
rect 349798 275408 349804 275460
rect 349856 275448 349862 275460
rect 361390 275448 361396 275460
rect 349856 275420 361396 275448
rect 349856 275408 349862 275420
rect 361390 275408 361396 275420
rect 361448 275408 361454 275460
rect 362954 275408 362960 275460
rect 363012 275448 363018 275460
rect 367278 275448 367284 275460
rect 363012 275420 367284 275448
rect 363012 275408 363018 275420
rect 367278 275408 367284 275420
rect 367336 275408 367342 275460
rect 376662 275408 376668 275460
rect 376720 275448 376726 275460
rect 393314 275448 393320 275460
rect 376720 275420 393320 275448
rect 376720 275408 376726 275420
rect 393314 275408 393320 275420
rect 393372 275408 393378 275460
rect 395430 275408 395436 275460
rect 395488 275448 395494 275460
rect 403986 275448 403992 275460
rect 395488 275420 403992 275448
rect 395488 275408 395494 275420
rect 403986 275408 403992 275420
rect 404044 275408 404050 275460
rect 407758 275408 407764 275460
rect 407816 275448 407822 275460
rect 432322 275448 432328 275460
rect 407816 275420 432328 275448
rect 407816 275408 407822 275420
rect 432322 275408 432328 275420
rect 432380 275408 432386 275460
rect 438854 275408 438860 275460
rect 438912 275448 438918 275460
rect 446490 275448 446496 275460
rect 438912 275420 446496 275448
rect 438912 275408 438918 275420
rect 446490 275408 446496 275420
rect 446548 275408 446554 275460
rect 450538 275408 450544 275460
rect 450596 275448 450602 275460
rect 509142 275448 509148 275460
rect 450596 275420 509148 275448
rect 450596 275408 450602 275420
rect 509142 275408 509148 275420
rect 509200 275408 509206 275460
rect 512178 275408 512184 275460
rect 512236 275448 512242 275460
rect 533982 275448 533988 275460
rect 512236 275420 533988 275448
rect 512236 275408 512242 275420
rect 533982 275408 533988 275420
rect 534040 275408 534046 275460
rect 535730 275408 535736 275460
rect 535788 275448 535794 275460
rect 633342 275448 633348 275460
rect 535788 275420 633348 275448
rect 535788 275408 535794 275420
rect 633342 275408 633348 275420
rect 633400 275408 633406 275460
rect 70578 275272 70584 275324
rect 70636 275312 70642 275324
rect 140130 275312 140136 275324
rect 70636 275284 140136 275312
rect 70636 275272 70642 275284
rect 140130 275272 140136 275284
rect 140188 275272 140194 275324
rect 156874 275272 156880 275324
rect 156932 275312 156938 275324
rect 199286 275312 199292 275324
rect 156932 275284 199292 275312
rect 156932 275272 156938 275284
rect 199286 275272 199292 275284
rect 199344 275272 199350 275324
rect 211246 275272 211252 275324
rect 211304 275312 211310 275324
rect 232682 275312 232688 275324
rect 211304 275284 232688 275312
rect 211304 275272 211310 275284
rect 232682 275272 232688 275284
rect 232740 275272 232746 275324
rect 246758 275272 246764 275324
rect 246816 275312 246822 275324
rect 256694 275312 256700 275324
rect 246816 275284 256700 275312
rect 246816 275272 246822 275284
rect 256694 275272 256700 275284
rect 256752 275272 256758 275324
rect 260926 275272 260932 275324
rect 260984 275312 260990 275324
rect 273530 275312 273536 275324
rect 260984 275284 273536 275312
rect 260984 275272 260990 275284
rect 273530 275272 273536 275284
rect 273588 275272 273594 275324
rect 273898 275272 273904 275324
rect 273956 275312 273962 275324
rect 283282 275312 283288 275324
rect 273956 275284 283288 275312
rect 273956 275272 273962 275284
rect 283282 275272 283288 275284
rect 283340 275272 283346 275324
rect 328270 275272 328276 275324
rect 328328 275312 328334 275324
rect 335354 275312 335360 275324
rect 328328 275284 335360 275312
rect 328328 275272 328334 275284
rect 335354 275272 335360 275284
rect 335412 275272 335418 275324
rect 347038 275272 347044 275324
rect 347096 275312 347102 275324
rect 356698 275312 356704 275324
rect 347096 275284 356704 275312
rect 347096 275272 347102 275284
rect 356698 275272 356704 275284
rect 356756 275272 356762 275324
rect 359458 275272 359464 275324
rect 359516 275312 359522 275324
rect 370866 275312 370872 275324
rect 359516 275284 370872 275312
rect 359516 275272 359522 275284
rect 370866 275272 370872 275284
rect 370924 275272 370930 275324
rect 377398 275272 377404 275324
rect 377456 275312 377462 275324
rect 396902 275312 396908 275324
rect 377456 275284 396908 275312
rect 377456 275272 377462 275284
rect 396902 275272 396908 275284
rect 396960 275272 396966 275324
rect 400398 275272 400404 275324
rect 400456 275312 400462 275324
rect 425238 275312 425244 275324
rect 400456 275284 425244 275312
rect 400456 275272 400462 275284
rect 425238 275272 425244 275284
rect 425296 275272 425302 275324
rect 427814 275272 427820 275324
rect 427872 275312 427878 275324
rect 442994 275312 443000 275324
rect 427872 275284 443000 275312
rect 427872 275272 427878 275284
rect 442994 275272 443000 275284
rect 443052 275272 443058 275324
rect 453758 275272 453764 275324
rect 453816 275312 453822 275324
rect 516226 275312 516232 275324
rect 453816 275284 516232 275312
rect 453816 275272 453822 275284
rect 516226 275272 516232 275284
rect 516284 275272 516290 275324
rect 523678 275272 523684 275324
rect 523736 275312 523742 275324
rect 545850 275312 545856 275324
rect 523736 275284 545856 275312
rect 523736 275272 523742 275284
rect 545850 275272 545856 275284
rect 545908 275272 545914 275324
rect 546034 275272 546040 275324
rect 546092 275312 546098 275324
rect 552934 275312 552940 275324
rect 546092 275284 552940 275312
rect 546092 275272 546098 275284
rect 552934 275272 552940 275284
rect 552992 275272 552998 275324
rect 553118 275272 553124 275324
rect 553176 275312 553182 275324
rect 574186 275312 574192 275324
rect 553176 275284 574192 275312
rect 553176 275272 553182 275284
rect 574186 275272 574192 275284
rect 574244 275272 574250 275324
rect 110782 275136 110788 275188
rect 110840 275176 110846 275188
rect 164970 275176 164976 275188
rect 110840 275148 164976 275176
rect 110840 275136 110846 275148
rect 164970 275136 164976 275148
rect 165028 275136 165034 275188
rect 171042 275136 171048 275188
rect 171100 275176 171106 275188
rect 191006 275176 191012 275188
rect 171100 275148 191012 275176
rect 171100 275136 171106 275148
rect 191006 275136 191012 275148
rect 191064 275136 191070 275188
rect 428918 275136 428924 275188
rect 428976 275176 428982 275188
rect 428976 275148 480254 275176
rect 428976 275136 428982 275148
rect 135622 275000 135628 275052
rect 135680 275040 135686 275052
rect 167638 275040 167644 275052
rect 135680 275012 167644 275040
rect 135680 275000 135686 275012
rect 167638 275000 167644 275012
rect 167696 275000 167702 275052
rect 290458 275000 290464 275052
rect 290516 275040 290522 275052
rect 294322 275040 294328 275052
rect 290516 275012 294328 275040
rect 290516 275000 290522 275012
rect 294322 275000 294328 275012
rect 294380 275000 294386 275052
rect 366358 275000 366364 275052
rect 366416 275040 366422 275052
rect 369670 275040 369676 275052
rect 366416 275012 369676 275040
rect 366416 275000 366422 275012
rect 369670 275000 369676 275012
rect 369728 275000 369734 275052
rect 426250 275000 426256 275052
rect 426308 275040 426314 275052
rect 477218 275040 477224 275052
rect 426308 275012 477224 275040
rect 426308 275000 426314 275012
rect 477218 275000 477224 275012
rect 477276 275000 477282 275052
rect 480226 275040 480254 275148
rect 481542 275136 481548 275188
rect 481600 275176 481606 275188
rect 544654 275176 544660 275188
rect 481600 275148 544660 275176
rect 481600 275136 481606 275148
rect 544654 275136 544660 275148
rect 544712 275136 544718 275188
rect 552658 275136 552664 275188
rect 552716 275176 552722 275188
rect 560018 275176 560024 275188
rect 552716 275148 560024 275176
rect 552716 275136 552722 275148
rect 560018 275136 560024 275148
rect 560076 275136 560082 275188
rect 480806 275040 480812 275052
rect 480226 275012 480812 275040
rect 480806 275000 480812 275012
rect 480864 275000 480870 275052
rect 487798 275000 487804 275052
rect 487856 275040 487862 275052
rect 530486 275040 530492 275052
rect 487856 275012 530492 275040
rect 487856 275000 487862 275012
rect 530486 275000 530492 275012
rect 530544 275000 530550 275052
rect 530670 275000 530676 275052
rect 530728 275040 530734 275052
rect 541066 275040 541072 275052
rect 530728 275012 541072 275040
rect 530728 275000 530734 275012
rect 541066 275000 541072 275012
rect 541124 275000 541130 275052
rect 542262 275000 542268 275052
rect 542320 275040 542326 275052
rect 549346 275040 549352 275052
rect 542320 275012 549352 275040
rect 542320 275000 542326 275012
rect 549346 275000 549352 275012
rect 549404 275000 549410 275052
rect 551554 275000 551560 275052
rect 551612 275040 551618 275052
rect 553118 275040 553124 275052
rect 551612 275012 553124 275040
rect 551612 275000 551618 275012
rect 553118 275000 553124 275012
rect 553176 275000 553182 275052
rect 559558 275000 559564 275052
rect 559616 275040 559622 275052
rect 567102 275040 567108 275052
rect 559616 275012 567108 275040
rect 559616 275000 559622 275012
rect 567102 275000 567108 275012
rect 567160 275000 567166 275052
rect 81250 274932 81256 274984
rect 81308 274972 81314 274984
rect 86218 274972 86224 274984
rect 81308 274944 86224 274972
rect 81308 274932 81314 274944
rect 86218 274932 86224 274944
rect 86276 274932 86282 274984
rect 129642 274864 129648 274916
rect 129700 274904 129706 274916
rect 136082 274904 136088 274916
rect 129700 274876 136088 274904
rect 129700 274864 129706 274876
rect 136082 274864 136088 274876
rect 136140 274864 136146 274916
rect 142706 274864 142712 274916
rect 142764 274904 142770 274916
rect 166258 274904 166264 274916
rect 142764 274876 166264 274904
rect 142764 274864 142770 274876
rect 166258 274864 166264 274876
rect 166316 274864 166322 274916
rect 469398 274864 469404 274916
rect 469456 274904 469462 274916
rect 483198 274904 483204 274916
rect 469456 274876 483204 274904
rect 469456 274864 469462 274876
rect 483198 274864 483204 274876
rect 483256 274864 483262 274916
rect 490558 274864 490564 274916
rect 490616 274904 490622 274916
rect 526898 274904 526904 274916
rect 490616 274876 526904 274904
rect 490616 274864 490622 274876
rect 526898 274864 526904 274876
rect 526956 274864 526962 274916
rect 543274 274864 543280 274916
rect 543332 274904 543338 274916
rect 645118 274904 645124 274916
rect 543332 274876 645124 274904
rect 543332 274864 543338 274876
rect 645118 274864 645124 274876
rect 645176 274864 645182 274916
rect 199470 274796 199476 274848
rect 199528 274836 199534 274848
rect 202230 274836 202236 274848
rect 199528 274808 202236 274836
rect 199528 274796 199534 274808
rect 202230 274796 202236 274808
rect 202288 274796 202294 274848
rect 208854 274796 208860 274848
rect 208912 274836 208918 274848
rect 211062 274836 211068 274848
rect 208912 274808 211068 274836
rect 208912 274796 208918 274808
rect 211062 274796 211068 274808
rect 211120 274796 211126 274848
rect 257338 274796 257344 274848
rect 257396 274836 257402 274848
rect 259914 274836 259920 274848
rect 257396 274808 259920 274836
rect 257396 274796 257402 274808
rect 259914 274796 259920 274808
rect 259972 274796 259978 274848
rect 357250 274796 357256 274848
rect 357308 274836 357314 274848
rect 360194 274836 360200 274848
rect 357308 274808 360200 274836
rect 357308 274796 357314 274808
rect 360194 274796 360200 274808
rect 360252 274796 360258 274848
rect 369854 274796 369860 274848
rect 369912 274836 369918 274848
rect 375558 274836 375564 274848
rect 369912 274808 375564 274836
rect 369912 274796 369918 274808
rect 375558 274796 375564 274808
rect 375616 274796 375622 274848
rect 146202 274728 146208 274780
rect 146260 274768 146266 274780
rect 149698 274768 149704 274780
rect 146260 274740 149704 274768
rect 146260 274728 146266 274740
rect 149698 274728 149704 274740
rect 149756 274728 149762 274780
rect 150986 274728 150992 274780
rect 151044 274768 151050 274780
rect 152734 274768 152740 274780
rect 151044 274740 152740 274768
rect 151044 274728 151050 274740
rect 152734 274728 152740 274740
rect 152792 274728 152798 274780
rect 163958 274728 163964 274780
rect 164016 274768 164022 274780
rect 170398 274768 170404 274780
rect 164016 274740 170404 274768
rect 164016 274728 164022 274740
rect 170398 274728 170404 274740
rect 170456 274728 170462 274780
rect 172238 274728 172244 274780
rect 172296 274768 172302 274780
rect 174354 274768 174360 274780
rect 172296 274740 174360 274768
rect 172296 274728 172302 274740
rect 174354 274728 174360 274740
rect 174412 274728 174418 274780
rect 387702 274728 387708 274780
rect 387760 274768 387766 274780
rect 394510 274768 394516 274780
rect 387760 274740 394516 274768
rect 387760 274728 387766 274740
rect 394510 274728 394516 274740
rect 394568 274728 394574 274780
rect 397086 274728 397092 274780
rect 397144 274768 397150 274780
rect 401502 274768 401508 274780
rect 397144 274740 401508 274768
rect 397144 274728 397150 274740
rect 401502 274728 401508 274740
rect 401560 274728 401566 274780
rect 415210 274728 415216 274780
rect 415268 274768 415274 274780
rect 419350 274768 419356 274780
rect 415268 274740 419356 274768
rect 415268 274728 415274 274740
rect 419350 274728 419356 274740
rect 419408 274728 419414 274780
rect 446398 274728 446404 274780
rect 446456 274768 446462 274780
rect 453574 274768 453580 274780
rect 446456 274740 453580 274768
rect 446456 274728 446462 274740
rect 453574 274728 453580 274740
rect 453632 274728 453638 274780
rect 483658 274728 483664 274780
rect 483716 274768 483722 274780
rect 493870 274768 493876 274780
rect 483716 274740 493876 274768
rect 483716 274728 483722 274740
rect 493870 274728 493876 274740
rect 493928 274728 493934 274780
rect 498470 274728 498476 274780
rect 498528 274768 498534 274780
rect 499758 274768 499764 274780
rect 498528 274740 499764 274768
rect 498528 274728 498534 274740
rect 499758 274728 499764 274740
rect 499816 274728 499822 274780
rect 501598 274728 501604 274780
rect 501656 274768 501662 274780
rect 505646 274768 505652 274780
rect 501656 274740 505652 274768
rect 501656 274728 501662 274740
rect 505646 274728 505652 274740
rect 505704 274728 505710 274780
rect 506474 274728 506480 274780
rect 506532 274768 506538 274780
rect 510338 274768 510344 274780
rect 506532 274740 510344 274768
rect 506532 274728 506538 274740
rect 510338 274728 510344 274740
rect 510396 274728 510402 274780
rect 510522 274728 510528 274780
rect 510580 274768 510586 274780
rect 537294 274768 537300 274780
rect 510580 274740 537300 274768
rect 510580 274728 510586 274740
rect 537294 274728 537300 274740
rect 537352 274728 537358 274780
rect 537662 274728 537668 274780
rect 537720 274768 537726 274780
rect 538766 274768 538772 274780
rect 537720 274740 538772 274768
rect 537720 274728 537726 274740
rect 538766 274728 538772 274740
rect 538824 274728 538830 274780
rect 539502 274728 539508 274780
rect 539560 274768 539566 274780
rect 542078 274768 542084 274780
rect 539560 274740 542084 274768
rect 539560 274728 539566 274740
rect 542078 274728 542084 274740
rect 542136 274728 542142 274780
rect 71774 274660 71780 274712
rect 71832 274700 71838 274712
rect 73798 274700 73804 274712
rect 71832 274672 73804 274700
rect 71832 274660 71838 274672
rect 73798 274660 73804 274672
rect 73856 274660 73862 274712
rect 74074 274660 74080 274712
rect 74132 274700 74138 274712
rect 77202 274700 77208 274712
rect 74132 274672 77208 274700
rect 74132 274660 74138 274672
rect 77202 274660 77208 274672
rect 77260 274660 77266 274712
rect 210050 274660 210056 274712
rect 210108 274700 210114 274712
rect 212258 274700 212264 274712
rect 210108 274672 212264 274700
rect 210108 274660 210114 274672
rect 212258 274660 212264 274672
rect 212316 274660 212322 274712
rect 243170 274660 243176 274712
rect 243228 274700 243234 274712
rect 249058 274700 249064 274712
rect 243228 274672 249064 274700
rect 243228 274660 243234 274672
rect 249058 274660 249064 274672
rect 249116 274660 249122 274712
rect 289262 274660 289268 274712
rect 289320 274700 289326 274712
rect 292758 274700 292764 274712
rect 289320 274672 292764 274700
rect 289320 274660 289326 274672
rect 292758 274660 292764 274672
rect 292816 274660 292822 274712
rect 296346 274660 296352 274712
rect 296404 274700 296410 274712
rect 298370 274700 298376 274712
rect 296404 274672 298376 274700
rect 296404 274660 296410 274672
rect 298370 274660 298376 274672
rect 298428 274660 298434 274712
rect 298738 274660 298744 274712
rect 298796 274700 298802 274712
rect 300118 274700 300124 274712
rect 298796 274672 300124 274700
rect 298796 274660 298802 274672
rect 300118 274660 300124 274672
rect 300176 274660 300182 274712
rect 324958 274660 324964 274712
rect 325016 274700 325022 274712
rect 327074 274700 327080 274712
rect 325016 274672 327080 274700
rect 325016 274660 325022 274672
rect 327074 274660 327080 274672
rect 327132 274660 327138 274712
rect 338022 274660 338028 274712
rect 338080 274700 338086 274712
rect 343634 274700 343640 274712
rect 338080 274672 343640 274700
rect 338080 274660 338086 274672
rect 343634 274660 343640 274672
rect 343692 274660 343698 274712
rect 344278 274660 344284 274712
rect 344336 274700 344342 274712
rect 347222 274700 347228 274712
rect 344336 274672 347228 274700
rect 344336 274660 344342 274672
rect 347222 274660 347228 274672
rect 347280 274660 347286 274712
rect 347406 274660 347412 274712
rect 347464 274700 347470 274712
rect 349614 274700 349620 274712
rect 347464 274672 349620 274700
rect 347464 274660 347470 274672
rect 349614 274660 349620 274672
rect 349672 274660 349678 274712
rect 360194 274660 360200 274712
rect 360252 274700 360258 274712
rect 363782 274700 363788 274712
rect 360252 274672 363788 274700
rect 360252 274660 360258 274672
rect 363782 274660 363788 274672
rect 363840 274660 363846 274712
rect 478966 274660 478972 274712
rect 479024 274700 479030 274712
rect 482002 274700 482008 274712
rect 479024 274672 482008 274700
rect 479024 274660 479030 274672
rect 482002 274660 482008 274672
rect 482060 274660 482066 274712
rect 619174 274660 619180 274712
rect 619232 274700 619238 274712
rect 623866 274700 623872 274712
rect 619232 274672 623872 274700
rect 619232 274660 619238 274672
rect 623866 274660 623872 274672
rect 623924 274660 623930 274712
rect 120258 274592 120264 274644
rect 120316 274632 120322 274644
rect 175274 274632 175280 274644
rect 120316 274604 175280 274632
rect 120316 274592 120322 274604
rect 175274 274592 175280 274604
rect 175332 274592 175338 274644
rect 384942 274592 384948 274644
rect 385000 274632 385006 274644
rect 400214 274632 400220 274644
rect 385000 274604 400220 274632
rect 385000 274592 385006 274604
rect 400214 274592 400220 274604
rect 400272 274592 400278 274644
rect 403986 274592 403992 274644
rect 404044 274632 404050 274644
rect 438854 274632 438860 274644
rect 404044 274604 438860 274632
rect 404044 274592 404050 274604
rect 438854 274592 438860 274604
rect 438912 274592 438918 274644
rect 445018 274592 445024 274644
rect 445076 274632 445082 274644
rect 478414 274632 478420 274644
rect 445076 274604 478420 274632
rect 445076 274592 445082 274604
rect 478414 274592 478420 274604
rect 478472 274592 478478 274644
rect 482186 274592 482192 274644
rect 482244 274632 482250 274644
rect 556430 274632 556436 274644
rect 482244 274604 556436 274632
rect 482244 274592 482250 274604
rect 556430 274592 556436 274604
rect 556488 274592 556494 274644
rect 559742 274592 559748 274644
rect 559800 274632 559806 274644
rect 587158 274632 587164 274644
rect 559800 274604 587164 274632
rect 559800 274592 559806 274604
rect 587158 274592 587164 274604
rect 587216 274592 587222 274644
rect 114278 274456 114284 274508
rect 114336 274496 114342 274508
rect 171594 274496 171600 274508
rect 114336 274468 171600 274496
rect 114336 274456 114342 274468
rect 171594 274456 171600 274468
rect 171652 274456 171658 274508
rect 179322 274456 179328 274508
rect 179380 274496 179386 274508
rect 213178 274496 213184 274508
rect 179380 274468 213184 274496
rect 179380 274456 179386 274468
rect 213178 274456 213184 274468
rect 213236 274456 213242 274508
rect 213638 274456 213644 274508
rect 213696 274496 213702 274508
rect 240410 274496 240416 274508
rect 213696 274468 240416 274496
rect 213696 274456 213702 274468
rect 240410 274456 240416 274468
rect 240468 274456 240474 274508
rect 378778 274456 378784 274508
rect 378836 274496 378842 274508
rect 378836 274468 393314 274496
rect 378836 274456 378842 274468
rect 93026 274320 93032 274372
rect 93084 274360 93090 274372
rect 95878 274360 95884 274372
rect 93084 274332 95884 274360
rect 93084 274320 93090 274332
rect 95878 274320 95884 274332
rect 95936 274320 95942 274372
rect 97718 274320 97724 274372
rect 97776 274360 97782 274372
rect 158806 274360 158812 274372
rect 97776 274332 158812 274360
rect 97776 274320 97782 274332
rect 158806 274320 158812 274332
rect 158864 274320 158870 274372
rect 180518 274320 180524 274372
rect 180576 274360 180582 274372
rect 216950 274360 216956 274372
rect 180576 274332 216956 274360
rect 180576 274320 180582 274332
rect 216950 274320 216956 274332
rect 217008 274320 217014 274372
rect 368290 274320 368296 274372
rect 368348 274360 368354 274372
rect 387702 274360 387708 274372
rect 368348 274332 387708 274360
rect 368348 274320 368354 274332
rect 387702 274320 387708 274332
rect 387760 274320 387766 274372
rect 95418 274184 95424 274236
rect 95476 274224 95482 274236
rect 157610 274224 157616 274236
rect 95476 274196 157616 274224
rect 95476 274184 95482 274196
rect 157610 274184 157616 274196
rect 157668 274184 157674 274236
rect 165614 274184 165620 274236
rect 165672 274224 165678 274236
rect 205726 274224 205732 274236
rect 165672 274196 205732 274224
rect 165672 274184 165678 274196
rect 205726 274184 205732 274196
rect 205784 274184 205790 274236
rect 206554 274184 206560 274236
rect 206612 274224 206618 274236
rect 234614 274224 234620 274236
rect 206612 274196 234620 274224
rect 206612 274184 206618 274196
rect 234614 274184 234620 274196
rect 234672 274184 234678 274236
rect 245654 274184 245660 274236
rect 245712 274224 245718 274236
rect 254026 274224 254032 274236
rect 245712 274196 254032 274224
rect 245712 274184 245718 274196
rect 254026 274184 254032 274196
rect 254084 274184 254090 274236
rect 351178 274184 351184 274236
rect 351236 274224 351242 274236
rect 362586 274224 362592 274236
rect 351236 274196 362592 274224
rect 351236 274184 351242 274196
rect 362586 274184 362592 274196
rect 362644 274184 362650 274236
rect 386230 274224 386236 274236
rect 373966 274196 386236 274224
rect 77662 274048 77668 274100
rect 77720 274088 77726 274100
rect 145098 274088 145104 274100
rect 77720 274060 145104 274088
rect 77720 274048 77726 274060
rect 145098 274048 145104 274060
rect 145156 274048 145162 274100
rect 145282 274048 145288 274100
rect 145340 274088 145346 274100
rect 189810 274088 189816 274100
rect 145340 274060 189816 274088
rect 145340 274048 145346 274060
rect 189810 274048 189816 274060
rect 189868 274048 189874 274100
rect 191190 274048 191196 274100
rect 191248 274088 191254 274100
rect 224770 274088 224776 274100
rect 191248 274060 224776 274088
rect 191248 274048 191254 274060
rect 224770 274048 224776 274060
rect 224828 274048 224834 274100
rect 224954 274048 224960 274100
rect 225012 274088 225018 274100
rect 245746 274088 245752 274100
rect 225012 274060 245752 274088
rect 225012 274048 225018 274060
rect 245746 274048 245752 274060
rect 245804 274048 245810 274100
rect 253474 274048 253480 274100
rect 253532 274088 253538 274100
rect 265250 274088 265256 274100
rect 253532 274060 265256 274088
rect 253532 274048 253538 274060
rect 265250 274048 265256 274060
rect 265308 274048 265314 274100
rect 339126 274048 339132 274100
rect 339184 274088 339190 274100
rect 353110 274088 353116 274100
rect 339184 274060 353116 274088
rect 339184 274048 339190 274060
rect 353110 274048 353116 274060
rect 353168 274048 353174 274100
rect 362770 274048 362776 274100
rect 362828 274088 362834 274100
rect 373966 274088 373994 274196
rect 386230 274184 386236 274196
rect 386288 274184 386294 274236
rect 393286 274224 393314 274468
rect 400122 274456 400128 274508
rect 400180 274496 400186 274508
rect 419534 274496 419540 274508
rect 400180 274468 419540 274496
rect 400180 274456 400186 274468
rect 419534 274456 419540 274468
rect 419592 274456 419598 274508
rect 420730 274456 420736 274508
rect 420788 274496 420794 274508
rect 470134 274496 470140 274508
rect 420788 274468 470140 274496
rect 420788 274456 420794 274468
rect 470134 274456 470140 274468
rect 470192 274456 470198 274508
rect 474366 274456 474372 274508
rect 474424 274496 474430 274508
rect 523678 274496 523684 274508
rect 474424 274468 523684 274496
rect 474424 274456 474430 274468
rect 523678 274456 523684 274468
rect 523736 274456 523742 274508
rect 537478 274456 537484 274508
rect 537536 274496 537542 274508
rect 613194 274496 613200 274508
rect 537536 274468 613200 274496
rect 537536 274456 537542 274468
rect 613194 274456 613200 274468
rect 613252 274456 613258 274508
rect 397270 274320 397276 274372
rect 397328 274360 397334 274372
rect 418338 274360 418344 274372
rect 397328 274332 418344 274360
rect 397328 274320 397334 274332
rect 418338 274320 418344 274332
rect 418396 274320 418402 274372
rect 419166 274320 419172 274372
rect 419224 274360 419230 274372
rect 467834 274360 467840 274372
rect 419224 274332 467840 274360
rect 419224 274320 419230 274332
rect 467834 274320 467840 274332
rect 467892 274320 467898 274372
rect 479334 274360 479340 274372
rect 470566 274332 479340 274360
rect 408678 274224 408684 274236
rect 393286 274196 408684 274224
rect 408678 274184 408684 274196
rect 408736 274184 408742 274236
rect 427446 274184 427452 274236
rect 427504 274224 427510 274236
rect 470566 274224 470594 274332
rect 479334 274320 479340 274332
rect 479392 274320 479398 274372
rect 479518 274320 479524 274372
rect 479576 274360 479582 274372
rect 481542 274360 481548 274372
rect 479576 274332 481548 274360
rect 479576 274320 479582 274332
rect 481542 274320 481548 274332
rect 481600 274320 481606 274372
rect 487062 274320 487068 274372
rect 487120 274360 487126 274372
rect 563514 274360 563520 274372
rect 487120 274332 563520 274360
rect 487120 274320 487126 274332
rect 563514 274320 563520 274332
rect 563572 274320 563578 274372
rect 563698 274320 563704 274372
rect 563756 274360 563762 274372
rect 611998 274360 612004 274372
rect 563756 274332 612004 274360
rect 563756 274320 563762 274332
rect 611998 274320 612004 274332
rect 612056 274320 612062 274372
rect 427504 274196 470594 274224
rect 427504 274184 427510 274196
rect 471974 274184 471980 274236
rect 472032 274224 472038 274236
rect 472032 274196 480254 274224
rect 472032 274184 472038 274196
rect 362828 274060 373994 274088
rect 362828 274048 362834 274060
rect 385678 274048 385684 274100
rect 385736 274088 385742 274100
rect 395154 274088 395160 274100
rect 385736 274060 395160 274088
rect 385736 274048 385742 274060
rect 395154 274048 395160 274060
rect 395212 274048 395218 274100
rect 395614 274048 395620 274100
rect 395672 274088 395678 274100
rect 426434 274088 426440 274100
rect 395672 274060 426440 274088
rect 395672 274048 395678 274060
rect 426434 274048 426440 274060
rect 426492 274048 426498 274100
rect 446582 274048 446588 274100
rect 446640 274088 446646 274100
rect 468938 274088 468944 274100
rect 446640 274060 468944 274088
rect 446640 274048 446646 274060
rect 468938 274048 468944 274060
rect 468996 274048 469002 274100
rect 469122 274048 469128 274100
rect 469180 274088 469186 274100
rect 469180 274060 475424 274088
rect 469180 274048 469186 274060
rect 75270 273912 75276 273964
rect 75328 273952 75334 273964
rect 142154 273952 142160 273964
rect 75328 273924 142160 273952
rect 75328 273912 75334 273924
rect 142154 273912 142160 273924
rect 142212 273912 142218 273964
rect 147398 273912 147404 273964
rect 147456 273952 147462 273964
rect 193306 273952 193312 273964
rect 147456 273924 193312 273952
rect 147456 273912 147462 273924
rect 193306 273912 193312 273924
rect 193364 273912 193370 273964
rect 193490 273912 193496 273964
rect 193548 273952 193554 273964
rect 222838 273952 222844 273964
rect 193548 273924 222844 273952
rect 193548 273912 193554 273924
rect 222838 273912 222844 273924
rect 222896 273912 222902 273964
rect 223114 273912 223120 273964
rect 223172 273952 223178 273964
rect 223172 273924 238754 273952
rect 223172 273912 223178 273924
rect 130838 273776 130844 273828
rect 130896 273816 130902 273828
rect 181438 273816 181444 273828
rect 130896 273788 181444 273816
rect 130896 273776 130902 273788
rect 181438 273776 181444 273788
rect 181496 273776 181502 273828
rect 238726 273816 238754 273924
rect 247034 273912 247040 273964
rect 247092 273952 247098 273964
rect 262214 273952 262220 273964
rect 247092 273924 262220 273952
rect 247092 273912 247098 273924
rect 262214 273912 262220 273924
rect 262272 273912 262278 273964
rect 265618 273912 265624 273964
rect 265676 273952 265682 273964
rect 276842 273952 276848 273964
rect 265676 273924 276848 273952
rect 265676 273912 265682 273924
rect 276842 273912 276848 273924
rect 276900 273912 276906 273964
rect 322750 273912 322756 273964
rect 322808 273952 322814 273964
rect 330662 273952 330668 273964
rect 322808 273924 330668 273952
rect 322808 273912 322814 273924
rect 330662 273912 330668 273924
rect 330720 273912 330726 273964
rect 333790 273912 333796 273964
rect 333848 273952 333854 273964
rect 344830 273952 344836 273964
rect 333848 273924 344836 273952
rect 333848 273912 333854 273924
rect 344830 273912 344836 273924
rect 344888 273912 344894 273964
rect 366358 273952 366364 273964
rect 354646 273924 366364 273952
rect 247034 273816 247040 273828
rect 238726 273788 247040 273816
rect 247034 273776 247040 273788
rect 247092 273776 247098 273828
rect 344646 273776 344652 273828
rect 344704 273816 344710 273828
rect 349798 273816 349804 273828
rect 344704 273788 349804 273816
rect 344704 273776 344710 273788
rect 349798 273776 349804 273788
rect 349856 273776 349862 273828
rect 350350 273776 350356 273828
rect 350408 273816 350414 273828
rect 354646 273816 354674 273924
rect 366358 273912 366364 273924
rect 366416 273912 366422 273964
rect 367002 273912 367008 273964
rect 367060 273952 367066 273964
rect 376662 273952 376668 273964
rect 367060 273924 376668 273952
rect 367060 273912 367066 273924
rect 376662 273912 376668 273924
rect 376720 273912 376726 273964
rect 407482 273952 407488 273964
rect 383626 273924 407488 273952
rect 350408 273788 354674 273816
rect 350408 273776 350414 273788
rect 376570 273776 376576 273828
rect 376628 273816 376634 273828
rect 383626 273816 383654 273924
rect 407482 273912 407488 273924
rect 407540 273912 407546 273964
rect 409230 273912 409236 273964
rect 409288 273952 409294 273964
rect 446398 273952 446404 273964
rect 409288 273924 446404 273952
rect 409288 273912 409294 273924
rect 446398 273912 446404 273924
rect 446456 273912 446462 273964
rect 468478 273912 468484 273964
rect 468536 273952 468542 273964
rect 471974 273952 471980 273964
rect 468536 273924 471980 273952
rect 468536 273912 468542 273924
rect 471974 273912 471980 273924
rect 472032 273912 472038 273964
rect 475396 273952 475424 274060
rect 475562 274048 475568 274100
rect 475620 274088 475626 274100
rect 479518 274088 479524 274100
rect 475620 274060 479524 274088
rect 475620 274048 475626 274060
rect 479518 274048 479524 274060
rect 479576 274048 479582 274100
rect 480226 274088 480254 274196
rect 481358 274184 481364 274236
rect 481416 274224 481422 274236
rect 482186 274224 482192 274236
rect 481416 274196 482192 274224
rect 481416 274184 481422 274196
rect 482186 274184 482192 274196
rect 482244 274184 482250 274236
rect 500862 274184 500868 274236
rect 500920 274224 500926 274236
rect 583662 274224 583668 274236
rect 500920 274196 583668 274224
rect 500920 274184 500926 274196
rect 583662 274184 583668 274196
rect 583720 274184 583726 274236
rect 494974 274088 494980 274100
rect 480226 274060 494980 274088
rect 494974 274048 494980 274060
rect 495032 274048 495038 274100
rect 533430 274048 533436 274100
rect 533488 274088 533494 274100
rect 630950 274088 630956 274100
rect 533488 274060 630956 274088
rect 533488 274048 533494 274060
rect 630950 274048 630956 274060
rect 631008 274048 631014 274100
rect 532786 273952 532792 273964
rect 475396 273924 532792 273952
rect 532786 273912 532792 273924
rect 532844 273912 532850 273964
rect 542078 273912 542084 273964
rect 542136 273952 542142 273964
rect 642726 273952 642732 273964
rect 542136 273924 642732 273952
rect 542136 273912 542142 273924
rect 642726 273912 642732 273924
rect 642784 273912 642790 273964
rect 376628 273788 383654 273816
rect 376628 273776 376634 273788
rect 431678 273776 431684 273828
rect 431736 273816 431742 273828
rect 485498 273816 485504 273828
rect 431736 273788 485504 273816
rect 431736 273776 431742 273788
rect 485498 273776 485504 273788
rect 485556 273776 485562 273828
rect 488350 273776 488356 273828
rect 488408 273816 488414 273828
rect 559558 273816 559564 273828
rect 488408 273788 559564 273816
rect 488408 273776 488414 273788
rect 559558 273776 559564 273788
rect 559616 273776 559622 273828
rect 124950 273640 124956 273692
rect 125008 273680 125014 273692
rect 148410 273680 148416 273692
rect 125008 273652 148416 273680
rect 125008 273640 125014 273652
rect 148410 273640 148416 273652
rect 148468 273640 148474 273692
rect 155678 273640 155684 273692
rect 155736 273680 155742 273692
rect 198090 273680 198096 273692
rect 155736 273652 198096 273680
rect 155736 273640 155742 273652
rect 198090 273640 198096 273652
rect 198148 273640 198154 273692
rect 457438 273640 457444 273692
rect 457496 273680 457502 273692
rect 484302 273680 484308 273692
rect 457496 273652 484308 273680
rect 457496 273640 457502 273652
rect 484302 273640 484308 273652
rect 484360 273640 484366 273692
rect 484486 273640 484492 273692
rect 484544 273680 484550 273692
rect 552658 273680 552664 273692
rect 484544 273652 552664 273680
rect 484544 273640 484550 273652
rect 552658 273640 552664 273652
rect 552716 273640 552722 273692
rect 439314 273504 439320 273556
rect 439372 273544 439378 273556
rect 471330 273544 471336 273556
rect 439372 273516 471336 273544
rect 439372 273504 439378 273516
rect 471330 273504 471336 273516
rect 471388 273504 471394 273556
rect 473078 273504 473084 273556
rect 473136 273544 473142 273556
rect 475562 273544 475568 273556
rect 473136 273516 475568 273544
rect 473136 273504 473142 273516
rect 475562 273504 475568 273516
rect 475620 273504 475626 273556
rect 478782 273504 478788 273556
rect 478840 273544 478846 273556
rect 546034 273544 546040 273556
rect 478840 273516 546040 273544
rect 478840 273504 478846 273516
rect 546034 273504 546040 273516
rect 546092 273504 546098 273556
rect 552658 273504 552664 273556
rect 552716 273544 552722 273556
rect 580074 273544 580080 273556
rect 552716 273516 580080 273544
rect 552716 273504 552722 273516
rect 580074 273504 580080 273516
rect 580132 273504 580138 273556
rect 464798 273368 464804 273420
rect 464856 273408 464862 273420
rect 469122 273408 469128 273420
rect 464856 273380 469128 273408
rect 464856 273368 464862 273380
rect 469122 273368 469128 273380
rect 469180 273368 469186 273420
rect 475930 273368 475936 273420
rect 475988 273408 475994 273420
rect 542262 273408 542268 273420
rect 475988 273380 542268 273408
rect 475988 273368 475994 273380
rect 542262 273368 542268 273380
rect 542320 273368 542326 273420
rect 330478 273232 330484 273284
rect 330536 273272 330542 273284
rect 333054 273272 333060 273284
rect 330536 273244 333060 273272
rect 330536 273232 330542 273244
rect 333054 273232 333060 273244
rect 333112 273232 333118 273284
rect 127342 273164 127348 273216
rect 127400 273204 127406 273216
rect 179874 273204 179880 273216
rect 127400 273176 179880 273204
rect 127400 273164 127406 273176
rect 179874 273164 179880 273176
rect 179932 273164 179938 273216
rect 401502 273164 401508 273216
rect 401560 273204 401566 273216
rect 427814 273204 427820 273216
rect 401560 273176 427820 273204
rect 401560 273164 401566 273176
rect 427814 273164 427820 273176
rect 427872 273164 427878 273216
rect 438118 273164 438124 273216
rect 438176 273204 438182 273216
rect 464246 273204 464252 273216
rect 438176 273176 464252 273204
rect 438176 273164 438182 273176
rect 464246 273164 464252 273176
rect 464304 273164 464310 273216
rect 471606 273164 471612 273216
rect 471664 273204 471670 273216
rect 543458 273204 543464 273216
rect 471664 273176 543464 273204
rect 471664 273164 471670 273176
rect 543458 273164 543464 273176
rect 543516 273164 543522 273216
rect 111978 273028 111984 273080
rect 112036 273068 112042 273080
rect 168374 273068 168380 273080
rect 112036 273040 168380 273068
rect 112036 273028 112042 273040
rect 168374 273028 168380 273040
rect 168432 273028 168438 273080
rect 182082 273028 182088 273080
rect 182140 273068 182146 273080
rect 207290 273068 207296 273080
rect 182140 273040 207296 273068
rect 182140 273028 182146 273040
rect 207290 273028 207296 273040
rect 207348 273028 207354 273080
rect 381998 273028 382004 273080
rect 382056 273068 382062 273080
rect 414566 273068 414572 273080
rect 382056 273040 414572 273068
rect 382056 273028 382062 273040
rect 414566 273028 414572 273040
rect 414624 273028 414630 273080
rect 429838 273028 429844 273080
rect 429896 273068 429902 273080
rect 447686 273068 447692 273080
rect 429896 273040 447692 273068
rect 429896 273028 429902 273040
rect 447686 273028 447692 273040
rect 447744 273028 447750 273080
rect 451090 273028 451096 273080
rect 451148 273068 451154 273080
rect 513926 273068 513932 273080
rect 451148 273040 513932 273068
rect 451148 273028 451154 273040
rect 513926 273028 513932 273040
rect 513984 273028 513990 273080
rect 520090 273028 520096 273080
rect 520148 273068 520154 273080
rect 610802 273068 610808 273080
rect 520148 273040 610808 273068
rect 520148 273028 520154 273040
rect 610802 273028 610808 273040
rect 610860 273028 610866 273080
rect 102502 272892 102508 272944
rect 102560 272932 102566 272944
rect 162118 272932 162124 272944
rect 102560 272904 162124 272932
rect 102560 272892 102566 272904
rect 162118 272892 162124 272904
rect 162176 272892 162182 272944
rect 189994 272892 190000 272944
rect 190052 272932 190058 272944
rect 190052 272904 213592 272932
rect 190052 272892 190058 272904
rect 94222 272756 94228 272808
rect 94280 272796 94286 272808
rect 155954 272796 155960 272808
rect 94280 272768 155960 272796
rect 94280 272756 94286 272768
rect 155954 272756 155960 272768
rect 156012 272756 156018 272808
rect 187602 272756 187608 272808
rect 187660 272796 187666 272808
rect 212534 272796 212540 272808
rect 187660 272768 212540 272796
rect 187660 272756 187666 272768
rect 212534 272756 212540 272768
rect 212592 272756 212598 272808
rect 213564 272796 213592 272904
rect 217134 272892 217140 272944
rect 217192 272932 217198 272944
rect 242986 272932 242992 272944
rect 217192 272904 242992 272932
rect 217192 272892 217198 272904
rect 242986 272892 242992 272904
rect 243044 272892 243050 272944
rect 286870 272892 286876 272944
rect 286928 272932 286934 272944
rect 287698 272932 287704 272944
rect 286928 272904 287704 272932
rect 286928 272892 286934 272904
rect 287698 272892 287704 272904
rect 287756 272892 287762 272944
rect 388806 272892 388812 272944
rect 388864 272932 388870 272944
rect 400398 272932 400404 272944
rect 388864 272904 400404 272932
rect 388864 272892 388870 272904
rect 400398 272892 400404 272904
rect 400456 272892 400462 272944
rect 406838 272892 406844 272944
rect 406896 272932 406902 272944
rect 450078 272932 450084 272944
rect 406896 272904 450084 272932
rect 406896 272892 406902 272904
rect 450078 272892 450084 272904
rect 450136 272892 450142 272944
rect 457990 272892 457996 272944
rect 458048 272932 458054 272944
rect 522206 272932 522212 272944
rect 458048 272904 522212 272932
rect 458048 272892 458054 272904
rect 522206 272892 522212 272904
rect 522264 272892 522270 272944
rect 524046 272892 524052 272944
rect 524104 272932 524110 272944
rect 617978 272932 617984 272944
rect 524104 272904 617984 272932
rect 524104 272892 524110 272904
rect 617978 272892 617984 272904
rect 618036 272892 618042 272944
rect 217410 272796 217416 272808
rect 213564 272768 217416 272796
rect 217410 272756 217416 272768
rect 217468 272756 217474 272808
rect 219894 272756 219900 272808
rect 219952 272796 219958 272808
rect 239214 272796 239220 272808
rect 219952 272768 239220 272796
rect 219952 272756 219958 272768
rect 239214 272756 239220 272768
rect 239272 272756 239278 272808
rect 252646 272756 252652 272808
rect 252704 272796 252710 272808
rect 267826 272796 267832 272808
rect 252704 272768 267832 272796
rect 252704 272756 252710 272768
rect 267826 272756 267832 272768
rect 267884 272756 267890 272808
rect 343542 272756 343548 272808
rect 343600 272796 343606 272808
rect 358998 272796 359004 272808
rect 343600 272768 359004 272796
rect 343600 272756 343606 272768
rect 358998 272756 359004 272768
rect 359056 272756 359062 272808
rect 360838 272756 360844 272808
rect 360896 272796 360902 272808
rect 381538 272796 381544 272808
rect 360896 272768 381544 272796
rect 360896 272756 360902 272768
rect 381538 272756 381544 272768
rect 381596 272756 381602 272808
rect 394326 272756 394332 272808
rect 394384 272796 394390 272808
rect 407758 272796 407764 272808
rect 394384 272768 407764 272796
rect 394384 272756 394390 272768
rect 407758 272756 407764 272768
rect 407816 272756 407822 272808
rect 408402 272756 408408 272808
rect 408460 272796 408466 272808
rect 452102 272796 452108 272808
rect 408460 272768 452108 272796
rect 408460 272756 408466 272768
rect 452102 272756 452108 272768
rect 452160 272756 452166 272808
rect 452286 272756 452292 272808
rect 452344 272796 452350 272808
rect 515122 272796 515128 272808
rect 452344 272768 515128 272796
rect 452344 272756 452350 272768
rect 515122 272756 515128 272768
rect 515180 272756 515186 272808
rect 517330 272756 517336 272808
rect 517388 272796 517394 272808
rect 525794 272796 525800 272808
rect 517388 272768 525800 272796
rect 517388 272756 517394 272768
rect 525794 272756 525800 272768
rect 525852 272756 525858 272808
rect 526806 272756 526812 272808
rect 526864 272796 526870 272808
rect 621474 272796 621480 272808
rect 526864 272768 621480 272796
rect 526864 272756 526870 272768
rect 621474 272756 621480 272768
rect 621532 272756 621538 272808
rect 82354 272620 82360 272672
rect 82412 272660 82418 272672
rect 148226 272660 148232 272672
rect 82412 272632 148232 272660
rect 82412 272620 82418 272632
rect 148226 272620 148232 272632
rect 148284 272620 148290 272672
rect 161566 272620 161572 272672
rect 161624 272660 161630 272672
rect 203058 272660 203064 272672
rect 161624 272632 203064 272660
rect 161624 272620 161630 272632
rect 203058 272620 203064 272632
rect 203116 272620 203122 272672
rect 203242 272620 203248 272672
rect 203300 272660 203306 272672
rect 233234 272660 233240 272672
rect 203300 272632 233240 272660
rect 203300 272620 203306 272632
rect 233234 272620 233240 272632
rect 233292 272620 233298 272672
rect 239582 272620 239588 272672
rect 239640 272660 239646 272672
rect 254578 272660 254584 272672
rect 239640 272632 254584 272660
rect 239640 272620 239646 272632
rect 254578 272620 254584 272632
rect 254636 272620 254642 272672
rect 280982 272620 280988 272672
rect 281040 272660 281046 272672
rect 286318 272660 286324 272672
rect 281040 272632 286324 272660
rect 281040 272620 281046 272632
rect 286318 272620 286324 272632
rect 286376 272620 286382 272672
rect 349798 272620 349804 272672
rect 349856 272660 349862 272672
rect 366082 272660 366088 272672
rect 349856 272632 366088 272660
rect 349856 272620 349862 272632
rect 366082 272620 366088 272632
rect 366140 272620 366146 272672
rect 370958 272620 370964 272672
rect 371016 272660 371022 272672
rect 399202 272660 399208 272672
rect 371016 272632 399208 272660
rect 371016 272620 371022 272632
rect 399202 272620 399208 272632
rect 399260 272620 399266 272672
rect 412266 272620 412272 272672
rect 412324 272660 412330 272672
rect 457162 272660 457168 272672
rect 412324 272632 457168 272660
rect 412324 272620 412330 272632
rect 457162 272620 457168 272632
rect 457220 272620 457226 272672
rect 461946 272620 461952 272672
rect 462004 272660 462010 272672
rect 529290 272660 529296 272672
rect 462004 272632 529296 272660
rect 462004 272620 462010 272632
rect 529290 272620 529296 272632
rect 529348 272620 529354 272672
rect 529750 272620 529756 272672
rect 529808 272660 529814 272672
rect 625062 272660 625068 272672
rect 529808 272632 625068 272660
rect 529808 272620 529814 272632
rect 625062 272620 625068 272632
rect 625120 272620 625126 272672
rect 65886 272484 65892 272536
rect 65944 272524 65950 272536
rect 136818 272524 136824 272536
rect 65944 272496 136824 272524
rect 65944 272484 65950 272496
rect 136818 272484 136824 272496
rect 136876 272484 136882 272536
rect 137922 272484 137928 272536
rect 137980 272524 137986 272536
rect 187694 272524 187700 272536
rect 137980 272496 187700 272524
rect 137980 272484 137986 272496
rect 187694 272484 187700 272496
rect 187752 272484 187758 272536
rect 192294 272484 192300 272536
rect 192352 272524 192358 272536
rect 225506 272524 225512 272536
rect 192352 272496 225512 272524
rect 192352 272484 192358 272496
rect 225506 272484 225512 272496
rect 225564 272484 225570 272536
rect 236086 272484 236092 272536
rect 236144 272524 236150 272536
rect 253198 272524 253204 272536
rect 236144 272496 253204 272524
rect 236144 272484 236150 272496
rect 253198 272484 253204 272496
rect 253256 272484 253262 272536
rect 255038 272484 255044 272536
rect 255096 272524 255102 272536
rect 269298 272524 269304 272536
rect 255096 272496 269304 272524
rect 255096 272484 255102 272496
rect 269298 272484 269304 272496
rect 269356 272484 269362 272536
rect 270218 272484 270224 272536
rect 270276 272524 270282 272536
rect 280338 272524 280344 272536
rect 270276 272496 280344 272524
rect 270276 272484 270282 272496
rect 280338 272484 280344 272496
rect 280396 272484 280402 272536
rect 331030 272484 331036 272536
rect 331088 272524 331094 272536
rect 342438 272524 342444 272536
rect 331088 272496 342444 272524
rect 331088 272484 331094 272496
rect 342438 272484 342444 272496
rect 342496 272484 342502 272536
rect 356882 272484 356888 272536
rect 356940 272524 356946 272536
rect 376846 272524 376852 272536
rect 356940 272496 376852 272524
rect 356940 272484 356946 272496
rect 376846 272484 376852 272496
rect 376904 272484 376910 272536
rect 380802 272484 380808 272536
rect 380860 272524 380866 272536
rect 411990 272524 411996 272536
rect 380860 272496 411996 272524
rect 380860 272484 380866 272496
rect 411990 272484 411996 272496
rect 412048 272484 412054 272536
rect 413922 272484 413928 272536
rect 413980 272524 413986 272536
rect 460658 272524 460664 272536
rect 413980 272496 460664 272524
rect 413980 272484 413986 272496
rect 460658 272484 460664 272496
rect 460716 272484 460722 272536
rect 467742 272484 467748 272536
rect 467800 272524 467806 272536
rect 536374 272524 536380 272536
rect 467800 272496 536380 272524
rect 467800 272484 467806 272496
rect 536374 272484 536380 272496
rect 536432 272484 536438 272536
rect 539318 272484 539324 272536
rect 539376 272524 539382 272536
rect 639230 272524 639236 272536
rect 539376 272496 639236 272524
rect 539376 272484 539382 272496
rect 639230 272484 639236 272496
rect 639288 272484 639294 272536
rect 128538 272348 128544 272400
rect 128596 272388 128602 272400
rect 181254 272388 181260 272400
rect 128596 272360 181260 272388
rect 128596 272348 128602 272360
rect 181254 272348 181260 272360
rect 181312 272348 181318 272400
rect 212534 272348 212540 272400
rect 212592 272388 212598 272400
rect 218790 272388 218796 272400
rect 212592 272360 218796 272388
rect 212592 272348 212598 272360
rect 218790 272348 218796 272360
rect 218848 272348 218854 272400
rect 457806 272348 457812 272400
rect 457864 272388 457870 272400
rect 466822 272388 466828 272400
rect 457864 272360 466828 272388
rect 457864 272348 457870 272360
rect 466822 272348 466828 272360
rect 466880 272348 466886 272400
rect 470502 272348 470508 272400
rect 470560 272388 470566 272400
rect 539870 272388 539876 272400
rect 470560 272360 539876 272388
rect 470560 272348 470566 272360
rect 539870 272348 539876 272360
rect 539928 272348 539934 272400
rect 541618 272348 541624 272400
rect 541676 272388 541682 272400
rect 603718 272388 603724 272400
rect 541676 272360 603724 272388
rect 541676 272348 541682 272360
rect 603718 272348 603724 272360
rect 603776 272348 603782 272400
rect 116670 272212 116676 272264
rect 116728 272252 116734 272264
rect 166074 272252 166080 272264
rect 116728 272224 166080 272252
rect 116728 272212 116734 272224
rect 166074 272212 166080 272224
rect 166132 272212 166138 272264
rect 166258 272212 166264 272264
rect 166316 272252 166322 272264
rect 191834 272252 191840 272264
rect 166316 272224 191840 272252
rect 166316 272212 166322 272224
rect 191834 272212 191840 272224
rect 191892 272212 191898 272264
rect 424962 272212 424968 272264
rect 425020 272252 425026 272264
rect 474918 272252 474924 272264
rect 425020 272224 474924 272252
rect 425020 272212 425026 272224
rect 474918 272212 474924 272224
rect 474976 272212 474982 272264
rect 479702 272212 479708 272264
rect 479760 272252 479766 272264
rect 548150 272252 548156 272264
rect 479760 272224 548156 272252
rect 479760 272212 479766 272224
rect 548150 272212 548156 272224
rect 548208 272212 548214 272264
rect 152182 272076 152188 272128
rect 152240 272116 152246 272128
rect 192478 272116 192484 272128
rect 152240 272088 192484 272116
rect 152240 272076 152246 272088
rect 192478 272076 192484 272088
rect 192536 272076 192542 272128
rect 447778 272076 447784 272128
rect 447836 272116 447842 272128
rect 506842 272116 506848 272128
rect 447836 272088 506848 272116
rect 447836 272076 447842 272088
rect 506842 272076 506848 272088
rect 506900 272076 506906 272128
rect 514018 272076 514024 272128
rect 514076 272116 514082 272128
rect 565906 272116 565912 272128
rect 514076 272088 565912 272116
rect 514076 272076 514082 272088
rect 565906 272076 565912 272088
rect 565964 272076 565970 272128
rect 121362 271804 121368 271856
rect 121420 271844 121426 271856
rect 176746 271844 176752 271856
rect 121420 271816 176752 271844
rect 121420 271804 121426 271816
rect 176746 271804 176752 271816
rect 176804 271804 176810 271856
rect 185210 271804 185216 271856
rect 185268 271844 185274 271856
rect 186958 271844 186964 271856
rect 185268 271816 186964 271844
rect 185268 271804 185274 271816
rect 186958 271804 186964 271816
rect 187016 271804 187022 271856
rect 187878 271804 187884 271856
rect 187936 271844 187942 271856
rect 196434 271844 196440 271856
rect 187936 271816 196440 271844
rect 187936 271804 187942 271816
rect 196434 271804 196440 271816
rect 196492 271804 196498 271856
rect 276290 271804 276296 271856
rect 276348 271844 276354 271856
rect 278038 271844 278044 271856
rect 276348 271816 278044 271844
rect 276348 271804 276354 271816
rect 278038 271804 278044 271816
rect 278096 271804 278102 271856
rect 288066 271804 288072 271856
rect 288124 271844 288130 271856
rect 292942 271844 292948 271856
rect 288124 271816 292948 271844
rect 288124 271804 288130 271816
rect 292942 271804 292948 271816
rect 293000 271804 293006 271856
rect 293218 271804 293224 271856
rect 293276 271844 293282 271856
rect 295794 271844 295800 271856
rect 293276 271816 295800 271844
rect 293276 271804 293282 271816
rect 295794 271804 295800 271816
rect 295852 271804 295858 271856
rect 375282 271804 375288 271856
rect 375340 271844 375346 271856
rect 395430 271844 395436 271856
rect 375340 271816 395436 271844
rect 375340 271804 375346 271816
rect 395430 271804 395436 271816
rect 395488 271804 395494 271856
rect 434438 271804 434444 271856
rect 434496 271844 434502 271856
rect 490282 271844 490288 271856
rect 434496 271816 490288 271844
rect 434496 271804 434502 271816
rect 490282 271804 490288 271816
rect 490340 271804 490346 271856
rect 496538 271804 496544 271856
rect 496596 271844 496602 271856
rect 578878 271844 578884 271856
rect 496596 271816 578884 271844
rect 496596 271804 496602 271816
rect 578878 271804 578884 271816
rect 578936 271804 578942 271856
rect 318610 271736 318616 271788
rect 318668 271776 318674 271788
rect 324774 271776 324780 271788
rect 318668 271748 324780 271776
rect 318668 271736 318674 271748
rect 324774 271736 324780 271748
rect 324832 271736 324838 271788
rect 104894 271668 104900 271720
rect 104952 271708 104958 271720
rect 163314 271708 163320 271720
rect 104952 271680 163320 271708
rect 104952 271668 104958 271680
rect 163314 271668 163320 271680
rect 163372 271668 163378 271720
rect 164142 271668 164148 271720
rect 164200 271708 164206 271720
rect 194778 271708 194784 271720
rect 164200 271680 194784 271708
rect 164200 271668 164206 271680
rect 194778 271668 194784 271680
rect 194836 271668 194842 271720
rect 197078 271668 197084 271720
rect 197136 271708 197142 271720
rect 224218 271708 224224 271720
rect 197136 271680 224224 271708
rect 197136 271668 197142 271680
rect 224218 271668 224224 271680
rect 224276 271668 224282 271720
rect 224586 271668 224592 271720
rect 224644 271708 224650 271720
rect 247770 271708 247776 271720
rect 224644 271680 247776 271708
rect 224644 271668 224650 271680
rect 247770 271668 247776 271680
rect 247828 271668 247834 271720
rect 363598 271668 363604 271720
rect 363656 271708 363662 271720
rect 374362 271708 374368 271720
rect 363656 271680 374368 271708
rect 363656 271668 363662 271680
rect 374362 271668 374368 271680
rect 374420 271668 374426 271720
rect 384758 271668 384764 271720
rect 384816 271708 384822 271720
rect 415210 271708 415216 271720
rect 384816 271680 415216 271708
rect 384816 271668 384822 271680
rect 415210 271668 415216 271680
rect 415268 271668 415274 271720
rect 418798 271668 418804 271720
rect 418856 271708 418862 271720
rect 429654 271708 429660 271720
rect 418856 271680 429660 271708
rect 418856 271668 418862 271680
rect 429654 271668 429660 271680
rect 429712 271668 429718 271720
rect 437198 271668 437204 271720
rect 437256 271708 437262 271720
rect 493686 271708 493692 271720
rect 437256 271680 493692 271708
rect 437256 271668 437262 271680
rect 493686 271668 493692 271680
rect 493744 271668 493750 271720
rect 499482 271668 499488 271720
rect 499540 271708 499546 271720
rect 582466 271708 582472 271720
rect 499540 271680 582472 271708
rect 499540 271668 499546 271680
rect 582466 271668 582472 271680
rect 582524 271668 582530 271720
rect 105998 271532 106004 271584
rect 106056 271572 106062 271584
rect 164786 271572 164792 271584
rect 106056 271544 164792 271572
rect 106056 271532 106062 271544
rect 164786 271532 164792 271544
rect 164844 271532 164850 271584
rect 178126 271532 178132 271584
rect 178184 271572 178190 271584
rect 184198 271572 184204 271584
rect 178184 271544 184204 271572
rect 178184 271532 178190 271544
rect 184198 271532 184204 271544
rect 184256 271532 184262 271584
rect 184474 271532 184480 271584
rect 184532 271572 184538 271584
rect 215938 271572 215944 271584
rect 184532 271544 215944 271572
rect 184532 271532 184538 271544
rect 215938 271532 215944 271544
rect 215996 271532 216002 271584
rect 216306 271532 216312 271584
rect 216364 271572 216370 271584
rect 242066 271572 242072 271584
rect 216364 271544 242072 271572
rect 216364 271532 216370 271544
rect 242066 271532 242072 271544
rect 242124 271532 242130 271584
rect 248414 271532 248420 271584
rect 248472 271572 248478 271584
rect 264330 271572 264336 271584
rect 248472 271544 264336 271572
rect 248472 271532 248478 271544
rect 264330 271532 264336 271544
rect 264388 271532 264394 271584
rect 340598 271532 340604 271584
rect 340656 271572 340662 271584
rect 355134 271572 355140 271584
rect 340656 271544 355140 271572
rect 340656 271532 340662 271544
rect 355134 271532 355140 271544
rect 355192 271532 355198 271584
rect 355318 271532 355324 271584
rect 355376 271572 355382 271584
rect 368474 271572 368480 271584
rect 355376 271544 368480 271572
rect 355376 271532 355382 271544
rect 368474 271532 368480 271544
rect 368532 271532 368538 271584
rect 369486 271532 369492 271584
rect 369544 271572 369550 271584
rect 377398 271572 377404 271584
rect 369544 271544 377404 271572
rect 369544 271532 369550 271544
rect 377398 271532 377404 271544
rect 377456 271532 377462 271584
rect 379330 271532 379336 271584
rect 379388 271572 379394 271584
rect 393774 271572 393780 271584
rect 379388 271544 393780 271572
rect 379388 271532 379394 271544
rect 393774 271532 393780 271544
rect 393832 271532 393838 271584
rect 395522 271532 395528 271584
rect 395580 271572 395586 271584
rect 427630 271572 427636 271584
rect 395580 271544 427636 271572
rect 395580 271532 395586 271544
rect 427630 271532 427636 271544
rect 427688 271532 427694 271584
rect 431926 271544 438164 271572
rect 89530 271396 89536 271448
rect 89588 271436 89594 271448
rect 152366 271436 152372 271448
rect 89588 271408 152372 271436
rect 89588 271396 89594 271408
rect 152366 271396 152372 271408
rect 152424 271396 152430 271448
rect 162762 271396 162768 271448
rect 162820 271436 162826 271448
rect 204714 271436 204720 271448
rect 162820 271408 204720 271436
rect 162820 271396 162826 271408
rect 204714 271396 204720 271408
rect 204772 271396 204778 271448
rect 205358 271396 205364 271448
rect 205416 271436 205422 271448
rect 234982 271436 234988 271448
rect 205416 271408 234988 271436
rect 205416 271396 205422 271408
rect 234982 271396 234988 271408
rect 235040 271396 235046 271448
rect 241882 271396 241888 271448
rect 241940 271436 241946 271448
rect 260282 271436 260288 271448
rect 241940 271408 260288 271436
rect 241940 271396 241946 271408
rect 260282 271396 260288 271408
rect 260340 271396 260346 271448
rect 334618 271396 334624 271448
rect 334676 271436 334682 271448
rect 341334 271436 341340 271448
rect 334676 271408 341340 271436
rect 334676 271396 334682 271408
rect 341334 271396 341340 271408
rect 341392 271396 341398 271448
rect 348878 271396 348884 271448
rect 348936 271436 348942 271448
rect 362954 271436 362960 271448
rect 348936 271408 362960 271436
rect 348936 271396 348942 271408
rect 362954 271396 362960 271408
rect 363012 271396 363018 271448
rect 366358 271396 366364 271448
rect 366416 271436 366422 271448
rect 379146 271436 379152 271448
rect 366416 271408 379152 271436
rect 366416 271396 366422 271408
rect 379146 271396 379152 271408
rect 379204 271396 379210 271448
rect 387610 271396 387616 271448
rect 387668 271436 387674 271448
rect 421650 271436 421656 271448
rect 387668 271408 421656 271436
rect 387668 271396 387674 271408
rect 421650 271396 421656 271408
rect 421708 271396 421714 271448
rect 425698 271396 425704 271448
rect 425756 271436 425762 271448
rect 431926 271436 431954 271544
rect 425756 271408 431954 271436
rect 425756 271396 425762 271408
rect 432966 271396 432972 271448
rect 433024 271436 433030 271448
rect 437934 271436 437940 271448
rect 433024 271408 437940 271436
rect 433024 271396 433030 271408
rect 437934 271396 437940 271408
rect 437992 271396 437998 271448
rect 68186 271260 68192 271312
rect 68244 271300 68250 271312
rect 138474 271300 138480 271312
rect 68244 271272 138480 271300
rect 68244 271260 68250 271272
rect 138474 271260 138480 271272
rect 138532 271260 138538 271312
rect 139118 271260 139124 271312
rect 139176 271300 139182 271312
rect 141602 271300 141608 271312
rect 139176 271272 141608 271300
rect 139176 271260 139182 271272
rect 141602 271260 141608 271272
rect 141660 271260 141666 271312
rect 141786 271260 141792 271312
rect 141844 271300 141850 271312
rect 189626 271300 189632 271312
rect 141844 271272 189632 271300
rect 141844 271260 141850 271272
rect 189626 271260 189632 271272
rect 189684 271260 189690 271312
rect 195698 271260 195704 271312
rect 195756 271300 195762 271312
rect 227898 271300 227904 271312
rect 195756 271272 227904 271300
rect 195756 271260 195762 271272
rect 227898 271260 227904 271272
rect 227956 271260 227962 271312
rect 228818 271260 228824 271312
rect 228876 271300 228882 271312
rect 236822 271300 236828 271312
rect 228876 271272 236828 271300
rect 228876 271260 228882 271272
rect 236822 271260 236828 271272
rect 236880 271260 236886 271312
rect 237282 271260 237288 271312
rect 237340 271300 237346 271312
rect 256970 271300 256976 271312
rect 237340 271272 256976 271300
rect 237340 271260 237346 271272
rect 256970 271260 256976 271272
rect 257028 271260 257034 271312
rect 259914 271260 259920 271312
rect 259972 271300 259978 271312
rect 270954 271300 270960 271312
rect 259972 271272 270960 271300
rect 259972 271260 259978 271272
rect 270954 271260 270960 271272
rect 271012 271260 271018 271312
rect 271506 271260 271512 271312
rect 271564 271300 271570 271312
rect 280890 271300 280896 271312
rect 271564 271272 280896 271300
rect 271564 271260 271570 271272
rect 280890 271260 280896 271272
rect 280948 271260 280954 271312
rect 315758 271260 315764 271312
rect 315816 271300 315822 271312
rect 319990 271300 319996 271312
rect 315816 271272 319996 271300
rect 315816 271260 315822 271272
rect 319990 271260 319996 271272
rect 320048 271260 320054 271312
rect 329742 271260 329748 271312
rect 329800 271300 329806 271312
rect 338942 271300 338948 271312
rect 329800 271272 338948 271300
rect 329800 271260 329806 271272
rect 338942 271260 338948 271272
rect 339000 271260 339006 271312
rect 341518 271260 341524 271312
rect 341576 271300 341582 271312
rect 348418 271300 348424 271312
rect 341576 271272 348424 271300
rect 341576 271260 341582 271272
rect 348418 271260 348424 271272
rect 348476 271260 348482 271312
rect 354582 271260 354588 271312
rect 354640 271300 354646 271312
rect 369854 271300 369860 271312
rect 354640 271272 369860 271300
rect 354640 271260 354646 271272
rect 369854 271260 369860 271272
rect 369912 271260 369918 271312
rect 372522 271260 372528 271312
rect 372580 271300 372586 271312
rect 382458 271300 382464 271312
rect 372580 271272 382464 271300
rect 372580 271260 372586 271272
rect 382458 271260 382464 271272
rect 382516 271260 382522 271312
rect 383378 271260 383384 271312
rect 383436 271300 383442 271312
rect 416958 271300 416964 271312
rect 383436 271272 416964 271300
rect 383436 271260 383442 271272
rect 416958 271260 416964 271272
rect 417016 271260 417022 271312
rect 421558 271260 421564 271312
rect 421616 271300 421622 271312
rect 437014 271300 437020 271312
rect 421616 271272 437020 271300
rect 421616 271260 421622 271272
rect 437014 271260 437020 271272
rect 437072 271260 437078 271312
rect 438136 271300 438164 271544
rect 442902 271532 442908 271584
rect 442960 271572 442966 271584
rect 500494 271572 500500 271584
rect 442960 271544 500500 271572
rect 442960 271532 442966 271544
rect 500494 271532 500500 271544
rect 500552 271532 500558 271584
rect 501966 271532 501972 271584
rect 502024 271572 502030 271584
rect 585594 271572 585600 271584
rect 502024 271544 585600 271572
rect 502024 271532 502030 271544
rect 585594 271532 585600 271544
rect 585652 271532 585658 271584
rect 585778 271532 585784 271584
rect 585836 271572 585842 271584
rect 608502 271572 608508 271584
rect 585836 271544 608508 271572
rect 585836 271532 585842 271544
rect 608502 271532 608508 271544
rect 608560 271532 608566 271584
rect 439958 271396 439964 271448
rect 440016 271436 440022 271448
rect 496998 271436 497004 271448
rect 440016 271408 497004 271436
rect 440016 271396 440022 271408
rect 496998 271396 497004 271408
rect 497056 271396 497062 271448
rect 504910 271396 504916 271448
rect 504968 271436 504974 271448
rect 589550 271436 589556 271448
rect 504968 271408 589556 271436
rect 504968 271396 504974 271408
rect 589550 271396 589556 271408
rect 589608 271396 589614 271448
rect 592678 271396 592684 271448
rect 592736 271436 592742 271448
rect 622670 271436 622676 271448
rect 592736 271408 622676 271436
rect 592736 271396 592742 271408
rect 622670 271396 622676 271408
rect 622728 271396 622734 271448
rect 438136 271272 441614 271300
rect 72970 271124 72976 271176
rect 73028 271164 73034 271176
rect 142338 271164 142344 271176
rect 73028 271136 142344 271164
rect 73028 271124 73034 271136
rect 142338 271124 142344 271136
rect 142396 271124 142402 271176
rect 143258 271124 143264 271176
rect 143316 271164 143322 271176
rect 144362 271164 144368 271176
rect 143316 271136 144368 271164
rect 143316 271124 143322 271136
rect 144362 271124 144368 271136
rect 144420 271124 144426 271176
rect 154298 271124 154304 271176
rect 154356 271164 154362 271176
rect 197906 271164 197912 271176
rect 154356 271136 197912 271164
rect 154356 271124 154362 271136
rect 197906 271124 197912 271136
rect 197964 271124 197970 271176
rect 198274 271124 198280 271176
rect 198332 271164 198338 271176
rect 229554 271164 229560 271176
rect 198332 271136 229560 271164
rect 198332 271124 198338 271136
rect 229554 271124 229560 271136
rect 229612 271124 229618 271176
rect 231394 271124 231400 271176
rect 231452 271164 231458 271176
rect 252738 271164 252744 271176
rect 231452 271136 252744 271164
rect 231452 271124 231458 271136
rect 252738 271124 252744 271136
rect 252796 271124 252802 271176
rect 263226 271124 263232 271176
rect 263284 271164 263290 271176
rect 275278 271164 275284 271176
rect 263284 271136 275284 271164
rect 263284 271124 263290 271136
rect 275278 271124 275284 271136
rect 275336 271124 275342 271176
rect 279786 271124 279792 271176
rect 279844 271164 279850 271176
rect 287146 271164 287152 271176
rect 279844 271136 287152 271164
rect 279844 271124 279850 271136
rect 287146 271124 287152 271136
rect 287204 271124 287210 271176
rect 325510 271124 325516 271176
rect 325568 271164 325574 271176
rect 334158 271164 334164 271176
rect 325568 271136 334164 271164
rect 325568 271124 325574 271136
rect 334158 271124 334164 271136
rect 334216 271124 334222 271176
rect 339310 271124 339316 271176
rect 339368 271164 339374 271176
rect 354306 271164 354312 271176
rect 339368 271136 354312 271164
rect 339368 271124 339374 271136
rect 354306 271124 354312 271136
rect 354364 271124 354370 271176
rect 362678 271124 362684 271176
rect 362736 271164 362742 271176
rect 387150 271164 387156 271176
rect 362736 271136 387156 271164
rect 362736 271124 362742 271136
rect 387150 271124 387156 271136
rect 387208 271124 387214 271176
rect 391750 271124 391756 271176
rect 391808 271164 391814 271176
rect 403434 271164 403440 271176
rect 391808 271136 403440 271164
rect 391808 271124 391814 271136
rect 403434 271124 403440 271136
rect 403492 271124 403498 271176
rect 404998 271124 405004 271176
rect 405056 271164 405062 271176
rect 441586 271164 441614 271272
rect 445662 271260 445668 271312
rect 445720 271300 445726 271312
rect 504450 271300 504456 271312
rect 445720 271272 504456 271300
rect 445720 271260 445726 271272
rect 504450 271260 504456 271272
rect 504508 271260 504514 271312
rect 509142 271260 509148 271312
rect 509200 271300 509206 271312
rect 596634 271300 596640 271312
rect 509200 271272 596640 271300
rect 509200 271260 509206 271272
rect 596634 271260 596640 271272
rect 596692 271260 596698 271312
rect 596818 271260 596824 271312
rect 596876 271300 596882 271312
rect 629754 271300 629760 271312
rect 596876 271272 629760 271300
rect 596876 271260 596882 271272
rect 629754 271260 629760 271272
rect 629812 271260 629818 271312
rect 448882 271164 448888 271176
rect 405056 271136 431954 271164
rect 441586 271136 448888 271164
rect 405056 271124 405062 271136
rect 83550 270988 83556 271040
rect 83608 271028 83614 271040
rect 123478 271028 123484 271040
rect 83608 271000 123484 271028
rect 83608 270988 83614 271000
rect 123478 270988 123484 271000
rect 123536 270988 123542 271040
rect 123754 270988 123760 271040
rect 123812 271028 123818 271040
rect 177482 271028 177488 271040
rect 123812 271000 177488 271028
rect 123812 270988 123818 271000
rect 177482 270988 177488 271000
rect 177540 270988 177546 271040
rect 431926 271028 431954 271136
rect 448882 271124 448888 271136
rect 448940 271124 448946 271176
rect 449802 271124 449808 271176
rect 449860 271164 449866 271176
rect 511534 271164 511540 271176
rect 449860 271136 511540 271164
rect 449860 271124 449866 271136
rect 511534 271124 511540 271136
rect 511592 271124 511598 271176
rect 511902 271124 511908 271176
rect 511960 271164 511966 271176
rect 600222 271164 600228 271176
rect 511960 271136 600228 271164
rect 511960 271124 511966 271136
rect 600222 271124 600228 271136
rect 600280 271124 600286 271176
rect 602338 271124 602344 271176
rect 602396 271164 602402 271176
rect 643922 271164 643928 271176
rect 602396 271136 643928 271164
rect 602396 271124 602402 271136
rect 643922 271124 643928 271136
rect 643980 271124 643986 271176
rect 434714 271028 434720 271040
rect 431926 271000 434720 271028
rect 434714 270988 434720 271000
rect 434772 270988 434778 271040
rect 434898 270988 434904 271040
rect 434956 271028 434962 271040
rect 486694 271028 486700 271040
rect 434956 271000 486700 271028
rect 434956 270988 434962 271000
rect 486694 270988 486700 271000
rect 486752 270988 486758 271040
rect 495250 270988 495256 271040
rect 495308 271028 495314 271040
rect 575382 271028 575388 271040
rect 495308 271000 575388 271028
rect 495308 270988 495314 271000
rect 575382 270988 575388 271000
rect 575440 270988 575446 271040
rect 576118 270988 576124 271040
rect 576176 271028 576182 271040
rect 594334 271028 594340 271040
rect 576176 271000 594340 271028
rect 576176 270988 576182 271000
rect 594334 270988 594340 271000
rect 594392 270988 594398 271040
rect 134426 270852 134432 270904
rect 134484 270892 134490 270904
rect 184934 270892 184940 270904
rect 134484 270864 184940 270892
rect 134484 270852 134490 270864
rect 184934 270852 184940 270864
rect 184992 270852 184998 270904
rect 418062 270852 418068 270904
rect 418120 270892 418126 270904
rect 456058 270892 456064 270904
rect 418120 270864 456064 270892
rect 418120 270852 418126 270864
rect 456058 270852 456064 270864
rect 456116 270852 456122 270904
rect 492582 270852 492588 270904
rect 492640 270892 492646 270904
rect 571794 270892 571800 270904
rect 492640 270864 571800 270892
rect 492640 270852 492646 270864
rect 571794 270852 571800 270864
rect 571852 270852 571858 270904
rect 113174 270716 113180 270768
rect 113232 270756 113238 270768
rect 154022 270756 154028 270768
rect 113232 270728 154028 270756
rect 113232 270716 113238 270728
rect 154022 270716 154028 270728
rect 154080 270716 154086 270768
rect 175826 270716 175832 270768
rect 175884 270756 175890 270768
rect 206278 270756 206284 270768
rect 175884 270728 206284 270756
rect 175884 270716 175890 270728
rect 206278 270716 206284 270728
rect 206336 270716 206342 270768
rect 404170 270716 404176 270768
rect 404228 270756 404234 270768
rect 445294 270756 445300 270768
rect 404228 270728 445300 270756
rect 404228 270716 404234 270728
rect 445294 270716 445300 270728
rect 445352 270716 445358 270768
rect 459186 270716 459192 270768
rect 459244 270756 459250 270768
rect 523034 270756 523040 270768
rect 459244 270728 523040 270756
rect 459244 270716 459250 270728
rect 523034 270716 523040 270728
rect 523092 270716 523098 270768
rect 526438 270716 526444 270768
rect 526496 270756 526502 270768
rect 576578 270756 576584 270768
rect 526496 270728 576584 270756
rect 526496 270716 526502 270728
rect 576578 270716 576584 270728
rect 576636 270716 576642 270768
rect 414474 270580 414480 270632
rect 414532 270620 414538 270632
rect 432966 270620 432972 270632
rect 414532 270592 432972 270620
rect 414532 270580 414538 270592
rect 432966 270580 432972 270592
rect 433024 270580 433030 270632
rect 433150 270580 433156 270632
rect 433208 270620 433214 270632
rect 434898 270620 434904 270632
rect 433208 270592 434904 270620
rect 433208 270580 433214 270592
rect 434898 270580 434904 270592
rect 434956 270580 434962 270632
rect 456058 270580 456064 270632
rect 456116 270620 456122 270632
rect 507946 270620 507952 270632
rect 456116 270592 507952 270620
rect 456116 270580 456122 270592
rect 507946 270580 507952 270592
rect 508004 270580 508010 270632
rect 509694 270580 509700 270632
rect 509752 270620 509758 270632
rect 510522 270620 510528 270632
rect 509752 270592 510528 270620
rect 509752 270580 509758 270592
rect 510522 270580 510528 270592
rect 510580 270580 510586 270632
rect 100662 270444 100668 270496
rect 100720 270484 100726 270496
rect 119798 270484 119804 270496
rect 100720 270456 119804 270484
rect 100720 270444 100726 270456
rect 119798 270444 119804 270456
rect 119856 270444 119862 270496
rect 122742 270444 122748 270496
rect 122800 270484 122806 270496
rect 176194 270484 176200 270496
rect 122800 270456 176200 270484
rect 122800 270444 122806 270456
rect 176194 270444 176200 270456
rect 176252 270444 176258 270496
rect 176930 270444 176936 270496
rect 176988 270484 176994 270496
rect 214742 270484 214748 270496
rect 176988 270456 214748 270484
rect 176988 270444 176994 270456
rect 214742 270444 214748 270456
rect 214800 270444 214806 270496
rect 219526 270444 219532 270496
rect 219584 270484 219590 270496
rect 219584 270456 229094 270484
rect 219584 270444 219590 270456
rect 78858 270308 78864 270360
rect 78916 270348 78922 270360
rect 132586 270348 132592 270360
rect 78916 270320 132592 270348
rect 78916 270308 78922 270320
rect 132586 270308 132592 270320
rect 132644 270308 132650 270360
rect 133782 270308 133788 270360
rect 133840 270348 133846 270360
rect 183646 270348 183652 270360
rect 133840 270320 183652 270348
rect 133840 270308 133846 270320
rect 183646 270308 183652 270320
rect 183704 270308 183710 270360
rect 186406 270308 186412 270360
rect 186464 270348 186470 270360
rect 201586 270348 201592 270360
rect 186464 270320 201592 270348
rect 186464 270308 186470 270320
rect 201586 270308 201592 270320
rect 201644 270308 201650 270360
rect 204162 270308 204168 270360
rect 204220 270348 204226 270360
rect 220262 270348 220268 270360
rect 204220 270320 220268 270348
rect 204220 270308 204226 270320
rect 220262 270308 220268 270320
rect 220320 270308 220326 270360
rect 229066 270348 229094 270456
rect 230382 270444 230388 270496
rect 230440 270484 230446 270496
rect 252094 270484 252100 270496
rect 230440 270456 252100 270484
rect 230440 270444 230446 270456
rect 252094 270444 252100 270456
rect 252152 270444 252158 270496
rect 275094 270444 275100 270496
rect 275152 270484 275158 270496
rect 276014 270484 276020 270496
rect 275152 270456 276020 270484
rect 275152 270444 275158 270456
rect 276014 270444 276020 270456
rect 276072 270444 276078 270496
rect 278682 270444 278688 270496
rect 278740 270484 278746 270496
rect 285950 270484 285956 270496
rect 278740 270456 285956 270484
rect 278740 270444 278746 270456
rect 285950 270444 285956 270456
rect 286008 270444 286014 270496
rect 291654 270444 291660 270496
rect 291712 270484 291718 270496
rect 295518 270484 295524 270496
rect 291712 270456 295524 270484
rect 291712 270444 291718 270456
rect 295518 270444 295524 270456
rect 295576 270444 295582 270496
rect 297910 270444 297916 270496
rect 297968 270484 297974 270496
rect 299566 270484 299572 270496
rect 297968 270456 299572 270484
rect 297968 270444 297974 270456
rect 299566 270444 299572 270456
rect 299624 270444 299630 270496
rect 299934 270444 299940 270496
rect 299992 270484 299998 270496
rect 300854 270484 300860 270496
rect 299992 270456 300860 270484
rect 299992 270444 299998 270456
rect 300854 270444 300860 270456
rect 300912 270444 300918 270496
rect 327074 270444 327080 270496
rect 327132 270484 327138 270496
rect 328454 270484 328460 270496
rect 327132 270456 328460 270484
rect 327132 270444 327138 270456
rect 328454 270444 328460 270456
rect 328512 270444 328518 270496
rect 360194 270484 360200 270496
rect 354646 270456 360200 270484
rect 244918 270348 244924 270360
rect 229066 270320 244924 270348
rect 244918 270308 244924 270320
rect 244976 270308 244982 270360
rect 335998 270308 336004 270360
rect 336056 270348 336062 270360
rect 347406 270348 347412 270360
rect 336056 270320 347412 270348
rect 336056 270308 336062 270320
rect 347406 270308 347412 270320
rect 347464 270308 347470 270360
rect 85482 270172 85488 270224
rect 85540 270212 85546 270224
rect 149422 270212 149428 270224
rect 85540 270184 149428 270212
rect 85540 270172 85546 270184
rect 149422 270172 149428 270184
rect 149480 270172 149486 270224
rect 153286 270172 153292 270224
rect 153344 270212 153350 270224
rect 169846 270212 169852 270224
rect 153344 270184 169852 270212
rect 153344 270172 153350 270184
rect 169846 270172 169852 270184
rect 169904 270172 169910 270224
rect 170030 270172 170036 270224
rect 170088 270212 170094 270224
rect 210142 270212 210148 270224
rect 170088 270184 210148 270212
rect 170088 270172 170094 270184
rect 210142 270172 210148 270184
rect 210200 270172 210206 270224
rect 211062 270172 211068 270224
rect 211120 270212 211126 270224
rect 237466 270212 237472 270224
rect 211120 270184 237472 270212
rect 211120 270172 211126 270184
rect 237466 270172 237472 270184
rect 237524 270172 237530 270224
rect 258534 270172 258540 270224
rect 258592 270212 258598 270224
rect 268010 270212 268016 270224
rect 258592 270184 268016 270212
rect 258592 270172 258598 270184
rect 268010 270172 268016 270184
rect 268068 270172 268074 270224
rect 321094 270172 321100 270224
rect 321152 270212 321158 270224
rect 327442 270212 327448 270224
rect 321152 270184 327448 270212
rect 321152 270172 321158 270184
rect 327442 270172 327448 270184
rect 327500 270172 327506 270224
rect 345934 270172 345940 270224
rect 345992 270212 345998 270224
rect 354646 270212 354674 270456
rect 360194 270444 360200 270456
rect 360252 270444 360258 270496
rect 377030 270444 377036 270496
rect 377088 270484 377094 270496
rect 387886 270484 387892 270496
rect 377088 270456 387892 270484
rect 377088 270444 377094 270456
rect 387886 270444 387892 270456
rect 387944 270444 387950 270496
rect 400582 270444 400588 270496
rect 400640 270484 400646 270496
rect 441614 270484 441620 270496
rect 400640 270456 441620 270484
rect 400640 270444 400646 270456
rect 441614 270444 441620 270456
rect 441672 270444 441678 270496
rect 453850 270444 453856 270496
rect 453908 270484 453914 270496
rect 516594 270484 516600 270496
rect 453908 270456 516600 270484
rect 453908 270444 453914 270456
rect 516594 270444 516600 270456
rect 516652 270444 516658 270496
rect 517698 270444 517704 270496
rect 517756 270484 517762 270496
rect 597554 270484 597560 270496
rect 517756 270456 597560 270484
rect 517756 270444 517762 270456
rect 597554 270444 597560 270456
rect 597612 270444 597618 270496
rect 359182 270308 359188 270360
rect 359240 270348 359246 270360
rect 382274 270348 382280 270360
rect 359240 270320 382280 270348
rect 359240 270308 359246 270320
rect 382274 270308 382280 270320
rect 382332 270308 382338 270360
rect 390370 270308 390376 270360
rect 390428 270348 390434 270360
rect 405734 270348 405740 270360
rect 390428 270320 405740 270348
rect 390428 270308 390434 270320
rect 405734 270308 405740 270320
rect 405792 270308 405798 270360
rect 407206 270308 407212 270360
rect 407264 270348 407270 270360
rect 451458 270348 451464 270360
rect 407264 270320 451464 270348
rect 407264 270308 407270 270320
rect 451458 270308 451464 270320
rect 451516 270308 451522 270360
rect 456426 270308 456432 270360
rect 456484 270348 456490 270360
rect 520274 270348 520280 270360
rect 456484 270320 520280 270348
rect 456484 270308 456490 270320
rect 520274 270308 520280 270320
rect 520332 270308 520338 270360
rect 523126 270308 523132 270360
rect 523184 270348 523190 270360
rect 605098 270348 605104 270360
rect 523184 270320 605104 270348
rect 523184 270308 523190 270320
rect 605098 270308 605104 270320
rect 605156 270308 605162 270360
rect 345992 270184 354674 270212
rect 345992 270172 345998 270184
rect 360194 270172 360200 270224
rect 360252 270212 360258 270224
rect 383654 270212 383660 270224
rect 360252 270184 383660 270212
rect 360252 270172 360258 270184
rect 383654 270172 383660 270184
rect 383712 270172 383718 270224
rect 388162 270172 388168 270224
rect 388220 270212 388226 270224
rect 410058 270212 410064 270224
rect 388220 270184 410064 270212
rect 388220 270172 388226 270184
rect 410058 270172 410064 270184
rect 410116 270172 410122 270224
rect 410794 270172 410800 270224
rect 410852 270212 410858 270224
rect 455414 270212 455420 270224
rect 410852 270184 455420 270212
rect 410852 270172 410858 270184
rect 455414 270172 455420 270184
rect 455472 270172 455478 270224
rect 461394 270172 461400 270224
rect 461452 270212 461458 270224
rect 527174 270212 527180 270224
rect 461452 270184 527180 270212
rect 461452 270172 461458 270184
rect 527174 270172 527180 270184
rect 527232 270172 527238 270224
rect 528094 270172 528100 270224
rect 528152 270212 528158 270224
rect 619174 270212 619180 270224
rect 528152 270184 619180 270212
rect 528152 270172 528158 270184
rect 619174 270172 619180 270184
rect 619232 270172 619238 270224
rect 309778 270104 309784 270156
rect 309836 270144 309842 270156
rect 311342 270144 311348 270156
rect 309836 270116 311348 270144
rect 309836 270104 309842 270116
rect 311342 270104 311348 270116
rect 311400 270104 311406 270156
rect 67542 270036 67548 270088
rect 67600 270076 67606 270088
rect 75914 270076 75920 270088
rect 67600 270048 75920 270076
rect 67600 270036 67606 270048
rect 75914 270036 75920 270048
rect 75972 270036 75978 270088
rect 80054 270036 80060 270088
rect 80112 270076 80118 270088
rect 146386 270076 146392 270088
rect 80112 270048 146392 270076
rect 80112 270036 80118 270048
rect 146386 270036 146392 270048
rect 146444 270036 146450 270088
rect 158622 270036 158628 270088
rect 158680 270076 158686 270088
rect 201034 270076 201040 270088
rect 158680 270048 201040 270076
rect 158680 270036 158686 270048
rect 201034 270036 201040 270048
rect 201092 270036 201098 270088
rect 202230 270036 202236 270088
rect 202288 270076 202294 270088
rect 230842 270076 230848 270088
rect 202288 270048 230848 270076
rect 202288 270036 202294 270048
rect 230842 270036 230848 270048
rect 230900 270036 230906 270088
rect 233694 270036 233700 270088
rect 233752 270076 233758 270088
rect 242710 270076 242716 270088
rect 233752 270048 242716 270076
rect 233752 270036 233758 270048
rect 242710 270036 242716 270048
rect 242768 270036 242774 270088
rect 245470 270036 245476 270088
rect 245528 270076 245534 270088
rect 263134 270076 263140 270088
rect 245528 270048 263140 270076
rect 245528 270036 245534 270048
rect 263134 270036 263140 270048
rect 263192 270036 263198 270088
rect 266814 270036 266820 270088
rect 266872 270076 266878 270088
rect 274634 270076 274640 270088
rect 266872 270048 274640 270076
rect 266872 270036 266878 270048
rect 274634 270036 274640 270048
rect 274692 270036 274698 270088
rect 316954 270036 316960 270088
rect 317012 270076 317018 270088
rect 321554 270076 321560 270088
rect 317012 270048 321560 270076
rect 317012 270036 317018 270048
rect 321554 270036 321560 270048
rect 321612 270036 321618 270088
rect 323578 270036 323584 270088
rect 323636 270076 323642 270088
rect 331214 270076 331220 270088
rect 323636 270048 331220 270076
rect 323636 270036 323642 270048
rect 331214 270036 331220 270048
rect 331272 270036 331278 270088
rect 346762 270036 346768 270088
rect 346820 270076 346826 270088
rect 364334 270076 364340 270088
rect 346820 270048 364340 270076
rect 346820 270036 346826 270048
rect 364334 270036 364340 270048
rect 364392 270036 364398 270088
rect 364978 270036 364984 270088
rect 365036 270076 365042 270088
rect 390554 270076 390560 270088
rect 365036 270048 390560 270076
rect 365036 270036 365042 270048
rect 390554 270036 390560 270048
rect 390612 270036 390618 270088
rect 409690 270036 409696 270088
rect 409748 270076 409754 270088
rect 454034 270076 454040 270088
rect 409748 270048 454040 270076
rect 409748 270036 409754 270048
rect 454034 270036 454040 270048
rect 454092 270036 454098 270088
rect 455046 270036 455052 270088
rect 455104 270076 455110 270088
rect 473354 270076 473360 270088
rect 455104 270048 473360 270076
rect 455104 270036 455110 270048
rect 473354 270036 473360 270048
rect 473412 270036 473418 270088
rect 525610 270036 525616 270088
rect 525668 270076 525674 270088
rect 619634 270076 619640 270088
rect 525668 270048 619640 270076
rect 525668 270036 525674 270048
rect 619634 270036 619640 270048
rect 619692 270036 619698 270088
rect 77202 269900 77208 269952
rect 77260 269940 77266 269952
rect 143902 269940 143908 269952
rect 77260 269912 143908 269940
rect 77260 269900 77266 269912
rect 143902 269900 143908 269912
rect 143960 269900 143966 269952
rect 144086 269900 144092 269952
rect 144144 269940 144150 269952
rect 190822 269940 190828 269952
rect 144144 269912 190828 269940
rect 144144 269900 144150 269912
rect 190822 269900 190828 269912
rect 190880 269900 190886 269952
rect 201770 269900 201776 269952
rect 201828 269940 201834 269952
rect 232498 269940 232504 269952
rect 201828 269912 232504 269940
rect 201828 269900 201834 269912
rect 232498 269900 232504 269912
rect 232556 269900 232562 269952
rect 234798 269900 234804 269952
rect 234856 269940 234862 269952
rect 255682 269940 255688 269952
rect 234856 269912 255688 269940
rect 234856 269900 234862 269912
rect 255682 269900 255688 269912
rect 255740 269900 255746 269952
rect 262030 269900 262036 269952
rect 262088 269940 262094 269952
rect 272518 269940 272524 269952
rect 262088 269912 272524 269940
rect 262088 269900 262094 269912
rect 272518 269900 272524 269912
rect 272576 269900 272582 269952
rect 273070 269900 273076 269952
rect 273128 269940 273134 269952
rect 282178 269940 282184 269952
rect 273128 269912 282184 269940
rect 273128 269900 273134 269912
rect 282178 269900 282184 269912
rect 282236 269900 282242 269952
rect 285766 269900 285772 269952
rect 285824 269940 285830 269952
rect 291286 269940 291292 269952
rect 285824 269912 291292 269940
rect 285824 269900 285830 269912
rect 291286 269900 291292 269912
rect 291344 269900 291350 269952
rect 329374 269900 329380 269952
rect 329432 269940 329438 269952
rect 339494 269940 339500 269952
rect 329432 269912 339500 269940
rect 329432 269900 329438 269912
rect 339494 269900 339500 269912
rect 339552 269900 339558 269952
rect 341794 269900 341800 269952
rect 341852 269940 341858 269952
rect 357434 269940 357440 269952
rect 341852 269912 357440 269940
rect 341852 269900 341858 269912
rect 357434 269900 357440 269912
rect 357492 269900 357498 269952
rect 364150 269900 364156 269952
rect 364208 269940 364214 269952
rect 389174 269940 389180 269952
rect 364208 269912 389180 269940
rect 364208 269900 364214 269912
rect 389174 269900 389180 269912
rect 389232 269900 389238 269952
rect 390186 269900 390192 269952
rect 390244 269940 390250 269952
rect 412634 269940 412640 269952
rect 390244 269912 412640 269940
rect 390244 269900 390250 269912
rect 412634 269900 412640 269912
rect 412692 269900 412698 269952
rect 414658 269900 414664 269952
rect 414716 269940 414722 269952
rect 460934 269940 460940 269952
rect 414716 269912 460940 269940
rect 414716 269900 414722 269912
rect 460934 269900 460940 269912
rect 460992 269900 460998 269952
rect 463510 269900 463516 269952
rect 463568 269940 463574 269952
rect 531314 269940 531320 269952
rect 463568 269912 531320 269940
rect 463568 269900 463574 269912
rect 531314 269900 531320 269912
rect 531372 269900 531378 269952
rect 531682 269900 531688 269952
rect 531740 269940 531746 269952
rect 627914 269940 627920 269952
rect 531740 269912 627920 269940
rect 531740 269900 531746 269912
rect 627914 269900 627920 269912
rect 627972 269900 627978 269952
rect 69382 269764 69388 269816
rect 69440 269804 69446 269816
rect 139762 269804 139768 269816
rect 69440 269776 139768 269804
rect 69440 269764 69446 269776
rect 139762 269764 139768 269776
rect 139820 269764 139826 269816
rect 140682 269764 140688 269816
rect 140740 269804 140746 269816
rect 188614 269804 188620 269816
rect 140740 269776 188620 269804
rect 140740 269764 140746 269776
rect 188614 269764 188620 269776
rect 188672 269764 188678 269816
rect 194594 269764 194600 269816
rect 194652 269804 194658 269816
rect 227254 269804 227260 269816
rect 194652 269776 227260 269804
rect 194652 269764 194658 269776
rect 227254 269764 227260 269776
rect 227312 269764 227318 269816
rect 249886 269804 249892 269816
rect 229066 269776 249892 269804
rect 119062 269628 119068 269680
rect 119120 269668 119126 269680
rect 173342 269668 173348 269680
rect 119120 269640 173348 269668
rect 119120 269628 119126 269640
rect 173342 269628 173348 269640
rect 173400 269628 173406 269680
rect 174354 269628 174360 269680
rect 174412 269668 174418 269680
rect 210970 269668 210976 269680
rect 174412 269640 210976 269668
rect 174412 269628 174418 269640
rect 210970 269628 210976 269640
rect 211028 269628 211034 269680
rect 226610 269628 226616 269680
rect 226668 269668 226674 269680
rect 229066 269668 229094 269776
rect 249886 269764 249892 269776
rect 249944 269764 249950 269816
rect 250254 269764 250260 269816
rect 250312 269804 250318 269816
rect 266446 269804 266452 269816
rect 250312 269776 266452 269804
rect 250312 269764 250318 269776
rect 266446 269764 266452 269776
rect 266504 269764 266510 269816
rect 268194 269764 268200 269816
rect 268252 269804 268258 269816
rect 278866 269804 278872 269816
rect 268252 269776 278872 269804
rect 268252 269764 268258 269776
rect 278866 269764 278872 269776
rect 278924 269764 278930 269816
rect 314470 269764 314476 269816
rect 314528 269804 314534 269816
rect 318978 269804 318984 269816
rect 314528 269776 318984 269804
rect 314528 269764 314534 269776
rect 318978 269764 318984 269776
rect 319036 269764 319042 269816
rect 326890 269764 326896 269816
rect 326948 269804 326954 269816
rect 335538 269804 335544 269816
rect 326948 269776 335544 269804
rect 326948 269764 326954 269776
rect 335538 269764 335544 269776
rect 335596 269764 335602 269816
rect 336918 269764 336924 269816
rect 336976 269804 336982 269816
rect 350534 269804 350540 269816
rect 336976 269776 350540 269804
rect 336976 269764 336982 269776
rect 350534 269764 350540 269776
rect 350592 269764 350598 269816
rect 351730 269764 351736 269816
rect 351788 269804 351794 269816
rect 371234 269804 371240 269816
rect 351788 269776 371240 269804
rect 351788 269764 351794 269776
rect 371234 269764 371240 269776
rect 371292 269764 371298 269816
rect 374914 269764 374920 269816
rect 374972 269804 374978 269816
rect 404354 269804 404360 269816
rect 374972 269776 404360 269804
rect 374972 269764 374978 269776
rect 404354 269764 404360 269776
rect 404412 269764 404418 269816
rect 412450 269764 412456 269816
rect 412508 269804 412514 269816
rect 458174 269804 458180 269816
rect 412508 269776 458180 269804
rect 412508 269764 412514 269776
rect 458174 269764 458180 269776
rect 458232 269764 458238 269816
rect 458542 269764 458548 269816
rect 458600 269804 458606 269816
rect 524414 269804 524420 269816
rect 458600 269776 524420 269804
rect 458600 269764 458606 269776
rect 524414 269764 524420 269776
rect 524472 269764 524478 269816
rect 535546 269764 535552 269816
rect 535604 269804 535610 269816
rect 633526 269804 633532 269816
rect 535604 269776 633532 269804
rect 535604 269764 535610 269776
rect 633526 269764 633532 269776
rect 633584 269764 633590 269816
rect 226668 269640 229094 269668
rect 226668 269628 226674 269640
rect 387426 269628 387432 269680
rect 387484 269668 387490 269680
rect 401686 269668 401692 269680
rect 387484 269640 401692 269668
rect 387484 269628 387490 269640
rect 401686 269628 401692 269640
rect 401744 269628 401750 269680
rect 401870 269628 401876 269680
rect 401928 269668 401934 269680
rect 419718 269668 419724 269680
rect 401928 269640 419724 269668
rect 401928 269628 401934 269640
rect 419718 269628 419724 269640
rect 419776 269628 419782 269680
rect 422110 269628 422116 269680
rect 422168 269668 422174 269680
rect 472158 269668 472164 269680
rect 422168 269640 472164 269668
rect 422168 269628 422174 269640
rect 472158 269628 472164 269640
rect 472216 269628 472222 269680
rect 474642 269628 474648 269680
rect 474700 269668 474706 269680
rect 546494 269668 546500 269680
rect 474700 269640 546500 269668
rect 474700 269628 474706 269640
rect 546494 269628 546500 269640
rect 546552 269628 546558 269680
rect 126882 269492 126888 269544
rect 126940 269532 126946 269544
rect 178678 269532 178684 269544
rect 126940 269504 178684 269532
rect 126940 269492 126946 269504
rect 178678 269492 178684 269504
rect 178736 269492 178742 269544
rect 183462 269492 183468 269544
rect 183520 269532 183526 269544
rect 204162 269532 204168 269544
rect 183520 269504 204168 269532
rect 183520 269492 183526 269504
rect 204162 269492 204168 269504
rect 204220 269492 204226 269544
rect 383654 269492 383660 269544
rect 383712 269532 383718 269544
rect 391934 269532 391940 269544
rect 383712 269504 391940 269532
rect 383712 269492 383718 269504
rect 391934 269492 391940 269504
rect 391992 269492 391998 269544
rect 392118 269492 392124 269544
rect 392176 269532 392182 269544
rect 409874 269532 409880 269544
rect 392176 269504 409880 269532
rect 392176 269492 392182 269504
rect 409874 269492 409880 269504
rect 409932 269492 409938 269544
rect 424594 269492 424600 269544
rect 424652 269532 424658 269544
rect 476114 269532 476120 269544
rect 424652 269504 476120 269532
rect 424652 269492 424658 269504
rect 476114 269492 476120 269504
rect 476172 269492 476178 269544
rect 476758 269492 476764 269544
rect 476816 269532 476822 269544
rect 549898 269532 549904 269544
rect 476816 269504 549904 269532
rect 476816 269492 476822 269504
rect 549898 269492 549904 269504
rect 549956 269492 549962 269544
rect 136082 269356 136088 269408
rect 136140 269396 136146 269408
rect 180886 269396 180892 269408
rect 136140 269368 180892 269396
rect 136140 269356 136146 269368
rect 180886 269356 180892 269368
rect 180944 269356 180950 269408
rect 419810 269356 419816 269408
rect 419868 269396 419874 269408
rect 465074 269396 465080 269408
rect 419868 269368 465080 269396
rect 419868 269356 419874 269368
rect 465074 269356 465080 269368
rect 465132 269356 465138 269408
rect 507854 269356 507860 269408
rect 507912 269396 507918 269408
rect 560294 269396 560300 269408
rect 507912 269368 560300 269396
rect 507912 269356 507918 269368
rect 560294 269356 560300 269368
rect 560352 269356 560358 269408
rect 251450 269220 251456 269272
rect 251508 269260 251514 269272
rect 258074 269260 258080 269272
rect 251508 269232 258080 269260
rect 251508 269220 251514 269232
rect 258074 269220 258080 269232
rect 258132 269220 258138 269272
rect 294046 269220 294052 269272
rect 294104 269260 294110 269272
rect 297082 269260 297088 269272
rect 294104 269232 297088 269260
rect 294104 269220 294110 269232
rect 297082 269220 297088 269232
rect 297140 269220 297146 269272
rect 441614 269220 441620 269272
rect 441672 269260 441678 269272
rect 462314 269260 462320 269272
rect 441672 269232 462320 269260
rect 441672 269220 441678 269232
rect 462314 269220 462320 269232
rect 462372 269220 462378 269272
rect 465994 269220 466000 269272
rect 466052 269260 466058 269272
rect 534166 269260 534172 269272
rect 466052 269232 534172 269260
rect 466052 269220 466058 269232
rect 534166 269220 534172 269232
rect 534224 269220 534230 269272
rect 146938 269152 146944 269204
rect 146996 269192 147002 269204
rect 153838 269192 153844 269204
rect 146996 269164 153844 269192
rect 146996 269152 147002 269164
rect 153838 269152 153844 269164
rect 153896 269152 153902 269204
rect 282822 269084 282828 269136
rect 282880 269124 282886 269136
rect 288802 269124 288808 269136
rect 282880 269096 288808 269124
rect 282880 269084 282886 269096
rect 288802 269084 288808 269096
rect 288860 269084 288866 269136
rect 295334 269084 295340 269136
rect 295392 269124 295398 269136
rect 297910 269124 297916 269136
rect 295392 269096 297916 269124
rect 295392 269084 295398 269096
rect 297910 269084 297916 269096
rect 297968 269084 297974 269136
rect 319438 269084 319444 269136
rect 319496 269124 319502 269136
rect 325694 269124 325700 269136
rect 319496 269096 325700 269124
rect 319496 269084 319502 269096
rect 325694 269084 325700 269096
rect 325752 269084 325758 269136
rect 331858 269084 331864 269136
rect 331916 269124 331922 269136
rect 338022 269124 338028 269136
rect 331916 269096 338028 269124
rect 331916 269084 331922 269096
rect 338022 269084 338028 269096
rect 338080 269084 338086 269136
rect 342254 269084 342260 269136
rect 342312 269124 342318 269136
rect 345106 269124 345112 269136
rect 342312 269096 345112 269124
rect 342312 269084 342318 269096
rect 345106 269084 345112 269096
rect 345164 269084 345170 269136
rect 115842 269016 115848 269068
rect 115900 269056 115906 269068
rect 171226 269056 171232 269068
rect 115900 269028 171232 269056
rect 115900 269016 115906 269028
rect 171226 269016 171232 269028
rect 171284 269016 171290 269068
rect 413002 269016 413008 269068
rect 413060 269056 413066 269068
rect 459738 269056 459744 269068
rect 413060 269028 459744 269056
rect 413060 269016 413066 269028
rect 459738 269016 459744 269028
rect 459796 269016 459802 269068
rect 469214 269016 469220 269068
rect 469272 269056 469278 269068
rect 495434 269056 495440 269068
rect 469272 269028 495440 269056
rect 469272 269016 469278 269028
rect 495434 269016 495440 269028
rect 495492 269016 495498 269068
rect 495802 269016 495808 269068
rect 495860 269056 495866 269068
rect 576854 269056 576860 269068
rect 495860 269028 576860 269056
rect 495860 269016 495866 269028
rect 576854 269016 576860 269028
rect 576912 269016 576918 269068
rect 108942 268880 108948 268932
rect 109000 268920 109006 268932
rect 166258 268920 166264 268932
rect 109000 268892 166264 268920
rect 109000 268880 109006 268892
rect 166258 268880 166264 268892
rect 166316 268880 166322 268932
rect 172422 268880 172428 268932
rect 172480 268920 172486 268932
rect 204346 268920 204352 268932
rect 172480 268892 204352 268920
rect 172480 268880 172486 268892
rect 204346 268880 204352 268892
rect 204404 268880 204410 268932
rect 208394 268880 208400 268932
rect 208452 268920 208458 268932
rect 214282 268920 214288 268932
rect 208452 268892 214288 268920
rect 208452 268880 208458 268892
rect 214282 268880 214288 268892
rect 214340 268880 214346 268932
rect 428734 268880 428740 268932
rect 428792 268920 428798 268932
rect 478966 268920 478972 268932
rect 428792 268892 478972 268920
rect 428792 268880 428798 268892
rect 478966 268880 478972 268892
rect 479024 268880 479030 268932
rect 498286 268880 498292 268932
rect 498344 268920 498350 268932
rect 580994 268920 581000 268932
rect 498344 268892 581000 268920
rect 498344 268880 498350 268892
rect 580994 268880 581000 268892
rect 581052 268880 581058 268932
rect 582190 268880 582196 268932
rect 582248 268920 582254 268932
rect 600406 268920 600412 268932
rect 582248 268892 600412 268920
rect 582248 268880 582254 268892
rect 600406 268880 600412 268892
rect 600464 268880 600470 268932
rect 99282 268744 99288 268796
rect 99340 268784 99346 268796
rect 99340 268756 103514 268784
rect 99340 268744 99346 268756
rect 91002 268608 91008 268660
rect 91060 268648 91066 268660
rect 99282 268648 99288 268660
rect 91060 268620 99288 268648
rect 91060 268608 91066 268620
rect 99282 268608 99288 268620
rect 99340 268608 99346 268660
rect 103486 268648 103514 268756
rect 110230 268744 110236 268796
rect 110288 268784 110294 268796
rect 167914 268784 167920 268796
rect 110288 268756 167920 268784
rect 110288 268744 110294 268756
rect 167914 268744 167920 268756
rect 167972 268744 167978 268796
rect 173802 268744 173808 268796
rect 173860 268784 173866 268796
rect 212626 268784 212632 268796
rect 173860 268756 212632 268784
rect 173860 268744 173866 268756
rect 212626 268744 212632 268756
rect 212684 268744 212690 268796
rect 215202 268744 215208 268796
rect 215260 268784 215266 268796
rect 223482 268784 223488 268796
rect 215260 268756 223488 268784
rect 215260 268744 215266 268756
rect 223482 268744 223488 268756
rect 223540 268744 223546 268796
rect 227714 268744 227720 268796
rect 227772 268784 227778 268796
rect 250714 268784 250720 268796
rect 227772 268756 250720 268784
rect 227772 268744 227778 268756
rect 250714 268744 250720 268756
rect 250772 268744 250778 268796
rect 372338 268744 372344 268796
rect 372396 268784 372402 268796
rect 397086 268784 397092 268796
rect 372396 268756 397092 268784
rect 372396 268744 372402 268756
rect 397086 268744 397092 268756
rect 397144 268744 397150 268796
rect 398742 268744 398748 268796
rect 398800 268784 398806 268796
rect 422294 268784 422300 268796
rect 398800 268756 422300 268784
rect 398800 268744 398806 268756
rect 422294 268744 422300 268756
rect 422352 268744 422358 268796
rect 433702 268744 433708 268796
rect 433760 268784 433766 268796
rect 488534 268784 488540 268796
rect 433760 268756 488540 268784
rect 433760 268744 433766 268756
rect 488534 268744 488540 268756
rect 488592 268744 488598 268796
rect 500678 268744 500684 268796
rect 500736 268784 500742 268796
rect 584122 268784 584128 268796
rect 500736 268756 584128 268784
rect 500736 268744 500742 268756
rect 584122 268744 584128 268756
rect 584180 268744 584186 268796
rect 160462 268648 160468 268660
rect 103486 268620 160468 268648
rect 160462 268608 160468 268620
rect 160520 268608 160526 268660
rect 168650 268608 168656 268660
rect 168708 268648 168714 268660
rect 208486 268648 208492 268660
rect 168708 268620 208492 268648
rect 168708 268608 168714 268620
rect 208486 268608 208492 268620
rect 208544 268608 208550 268660
rect 212258 268608 212264 268660
rect 212316 268648 212322 268660
rect 238294 268648 238300 268660
rect 212316 268620 238300 268648
rect 212316 268608 212322 268620
rect 238294 268608 238300 268620
rect 238352 268608 238358 268660
rect 256694 268608 256700 268660
rect 256752 268648 256758 268660
rect 263962 268648 263968 268660
rect 256752 268620 263968 268648
rect 256752 268608 256758 268620
rect 263962 268608 263968 268620
rect 264020 268608 264026 268660
rect 326062 268608 326068 268660
rect 326120 268648 326126 268660
rect 328270 268648 328276 268660
rect 326120 268620 328276 268648
rect 326120 268608 326126 268620
rect 328270 268608 328276 268620
rect 328328 268608 328334 268660
rect 355870 268608 355876 268660
rect 355928 268648 355934 268660
rect 367830 268648 367836 268660
rect 355928 268620 367836 268648
rect 355928 268608 355934 268620
rect 367830 268608 367836 268620
rect 367888 268608 367894 268660
rect 382366 268608 382372 268660
rect 382424 268648 382430 268660
rect 415394 268648 415400 268660
rect 382424 268620 415400 268648
rect 382424 268608 382430 268620
rect 415394 268608 415400 268620
rect 415452 268608 415458 268660
rect 416682 268608 416688 268660
rect 416740 268648 416746 268660
rect 433334 268648 433340 268660
rect 416740 268620 433340 268648
rect 416740 268608 416746 268620
rect 433334 268608 433340 268620
rect 433392 268608 433398 268660
rect 436186 268608 436192 268660
rect 436244 268648 436250 268660
rect 491846 268648 491852 268660
rect 436244 268620 491852 268648
rect 436244 268608 436250 268620
rect 491846 268608 491852 268620
rect 491904 268608 491910 268660
rect 498470 268648 498476 268660
rect 492048 268620 498476 268648
rect 92382 268472 92388 268524
rect 92440 268512 92446 268524
rect 155494 268512 155500 268524
rect 92440 268484 155500 268512
rect 92440 268472 92446 268484
rect 155494 268472 155500 268484
rect 155552 268472 155558 268524
rect 160002 268472 160008 268524
rect 160060 268512 160066 268524
rect 200390 268512 200396 268524
rect 160060 268484 200396 268512
rect 160060 268472 160066 268484
rect 200390 268472 200396 268484
rect 200448 268472 200454 268524
rect 208210 268472 208216 268524
rect 208268 268512 208274 268524
rect 236638 268512 236644 268524
rect 208268 268484 236644 268512
rect 208268 268472 208274 268484
rect 236638 268472 236644 268484
rect 236696 268472 236702 268524
rect 241422 268472 241428 268524
rect 241480 268512 241486 268524
rect 256694 268512 256700 268524
rect 241480 268484 256700 268512
rect 241480 268472 241486 268484
rect 256694 268472 256700 268484
rect 256752 268472 256758 268524
rect 269114 268472 269120 268524
rect 269172 268512 269178 268524
rect 279694 268512 279700 268524
rect 269172 268484 279700 268512
rect 269172 268472 269178 268484
rect 279694 268472 279700 268484
rect 279752 268472 279758 268524
rect 343358 268472 343364 268524
rect 343416 268512 343422 268524
rect 357250 268512 357256 268524
rect 343416 268484 357256 268512
rect 343416 268472 343422 268484
rect 357250 268472 357256 268484
rect 357308 268472 357314 268524
rect 357526 268472 357532 268524
rect 357584 268512 357590 268524
rect 379514 268512 379520 268524
rect 357584 268484 379520 268512
rect 357584 268472 357590 268484
rect 379514 268472 379520 268484
rect 379572 268472 379578 268524
rect 393130 268472 393136 268524
rect 393188 268512 393194 268524
rect 430574 268512 430580 268524
rect 393188 268484 430580 268512
rect 393188 268472 393194 268484
rect 430574 268472 430580 268484
rect 430632 268472 430638 268524
rect 441154 268472 441160 268524
rect 441212 268512 441218 268524
rect 492048 268512 492076 268620
rect 498470 268608 498476 268620
rect 498528 268608 498534 268660
rect 503254 268608 503260 268660
rect 503312 268648 503318 268660
rect 587894 268648 587900 268660
rect 503312 268620 587900 268648
rect 503312 268608 503318 268620
rect 587894 268608 587900 268620
rect 587952 268608 587958 268660
rect 441212 268484 492076 268512
rect 441212 268472 441218 268484
rect 492214 268472 492220 268524
rect 492272 268512 492278 268524
rect 492272 268484 509234 268512
rect 492272 268472 492278 268484
rect 87138 268336 87144 268388
rect 87196 268376 87202 268388
rect 152182 268376 152188 268388
rect 87196 268348 152188 268376
rect 87196 268336 87202 268348
rect 152182 268336 152188 268348
rect 152240 268336 152246 268388
rect 152734 268336 152740 268388
rect 152792 268376 152798 268388
rect 196066 268376 196072 268388
rect 152792 268348 196072 268376
rect 152792 268336 152798 268348
rect 196066 268336 196072 268348
rect 196124 268336 196130 268388
rect 200574 268336 200580 268388
rect 200632 268376 200638 268388
rect 231670 268376 231676 268388
rect 200632 268348 231676 268376
rect 200632 268336 200638 268348
rect 231670 268336 231676 268348
rect 231728 268336 231734 268388
rect 238662 268336 238668 268388
rect 238720 268376 238726 268388
rect 256142 268376 256148 268388
rect 238720 268348 256148 268376
rect 238720 268336 238726 268348
rect 256142 268336 256148 268348
rect 256200 268336 256206 268388
rect 256510 268336 256516 268388
rect 256568 268376 256574 268388
rect 270586 268376 270592 268388
rect 256568 268348 270592 268376
rect 256568 268336 256574 268348
rect 270586 268336 270592 268348
rect 270644 268336 270650 268388
rect 327718 268336 327724 268388
rect 327776 268376 327782 268388
rect 336734 268376 336740 268388
rect 327776 268348 336740 268376
rect 327776 268336 327782 268348
rect 336734 268336 336740 268348
rect 336792 268336 336798 268388
rect 337654 268336 337660 268388
rect 337712 268376 337718 268388
rect 352098 268376 352104 268388
rect 337712 268348 352104 268376
rect 337712 268336 337718 268348
rect 352098 268336 352104 268348
rect 352156 268336 352162 268388
rect 352558 268336 352564 268388
rect 352616 268376 352622 268388
rect 368842 268376 368848 268388
rect 352616 268348 368848 268376
rect 352616 268336 352622 268348
rect 368842 268336 368848 268348
rect 368900 268336 368906 268388
rect 369946 268336 369952 268388
rect 370004 268376 370010 268388
rect 397454 268376 397460 268388
rect 370004 268348 397460 268376
rect 370004 268336 370010 268348
rect 397454 268336 397460 268348
rect 397512 268336 397518 268388
rect 399754 268336 399760 268388
rect 399812 268376 399818 268388
rect 440234 268376 440240 268388
rect 399812 268348 440240 268376
rect 399812 268336 399818 268348
rect 440234 268336 440240 268348
rect 440292 268336 440298 268388
rect 443638 268336 443644 268388
rect 443696 268376 443702 268388
rect 502334 268376 502340 268388
rect 443696 268348 502340 268376
rect 443696 268336 443702 268348
rect 502334 268336 502340 268348
rect 502392 268336 502398 268388
rect 509206 268376 509234 268484
rect 510706 268472 510712 268524
rect 510764 268512 510770 268524
rect 598934 268512 598940 268524
rect 510764 268484 598940 268512
rect 510764 268472 510770 268484
rect 598934 268472 598940 268484
rect 598992 268472 598998 268524
rect 517882 268376 517888 268388
rect 509206 268348 517888 268376
rect 517882 268336 517888 268348
rect 517940 268336 517946 268388
rect 534718 268336 534724 268388
rect 534776 268376 534782 268388
rect 535730 268376 535736 268388
rect 534776 268348 535736 268376
rect 534776 268336 534782 268348
rect 535730 268336 535736 268348
rect 535788 268336 535794 268388
rect 536374 268336 536380 268388
rect 536432 268376 536438 268388
rect 634814 268376 634820 268388
rect 536432 268348 634820 268376
rect 536432 268336 536438 268348
rect 634814 268336 634820 268348
rect 634872 268336 634878 268388
rect 118602 268200 118608 268252
rect 118660 268240 118666 268252
rect 174538 268240 174544 268252
rect 118660 268212 174544 268240
rect 118660 268200 118666 268212
rect 174538 268200 174544 268212
rect 174596 268200 174602 268252
rect 429562 268200 429568 268252
rect 429620 268240 429626 268252
rect 469398 268240 469404 268252
rect 429620 268212 469404 268240
rect 429620 268200 429626 268212
rect 469398 268200 469404 268212
rect 469456 268200 469462 268252
rect 492122 268240 492128 268252
rect 470566 268212 492128 268240
rect 137002 268064 137008 268116
rect 137060 268104 137066 268116
rect 183002 268104 183008 268116
rect 137060 268076 183008 268104
rect 137060 268064 137066 268076
rect 183002 268064 183008 268076
rect 183060 268064 183066 268116
rect 422294 268064 422300 268116
rect 422352 268104 422358 268116
rect 443270 268104 443276 268116
rect 422352 268076 443276 268104
rect 422352 268064 422358 268076
rect 443270 268064 443276 268076
rect 443328 268064 443334 268116
rect 459554 268064 459560 268116
rect 459612 268104 459618 268116
rect 470566 268104 470594 268212
rect 492122 268200 492128 268212
rect 492180 268200 492186 268252
rect 492306 268200 492312 268252
rect 492364 268240 492370 268252
rect 569954 268240 569960 268252
rect 492364 268212 569960 268240
rect 492364 268200 492370 268212
rect 569954 268200 569960 268212
rect 570012 268200 570018 268252
rect 567378 268104 567384 268116
rect 459612 268076 470594 268104
rect 489886 268076 567384 268104
rect 459612 268064 459618 268076
rect 489178 267928 489184 267980
rect 489236 267968 489242 267980
rect 489886 267968 489914 268076
rect 567378 268064 567384 268076
rect 567436 268064 567442 268116
rect 489236 267940 489914 267968
rect 489236 267928 489242 267940
rect 490834 267928 490840 267980
rect 490892 267968 490898 267980
rect 492306 267968 492312 267980
rect 490892 267940 492312 267968
rect 490892 267928 490898 267940
rect 492306 267928 492312 267940
rect 492364 267928 492370 267980
rect 493318 267928 493324 267980
rect 493376 267968 493382 267980
rect 551554 267968 551560 267980
rect 493376 267940 551560 267968
rect 493376 267928 493382 267940
rect 551554 267928 551560 267940
rect 551612 267928 551618 267980
rect 193122 267832 193128 267844
rect 192312 267804 193128 267832
rect 132402 267656 132408 267708
rect 132460 267696 132466 267708
rect 132460 267668 180794 267696
rect 132460 267656 132466 267668
rect 99282 267520 99288 267572
rect 99340 267560 99346 267572
rect 154666 267560 154672 267572
rect 99340 267532 154672 267560
rect 99340 267520 99346 267532
rect 154666 267520 154672 267532
rect 154724 267520 154730 267572
rect 160738 267520 160744 267572
rect 160796 267560 160802 267572
rect 164602 267560 164608 267572
rect 160796 267532 164608 267560
rect 160796 267520 160802 267532
rect 164602 267520 164608 267532
rect 164660 267520 164666 267572
rect 166442 267520 166448 267572
rect 166500 267560 166506 267572
rect 172882 267560 172888 267572
rect 166500 267532 172888 267560
rect 166500 267520 166506 267532
rect 172882 267520 172888 267532
rect 172940 267520 172946 267572
rect 180766 267560 180794 267668
rect 184198 267656 184204 267708
rect 184256 267696 184262 267708
rect 192312 267696 192340 267804
rect 193122 267792 193128 267804
rect 193180 267792 193186 267844
rect 448606 267792 448612 267844
rect 448664 267832 448670 267844
rect 506474 267832 506480 267844
rect 448664 267804 506480 267832
rect 448664 267792 448670 267804
rect 506474 267792 506480 267804
rect 506532 267792 506538 267844
rect 184256 267668 192340 267696
rect 184256 267656 184262 267668
rect 193122 267656 193128 267708
rect 193180 267656 193186 267708
rect 204162 267656 204168 267708
rect 204220 267696 204226 267708
rect 218422 267696 218428 267708
rect 204220 267668 218428 267696
rect 204220 267656 204226 267668
rect 218422 267656 218428 267668
rect 218480 267656 218486 267708
rect 218790 267656 218796 267708
rect 218848 267696 218854 267708
rect 222562 267696 222568 267708
rect 218848 267668 222568 267696
rect 218848 267656 218854 267668
rect 222562 267656 222568 267668
rect 222620 267656 222626 267708
rect 377766 267656 377772 267708
rect 377824 267696 377830 267708
rect 385678 267696 385684 267708
rect 377824 267668 385684 267696
rect 377824 267656 377830 267668
rect 385678 267656 385684 267668
rect 385736 267656 385742 267708
rect 387242 267656 387248 267708
rect 387300 267696 387306 267708
rect 398742 267696 398748 267708
rect 387300 267668 398748 267696
rect 387300 267656 387306 267668
rect 398742 267656 398748 267668
rect 398800 267656 398806 267708
rect 404722 267656 404728 267708
rect 404780 267696 404786 267708
rect 429838 267696 429844 267708
rect 404780 267668 429844 267696
rect 404780 267656 404786 267668
rect 429838 267656 429844 267668
rect 429896 267656 429902 267708
rect 436738 267656 436744 267708
rect 436796 267696 436802 267708
rect 441614 267696 441620 267708
rect 436796 267668 441620 267696
rect 436796 267656 436802 267668
rect 441614 267656 441620 267668
rect 441672 267656 441678 267708
rect 442718 267656 442724 267708
rect 442776 267696 442782 267708
rect 483658 267696 483664 267708
rect 442776 267668 483664 267696
rect 442776 267656 442782 267668
rect 483658 267656 483664 267668
rect 483716 267656 483722 267708
rect 483842 267656 483848 267708
rect 483900 267696 483906 267708
rect 483900 267668 489914 267696
rect 483900 267656 483906 267668
rect 184474 267560 184480 267572
rect 180766 267532 184480 267560
rect 184474 267520 184480 267532
rect 184532 267520 184538 267572
rect 186958 267520 186964 267572
rect 187016 267560 187022 267572
rect 193140 267560 193168 267656
rect 216766 267560 216772 267572
rect 187016 267532 193076 267560
rect 193140 267532 216772 267560
rect 187016 267520 187022 267532
rect 107654 267384 107660 267436
rect 107712 267424 107718 267436
rect 167086 267424 167092 267436
rect 107712 267396 167092 267424
rect 107712 267384 107718 267396
rect 167086 267384 167092 267396
rect 167144 267384 167150 267436
rect 167638 267384 167644 267436
rect 167696 267424 167702 267436
rect 186958 267424 186964 267436
rect 167696 267396 186964 267424
rect 167696 267384 167702 267396
rect 186958 267384 186964 267396
rect 187016 267384 187022 267436
rect 189902 267384 189908 267436
rect 189960 267424 189966 267436
rect 192754 267424 192760 267436
rect 189960 267396 192760 267424
rect 189960 267384 189966 267396
rect 192754 267384 192760 267396
rect 192812 267384 192818 267436
rect 193048 267424 193076 267532
rect 216766 267520 216772 267532
rect 216824 267520 216830 267572
rect 217410 267520 217416 267572
rect 217468 267560 217474 267572
rect 223022 267560 223028 267572
rect 217468 267532 223028 267560
rect 217468 267520 217474 267532
rect 223022 267520 223028 267532
rect 223080 267520 223086 267572
rect 224218 267520 224224 267572
rect 224276 267560 224282 267572
rect 229186 267560 229192 267572
rect 224276 267532 229192 267560
rect 224276 267520 224282 267532
rect 229186 267520 229192 267532
rect 229244 267520 229250 267572
rect 373258 267520 373264 267572
rect 373316 267560 373322 267572
rect 387426 267560 387432 267572
rect 373316 267532 387432 267560
rect 373316 267520 373322 267532
rect 387426 267520 387432 267532
rect 387484 267520 387490 267572
rect 402238 267520 402244 267572
rect 402296 267560 402302 267572
rect 422294 267560 422300 267572
rect 402296 267532 422300 267560
rect 402296 267520 402302 267532
rect 422294 267520 422300 267532
rect 422352 267520 422358 267572
rect 430390 267520 430396 267572
rect 430448 267560 430454 267572
rect 457438 267560 457444 267572
rect 430448 267532 457444 267560
rect 430448 267520 430454 267532
rect 457438 267520 457444 267532
rect 457496 267520 457502 267572
rect 462682 267520 462688 267572
rect 462740 267560 462746 267572
rect 468938 267560 468944 267572
rect 462740 267532 468944 267560
rect 462740 267520 462746 267532
rect 468938 267520 468944 267532
rect 468996 267520 469002 267572
rect 475102 267520 475108 267572
rect 475160 267560 475166 267572
rect 479702 267560 479708 267572
rect 475160 267532 479708 267560
rect 475160 267520 475166 267532
rect 479702 267520 479708 267532
rect 479760 267520 479766 267572
rect 484026 267520 484032 267572
rect 484084 267560 484090 267572
rect 487798 267560 487804 267572
rect 484084 267532 487804 267560
rect 484084 267520 484090 267532
rect 487798 267520 487804 267532
rect 487856 267520 487862 267572
rect 489886 267560 489914 267668
rect 490006 267656 490012 267708
rect 490064 267696 490070 267708
rect 497274 267696 497280 267708
rect 490064 267668 497280 267696
rect 490064 267656 490070 267668
rect 497274 267656 497280 267668
rect 497332 267656 497338 267708
rect 499666 267656 499672 267708
rect 499724 267696 499730 267708
rect 526438 267696 526444 267708
rect 499724 267668 526444 267696
rect 499724 267656 499730 267668
rect 526438 267656 526444 267668
rect 526496 267656 526502 267708
rect 527266 267656 527272 267708
rect 527324 267696 527330 267708
rect 592678 267696 592684 267708
rect 527324 267668 592684 267696
rect 527324 267656 527330 267668
rect 592678 267656 592684 267668
rect 592736 267656 592742 267708
rect 507854 267560 507860 267572
rect 489886 267532 507860 267560
rect 507854 267520 507860 267532
rect 507912 267520 507918 267572
rect 508222 267520 508228 267572
rect 508280 267560 508286 267572
rect 522390 267560 522396 267572
rect 508280 267532 522396 267560
rect 508280 267520 508286 267532
rect 522390 267520 522396 267532
rect 522448 267520 522454 267572
rect 523678 267520 523684 267572
rect 523736 267560 523742 267572
rect 530670 267560 530676 267572
rect 523736 267532 530676 267560
rect 523736 267520 523742 267532
rect 530670 267520 530676 267532
rect 530728 267520 530734 267572
rect 532234 267520 532240 267572
rect 532292 267560 532298 267572
rect 596818 267560 596824 267572
rect 532292 267532 596824 267560
rect 532292 267520 532298 267532
rect 596818 267520 596824 267532
rect 596876 267520 596882 267572
rect 221734 267424 221740 267436
rect 193048 267396 221740 267424
rect 221734 267384 221740 267396
rect 221792 267384 221798 267436
rect 232682 267384 232688 267436
rect 232740 267424 232746 267436
rect 239122 267424 239128 267436
rect 232740 267396 239128 267424
rect 232740 267384 232746 267396
rect 239122 267384 239128 267396
rect 239180 267384 239186 267436
rect 261478 267384 261484 267436
rect 261536 267424 261542 267436
rect 268930 267424 268936 267436
rect 261536 267396 268936 267424
rect 261536 267384 261542 267396
rect 268930 267384 268936 267396
rect 268988 267384 268994 267436
rect 340966 267384 340972 267436
rect 341024 267424 341030 267436
rect 347038 267424 347044 267436
rect 341024 267396 347044 267424
rect 341024 267384 341030 267396
rect 347038 267384 347044 267396
rect 347096 267384 347102 267436
rect 350902 267384 350908 267436
rect 350960 267424 350966 267436
rect 359458 267424 359464 267436
rect 350960 267396 359464 267424
rect 350960 267384 350966 267396
rect 359458 267384 359464 267396
rect 359516 267384 359522 267436
rect 361114 267384 361120 267436
rect 361172 267424 361178 267436
rect 373074 267424 373080 267436
rect 361172 267396 373080 267424
rect 361172 267384 361178 267396
rect 373074 267384 373080 267396
rect 373132 267384 373138 267436
rect 375742 267384 375748 267436
rect 375800 267424 375806 267436
rect 390370 267424 390376 267436
rect 375800 267396 390376 267424
rect 375800 267384 375806 267396
rect 390370 267384 390376 267396
rect 390428 267384 390434 267436
rect 390646 267384 390652 267436
rect 390704 267424 390710 267436
rect 395522 267424 395528 267436
rect 390704 267396 395528 267424
rect 390704 267384 390710 267396
rect 395522 267384 395528 267396
rect 395580 267384 395586 267436
rect 397086 267384 397092 267436
rect 397144 267424 397150 267436
rect 421558 267424 421564 267436
rect 397144 267396 421564 267424
rect 397144 267384 397150 267396
rect 421558 267384 421564 267396
rect 421616 267384 421622 267436
rect 436554 267384 436560 267436
rect 436612 267424 436618 267436
rect 445018 267424 445024 267436
rect 436612 267396 445024 267424
rect 436612 267384 436618 267396
rect 445018 267384 445024 267396
rect 445076 267384 445082 267436
rect 450262 267384 450268 267436
rect 450320 267424 450326 267436
rect 505830 267424 505836 267436
rect 450320 267396 505836 267424
rect 450320 267384 450326 267396
rect 505830 267384 505836 267396
rect 505888 267384 505894 267436
rect 507394 267384 507400 267436
rect 507452 267424 507458 267436
rect 576118 267424 576124 267436
rect 507452 267396 576124 267424
rect 507452 267384 507458 267396
rect 576118 267384 576124 267396
rect 576176 267384 576182 267436
rect 95878 267248 95884 267300
rect 95936 267288 95942 267300
rect 157150 267288 157156 267300
rect 95936 267260 157156 267288
rect 95936 267248 95942 267260
rect 157150 267248 157156 267260
rect 157208 267248 157214 267300
rect 170398 267248 170404 267300
rect 170456 267288 170462 267300
rect 170456 267260 206140 267288
rect 170456 267248 170462 267260
rect 86218 267112 86224 267164
rect 86276 267152 86282 267164
rect 148042 267152 148048 267164
rect 86276 267124 148048 267152
rect 86276 267112 86282 267124
rect 148042 267112 148048 267124
rect 148100 267112 148106 267164
rect 149698 267112 149704 267164
rect 149756 267152 149762 267164
rect 194410 267152 194416 267164
rect 149756 267124 194416 267152
rect 149756 267112 149762 267124
rect 194410 267112 194416 267124
rect 194468 267112 194474 267164
rect 198182 267112 198188 267164
rect 198240 267152 198246 267164
rect 200206 267152 200212 267164
rect 198240 267124 200212 267152
rect 198240 267112 198246 267124
rect 200206 267112 200212 267124
rect 200264 267112 200270 267164
rect 206112 267152 206140 267260
rect 206278 267248 206284 267300
rect 206336 267288 206342 267300
rect 213454 267288 213460 267300
rect 206336 267260 213460 267288
rect 206336 267248 206342 267260
rect 213454 267248 213460 267260
rect 213512 267248 213518 267300
rect 215938 267248 215944 267300
rect 215996 267288 216002 267300
rect 220078 267288 220084 267300
rect 215996 267260 220084 267288
rect 215996 267248 216002 267260
rect 220078 267248 220084 267260
rect 220136 267248 220142 267300
rect 220262 267248 220268 267300
rect 220320 267288 220326 267300
rect 234154 267288 234160 267300
rect 220320 267260 234160 267288
rect 220320 267248 220326 267260
rect 234154 267248 234160 267260
rect 234212 267248 234218 267300
rect 236822 267248 236828 267300
rect 236880 267288 236886 267300
rect 251542 267288 251548 267300
rect 236880 267260 251548 267288
rect 236880 267248 236886 267260
rect 251542 267248 251548 267260
rect 251600 267248 251606 267300
rect 286318 267248 286324 267300
rect 286376 267288 286382 267300
rect 287974 267288 287980 267300
rect 286376 267260 287980 267288
rect 286376 267248 286382 267260
rect 287974 267248 287980 267260
rect 288032 267248 288038 267300
rect 313642 267248 313648 267300
rect 313700 267288 313706 267300
rect 317414 267288 317420 267300
rect 313700 267260 317420 267288
rect 313700 267248 313706 267260
rect 317414 267248 317420 267260
rect 317472 267248 317478 267300
rect 335170 267248 335176 267300
rect 335228 267288 335234 267300
rect 341518 267288 341524 267300
rect 335228 267260 341524 267288
rect 335228 267248 335234 267260
rect 341518 267248 341524 267260
rect 341576 267248 341582 267300
rect 363322 267248 363328 267300
rect 363380 267288 363386 267300
rect 377030 267288 377036 267300
rect 363380 267260 377036 267288
rect 363380 267248 363386 267260
rect 377030 267248 377036 267260
rect 377088 267248 377094 267300
rect 394786 267248 394792 267300
rect 394844 267288 394850 267300
rect 416682 267288 416688 267300
rect 394844 267260 416688 267288
rect 394844 267248 394850 267260
rect 416682 267248 416688 267260
rect 416740 267248 416746 267300
rect 419626 267248 419632 267300
rect 419684 267288 419690 267300
rect 446582 267288 446588 267300
rect 419684 267260 446588 267288
rect 419684 267248 419690 267260
rect 446582 267248 446588 267260
rect 446640 267248 446646 267300
rect 455230 267248 455236 267300
rect 455288 267288 455294 267300
rect 507854 267288 507860 267300
rect 455288 267260 507860 267288
rect 455288 267248 455294 267260
rect 507854 267248 507860 267260
rect 507912 267248 507918 267300
rect 509878 267248 509884 267300
rect 509936 267288 509942 267300
rect 517698 267288 517704 267300
rect 509936 267260 517704 267288
rect 509936 267248 509942 267260
rect 517698 267248 517704 267260
rect 517756 267248 517762 267300
rect 582190 267288 582196 267300
rect 518866 267260 582196 267288
rect 206830 267152 206836 267164
rect 206112 267124 206836 267152
rect 206830 267112 206836 267124
rect 206888 267112 206894 267164
rect 207014 267112 207020 267164
rect 207072 267152 207078 267164
rect 220906 267152 220912 267164
rect 207072 267124 220912 267152
rect 207072 267112 207078 267124
rect 220906 267112 220912 267124
rect 220964 267112 220970 267164
rect 223482 267112 223488 267164
rect 223540 267152 223546 267164
rect 241606 267152 241612 267164
rect 223540 267124 241612 267152
rect 223540 267112 223546 267124
rect 241606 267112 241612 267124
rect 241664 267112 241670 267164
rect 242710 267112 242716 267164
rect 242768 267152 242774 267164
rect 254854 267152 254860 267164
rect 242768 267124 254860 267152
rect 242768 267112 242774 267124
rect 254854 267112 254860 267124
rect 254912 267112 254918 267164
rect 266998 267112 267004 267164
rect 267056 267152 267062 267164
rect 273070 267152 273076 267164
rect 267056 267124 273076 267152
rect 267056 267112 267062 267124
rect 273070 267112 273076 267124
rect 273128 267112 273134 267164
rect 276014 267112 276020 267164
rect 276072 267152 276078 267164
rect 283834 267152 283840 267164
rect 276072 267124 283840 267152
rect 276072 267112 276078 267124
rect 283834 267112 283840 267124
rect 283892 267112 283898 267164
rect 324406 267112 324412 267164
rect 324464 267152 324470 267164
rect 330478 267152 330484 267164
rect 324464 267124 330484 267152
rect 324464 267112 324470 267124
rect 330478 267112 330484 267124
rect 330536 267112 330542 267164
rect 334342 267112 334348 267164
rect 334400 267152 334406 267164
rect 344278 267152 344284 267164
rect 334400 267124 344284 267152
rect 334400 267112 334406 267124
rect 344278 267112 344284 267124
rect 344336 267112 344342 267164
rect 353386 267112 353392 267164
rect 353444 267152 353450 267164
rect 363598 267152 363604 267164
rect 353444 267124 363604 267152
rect 353444 267112 353450 267124
rect 363598 267112 363604 267124
rect 363656 267112 363662 267164
rect 365806 267112 365812 267164
rect 365864 267152 365870 267164
rect 365864 267124 378824 267152
rect 365864 267112 365870 267124
rect 73798 266976 73804 267028
rect 73856 267016 73862 267028
rect 141418 267016 141424 267028
rect 73856 266988 141424 267016
rect 73856 266976 73862 266988
rect 141418 266976 141424 266988
rect 141476 266976 141482 267028
rect 146938 266976 146944 267028
rect 146996 267016 147002 267028
rect 189442 267016 189448 267028
rect 146996 266988 189448 267016
rect 146996 266976 147002 266988
rect 189442 266976 189448 266988
rect 189500 266976 189506 267028
rect 191006 266976 191012 267028
rect 191064 267016 191070 267028
rect 211798 267016 211804 267028
rect 191064 266988 211804 267016
rect 191064 266976 191070 266988
rect 211798 266976 211804 266988
rect 211856 266976 211862 267028
rect 222010 266976 222016 267028
rect 222068 267016 222074 267028
rect 246574 267016 246580 267028
rect 222068 266988 246580 267016
rect 222068 266976 222074 266988
rect 246574 266976 246580 266988
rect 246632 266976 246638 267028
rect 249058 266976 249064 267028
rect 249116 267016 249122 267028
rect 261478 267016 261484 267028
rect 249116 266988 261484 267016
rect 249116 266976 249122 266988
rect 261478 266976 261484 266988
rect 261536 266976 261542 267028
rect 264974 266976 264980 267028
rect 265032 267016 265038 267028
rect 276382 267016 276388 267028
rect 265032 266988 276388 267016
rect 265032 266976 265038 266988
rect 276382 266976 276388 266988
rect 276440 266976 276446 267028
rect 278038 266976 278044 267028
rect 278096 267016 278102 267028
rect 284662 267016 284668 267028
rect 278096 266988 284668 267016
rect 278096 266976 278102 266988
rect 284662 266976 284668 266988
rect 284720 266976 284726 267028
rect 333514 266976 333520 267028
rect 333572 267016 333578 267028
rect 342254 267016 342260 267028
rect 333572 266988 342260 267016
rect 333572 266976 333578 266988
rect 342254 266976 342260 266988
rect 342312 266976 342318 267028
rect 368106 266976 368112 267028
rect 368164 267016 368170 267028
rect 377766 267016 377772 267028
rect 368164 266988 377772 267016
rect 368164 266976 368170 266988
rect 377766 266976 377772 266988
rect 377824 266976 377830 267028
rect 119798 266840 119804 266892
rect 119856 266880 119862 266892
rect 161750 266880 161756 266892
rect 119856 266852 161756 266880
rect 119856 266840 119862 266852
rect 161750 266840 161756 266852
rect 161808 266840 161814 266892
rect 169846 266840 169852 266892
rect 169904 266880 169910 266892
rect 199102 266880 199108 266892
rect 169904 266852 199108 266880
rect 169904 266840 169910 266852
rect 199102 266840 199108 266852
rect 199160 266840 199166 266892
rect 199286 266840 199292 266892
rect 199344 266880 199350 266892
rect 201862 266880 201868 266892
rect 199344 266852 201868 266880
rect 199344 266840 199350 266852
rect 201862 266840 201868 266852
rect 201920 266840 201926 266892
rect 243538 266840 243544 266892
rect 243596 266880 243602 266892
rect 249058 266880 249064 266892
rect 243596 266852 249064 266880
rect 243596 266840 243602 266852
rect 249058 266840 249064 266852
rect 249116 266840 249122 266892
rect 254578 266840 254584 266892
rect 254636 266880 254642 266892
rect 258994 266880 259000 266892
rect 254636 266852 259000 266880
rect 254636 266840 254642 266852
rect 258994 266840 259000 266852
rect 259052 266840 259058 266892
rect 274634 266840 274640 266892
rect 274692 266880 274698 266892
rect 278038 266880 278044 266892
rect 274692 266852 278044 266880
rect 274692 266840 274698 266852
rect 278038 266840 278044 266852
rect 278096 266840 278102 266892
rect 317782 266840 317788 266892
rect 317840 266880 317846 266892
rect 322934 266880 322940 266892
rect 317840 266852 322940 266880
rect 317840 266840 317846 266852
rect 322934 266840 322940 266852
rect 322992 266840 322998 266892
rect 349246 266840 349252 266892
rect 349304 266880 349310 266892
rect 355318 266880 355324 266892
rect 349304 266852 355324 266880
rect 349304 266840 349310 266852
rect 355318 266840 355324 266852
rect 355376 266840 355382 266892
rect 356698 266840 356704 266892
rect 356756 266880 356762 266892
rect 366358 266880 366364 266892
rect 356756 266852 366364 266880
rect 356756 266840 356762 266852
rect 366358 266840 366364 266852
rect 366416 266840 366422 266892
rect 132586 266704 132592 266756
rect 132644 266744 132650 266756
rect 147214 266744 147220 266756
rect 132644 266716 147220 266744
rect 132644 266704 132650 266716
rect 147214 266704 147220 266716
rect 147272 266704 147278 266756
rect 148502 266704 148508 266756
rect 148560 266744 148566 266756
rect 179506 266744 179512 266756
rect 148560 266716 179512 266744
rect 148560 266704 148566 266716
rect 179506 266704 179512 266716
rect 179564 266704 179570 266756
rect 201586 266704 201592 266756
rect 201644 266744 201650 266756
rect 207014 266744 207020 266756
rect 201644 266716 207020 266744
rect 201644 266704 201650 266716
rect 207014 266704 207020 266716
rect 207072 266704 207078 266756
rect 321922 266704 321928 266756
rect 321980 266744 321986 266756
rect 327074 266744 327080 266756
rect 321980 266716 327080 266744
rect 321980 266704 321986 266716
rect 327074 266704 327080 266716
rect 327132 266704 327138 266756
rect 378796 266744 378824 267124
rect 385678 267112 385684 267164
rect 385736 267152 385742 267164
rect 401870 267152 401876 267164
rect 385736 267124 401876 267152
rect 385736 267112 385742 267124
rect 401870 267112 401876 267124
rect 401928 267112 401934 267164
rect 415486 267112 415492 267164
rect 415544 267152 415550 267164
rect 436738 267152 436744 267164
rect 415544 267124 436744 267152
rect 415544 267112 415550 267124
rect 436738 267112 436744 267124
rect 436796 267112 436802 267164
rect 445294 267112 445300 267164
rect 445352 267152 445358 267164
rect 450722 267152 450728 267164
rect 445352 267124 450728 267152
rect 445352 267112 445358 267124
rect 450722 267112 450728 267124
rect 450780 267112 450786 267164
rect 452562 267112 452568 267164
rect 452620 267152 452626 267164
rect 456058 267152 456064 267164
rect 452620 267124 456064 267152
rect 452620 267112 452626 267124
rect 456058 267112 456064 267124
rect 456116 267112 456122 267164
rect 469122 267152 469128 267164
rect 464632 267124 469128 267152
rect 378962 266976 378968 267028
rect 379020 267016 379026 267028
rect 392118 267016 392124 267028
rect 379020 266988 392124 267016
rect 379020 266976 379026 266988
rect 392118 266976 392124 266988
rect 392176 266976 392182 267028
rect 392302 266976 392308 267028
rect 392360 267016 392366 267028
rect 418798 267016 418804 267028
rect 392360 266988 418804 267016
rect 392360 266976 392366 266988
rect 418798 266976 418804 266988
rect 418856 266976 418862 267028
rect 422938 266976 422944 267028
rect 422996 267016 423002 267028
rect 455046 267016 455052 267028
rect 422996 266988 455052 267016
rect 422996 266976 423002 266988
rect 455046 266976 455052 266988
rect 455104 266976 455110 267028
rect 455414 266976 455420 267028
rect 455472 267016 455478 267028
rect 459554 267016 459560 267028
rect 455472 266988 459560 267016
rect 455472 266976 455478 266988
rect 459554 266976 459560 266988
rect 459612 266976 459618 267028
rect 380618 266840 380624 266892
rect 380676 266880 380682 266892
rect 390186 266880 390192 266892
rect 380676 266852 390192 266880
rect 380676 266840 380682 266852
rect 390186 266840 390192 266852
rect 390244 266840 390250 266892
rect 405550 266840 405556 266892
rect 405608 266880 405614 266892
rect 425698 266880 425704 266892
rect 405608 266852 425704 266880
rect 405608 266840 405614 266852
rect 425698 266840 425704 266852
rect 425756 266840 425762 266892
rect 426066 266840 426072 266892
rect 426124 266880 426130 266892
rect 436554 266880 436560 266892
rect 426124 266852 436560 266880
rect 426124 266840 426130 266852
rect 436554 266840 436560 266852
rect 436612 266840 436618 266892
rect 438670 266840 438676 266892
rect 438728 266880 438734 266892
rect 464632 266880 464660 267124
rect 469122 267112 469128 267124
rect 469180 267112 469186 267164
rect 469306 267112 469312 267164
rect 469364 267152 469370 267164
rect 470502 267152 470508 267164
rect 469364 267124 470508 267152
rect 469364 267112 469370 267124
rect 470502 267112 470508 267124
rect 470560 267112 470566 267164
rect 473262 267112 473268 267164
rect 473320 267152 473326 267164
rect 512178 267152 512184 267164
rect 473320 267124 512184 267152
rect 473320 267112 473326 267124
rect 512178 267112 512184 267124
rect 512236 267112 512242 267164
rect 512362 267112 512368 267164
rect 512420 267152 512426 267164
rect 518866 267152 518894 267260
rect 582190 267248 582196 267260
rect 582248 267248 582254 267300
rect 512420 267124 518894 267152
rect 512420 267112 512426 267124
rect 520642 267112 520648 267164
rect 520700 267152 520706 267164
rect 524230 267152 524236 267164
rect 520700 267124 524236 267152
rect 520700 267112 520706 267124
rect 524230 267112 524236 267124
rect 524288 267112 524294 267164
rect 615494 267152 615500 267164
rect 528526 267124 615500 267152
rect 468478 267016 468484 267028
rect 438728 266852 464660 266880
rect 464724 266988 468484 267016
rect 438728 266840 438734 266852
rect 383654 266744 383660 266756
rect 378796 266716 383660 266744
rect 383654 266704 383660 266716
rect 383712 266704 383718 266756
rect 398098 266704 398104 266756
rect 398156 266744 398162 266756
rect 414474 266744 414480 266756
rect 398156 266716 414480 266744
rect 398156 266704 398162 266716
rect 414474 266704 414480 266716
rect 414532 266704 414538 266756
rect 423766 266704 423772 266756
rect 423824 266744 423830 266756
rect 424962 266744 424968 266756
rect 423824 266716 424968 266744
rect 423824 266704 423830 266716
rect 424962 266704 424968 266716
rect 425020 266704 425026 266756
rect 425422 266704 425428 266756
rect 425480 266744 425486 266756
rect 426250 266744 426256 266756
rect 425480 266716 426256 266744
rect 425480 266704 425486 266716
rect 426250 266704 426256 266716
rect 426308 266704 426314 266756
rect 427906 266704 427912 266756
rect 427964 266744 427970 266756
rect 428918 266744 428924 266756
rect 427964 266716 428924 266744
rect 427964 266704 427970 266716
rect 428918 266704 428924 266716
rect 428976 266704 428982 266756
rect 437842 266704 437848 266756
rect 437900 266744 437906 266756
rect 464724 266744 464752 266988
rect 468478 266976 468484 266988
rect 468536 266976 468542 267028
rect 468938 266976 468944 267028
rect 468996 267016 469002 267028
rect 484026 267016 484032 267028
rect 468996 266988 484032 267016
rect 468996 266976 469002 266988
rect 484026 266976 484032 266988
rect 484084 266976 484090 267028
rect 523678 267016 523684 267028
rect 485056 266988 523684 267016
rect 465166 266840 465172 266892
rect 465224 266880 465230 266892
rect 465224 266852 467972 266880
rect 465224 266840 465230 266852
rect 437900 266716 464752 266744
rect 437900 266704 437906 266716
rect 466822 266704 466828 266756
rect 466880 266744 466886 266756
rect 467742 266744 467748 266756
rect 466880 266716 467748 266744
rect 466880 266704 466886 266716
rect 467742 266704 467748 266716
rect 467800 266704 467806 266756
rect 467944 266744 467972 266852
rect 470134 266840 470140 266892
rect 470192 266880 470198 266892
rect 485056 266880 485084 266988
rect 523678 266976 523684 266988
rect 523736 266976 523742 267028
rect 528526 267016 528554 267124
rect 615494 267112 615500 267124
rect 615552 267112 615558 267164
rect 523880 266988 528554 267016
rect 528756 266988 530072 267016
rect 470192 266852 485084 266880
rect 470192 266840 470198 266852
rect 487522 266840 487528 266892
rect 487580 266880 487586 266892
rect 514018 266880 514024 266892
rect 487580 266852 514024 266880
rect 487580 266840 487586 266852
rect 514018 266840 514024 266852
rect 514076 266840 514082 266892
rect 514386 266840 514392 266892
rect 514444 266880 514450 266892
rect 517514 266880 517520 266892
rect 514444 266852 517520 266880
rect 514444 266840 514450 266852
rect 517514 266840 517520 266852
rect 517572 266840 517578 266892
rect 518986 266840 518992 266892
rect 519044 266880 519050 266892
rect 520090 266880 520096 266892
rect 519044 266852 520096 266880
rect 519044 266840 519050 266852
rect 520090 266840 520096 266852
rect 520148 266840 520154 266892
rect 522298 266840 522304 266892
rect 522356 266880 522362 266892
rect 523880 266880 523908 266988
rect 522356 266852 523908 266880
rect 522356 266840 522362 266852
rect 524230 266840 524236 266892
rect 524288 266880 524294 266892
rect 528756 266880 528784 266988
rect 524288 266852 528784 266880
rect 524288 266840 524294 266852
rect 528922 266840 528928 266892
rect 528980 266880 528986 266892
rect 529750 266880 529756 266892
rect 528980 266852 529756 266880
rect 528980 266840 528986 266852
rect 529750 266840 529756 266852
rect 529808 266840 529814 266892
rect 530044 266880 530072 266988
rect 537202 266976 537208 267028
rect 537260 267016 537266 267028
rect 636194 267016 636200 267028
rect 537260 266988 636200 267016
rect 537260 266976 537266 266988
rect 636194 266976 636200 266988
rect 636252 266976 636258 267028
rect 537478 266880 537484 266892
rect 530044 266852 537484 266880
rect 537478 266840 537484 266852
rect 537536 266840 537542 266892
rect 540974 266840 540980 266892
rect 541032 266880 541038 266892
rect 541618 266880 541624 266892
rect 541032 266852 541624 266880
rect 541032 266840 541038 266852
rect 541618 266840 541624 266852
rect 541676 266840 541682 266892
rect 541894 266840 541900 266892
rect 541952 266880 541958 266892
rect 602338 266880 602344 266892
rect 541952 266852 602344 266880
rect 541952 266840 541958 266852
rect 602338 266840 602344 266852
rect 602396 266840 602402 266892
rect 473262 266744 473268 266756
rect 467944 266716 473268 266744
rect 473262 266704 473268 266716
rect 473320 266704 473326 266756
rect 473446 266704 473452 266756
rect 473504 266744 473510 266756
rect 474366 266744 474372 266756
rect 473504 266716 474372 266744
rect 473504 266704 473510 266716
rect 474366 266704 474372 266716
rect 474424 266704 474430 266756
rect 477586 266704 477592 266756
rect 477644 266744 477650 266756
rect 478598 266744 478604 266756
rect 477644 266716 478604 266744
rect 477644 266704 477650 266716
rect 478598 266704 478604 266716
rect 478656 266704 478662 266756
rect 483382 266704 483388 266756
rect 483440 266744 483446 266756
rect 484302 266744 484308 266756
rect 483440 266716 484308 266744
rect 483440 266704 483446 266716
rect 484302 266704 484308 266716
rect 484360 266704 484366 266756
rect 485866 266704 485872 266756
rect 485924 266744 485930 266756
rect 487062 266744 487068 266756
rect 485924 266716 487068 266744
rect 485924 266704 485930 266716
rect 487062 266704 487068 266716
rect 487120 266704 487126 266756
rect 494974 266704 494980 266756
rect 495032 266744 495038 266756
rect 499666 266744 499672 266756
rect 495032 266716 499672 266744
rect 495032 266704 495038 266716
rect 499666 266704 499672 266716
rect 499724 266704 499730 266756
rect 499850 266704 499856 266756
rect 499908 266744 499914 266756
rect 501598 266744 501604 266756
rect 499908 266716 501604 266744
rect 499908 266704 499914 266716
rect 501598 266704 501604 266716
rect 501656 266704 501662 266756
rect 502426 266704 502432 266756
rect 502484 266744 502490 266756
rect 559742 266744 559748 266756
rect 502484 266716 559748 266744
rect 502484 266704 502490 266716
rect 559742 266704 559748 266716
rect 559800 266704 559806 266756
rect 258074 266636 258080 266688
rect 258132 266676 258138 266688
rect 267274 266676 267280 266688
rect 258132 266648 267280 266676
rect 258132 266636 258138 266648
rect 267274 266636 267280 266648
rect 267332 266636 267338 266688
rect 312814 266636 312820 266688
rect 312872 266676 312878 266688
rect 316402 266676 316408 266688
rect 312872 266648 316408 266676
rect 312872 266636 312878 266648
rect 316402 266636 316408 266648
rect 316460 266636 316466 266688
rect 389818 266636 389824 266688
rect 389876 266676 389882 266688
rect 395338 266676 395344 266688
rect 389876 266648 395344 266676
rect 389876 266636 389882 266648
rect 395338 266636 395344 266648
rect 395396 266636 395402 266688
rect 123478 266568 123484 266620
rect 123536 266608 123542 266620
rect 150526 266608 150532 266620
rect 123536 266580 150532 266608
rect 123536 266568 123542 266580
rect 150526 266568 150532 266580
rect 150584 266568 150590 266620
rect 154022 266568 154028 266620
rect 154080 266608 154086 266620
rect 170398 266608 170404 266620
rect 154080 266580 170404 266608
rect 154080 266568 154086 266580
rect 170398 266568 170404 266580
rect 170456 266568 170462 266620
rect 416314 266568 416320 266620
rect 416372 266608 416378 266620
rect 438118 266608 438124 266620
rect 416372 266580 438124 266608
rect 416372 266568 416378 266580
rect 438118 266568 438124 266580
rect 438176 266568 438182 266620
rect 446950 266568 446956 266620
rect 447008 266608 447014 266620
rect 452562 266608 452568 266620
rect 447008 266580 452568 266608
rect 447008 266568 447014 266580
rect 452562 266568 452568 266580
rect 452620 266568 452626 266620
rect 452746 266568 452752 266620
rect 452804 266608 452810 266620
rect 453666 266608 453672 266620
rect 452804 266580 453672 266608
rect 452804 266568 452810 266580
rect 453666 266568 453672 266580
rect 453724 266568 453730 266620
rect 454402 266568 454408 266620
rect 454460 266608 454466 266620
rect 455414 266608 455420 266620
rect 454460 266580 455420 266608
rect 454460 266568 454466 266580
rect 455414 266568 455420 266580
rect 455472 266568 455478 266620
rect 456886 266568 456892 266620
rect 456944 266608 456950 266620
rect 457990 266608 457996 266620
rect 456944 266580 457996 266608
rect 456944 266568 456950 266580
rect 457990 266568 457996 266580
rect 458048 266568 458054 266620
rect 460198 266568 460204 266620
rect 460256 266608 460262 266620
rect 490558 266608 490564 266620
rect 460256 266580 490564 266608
rect 460256 266568 460262 266580
rect 490558 266568 490564 266580
rect 490616 266568 490622 266620
rect 491662 266568 491668 266620
rect 491720 266608 491726 266620
rect 492582 266608 492588 266620
rect 491720 266580 492588 266608
rect 491720 266568 491726 266580
rect 492582 266568 492588 266580
rect 492640 266568 492646 266620
rect 494146 266568 494152 266620
rect 494204 266608 494210 266620
rect 495250 266608 495256 266620
rect 494204 266580 495256 266608
rect 494204 266568 494210 266580
rect 495250 266568 495256 266580
rect 495308 266568 495314 266620
rect 497458 266568 497464 266620
rect 497516 266608 497522 266620
rect 552658 266608 552664 266620
rect 497516 266580 552664 266608
rect 497516 266568 497522 266580
rect 552658 266568 552664 266580
rect 552716 266568 552722 266620
rect 222838 266500 222844 266552
rect 222896 266540 222902 266552
rect 226702 266540 226708 266552
rect 222896 266512 226708 266540
rect 222896 266500 222902 266512
rect 226702 266500 226708 266512
rect 226760 266500 226766 266552
rect 253198 266500 253204 266552
rect 253256 266540 253262 266552
rect 256510 266540 256516 266552
rect 253256 266512 256516 266540
rect 253256 266500 253262 266512
rect 256510 266500 256516 266512
rect 256568 266500 256574 266552
rect 256694 266500 256700 266552
rect 256752 266540 256758 266552
rect 259822 266540 259828 266552
rect 256752 266512 259828 266540
rect 256752 266500 256758 266512
rect 259822 266500 259828 266512
rect 259880 266500 259886 266552
rect 308674 266500 308680 266552
rect 308732 266540 308738 266552
rect 310882 266540 310888 266552
rect 308732 266512 310888 266540
rect 308732 266500 308738 266512
rect 310882 266500 310888 266512
rect 310940 266500 310946 266552
rect 311158 266500 311164 266552
rect 311216 266540 311222 266552
rect 313274 266540 313280 266552
rect 311216 266512 313280 266540
rect 311216 266500 311222 266512
rect 313274 266500 313280 266512
rect 313332 266500 313338 266552
rect 320266 266500 320272 266552
rect 320324 266540 320330 266552
rect 324958 266540 324964 266552
rect 320324 266512 324964 266540
rect 320324 266500 320330 266512
rect 324958 266500 324964 266512
rect 325016 266500 325022 266552
rect 330202 266500 330208 266552
rect 330260 266540 330266 266552
rect 334618 266540 334624 266552
rect 330260 266512 334624 266540
rect 330260 266500 330266 266512
rect 334618 266500 334624 266512
rect 334676 266500 334682 266552
rect 345106 266500 345112 266552
rect 345164 266540 345170 266552
rect 351178 266540 351184 266552
rect 345164 266512 351184 266540
rect 345164 266500 345170 266512
rect 351178 266500 351184 266512
rect 351236 266500 351242 266552
rect 395614 266500 395620 266552
rect 395672 266540 395678 266552
rect 404998 266540 405004 266552
rect 395672 266512 405004 266540
rect 395672 266500 395678 266512
rect 404998 266500 405004 266512
rect 405056 266500 405062 266552
rect 141602 266432 141608 266484
rect 141660 266472 141666 266484
rect 146938 266472 146944 266484
rect 141660 266444 146944 266472
rect 141660 266432 141666 266444
rect 146938 266432 146944 266444
rect 146996 266432 147002 266484
rect 421282 266432 421288 266484
rect 421340 266472 421346 266484
rect 421340 266444 431954 266472
rect 421340 266432 421346 266444
rect 156598 266364 156604 266416
rect 156656 266404 156662 266416
rect 159634 266404 159640 266416
rect 156656 266376 159640 266404
rect 156656 266364 156662 266376
rect 159634 266364 159640 266376
rect 159692 266364 159698 266416
rect 162118 266364 162124 266416
rect 162176 266404 162182 266416
rect 162946 266404 162952 266416
rect 162176 266376 162952 266404
rect 162176 266364 162182 266376
rect 162946 266364 162952 266376
rect 163004 266364 163010 266416
rect 165062 266364 165068 266416
rect 165120 266404 165126 266416
rect 169570 266404 169576 266416
rect 165120 266376 169576 266404
rect 165120 266364 165126 266376
rect 169570 266364 169576 266376
rect 169628 266364 169634 266416
rect 181530 266364 181536 266416
rect 181588 266404 181594 266416
rect 182818 266404 182824 266416
rect 181588 266376 182824 266404
rect 181588 266364 181594 266376
rect 182818 266364 182824 266376
rect 182876 266364 182882 266416
rect 183002 266364 183008 266416
rect 183060 266404 183066 266416
rect 186130 266404 186136 266416
rect 183060 266376 186136 266404
rect 183060 266364 183066 266376
rect 186130 266364 186136 266376
rect 186188 266364 186194 266416
rect 192478 266364 192484 266416
rect 192536 266404 192542 266416
rect 197722 266404 197728 266416
rect 192536 266376 197728 266404
rect 192536 266364 192542 266376
rect 197722 266364 197728 266376
rect 197780 266364 197786 266416
rect 200390 266364 200396 266416
rect 200448 266404 200454 266416
rect 202690 266404 202696 266416
rect 200448 266376 202696 266404
rect 200448 266364 200454 266376
rect 202690 266364 202696 266376
rect 202748 266364 202754 266416
rect 213178 266364 213184 266416
rect 213236 266404 213242 266416
rect 215938 266404 215944 266416
rect 213236 266376 215944 266404
rect 213236 266364 213242 266376
rect 215938 266364 215944 266376
rect 215996 266364 216002 266416
rect 221458 266364 221464 266416
rect 221516 266404 221522 266416
rect 224218 266404 224224 266416
rect 221516 266376 224224 266404
rect 221516 266364 221522 266376
rect 224218 266364 224224 266376
rect 224276 266364 224282 266416
rect 239490 266364 239496 266416
rect 239548 266404 239554 266416
rect 244090 266404 244096 266416
rect 239548 266376 244096 266404
rect 239548 266364 239554 266376
rect 244090 266364 244096 266376
rect 244148 266364 244154 266416
rect 256142 266364 256148 266416
rect 256200 266404 256206 266416
rect 258166 266404 258172 266416
rect 256200 266376 258172 266404
rect 256200 266364 256206 266376
rect 258166 266364 258172 266376
rect 258224 266364 258230 266416
rect 268010 266364 268016 266416
rect 268068 266404 268074 266416
rect 272242 266404 272248 266416
rect 268068 266376 272248 266404
rect 268068 266364 268074 266376
rect 272242 266364 272248 266376
rect 272300 266364 272306 266416
rect 272518 266364 272524 266416
rect 272576 266404 272582 266416
rect 274726 266404 274732 266416
rect 272576 266376 274732 266404
rect 272576 266364 272582 266376
rect 274726 266364 274732 266376
rect 274784 266364 274790 266416
rect 287698 266364 287704 266416
rect 287756 266404 287762 266416
rect 292114 266404 292120 266416
rect 287756 266376 292120 266404
rect 287756 266364 287762 266376
rect 292114 266364 292120 266376
rect 292172 266364 292178 266416
rect 301038 266364 301044 266416
rect 301096 266404 301102 266416
rect 302050 266404 302056 266416
rect 301096 266376 302056 266404
rect 301096 266364 301102 266376
rect 302050 266364 302056 266376
rect 302108 266364 302114 266416
rect 307846 266364 307852 266416
rect 307904 266404 307910 266416
rect 309502 266404 309508 266416
rect 307904 266376 309508 266404
rect 307904 266364 307910 266376
rect 309502 266364 309508 266376
rect 309560 266364 309566 266416
rect 310330 266364 310336 266416
rect 310388 266404 310394 266416
rect 311894 266404 311900 266416
rect 310388 266376 311900 266404
rect 310388 266364 310394 266376
rect 311894 266364 311900 266376
rect 311952 266364 311958 266416
rect 312354 266364 312360 266416
rect 312412 266404 312418 266416
rect 314654 266404 314660 266416
rect 312412 266376 314660 266404
rect 312412 266364 312418 266376
rect 314654 266364 314660 266376
rect 314712 266364 314718 266416
rect 316126 266364 316132 266416
rect 316184 266404 316190 266416
rect 320542 266404 320548 266416
rect 316184 266376 320548 266404
rect 316184 266364 316190 266376
rect 320542 266364 320548 266376
rect 320600 266364 320606 266416
rect 328546 266364 328552 266416
rect 328604 266404 328610 266416
rect 329742 266404 329748 266416
rect 328604 266376 329748 266404
rect 328604 266364 328610 266376
rect 329742 266364 329748 266376
rect 329800 266364 329806 266416
rect 332686 266364 332692 266416
rect 332744 266404 332750 266416
rect 333790 266404 333796 266416
rect 332744 266376 333796 266404
rect 332744 266364 332750 266376
rect 333790 266364 333796 266376
rect 333848 266364 333854 266416
rect 342622 266364 342628 266416
rect 342680 266404 342686 266416
rect 343542 266404 343548 266416
rect 342680 266376 343548 266404
rect 342680 266364 342686 266376
rect 343542 266364 343548 266376
rect 343600 266364 343606 266416
rect 347590 266364 347596 266416
rect 347648 266404 347654 266416
rect 349798 266404 349804 266416
rect 347648 266376 349804 266404
rect 347648 266364 347654 266376
rect 349798 266364 349804 266376
rect 349856 266364 349862 266416
rect 355042 266364 355048 266416
rect 355100 266404 355106 266416
rect 356882 266404 356888 266416
rect 355100 266376 356888 266404
rect 355100 266364 355106 266376
rect 356882 266364 356888 266376
rect 356940 266364 356946 266416
rect 358354 266364 358360 266416
rect 358412 266404 358418 266416
rect 360838 266404 360844 266416
rect 358412 266376 360844 266404
rect 358412 266364 358418 266376
rect 360838 266364 360844 266376
rect 360896 266364 360902 266416
rect 361666 266364 361672 266416
rect 361724 266404 361730 266416
rect 362862 266404 362868 266416
rect 361724 266376 362868 266404
rect 361724 266364 361730 266376
rect 362862 266364 362868 266376
rect 362920 266364 362926 266416
rect 367462 266364 367468 266416
rect 367520 266404 367526 266416
rect 368290 266404 368296 266416
rect 367520 266376 368296 266404
rect 367520 266364 367526 266376
rect 368290 266364 368296 266376
rect 368348 266364 368354 266416
rect 371602 266364 371608 266416
rect 371660 266404 371666 266416
rect 372522 266404 372528 266416
rect 371660 266376 372528 266404
rect 371660 266364 371666 266376
rect 372522 266364 372528 266376
rect 372580 266364 372586 266416
rect 374086 266364 374092 266416
rect 374144 266404 374150 266416
rect 375282 266404 375288 266416
rect 374144 266376 375288 266404
rect 374144 266364 374150 266376
rect 375282 266364 375288 266376
rect 375340 266364 375346 266416
rect 377398 266364 377404 266416
rect 377456 266404 377462 266416
rect 378778 266404 378784 266416
rect 377456 266376 378784 266404
rect 377456 266364 377462 266376
rect 378778 266364 378784 266376
rect 378836 266364 378842 266416
rect 379882 266364 379888 266416
rect 379940 266404 379946 266416
rect 380802 266404 380808 266416
rect 379940 266376 380808 266404
rect 379940 266364 379946 266376
rect 380802 266364 380808 266376
rect 380860 266364 380866 266416
rect 384022 266364 384028 266416
rect 384080 266404 384086 266416
rect 384942 266404 384948 266416
rect 384080 266376 384948 266404
rect 384080 266364 384086 266376
rect 384942 266364 384948 266376
rect 385000 266364 385006 266416
rect 386506 266364 386512 266416
rect 386564 266404 386570 266416
rect 387610 266404 387616 266416
rect 386564 266376 387616 266404
rect 386564 266364 386570 266376
rect 387610 266364 387616 266376
rect 387668 266364 387674 266416
rect 396442 266364 396448 266416
rect 396500 266404 396506 266416
rect 397270 266404 397276 266416
rect 396500 266376 397276 266404
rect 396500 266364 396506 266376
rect 397270 266364 397276 266376
rect 397328 266364 397334 266416
rect 398926 266364 398932 266416
rect 398984 266404 398990 266416
rect 400122 266404 400128 266416
rect 398984 266376 400128 266404
rect 398984 266364 398990 266376
rect 400122 266364 400128 266376
rect 400180 266364 400186 266416
rect 403066 266364 403072 266416
rect 403124 266404 403130 266416
rect 404170 266404 404176 266416
rect 403124 266376 404176 266404
rect 403124 266364 403130 266376
rect 404170 266364 404176 266376
rect 404228 266364 404234 266416
rect 411346 266364 411352 266416
rect 411404 266404 411410 266416
rect 412266 266404 412272 266416
rect 411404 266376 412272 266404
rect 411404 266364 411410 266376
rect 412266 266364 412272 266376
rect 412324 266364 412330 266416
rect 417142 266364 417148 266416
rect 417200 266404 417206 266416
rect 419810 266404 419816 266416
rect 417200 266376 419816 266404
rect 417200 266364 417206 266376
rect 419810 266364 419816 266376
rect 419868 266364 419874 266416
rect 431926 266268 431954 266444
rect 450722 266432 450728 266484
rect 450780 266472 450786 266484
rect 499758 266472 499764 266484
rect 450780 266444 499764 266472
rect 450780 266432 450786 266444
rect 499758 266432 499764 266444
rect 499816 266432 499822 266484
rect 499942 266432 499948 266484
rect 500000 266472 500006 266484
rect 500862 266472 500868 266484
rect 500000 266444 500868 266472
rect 500000 266432 500006 266444
rect 500862 266432 500868 266444
rect 500920 266432 500926 266484
rect 504082 266432 504088 266484
rect 504140 266472 504146 266484
rect 504910 266472 504916 266484
rect 504140 266444 504916 266472
rect 504140 266432 504146 266444
rect 504910 266432 504916 266444
rect 504968 266432 504974 266484
rect 506566 266432 506572 266484
rect 506624 266472 506630 266484
rect 507670 266472 507676 266484
rect 506624 266444 507676 266472
rect 506624 266432 506630 266444
rect 507670 266432 507676 266444
rect 507728 266432 507734 266484
rect 507854 266432 507860 266484
rect 507912 266472 507918 266484
rect 510062 266472 510068 266484
rect 507912 266444 510068 266472
rect 507912 266432 507918 266444
rect 510062 266432 510068 266444
rect 510120 266432 510126 266484
rect 514846 266432 514852 266484
rect 514904 266472 514910 266484
rect 516042 266472 516048 266484
rect 514904 266444 516048 266472
rect 514904 266432 514910 266444
rect 516042 266432 516048 266444
rect 516100 266432 516106 266484
rect 516502 266432 516508 266484
rect 516560 266472 516566 266484
rect 517330 266472 517336 266484
rect 516560 266444 517336 266472
rect 516560 266432 516566 266444
rect 517330 266432 517336 266444
rect 517388 266432 517394 266484
rect 517514 266432 517520 266484
rect 517572 266472 517578 266484
rect 540974 266472 540980 266484
rect 517572 266444 540980 266472
rect 517572 266432 517578 266444
rect 540974 266432 540980 266444
rect 541032 266432 541038 266484
rect 541342 266432 541348 266484
rect 541400 266472 541406 266484
rect 542078 266472 542084 266484
rect 541400 266444 542084 266472
rect 541400 266432 541406 266444
rect 542078 266432 542084 266444
rect 542136 266432 542142 266484
rect 432046 266364 432052 266416
rect 432104 266404 432110 266416
rect 433150 266404 433156 266416
rect 432104 266376 433156 266404
rect 432104 266364 432110 266376
rect 433150 266364 433156 266376
rect 433208 266364 433214 266416
rect 439314 266404 439320 266416
rect 433352 266376 439320 266404
rect 433352 266268 433380 266376
rect 439314 266364 439320 266376
rect 439372 266364 439378 266416
rect 440326 266364 440332 266416
rect 440384 266404 440390 266416
rect 441338 266404 441344 266416
rect 440384 266376 441344 266404
rect 440384 266364 440390 266376
rect 441338 266364 441344 266376
rect 441396 266364 441402 266416
rect 441982 266364 441988 266416
rect 442040 266404 442046 266416
rect 442902 266404 442908 266416
rect 442040 266376 442908 266404
rect 442040 266364 442046 266376
rect 442902 266364 442908 266376
rect 442960 266364 442966 266416
rect 444466 266364 444472 266416
rect 444524 266404 444530 266416
rect 445662 266404 445668 266416
rect 444524 266376 445668 266404
rect 444524 266364 444530 266376
rect 445662 266364 445668 266376
rect 445720 266364 445726 266416
rect 446122 266364 446128 266416
rect 446180 266404 446186 266416
rect 447778 266404 447784 266416
rect 446180 266376 447784 266404
rect 446180 266364 446186 266376
rect 447778 266364 447784 266376
rect 447836 266364 447842 266416
rect 448146 266364 448152 266416
rect 448204 266404 448210 266416
rect 450538 266404 450544 266416
rect 448204 266376 450544 266404
rect 448204 266364 448210 266376
rect 450538 266364 450544 266376
rect 450596 266364 450602 266416
rect 480070 266296 480076 266348
rect 480128 266336 480134 266348
rect 554774 266336 554780 266348
rect 480128 266308 554780 266336
rect 480128 266296 480134 266308
rect 554774 266296 554780 266308
rect 554832 266296 554838 266348
rect 431926 266240 433380 266268
rect 485038 266160 485044 266212
rect 485096 266200 485102 266212
rect 561674 266200 561680 266212
rect 485096 266172 561680 266200
rect 485096 266160 485102 266172
rect 561674 266160 561680 266172
rect 561732 266160 561738 266212
rect 486694 266024 486700 266076
rect 486752 266064 486758 266076
rect 564434 266064 564440 266076
rect 486752 266036 564440 266064
rect 486752 266024 486758 266036
rect 564434 266024 564440 266036
rect 564492 266024 564498 266076
rect 142154 265888 142160 265940
rect 142212 265928 142218 265940
rect 142798 265928 142804 265940
rect 142212 265900 142804 265928
rect 142212 265888 142218 265900
rect 142798 265888 142804 265900
rect 142856 265888 142862 265940
rect 234614 265888 234620 265940
rect 234672 265928 234678 265940
rect 235534 265928 235540 265940
rect 234672 265900 235540 265928
rect 234672 265888 234678 265900
rect 235534 265888 235540 265900
rect 235592 265888 235598 265940
rect 292758 265888 292764 265940
rect 292816 265928 292822 265940
rect 293494 265928 293500 265940
rect 292816 265900 293500 265928
rect 292816 265888 292822 265900
rect 293494 265888 293500 265900
rect 293552 265888 293558 265940
rect 492490 265888 492496 265940
rect 492548 265928 492554 265940
rect 572714 265928 572720 265940
rect 492548 265900 572720 265928
rect 492548 265888 492554 265900
rect 572714 265888 572720 265900
rect 572772 265888 572778 265940
rect 515674 265752 515680 265804
rect 515732 265792 515738 265804
rect 605834 265792 605840 265804
rect 515732 265764 605840 265792
rect 515732 265752 515738 265764
rect 605834 265752 605840 265764
rect 605892 265752 605898 265804
rect 518158 265616 518164 265668
rect 518216 265656 518222 265668
rect 608686 265656 608692 265668
rect 518216 265628 608692 265656
rect 518216 265616 518222 265628
rect 608686 265616 608692 265628
rect 608744 265616 608750 265668
rect 481726 265480 481732 265532
rect 481784 265520 481790 265532
rect 557534 265520 557540 265532
rect 481784 265492 557540 265520
rect 481784 265480 481790 265492
rect 557534 265480 557540 265492
rect 557592 265480 557598 265532
rect 479242 265344 479248 265396
rect 479300 265384 479306 265396
rect 553394 265384 553400 265396
rect 479300 265356 553400 265384
rect 479300 265344 479306 265356
rect 553394 265344 553400 265356
rect 553452 265344 553458 265396
rect 577498 261604 577504 261656
rect 577556 261644 577562 261656
rect 648614 261644 648620 261656
rect 577556 261616 648620 261644
rect 577556 261604 577562 261616
rect 648614 261604 648620 261616
rect 648672 261604 648678 261656
rect 570598 261468 570604 261520
rect 570656 261508 570662 261520
rect 645854 261508 645860 261520
rect 570656 261480 645860 261508
rect 570656 261468 570662 261480
rect 645854 261468 645860 261480
rect 645912 261468 645918 261520
rect 554406 260856 554412 260908
rect 554464 260896 554470 260908
rect 568574 260896 568580 260908
rect 554464 260868 568580 260896
rect 554464 260856 554470 260868
rect 568574 260856 568580 260868
rect 568632 260856 568638 260908
rect 675846 260176 675852 260228
rect 675904 260216 675910 260228
rect 676398 260216 676404 260228
rect 675904 260188 676404 260216
rect 675904 260176 675910 260188
rect 676398 260176 676404 260188
rect 676456 260176 676462 260228
rect 554314 259428 554320 259480
rect 554372 259468 554378 259480
rect 560938 259468 560944 259480
rect 554372 259440 560944 259468
rect 554372 259428 554378 259440
rect 560938 259428 560944 259440
rect 560996 259428 561002 259480
rect 553946 256708 553952 256760
rect 554004 256748 554010 256760
rect 559558 256748 559564 256760
rect 554004 256720 559564 256748
rect 554004 256708 554010 256720
rect 559558 256708 559564 256720
rect 559616 256708 559622 256760
rect 35802 252696 35808 252748
rect 35860 252736 35866 252748
rect 41690 252736 41696 252748
rect 35860 252708 41696 252736
rect 35860 252696 35866 252708
rect 41690 252696 41696 252708
rect 41748 252696 41754 252748
rect 35618 252560 35624 252612
rect 35676 252600 35682 252612
rect 40678 252600 40684 252612
rect 35676 252572 40684 252600
rect 35676 252560 35682 252572
rect 40678 252560 40684 252572
rect 40736 252560 40742 252612
rect 554406 252560 554412 252612
rect 554464 252600 554470 252612
rect 562318 252600 562324 252612
rect 554464 252572 562324 252600
rect 554464 252560 554470 252572
rect 562318 252560 562324 252572
rect 562376 252560 562382 252612
rect 675846 252220 675852 252272
rect 675904 252260 675910 252272
rect 678238 252260 678244 252272
rect 675904 252232 678244 252260
rect 675904 252220 675910 252232
rect 678238 252220 678244 252232
rect 678296 252220 678302 252272
rect 35802 251200 35808 251252
rect 35860 251240 35866 251252
rect 37918 251240 37924 251252
rect 35860 251212 37924 251240
rect 35860 251200 35866 251212
rect 37918 251200 37924 251212
rect 37976 251200 37982 251252
rect 554130 251200 554136 251252
rect 554188 251240 554194 251252
rect 556798 251240 556804 251252
rect 554188 251212 556804 251240
rect 554188 251200 554194 251212
rect 556798 251200 556804 251212
rect 556856 251200 556862 251252
rect 675478 251200 675484 251252
rect 675536 251200 675542 251252
rect 675496 250980 675524 251200
rect 675478 250928 675484 250980
rect 675536 250928 675542 250980
rect 553486 249024 553492 249076
rect 553544 249064 553550 249076
rect 571334 249064 571340 249076
rect 553544 249036 571340 249064
rect 553544 249024 553550 249036
rect 571334 249024 571340 249036
rect 571392 249024 571398 249076
rect 553854 246304 553860 246356
rect 553912 246344 553918 246356
rect 632698 246344 632704 246356
rect 553912 246316 632704 246344
rect 553912 246304 553918 246316
rect 632698 246304 632704 246316
rect 632756 246304 632762 246356
rect 554406 245624 554412 245676
rect 554464 245664 554470 245676
rect 592678 245664 592684 245676
rect 554464 245636 592684 245664
rect 554464 245624 554470 245636
rect 592678 245624 592684 245636
rect 592736 245624 592742 245676
rect 553394 244264 553400 244316
rect 553452 244304 553458 244316
rect 555418 244304 555424 244316
rect 553452 244276 555424 244304
rect 553452 244264 553458 244276
rect 555418 244264 555424 244276
rect 555476 244264 555482 244316
rect 37918 242836 37924 242888
rect 37976 242876 37982 242888
rect 41690 242876 41696 242888
rect 37976 242848 41696 242876
rect 37976 242836 37982 242848
rect 41690 242836 41696 242848
rect 41748 242836 41754 242888
rect 34422 242156 34428 242208
rect 34480 242196 34486 242208
rect 41690 242196 41696 242208
rect 34480 242168 41696 242196
rect 34480 242156 34486 242168
rect 41690 242156 41696 242168
rect 41748 242156 41754 242208
rect 558178 242156 558184 242208
rect 558236 242196 558242 242208
rect 647234 242196 647240 242208
rect 558236 242168 647240 242196
rect 558236 242156 558242 242168
rect 647234 242156 647240 242168
rect 647292 242156 647298 242208
rect 553946 241476 553952 241528
rect 554004 241516 554010 241528
rect 621658 241516 621664 241528
rect 554004 241488 621664 241516
rect 554004 241476 554010 241488
rect 621658 241476 621664 241488
rect 621716 241476 621722 241528
rect 554314 238688 554320 238740
rect 554372 238728 554378 238740
rect 577498 238728 577504 238740
rect 554372 238700 577504 238728
rect 554372 238688 554378 238700
rect 577498 238688 577504 238700
rect 577556 238688 577562 238740
rect 671062 237804 671068 237856
rect 671120 237844 671126 237856
rect 672756 237844 672784 238102
rect 671120 237816 672784 237844
rect 671120 237804 671126 237816
rect 671706 237532 671712 237584
rect 671764 237572 671770 237584
rect 672874 237572 672902 237898
rect 671764 237544 672902 237572
rect 671764 237532 671770 237544
rect 668762 237396 668768 237448
rect 668820 237436 668826 237448
rect 672966 237436 672994 237694
rect 668820 237408 672994 237436
rect 668820 237396 668826 237408
rect 671338 237124 671344 237176
rect 671396 237164 671402 237176
rect 673104 237164 673132 237490
rect 671396 237136 673132 237164
rect 671396 237124 671402 237136
rect 671522 236988 671528 237040
rect 671580 237028 671586 237040
rect 673196 237028 673224 237286
rect 671580 237000 673224 237028
rect 671580 236988 671586 237000
rect 673086 236716 673092 236768
rect 673144 236756 673150 236768
rect 673316 236756 673344 237082
rect 673414 236904 673466 236910
rect 673414 236846 673466 236852
rect 673528 236904 673580 236910
rect 673528 236846 673580 236852
rect 673144 236728 673344 236756
rect 673144 236716 673150 236728
rect 672534 236444 672540 236496
rect 672592 236484 672598 236496
rect 672592 236456 673670 236484
rect 672592 236444 672598 236456
rect 673752 236292 673804 236298
rect 673752 236234 673804 236240
rect 673454 236104 673460 236156
rect 673512 236144 673518 236156
rect 673512 236116 673900 236144
rect 673512 236104 673518 236116
rect 554498 236036 554504 236088
rect 554556 236076 554562 236088
rect 558178 236076 558184 236088
rect 554556 236048 558184 236076
rect 554556 236036 554562 236048
rect 558178 236036 558184 236048
rect 558236 236036 558242 236088
rect 673454 235900 673460 235952
rect 673512 235940 673518 235952
rect 673512 235912 673992 235940
rect 673512 235900 673518 235912
rect 674082 235628 674088 235680
rect 674140 235628 674146 235680
rect 673362 235492 673368 235544
rect 673420 235532 673426 235544
rect 673420 235504 674222 235532
rect 673420 235492 673426 235504
rect 674098 235124 674104 235136
rect 672552 235096 674104 235124
rect 672552 235000 672580 235096
rect 674098 235084 674104 235096
rect 674156 235084 674162 235136
rect 672534 234948 672540 235000
rect 672592 234948 672598 235000
rect 674324 234988 674352 235314
rect 673426 234960 674352 234988
rect 554406 234540 554412 234592
rect 554464 234580 554470 234592
rect 570598 234580 570604 234592
rect 554464 234552 570604 234580
rect 554464 234540 554470 234552
rect 570598 234540 570604 234552
rect 570656 234540 570662 234592
rect 668118 234540 668124 234592
rect 668176 234580 668182 234592
rect 673426 234580 673454 234960
rect 674190 234812 674196 234864
rect 674248 234852 674254 234864
rect 674438 234852 674466 235110
rect 674536 235000 674588 235006
rect 674536 234942 674588 234948
rect 674248 234824 674466 234852
rect 674248 234812 674254 234824
rect 668176 234552 673454 234580
rect 668176 234540 668182 234552
rect 669590 234336 669596 234388
rect 669648 234376 669654 234388
rect 674668 234376 674696 234702
rect 669648 234348 674696 234376
rect 669648 234336 669654 234348
rect 674760 234308 674788 234498
rect 675846 234336 675852 234388
rect 675904 234376 675910 234388
rect 680998 234376 681004 234388
rect 675904 234348 681004 234376
rect 675904 234336 675910 234348
rect 680998 234336 681004 234348
rect 681056 234336 681062 234388
rect 674744 234280 674788 234308
rect 673822 234200 673828 234252
rect 673880 234240 673886 234252
rect 674744 234240 674772 234280
rect 673880 234212 674772 234240
rect 673880 234200 673886 234212
rect 674898 234172 674926 234294
rect 674852 234144 674926 234172
rect 674852 234104 674880 234144
rect 674760 234076 674880 234104
rect 671706 233996 671712 234048
rect 671764 234036 671770 234048
rect 674760 234036 674788 234076
rect 671764 234008 674788 234036
rect 671764 233996 671770 234008
rect 674990 233968 675018 234090
rect 674898 233940 675018 233968
rect 670970 233860 670976 233912
rect 671028 233900 671034 233912
rect 674742 233900 674748 233912
rect 671028 233872 674748 233900
rect 671028 233860 671034 233872
rect 674742 233860 674748 233872
rect 674800 233860 674806 233912
rect 674898 233832 674926 233940
rect 675096 233912 675148 233918
rect 675096 233854 675148 233860
rect 675236 233912 675288 233918
rect 675236 233854 675288 233860
rect 674898 233804 675018 233832
rect 672948 233656 672954 233708
rect 673006 233696 673012 233708
rect 674834 233696 674840 233708
rect 673006 233668 674840 233696
rect 673006 233656 673012 233668
rect 674834 233656 674840 233668
rect 674892 233656 674898 233708
rect 674990 233628 675018 233804
rect 675846 233724 675852 233776
rect 675904 233764 675910 233776
rect 675904 233736 678974 233764
rect 675904 233724 675910 233736
rect 675110 233628 675116 233640
rect 674990 233600 675116 233628
rect 675110 233588 675116 233600
rect 675168 233588 675174 233640
rect 675846 233588 675852 233640
rect 675904 233628 675910 233640
rect 677686 233628 677692 233640
rect 675904 233600 677692 233628
rect 675904 233588 675910 233600
rect 677686 233588 677692 233600
rect 677744 233588 677750 233640
rect 670786 233316 670792 233368
rect 670844 233356 670850 233368
rect 675358 233356 675386 233478
rect 675846 233452 675852 233504
rect 675904 233492 675910 233504
rect 675904 233464 678100 233492
rect 675904 233452 675910 233464
rect 670844 233328 675386 233356
rect 670844 233316 670850 233328
rect 676030 233316 676036 233368
rect 676088 233356 676094 233368
rect 677870 233356 677876 233368
rect 676088 233328 677876 233356
rect 676088 233316 676094 233328
rect 677870 233316 677876 233328
rect 677928 233316 677934 233368
rect 678072 233288 678100 233464
rect 678946 233424 678974 233736
rect 683114 233424 683120 233436
rect 678946 233396 683120 233424
rect 683114 233384 683120 233396
rect 683172 233384 683178 233436
rect 684494 233288 684500 233300
rect 678072 233260 684500 233288
rect 684494 233248 684500 233260
rect 684552 233248 684558 233300
rect 672994 233180 673000 233232
rect 673052 233220 673058 233232
rect 673942 233220 673948 233232
rect 673052 233192 673948 233220
rect 673052 233180 673058 233192
rect 673942 233180 673948 233192
rect 674000 233180 674006 233232
rect 669038 232976 669044 233028
rect 669096 233016 669102 233028
rect 670234 233016 670240 233028
rect 669096 232988 670240 233016
rect 669096 232976 669102 232988
rect 670234 232976 670240 232988
rect 670292 232976 670298 233028
rect 669774 232840 669780 232892
rect 669832 232880 669838 232892
rect 673362 232880 673368 232892
rect 669832 232852 673368 232880
rect 669832 232840 669838 232852
rect 673362 232840 673368 232852
rect 673420 232840 673426 232892
rect 661862 232500 661868 232552
rect 661920 232540 661926 232552
rect 661920 232512 663794 232540
rect 661920 232500 661926 232512
rect 663766 232472 663794 232512
rect 675846 232500 675852 232552
rect 675904 232540 675910 232552
rect 683482 232540 683488 232552
rect 675904 232512 683488 232540
rect 675904 232500 675910 232512
rect 683482 232500 683488 232512
rect 683540 232500 683546 232552
rect 675478 232472 675484 232484
rect 663766 232444 675484 232472
rect 675478 232432 675484 232444
rect 675536 232432 675542 232484
rect 665082 232160 665088 232212
rect 665140 232200 665146 232212
rect 665140 232172 675556 232200
rect 665140 232160 665146 232172
rect 673454 231956 673460 232008
rect 673512 231996 673518 232008
rect 673512 231968 675372 231996
rect 673512 231956 673518 231968
rect 675180 231736 675232 231742
rect 675180 231678 675232 231684
rect 674166 231616 674172 231668
rect 674224 231656 674230 231668
rect 674466 231656 674472 231668
rect 674224 231628 674472 231656
rect 674224 231616 674230 231628
rect 674466 231616 674472 231628
rect 674524 231616 674530 231668
rect 675070 231532 675122 231538
rect 675070 231474 675122 231480
rect 674956 231328 675008 231334
rect 673454 231316 673460 231328
rect 663766 231288 673460 231316
rect 662230 231072 662236 231124
rect 662288 231112 662294 231124
rect 663766 231112 663794 231288
rect 673454 231276 673460 231288
rect 673512 231276 673518 231328
rect 674956 231270 675008 231276
rect 667934 231140 667940 231192
rect 667992 231180 667998 231192
rect 667992 231152 674866 231180
rect 667992 231140 667998 231152
rect 662288 231084 663794 231112
rect 662288 231072 662294 231084
rect 675846 231072 675852 231124
rect 675904 231112 675910 231124
rect 678606 231112 678612 231124
rect 675904 231084 678612 231112
rect 675904 231072 675910 231084
rect 678606 231072 678612 231084
rect 678664 231072 678670 231124
rect 674732 230920 674784 230926
rect 129642 230868 129648 230920
rect 129700 230908 129706 230920
rect 199102 230908 199108 230920
rect 129700 230880 199108 230908
rect 129700 230868 129706 230880
rect 199102 230868 199108 230880
rect 199160 230868 199166 230920
rect 674732 230862 674784 230868
rect 674466 230840 674472 230852
rect 674300 230812 674472 230840
rect 104802 230732 104808 230784
rect 104860 230772 104866 230784
rect 179138 230772 179144 230784
rect 104860 230744 179144 230772
rect 104860 230732 104866 230744
rect 179138 230732 179144 230744
rect 179196 230732 179202 230784
rect 97902 230596 97908 230648
rect 97960 230636 97966 230648
rect 173986 230636 173992 230648
rect 97960 230608 173992 230636
rect 97960 230596 97966 230608
rect 173986 230596 173992 230608
rect 174044 230596 174050 230648
rect 91002 230460 91008 230512
rect 91060 230500 91066 230512
rect 168834 230500 168840 230512
rect 91060 230472 168840 230500
rect 91060 230460 91066 230472
rect 168834 230460 168840 230472
rect 168892 230460 168898 230512
rect 511810 230460 511816 230512
rect 511868 230500 511874 230512
rect 511868 230472 512040 230500
rect 511868 230460 511874 230472
rect 196066 230392 196072 230444
rect 196124 230432 196130 230444
rect 198458 230432 198464 230444
rect 196124 230404 198464 230432
rect 196124 230392 196130 230404
rect 198458 230392 198464 230404
rect 198516 230392 198522 230444
rect 207658 230392 207664 230444
rect 207716 230432 207722 230444
rect 251266 230432 251272 230444
rect 207716 230404 251272 230432
rect 207716 230392 207722 230404
rect 251266 230392 251272 230404
rect 251324 230392 251330 230444
rect 256602 230392 256608 230444
rect 256660 230432 256666 230444
rect 297634 230432 297640 230444
rect 256660 230404 297640 230432
rect 256660 230392 256666 230404
rect 297634 230392 297640 230404
rect 297692 230392 297698 230444
rect 311894 230392 311900 230444
rect 311952 230432 311958 230444
rect 340138 230432 340144 230444
rect 311952 230404 340144 230432
rect 311952 230392 311958 230404
rect 340138 230392 340144 230404
rect 340196 230392 340202 230444
rect 441890 230392 441896 230444
rect 441948 230432 441954 230444
rect 443546 230432 443552 230444
rect 441948 230404 443552 230432
rect 441948 230392 441954 230404
rect 443546 230392 443552 230404
rect 443604 230392 443610 230444
rect 444466 230392 444472 230444
rect 444524 230432 444530 230444
rect 447594 230432 447600 230444
rect 444524 230404 447600 230432
rect 444524 230392 444530 230404
rect 447594 230392 447600 230404
rect 447652 230392 447658 230444
rect 476114 230392 476120 230444
rect 476172 230432 476178 230444
rect 478598 230432 478604 230444
rect 476172 230404 478604 230432
rect 476172 230392 476178 230404
rect 478598 230392 478604 230404
rect 478656 230392 478662 230444
rect 387426 230324 387432 230376
rect 387484 230364 387490 230376
rect 388438 230364 388444 230376
rect 387484 230336 388444 230364
rect 387484 230324 387490 230336
rect 388438 230324 388444 230336
rect 388496 230324 388502 230376
rect 439314 230324 439320 230376
rect 439372 230364 439378 230376
rect 440326 230364 440332 230376
rect 439372 230336 440332 230364
rect 439372 230324 439378 230336
rect 440326 230324 440332 230336
rect 440384 230324 440390 230376
rect 449618 230324 449624 230376
rect 449676 230364 449682 230376
rect 450538 230364 450544 230376
rect 449676 230336 450544 230364
rect 449676 230324 449682 230336
rect 450538 230324 450544 230336
rect 450596 230324 450602 230376
rect 451550 230324 451556 230376
rect 451608 230364 451614 230376
rect 453298 230364 453304 230376
rect 451608 230336 453304 230364
rect 451608 230324 451614 230336
rect 453298 230324 453304 230336
rect 453356 230324 453362 230376
rect 455414 230324 455420 230376
rect 455472 230364 455478 230376
rect 457162 230364 457168 230376
rect 455472 230336 457168 230364
rect 455472 230324 455478 230336
rect 457162 230324 457168 230336
rect 457220 230324 457226 230376
rect 463786 230324 463792 230376
rect 463844 230364 463850 230376
rect 465718 230364 465724 230376
rect 463844 230336 465724 230364
rect 463844 230324 463850 230336
rect 465718 230324 465724 230336
rect 465776 230324 465782 230376
rect 481818 230324 481824 230376
rect 481876 230364 481882 230376
rect 486510 230364 486516 230376
rect 481876 230336 486516 230364
rect 481876 230324 481882 230336
rect 486510 230324 486516 230336
rect 486568 230324 486574 230376
rect 503714 230324 503720 230376
rect 503772 230364 503778 230376
rect 507118 230364 507124 230376
rect 503772 230336 507124 230364
rect 503772 230324 503778 230336
rect 507118 230324 507124 230336
rect 507176 230324 507182 230376
rect 510798 230324 510804 230376
rect 510856 230364 510862 230376
rect 511810 230364 511816 230376
rect 510856 230336 511816 230364
rect 510856 230324 510862 230336
rect 511810 230324 511816 230336
rect 511868 230324 511874 230376
rect 133690 230256 133696 230308
rect 133748 230296 133754 230308
rect 202322 230296 202328 230308
rect 133748 230268 202328 230296
rect 133748 230256 133754 230268
rect 202322 230256 202328 230268
rect 202380 230256 202386 230308
rect 240962 230296 240968 230308
rect 209746 230268 240968 230296
rect 126882 230120 126888 230172
rect 126940 230160 126946 230172
rect 197170 230160 197176 230172
rect 126940 230132 197176 230160
rect 126940 230120 126946 230132
rect 197170 230120 197176 230132
rect 197228 230120 197234 230172
rect 197446 230120 197452 230172
rect 197504 230160 197510 230172
rect 201034 230160 201040 230172
rect 197504 230132 201040 230160
rect 197504 230120 197510 230132
rect 201034 230120 201040 230132
rect 201092 230120 201098 230172
rect 202138 230120 202144 230172
rect 202196 230160 202202 230172
rect 209746 230160 209774 230268
rect 240962 230256 240968 230268
rect 241020 230256 241026 230308
rect 242526 230256 242532 230308
rect 242584 230296 242590 230308
rect 287330 230296 287336 230308
rect 242584 230268 287336 230296
rect 242584 230256 242590 230268
rect 287330 230256 287336 230268
rect 287388 230256 287394 230308
rect 305638 230256 305644 230308
rect 305696 230296 305702 230308
rect 334986 230296 334992 230308
rect 305696 230268 334992 230296
rect 305696 230256 305702 230268
rect 334986 230256 334992 230268
rect 335044 230256 335050 230308
rect 376018 230256 376024 230308
rect 376076 230296 376082 230308
rect 380710 230296 380716 230308
rect 376076 230268 380716 230296
rect 376076 230256 376082 230268
rect 380710 230256 380716 230268
rect 380768 230256 380774 230308
rect 512012 230296 512040 230472
rect 531130 230460 531136 230512
rect 531188 230500 531194 230512
rect 531188 230472 531452 230500
rect 531188 230460 531194 230472
rect 526898 230392 526904 230444
rect 526956 230432 526962 230444
rect 526956 230404 528554 230432
rect 526956 230392 526962 230404
rect 520458 230324 520464 230376
rect 520516 230364 520522 230376
rect 521562 230364 521568 230376
rect 520516 230336 521568 230364
rect 520516 230324 520522 230336
rect 521562 230324 521568 230336
rect 521620 230324 521626 230376
rect 518894 230296 518900 230308
rect 512012 230268 518900 230296
rect 518894 230256 518900 230268
rect 518952 230256 518958 230308
rect 413830 230188 413836 230240
rect 413888 230228 413894 230240
rect 419994 230228 420000 230240
rect 413888 230200 420000 230228
rect 413888 230188 413894 230200
rect 419994 230188 420000 230200
rect 420052 230188 420058 230240
rect 443822 230188 443828 230240
rect 443880 230228 443886 230240
rect 444650 230228 444656 230240
rect 443880 230200 444656 230228
rect 443880 230188 443886 230200
rect 444650 230188 444656 230200
rect 444708 230188 444714 230240
rect 452838 230188 452844 230240
rect 452896 230228 452902 230240
rect 454310 230228 454316 230240
rect 452896 230200 454316 230228
rect 452896 230188 452902 230200
rect 454310 230188 454316 230200
rect 454368 230188 454374 230240
rect 465442 230188 465448 230240
rect 465500 230228 465506 230240
rect 469398 230228 469404 230240
rect 465500 230200 469404 230228
rect 465500 230188 465506 230200
rect 469398 230188 469404 230200
rect 469456 230188 469462 230240
rect 477954 230188 477960 230240
rect 478012 230228 478018 230240
rect 478782 230228 478788 230240
rect 478012 230200 478788 230228
rect 478012 230188 478018 230200
rect 478782 230188 478788 230200
rect 478840 230188 478846 230240
rect 499850 230188 499856 230240
rect 499908 230228 499914 230240
rect 504358 230228 504364 230240
rect 499908 230200 504364 230228
rect 499908 230188 499914 230200
rect 504358 230188 504364 230200
rect 504416 230188 504422 230240
rect 528526 230228 528554 230404
rect 530118 230324 530124 230376
rect 530176 230364 530182 230376
rect 531222 230364 531228 230376
rect 530176 230336 531228 230364
rect 530176 230324 530182 230336
rect 531222 230324 531228 230336
rect 531280 230324 531286 230376
rect 531424 230364 531452 230472
rect 674300 230432 674328 230812
rect 674466 230800 674472 230812
rect 674524 230800 674530 230852
rect 674610 230716 674662 230722
rect 674610 230658 674662 230664
rect 674390 230596 674396 230648
rect 674448 230636 674454 230648
rect 674448 230608 674544 230636
rect 674448 230596 674454 230608
rect 674208 230404 674328 230432
rect 531424 230336 535040 230364
rect 534810 230228 534816 230240
rect 528526 230200 534816 230228
rect 534810 230188 534816 230200
rect 534868 230188 534874 230240
rect 202196 230132 209774 230160
rect 202196 230120 202202 230132
rect 230474 230120 230480 230172
rect 230532 230160 230538 230172
rect 277026 230160 277032 230172
rect 230532 230132 277032 230160
rect 230532 230120 230538 230132
rect 277026 230120 277032 230132
rect 277084 230120 277090 230172
rect 294598 230120 294604 230172
rect 294656 230160 294662 230172
rect 323394 230160 323400 230172
rect 294656 230132 323400 230160
rect 294656 230120 294662 230132
rect 323394 230120 323400 230132
rect 323452 230120 323458 230172
rect 323578 230120 323584 230172
rect 323636 230160 323642 230172
rect 324682 230160 324688 230172
rect 323636 230132 324688 230160
rect 323636 230120 323642 230132
rect 324682 230120 324688 230132
rect 324740 230120 324746 230172
rect 354858 230120 354864 230172
rect 354916 230160 354922 230172
rect 371050 230160 371056 230172
rect 354916 230132 371056 230160
rect 354916 230120 354922 230132
rect 371050 230120 371056 230132
rect 371108 230120 371114 230172
rect 505646 230120 505652 230172
rect 505704 230160 505710 230172
rect 513834 230160 513840 230172
rect 505704 230132 513840 230160
rect 505704 230120 505710 230132
rect 513834 230120 513840 230132
rect 513892 230120 513898 230172
rect 515306 230120 515312 230172
rect 515364 230160 515370 230172
rect 525150 230160 525156 230172
rect 515364 230132 525156 230160
rect 515364 230120 515370 230132
rect 525150 230120 525156 230132
rect 525208 230120 525214 230172
rect 535012 230160 535040 230336
rect 535454 230256 535460 230308
rect 535512 230296 535518 230308
rect 539594 230296 539600 230308
rect 535512 230268 539600 230296
rect 535512 230256 535518 230268
rect 539594 230256 539600 230268
rect 539652 230256 539658 230308
rect 668118 230256 668124 230308
rect 668176 230296 668182 230308
rect 673822 230296 673828 230308
rect 668176 230268 673828 230296
rect 668176 230256 668182 230268
rect 673822 230256 673828 230268
rect 673880 230256 673886 230308
rect 674208 230228 674236 230404
rect 674396 230308 674448 230314
rect 674396 230250 674448 230256
rect 674208 230200 674314 230228
rect 543642 230160 543648 230172
rect 535012 230132 543648 230160
rect 543642 230120 543648 230132
rect 543700 230120 543706 230172
rect 454126 230052 454132 230104
rect 454184 230092 454190 230104
rect 455322 230092 455328 230104
rect 454184 230064 455328 230092
rect 454184 230052 454190 230064
rect 455322 230052 455328 230064
rect 455380 230052 455386 230104
rect 86218 229984 86224 230036
rect 86276 230024 86282 230036
rect 155954 230024 155960 230036
rect 86276 229996 155960 230024
rect 86276 229984 86282 229996
rect 155954 229984 155960 229996
rect 156012 229984 156018 230036
rect 160186 229984 160192 230036
rect 160244 230024 160250 230036
rect 220354 230024 220360 230036
rect 160244 229996 220360 230024
rect 160244 229984 160250 229996
rect 220354 229984 220360 229996
rect 220412 229984 220418 230036
rect 224954 229984 224960 230036
rect 225012 230024 225018 230036
rect 271874 230024 271880 230036
rect 225012 229996 271880 230024
rect 225012 229984 225018 229996
rect 271874 229984 271880 229996
rect 271932 229984 271938 230036
rect 300118 229984 300124 230036
rect 300176 230024 300182 230036
rect 329834 230024 329840 230036
rect 300176 229996 329840 230024
rect 300176 229984 300182 229996
rect 329834 229984 329840 229996
rect 329892 229984 329898 230036
rect 337838 229984 337844 230036
rect 337896 230024 337902 230036
rect 360746 230024 360752 230036
rect 337896 229996 360752 230024
rect 337896 229984 337902 229996
rect 360746 229984 360752 229996
rect 360804 229984 360810 230036
rect 457346 229984 457352 230036
rect 457404 230024 457410 230036
rect 464062 230024 464068 230036
rect 457404 229996 464068 230024
rect 457404 229984 457410 229996
rect 464062 229984 464068 229996
rect 464120 229984 464126 230036
rect 476666 229984 476672 230036
rect 476724 230024 476730 230036
rect 480714 230024 480720 230036
rect 476724 229996 480720 230024
rect 476724 229984 476730 229996
rect 480714 229984 480720 229996
rect 480772 229984 480778 230036
rect 501782 229984 501788 230036
rect 501840 230024 501846 230036
rect 509878 230024 509884 230036
rect 501840 229996 509884 230024
rect 501840 229984 501846 229996
rect 509878 229984 509884 229996
rect 509936 229984 509942 230036
rect 519170 229984 519176 230036
rect 519228 230024 519234 230036
rect 528554 230024 528560 230036
rect 519228 229996 528560 230024
rect 519228 229984 519234 229996
rect 528554 229984 528560 229996
rect 528612 229984 528618 230036
rect 534626 229984 534632 230036
rect 534684 230024 534690 230036
rect 552750 230024 552756 230036
rect 534684 229996 552756 230024
rect 534684 229984 534690 229996
rect 552750 229984 552756 229996
rect 552808 229984 552814 230036
rect 559558 229984 559564 230036
rect 559616 230024 559622 230036
rect 567194 230024 567200 230036
rect 559616 229996 567200 230024
rect 559616 229984 559622 229996
rect 567194 229984 567200 229996
rect 567252 229984 567258 230036
rect 672150 229984 672156 230036
rect 672208 230024 672214 230036
rect 672534 230024 672540 230036
rect 672208 229996 672540 230024
rect 672208 229984 672214 229996
rect 672534 229984 672540 229996
rect 672592 229984 672598 230036
rect 673270 229984 673276 230036
rect 673328 230024 673334 230036
rect 673328 229996 674198 230024
rect 673328 229984 673334 229996
rect 675846 229984 675852 230036
rect 675904 230024 675910 230036
rect 676490 230024 676496 230036
rect 675904 229996 676496 230024
rect 675904 229984 675910 229996
rect 676490 229984 676496 229996
rect 676548 229984 676554 230036
rect 453482 229916 453488 229968
rect 453540 229956 453546 229968
rect 455782 229956 455788 229968
rect 453540 229928 455788 229956
rect 453540 229916 453546 229928
rect 455782 229916 455788 229928
rect 455840 229916 455846 229968
rect 117222 229848 117228 229900
rect 117280 229888 117286 229900
rect 189442 229888 189448 229900
rect 117280 229860 189448 229888
rect 117280 229848 117286 229860
rect 189442 229848 189448 229860
rect 189500 229848 189506 229900
rect 189718 229848 189724 229900
rect 189776 229888 189782 229900
rect 235810 229888 235816 229900
rect 189776 229860 235816 229888
rect 189776 229848 189782 229860
rect 235810 229848 235816 229860
rect 235868 229848 235874 229900
rect 283558 229848 283564 229900
rect 283616 229888 283622 229900
rect 318242 229888 318248 229900
rect 283616 229860 318248 229888
rect 283616 229848 283622 229860
rect 318242 229848 318248 229860
rect 318300 229848 318306 229900
rect 324958 229848 324964 229900
rect 325016 229888 325022 229900
rect 350442 229888 350448 229900
rect 325016 229860 350448 229888
rect 325016 229848 325022 229860
rect 350442 229848 350448 229860
rect 350500 229848 350506 229900
rect 361206 229848 361212 229900
rect 361264 229888 361270 229900
rect 378778 229888 378784 229900
rect 361264 229860 378784 229888
rect 361264 229848 361270 229860
rect 378778 229848 378784 229860
rect 378836 229848 378842 229900
rect 389910 229848 389916 229900
rect 389968 229888 389974 229900
rect 399386 229888 399392 229900
rect 389968 229860 399392 229888
rect 389968 229848 389974 229860
rect 399386 229848 399392 229860
rect 399444 229848 399450 229900
rect 410794 229848 410800 229900
rect 410852 229888 410858 229900
rect 417418 229888 417424 229900
rect 410852 229860 417424 229888
rect 410852 229848 410858 229860
rect 417418 229848 417424 229860
rect 417476 229848 417482 229900
rect 479242 229848 479248 229900
rect 479300 229888 479306 229900
rect 490558 229888 490564 229900
rect 479300 229860 490564 229888
rect 479300 229848 479306 229860
rect 490558 229848 490564 229860
rect 490616 229848 490622 229900
rect 494054 229848 494060 229900
rect 494112 229888 494118 229900
rect 506106 229888 506112 229900
rect 494112 229860 506112 229888
rect 494112 229848 494118 229860
rect 506106 229848 506112 229860
rect 506164 229848 506170 229900
rect 517238 229848 517244 229900
rect 517296 229888 517302 229900
rect 525978 229888 525984 229900
rect 517296 229860 525984 229888
rect 517296 229848 517302 229860
rect 525978 229848 525984 229860
rect 526036 229848 526042 229900
rect 528830 229848 528836 229900
rect 528888 229888 528894 229900
rect 535454 229888 535460 229900
rect 528888 229860 535460 229888
rect 528888 229848 528894 229860
rect 535454 229848 535460 229860
rect 535512 229848 535518 229900
rect 536558 229848 536564 229900
rect 536616 229888 536622 229900
rect 559742 229888 559748 229900
rect 536616 229860 559748 229888
rect 536616 229848 536622 229860
rect 559742 229848 559748 229860
rect 559800 229848 559806 229900
rect 433518 229780 433524 229832
rect 433576 229820 433582 229832
rect 434162 229820 434168 229832
rect 433576 229792 434168 229820
rect 433576 229780 433582 229792
rect 434162 229780 434168 229792
rect 434220 229780 434226 229832
rect 438670 229780 438676 229832
rect 438728 229820 438734 229832
rect 439314 229820 439320 229832
rect 438728 229792 439320 229820
rect 438728 229780 438734 229792
rect 439314 229780 439320 229792
rect 439372 229780 439378 229832
rect 673822 229780 673828 229832
rect 673880 229820 673886 229832
rect 673880 229792 674084 229820
rect 673880 229780 673886 229792
rect 110322 229712 110328 229764
rect 110380 229752 110386 229764
rect 184290 229752 184296 229764
rect 110380 229724 184296 229752
rect 110380 229712 110386 229724
rect 184290 229712 184296 229724
rect 184348 229712 184354 229764
rect 184474 229712 184480 229764
rect 184532 229752 184538 229764
rect 225506 229752 225512 229764
rect 184532 229724 225512 229752
rect 184532 229712 184538 229724
rect 225506 229712 225512 229724
rect 225564 229712 225570 229764
rect 270126 229712 270132 229764
rect 270184 229752 270190 229764
rect 307938 229752 307944 229764
rect 270184 229724 307944 229752
rect 270184 229712 270190 229724
rect 307938 229712 307944 229724
rect 307996 229712 308002 229764
rect 318058 229712 318064 229764
rect 318116 229752 318122 229764
rect 345290 229752 345296 229764
rect 318116 229724 345296 229752
rect 318116 229712 318122 229724
rect 345290 229712 345296 229724
rect 345348 229712 345354 229764
rect 345658 229712 345664 229764
rect 345716 229752 345722 229764
rect 355594 229752 355600 229764
rect 345716 229724 355600 229752
rect 345716 229712 345722 229724
rect 355594 229712 355600 229724
rect 355652 229712 355658 229764
rect 357066 229712 357072 229764
rect 357124 229752 357130 229764
rect 376202 229752 376208 229764
rect 357124 229724 376208 229752
rect 357124 229712 357130 229724
rect 376202 229712 376208 229724
rect 376260 229712 376266 229764
rect 380710 229712 380716 229764
rect 380768 229752 380774 229764
rect 394234 229752 394240 229764
rect 380768 229724 394240 229752
rect 380768 229712 380774 229724
rect 394234 229712 394240 229724
rect 394292 229712 394298 229764
rect 399846 229712 399852 229764
rect 399904 229752 399910 229764
rect 409690 229752 409696 229764
rect 399904 229724 409696 229752
rect 399904 229712 399910 229724
rect 409690 229712 409696 229724
rect 409748 229712 409754 229764
rect 469582 229712 469588 229764
rect 469640 229752 469646 229764
rect 476758 229752 476764 229764
rect 469640 229724 476764 229752
rect 469640 229712 469646 229724
rect 476758 229712 476764 229724
rect 476816 229712 476822 229764
rect 484762 229712 484768 229764
rect 484820 229752 484826 229764
rect 496814 229752 496820 229764
rect 484820 229724 496820 229752
rect 484820 229712 484826 229724
rect 496814 229712 496820 229724
rect 496872 229712 496878 229764
rect 507578 229712 507584 229764
rect 507636 229752 507642 229764
rect 516778 229752 516784 229764
rect 507636 229724 516784 229752
rect 507636 229712 507642 229724
rect 516778 229712 516784 229724
rect 516836 229712 516842 229764
rect 523034 229712 523040 229764
rect 523092 229752 523098 229764
rect 534626 229752 534632 229764
rect 523092 229724 534632 229752
rect 523092 229712 523098 229724
rect 534626 229712 534632 229724
rect 534684 229712 534690 229764
rect 538490 229712 538496 229764
rect 538548 229752 538554 229764
rect 565078 229752 565084 229764
rect 538548 229724 565084 229752
rect 538548 229712 538554 229724
rect 565078 229712 565084 229724
rect 565136 229712 565142 229764
rect 95234 229576 95240 229628
rect 95292 229616 95298 229628
rect 161106 229616 161112 229628
rect 95292 229588 161112 229616
rect 95292 229576 95298 229588
rect 161106 229576 161112 229588
rect 161164 229576 161170 229628
rect 161290 229576 161296 229628
rect 161348 229616 161354 229628
rect 217778 229616 217784 229628
rect 161348 229588 217784 229616
rect 161348 229576 161354 229588
rect 217778 229576 217784 229588
rect 217836 229576 217842 229628
rect 251726 229576 251732 229628
rect 251784 229616 251790 229628
rect 292482 229616 292488 229628
rect 251784 229588 292488 229616
rect 251784 229576 251790 229588
rect 292482 229576 292488 229588
rect 292540 229576 292546 229628
rect 490190 229576 490196 229628
rect 490248 229616 490254 229628
rect 493962 229616 493968 229628
rect 490248 229588 493968 229616
rect 490248 229576 490254 229588
rect 493962 229576 493968 229588
rect 494020 229576 494026 229628
rect 513650 229576 513656 229628
rect 513708 229616 513714 229628
rect 522482 229616 522488 229628
rect 513708 229588 522488 229616
rect 513708 229576 513714 229588
rect 522482 229576 522488 229588
rect 522540 229576 522546 229628
rect 676030 229576 676036 229628
rect 676088 229616 676094 229628
rect 677410 229616 677416 229628
rect 676088 229588 677416 229616
rect 676088 229576 676094 229588
rect 677410 229576 677416 229588
rect 677468 229576 677474 229628
rect 673948 229560 674000 229566
rect 673948 229502 674000 229508
rect 144178 229440 144184 229492
rect 144236 229480 144242 229492
rect 148870 229480 148876 229492
rect 144236 229452 148876 229480
rect 144236 229440 144242 229452
rect 148870 229440 148876 229452
rect 148928 229440 148934 229492
rect 150434 229440 150440 229492
rect 150492 229480 150498 229492
rect 215202 229480 215208 229492
rect 150492 229452 215208 229480
rect 150492 229440 150498 229452
rect 215202 229440 215208 229452
rect 215260 229440 215266 229492
rect 217318 229440 217324 229492
rect 217376 229480 217382 229492
rect 266722 229480 266728 229492
rect 217376 229452 266728 229480
rect 217376 229440 217382 229452
rect 266722 229440 266728 229452
rect 266780 229440 266786 229492
rect 276658 229440 276664 229492
rect 276716 229480 276722 229492
rect 302786 229480 302792 229492
rect 276716 229452 302792 229480
rect 276716 229440 276722 229452
rect 302786 229440 302792 229452
rect 302844 229440 302850 229492
rect 673454 229440 673460 229492
rect 673512 229480 673518 229492
rect 673512 229452 673854 229480
rect 673512 229440 673518 229452
rect 675846 229440 675852 229492
rect 675904 229480 675910 229492
rect 676674 229480 676680 229492
rect 675904 229452 676680 229480
rect 675904 229440 675910 229452
rect 676674 229440 676680 229452
rect 676732 229440 676738 229492
rect 448974 229372 448980 229424
rect 449032 229412 449038 229424
rect 451366 229412 451372 229424
rect 449032 229384 451372 229412
rect 449032 229372 449038 229384
rect 451366 229372 451372 229384
rect 451424 229372 451430 229424
rect 509510 229372 509516 229424
rect 509568 229412 509574 229424
rect 518158 229412 518164 229424
rect 509568 229384 518164 229412
rect 509568 229372 509574 229384
rect 518158 229372 518164 229384
rect 518216 229372 518222 229424
rect 133874 229304 133880 229356
rect 133932 229344 133938 229356
rect 146294 229344 146300 229356
rect 133932 229316 146300 229344
rect 133932 229304 133938 229316
rect 146294 229304 146300 229316
rect 146352 229304 146358 229356
rect 148686 229304 148692 229356
rect 148744 229344 148750 229356
rect 210050 229344 210056 229356
rect 148744 229316 210056 229344
rect 148744 229304 148750 229316
rect 210050 229304 210056 229316
rect 210108 229304 210114 229356
rect 210418 229304 210424 229356
rect 210476 229344 210482 229356
rect 261294 229344 261300 229356
rect 210476 229316 261300 229344
rect 210476 229304 210482 229316
rect 261294 229304 261300 229316
rect 261352 229304 261358 229356
rect 261478 229304 261484 229356
rect 261536 229344 261542 229356
rect 282178 229344 282184 229356
rect 261536 229316 282184 229344
rect 261536 229304 261542 229316
rect 282178 229304 282184 229316
rect 282236 229304 282242 229356
rect 288710 229304 288716 229356
rect 288768 229344 288774 229356
rect 313090 229344 313096 229356
rect 288768 229316 313096 229344
rect 288768 229304 288774 229316
rect 313090 229304 313096 229316
rect 313148 229304 313154 229356
rect 450262 229236 450268 229288
rect 450320 229276 450326 229288
rect 451826 229276 451832 229288
rect 450320 229248 451832 229276
rect 450320 229236 450326 229248
rect 451826 229236 451832 229248
rect 451884 229236 451890 229288
rect 493410 229236 493416 229288
rect 493468 229276 493474 229288
rect 500218 229276 500224 229288
rect 493468 229248 500224 229276
rect 493468 229236 493474 229248
rect 500218 229236 500224 229248
rect 500276 229236 500282 229288
rect 532694 229236 532700 229288
rect 532752 229276 532758 229288
rect 536742 229276 536748 229288
rect 532752 229248 536748 229276
rect 532752 229236 532758 229248
rect 536742 229236 536748 229248
rect 536800 229236 536806 229288
rect 673454 229236 673460 229288
rect 673512 229276 673518 229288
rect 673512 229248 673762 229276
rect 673512 229236 673518 229248
rect 94498 229168 94504 229220
rect 94556 229208 94562 229220
rect 145650 229208 145656 229220
rect 94556 229180 145656 229208
rect 94556 229168 94562 229180
rect 145650 229168 145656 229180
rect 145708 229168 145714 229220
rect 146202 229168 146208 229220
rect 146260 229208 146266 229220
rect 207474 229208 207480 229220
rect 146260 229180 207480 229208
rect 146260 229168 146266 229180
rect 207474 229168 207480 229180
rect 207532 229168 207538 229220
rect 213086 229168 213092 229220
rect 213144 229208 213150 229220
rect 256418 229208 256424 229220
rect 213144 229180 256424 229208
rect 213144 229168 213150 229180
rect 256418 229168 256424 229180
rect 256476 229168 256482 229220
rect 419626 229100 419632 229152
rect 419684 229140 419690 229152
rect 421926 229140 421932 229152
rect 419684 229112 421932 229140
rect 419684 229100 419690 229112
rect 421926 229100 421932 229112
rect 421984 229100 421990 229152
rect 423490 229100 423496 229152
rect 423548 229140 423554 229152
rect 427722 229140 427728 229152
rect 423548 229112 427728 229140
rect 423548 229100 423554 229112
rect 427722 229100 427728 229112
rect 427780 229100 427786 229152
rect 441246 229100 441252 229152
rect 441304 229140 441310 229152
rect 442074 229140 442080 229152
rect 441304 229112 442080 229140
rect 441304 229100 441310 229112
rect 442074 229100 442080 229112
rect 442132 229100 442138 229152
rect 446398 229100 446404 229152
rect 446456 229140 446462 229152
rect 446456 229112 448560 229140
rect 446456 229100 446462 229112
rect 126422 229032 126428 229084
rect 126480 229072 126486 229084
rect 195238 229072 195244 229084
rect 126480 229044 195244 229072
rect 126480 229032 126486 229044
rect 195238 229032 195244 229044
rect 195296 229032 195302 229084
rect 205266 229032 205272 229084
rect 205324 229072 205330 229084
rect 257062 229072 257068 229084
rect 205324 229044 257068 229072
rect 205324 229032 205330 229044
rect 257062 229032 257068 229044
rect 257120 229032 257126 229084
rect 265618 229032 265624 229084
rect 265676 229072 265682 229084
rect 274450 229072 274456 229084
rect 265676 229044 274456 229072
rect 265676 229032 265682 229044
rect 274450 229032 274456 229044
rect 274508 229032 274514 229084
rect 274634 229032 274640 229084
rect 274692 229072 274698 229084
rect 309226 229072 309232 229084
rect 274692 229044 309232 229072
rect 274692 229032 274698 229044
rect 309226 229032 309232 229044
rect 309284 229032 309290 229084
rect 309686 229032 309692 229084
rect 309744 229072 309750 229084
rect 320818 229072 320824 229084
rect 309744 229044 320824 229072
rect 309744 229032 309750 229044
rect 320818 229032 320824 229044
rect 320876 229032 320882 229084
rect 327718 229032 327724 229084
rect 327776 229072 327782 229084
rect 337562 229072 337568 229084
rect 327776 229044 337568 229072
rect 327776 229032 327782 229044
rect 337562 229032 337568 229044
rect 337620 229032 337626 229084
rect 448532 229016 448560 229112
rect 450906 229100 450912 229152
rect 450964 229140 450970 229152
rect 452746 229140 452752 229152
rect 450964 229112 452752 229140
rect 450964 229100 450970 229112
rect 452746 229100 452752 229112
rect 452804 229100 452810 229152
rect 497918 229100 497924 229152
rect 497976 229140 497982 229152
rect 497976 229112 502334 229140
rect 497976 229100 497982 229112
rect 502306 229072 502334 229112
rect 524966 229100 524972 229152
rect 525024 229140 525030 229152
rect 525024 229112 529980 229140
rect 525024 229100 525030 229112
rect 514846 229072 514852 229084
rect 502306 229044 514852 229072
rect 514846 229032 514852 229044
rect 514904 229032 514910 229084
rect 448514 228964 448520 229016
rect 448572 228964 448578 229016
rect 119798 228896 119804 228948
rect 119856 228936 119862 228948
rect 190086 228936 190092 228948
rect 119856 228908 190092 228936
rect 119856 228896 119862 228908
rect 190086 228896 190092 228908
rect 190144 228896 190150 228948
rect 193122 228896 193128 228948
rect 193180 228936 193186 228948
rect 246758 228936 246764 228948
rect 193180 228908 246764 228936
rect 193180 228896 193186 228908
rect 246758 228896 246764 228908
rect 246816 228896 246822 228948
rect 257798 228896 257804 228948
rect 257856 228936 257862 228948
rect 299566 228936 299572 228948
rect 257856 228908 299572 228936
rect 257856 228896 257862 228908
rect 299566 228896 299572 228908
rect 299624 228896 299630 228948
rect 312906 228896 312912 228948
rect 312964 228936 312970 228948
rect 340782 228936 340788 228948
rect 312964 228908 340788 228936
rect 312964 228896 312970 228908
rect 340782 228896 340788 228908
rect 340840 228896 340846 228948
rect 349982 228896 349988 228948
rect 350040 228936 350046 228948
rect 369118 228936 369124 228948
rect 350040 228908 369124 228936
rect 350040 228896 350046 228908
rect 369118 228896 369124 228908
rect 369176 228896 369182 228948
rect 377950 228896 377956 228948
rect 378008 228936 378014 228948
rect 390370 228936 390376 228948
rect 378008 228908 390376 228936
rect 378008 228896 378014 228908
rect 390370 228896 390376 228908
rect 390428 228896 390434 228948
rect 529952 228936 529980 229112
rect 673598 228948 673650 228954
rect 549530 228936 549536 228948
rect 529952 228908 549536 228936
rect 549530 228896 549536 228908
rect 549588 228896 549594 228948
rect 673598 228890 673650 228896
rect 465994 228828 466000 228880
rect 466052 228868 466058 228880
rect 469858 228868 469864 228880
rect 466052 228840 469864 228868
rect 466052 228828 466058 228840
rect 469858 228828 469864 228840
rect 469916 228828 469922 228880
rect 673362 228828 673368 228880
rect 673420 228868 673426 228880
rect 673420 228840 673532 228868
rect 673420 228828 673426 228840
rect 100662 228760 100668 228812
rect 100720 228800 100726 228812
rect 174630 228800 174636 228812
rect 100720 228772 174636 228800
rect 100720 228760 100726 228772
rect 174630 228760 174636 228772
rect 174688 228760 174694 228812
rect 176470 228760 176476 228812
rect 176528 228800 176534 228812
rect 233878 228800 233884 228812
rect 176528 228772 233884 228800
rect 176528 228760 176534 228772
rect 233878 228760 233884 228772
rect 233936 228760 233942 228812
rect 234522 228760 234528 228812
rect 234580 228800 234586 228812
rect 278314 228800 278320 228812
rect 234580 228772 278320 228800
rect 234580 228760 234586 228772
rect 278314 228760 278320 228772
rect 278372 228760 278378 228812
rect 285582 228760 285588 228812
rect 285640 228800 285646 228812
rect 318886 228800 318892 228812
rect 285640 228772 318892 228800
rect 285640 228760 285646 228772
rect 318886 228760 318892 228772
rect 318944 228760 318950 228812
rect 320818 228760 320824 228812
rect 320876 228800 320882 228812
rect 327258 228800 327264 228812
rect 320876 228772 327264 228800
rect 320876 228760 320882 228772
rect 327258 228760 327264 228772
rect 327316 228760 327322 228812
rect 335078 228760 335084 228812
rect 335136 228800 335142 228812
rect 356882 228800 356888 228812
rect 335136 228772 356888 228800
rect 335136 228760 335142 228772
rect 356882 228760 356888 228772
rect 356940 228760 356946 228812
rect 373810 228760 373816 228812
rect 373868 228800 373874 228812
rect 387150 228800 387156 228812
rect 373868 228772 387156 228800
rect 373868 228760 373874 228772
rect 387150 228760 387156 228772
rect 387208 228760 387214 228812
rect 447042 228760 447048 228812
rect 447100 228800 447106 228812
rect 450170 228800 450176 228812
rect 447100 228772 450176 228800
rect 447100 228760 447106 228772
rect 450170 228760 450176 228772
rect 450228 228760 450234 228812
rect 518526 228760 518532 228812
rect 518584 228800 518590 228812
rect 541250 228800 541256 228812
rect 518584 228772 541256 228800
rect 518584 228760 518590 228772
rect 541250 228760 541256 228772
rect 541308 228760 541314 228812
rect 106182 228624 106188 228676
rect 106240 228664 106246 228676
rect 179782 228664 179788 228676
rect 106240 228636 179788 228664
rect 106240 228624 106246 228636
rect 179782 228624 179788 228636
rect 179840 228624 179846 228676
rect 183462 228624 183468 228676
rect 183520 228664 183526 228676
rect 239030 228664 239036 228676
rect 183520 228636 239036 228664
rect 183520 228624 183526 228636
rect 239030 228624 239036 228636
rect 239088 228624 239094 228676
rect 246298 228624 246304 228676
rect 246356 228664 246362 228676
rect 289262 228664 289268 228676
rect 246356 228636 289268 228664
rect 246356 228624 246362 228636
rect 289262 228624 289268 228636
rect 289320 228624 289326 228676
rect 304902 228624 304908 228676
rect 304960 228664 304966 228676
rect 333698 228664 333704 228676
rect 304960 228636 333704 228664
rect 304960 228624 304966 228636
rect 333698 228624 333704 228636
rect 333756 228624 333762 228676
rect 340138 228624 340144 228676
rect 340196 228664 340202 228676
rect 362678 228664 362684 228676
rect 340196 228636 362684 228664
rect 340196 228624 340202 228636
rect 362678 228624 362684 228636
rect 362736 228624 362742 228676
rect 371050 228624 371056 228676
rect 371108 228664 371114 228676
rect 385218 228664 385224 228676
rect 371108 228636 385224 228664
rect 371108 228624 371114 228636
rect 385218 228624 385224 228636
rect 385276 228624 385282 228676
rect 403986 228624 403992 228676
rect 404044 228664 404050 228676
rect 411070 228664 411076 228676
rect 404044 228636 411076 228664
rect 404044 228624 404050 228636
rect 411070 228624 411076 228636
rect 411128 228624 411134 228676
rect 485038 228624 485044 228676
rect 485096 228664 485102 228676
rect 498838 228664 498844 228676
rect 485096 228636 498844 228664
rect 485096 228624 485102 228636
rect 498838 228624 498844 228636
rect 498896 228624 498902 228676
rect 514018 228624 514024 228676
rect 514076 228664 514082 228676
rect 535730 228664 535736 228676
rect 514076 228636 535736 228664
rect 514076 228624 514082 228636
rect 535730 228624 535736 228636
rect 535788 228624 535794 228676
rect 535914 228624 535920 228676
rect 535972 228664 535978 228676
rect 563054 228664 563060 228676
rect 535972 228636 563060 228664
rect 535972 228624 535978 228636
rect 563054 228624 563060 228636
rect 563112 228624 563118 228676
rect 673388 228540 673440 228546
rect 93762 228488 93768 228540
rect 93820 228528 93826 228540
rect 169478 228528 169484 228540
rect 93820 228500 169484 228528
rect 93820 228488 93826 228500
rect 169478 228488 169484 228500
rect 169536 228488 169542 228540
rect 169938 228488 169944 228540
rect 169996 228528 170002 228540
rect 228726 228528 228732 228540
rect 169996 228500 228732 228528
rect 169996 228488 170002 228500
rect 228726 228488 228732 228500
rect 228784 228488 228790 228540
rect 235718 228488 235724 228540
rect 235776 228528 235782 228540
rect 280246 228528 280252 228540
rect 235776 228500 280252 228528
rect 235776 228488 235782 228500
rect 280246 228488 280252 228500
rect 280304 228488 280310 228540
rect 288342 228488 288348 228540
rect 288400 228528 288406 228540
rect 322750 228528 322756 228540
rect 288400 228500 322756 228528
rect 288400 228488 288406 228500
rect 322750 228488 322756 228500
rect 322808 228488 322814 228540
rect 326798 228488 326804 228540
rect 326856 228528 326862 228540
rect 351086 228528 351092 228540
rect 326856 228500 351092 228528
rect 326856 228488 326862 228500
rect 351086 228488 351092 228500
rect 351144 228488 351150 228540
rect 362586 228488 362592 228540
rect 362644 228528 362650 228540
rect 379422 228528 379428 228540
rect 362644 228500 379428 228528
rect 362644 228488 362650 228500
rect 379422 228488 379428 228500
rect 379480 228488 379486 228540
rect 390186 228488 390192 228540
rect 390244 228528 390250 228540
rect 400030 228528 400036 228540
rect 390244 228500 400036 228528
rect 390244 228488 390250 228500
rect 400030 228488 400036 228500
rect 400088 228488 400094 228540
rect 407758 228528 407764 228540
rect 402946 228500 407764 228528
rect 57238 228352 57244 228404
rect 57296 228392 57302 228404
rect 141142 228392 141148 228404
rect 57296 228364 141148 228392
rect 57296 228352 57302 228364
rect 141142 228352 141148 228364
rect 141200 228352 141206 228404
rect 146018 228352 146024 228404
rect 146076 228392 146082 228404
rect 210694 228392 210700 228404
rect 146076 228364 210700 228392
rect 146076 228352 146082 228364
rect 210694 228352 210700 228364
rect 210752 228352 210758 228404
rect 215018 228352 215024 228404
rect 215076 228392 215082 228404
rect 266078 228392 266084 228404
rect 215076 228364 266084 228392
rect 215076 228352 215082 228364
rect 266078 228352 266084 228364
rect 266136 228352 266142 228404
rect 271782 228352 271788 228404
rect 271840 228392 271846 228404
rect 308582 228392 308588 228404
rect 271840 228364 308588 228392
rect 271840 228352 271846 228364
rect 308582 228352 308588 228364
rect 308640 228352 308646 228404
rect 309042 228352 309048 228404
rect 309100 228392 309106 228404
rect 336274 228392 336280 228404
rect 309100 228364 336280 228392
rect 309100 228352 309106 228364
rect 336274 228352 336280 228364
rect 336332 228352 336338 228404
rect 336642 228352 336648 228404
rect 336700 228392 336706 228404
rect 358814 228392 358820 228404
rect 336700 228364 358820 228392
rect 336700 228352 336706 228364
rect 358814 228352 358820 228364
rect 358872 228352 358878 228404
rect 359918 228352 359924 228404
rect 359976 228392 359982 228404
rect 376846 228392 376852 228404
rect 359976 228364 376852 228392
rect 359976 228352 359982 228364
rect 376846 228352 376852 228364
rect 376904 228352 376910 228404
rect 378962 228352 378968 228404
rect 379020 228392 379026 228404
rect 393590 228392 393596 228404
rect 379020 228364 393596 228392
rect 379020 228352 379026 228364
rect 393590 228352 393596 228364
rect 393648 228352 393654 228404
rect 400030 228352 400036 228404
rect 400088 228392 400094 228404
rect 402946 228392 402974 228500
rect 407758 228488 407764 228500
rect 407816 228488 407822 228540
rect 411070 228488 411076 228540
rect 411128 228528 411134 228540
rect 416130 228528 416136 228540
rect 411128 228500 416136 228528
rect 411128 228488 411134 228500
rect 416130 228488 416136 228500
rect 416188 228488 416194 228540
rect 478966 228488 478972 228540
rect 479024 228528 479030 228540
rect 490742 228528 490748 228540
rect 479024 228500 490748 228528
rect 479024 228488 479030 228500
rect 490742 228488 490748 228500
rect 490800 228488 490806 228540
rect 491478 228488 491484 228540
rect 491536 228528 491542 228540
rect 506474 228528 506480 228540
rect 491536 228500 506480 228528
rect 491536 228488 491542 228500
rect 506474 228488 506480 228500
rect 506532 228488 506538 228540
rect 510154 228488 510160 228540
rect 510212 228528 510218 228540
rect 530946 228528 530952 228540
rect 510212 228500 530952 228528
rect 510212 228488 510218 228500
rect 530946 228488 530952 228500
rect 531004 228488 531010 228540
rect 531406 228488 531412 228540
rect 531464 228528 531470 228540
rect 558362 228528 558368 228540
rect 531464 228500 558368 228528
rect 531464 228488 531470 228500
rect 558362 228488 558368 228500
rect 558420 228488 558426 228540
rect 673388 228482 673440 228488
rect 400088 228364 402974 228392
rect 400088 228352 400094 228364
rect 409598 228352 409604 228404
rect 409656 228392 409662 228404
rect 415486 228392 415492 228404
rect 409656 228364 415492 228392
rect 409656 228352 409662 228364
rect 415486 228352 415492 228364
rect 415544 228352 415550 228404
rect 470226 228352 470232 228404
rect 470284 228392 470290 228404
rect 479518 228392 479524 228404
rect 470284 228364 479524 228392
rect 470284 228352 470290 228364
rect 479518 228352 479524 228364
rect 479576 228352 479582 228404
rect 486970 228352 486976 228404
rect 487028 228392 487034 228404
rect 501322 228392 501328 228404
rect 487028 228364 501328 228392
rect 487028 228352 487034 228364
rect 501322 228352 501328 228364
rect 501380 228352 501386 228404
rect 502426 228352 502432 228404
rect 502484 228392 502490 228404
rect 521286 228392 521292 228404
rect 502484 228364 521292 228392
rect 502484 228352 502490 228364
rect 521286 228352 521292 228364
rect 521344 228352 521350 228404
rect 521746 228352 521752 228404
rect 521804 228392 521810 228404
rect 545758 228392 545764 228404
rect 521804 228364 545764 228392
rect 521804 228352 521810 228364
rect 545758 228352 545764 228364
rect 545816 228352 545822 228404
rect 554038 228352 554044 228404
rect 554096 228392 554102 228404
rect 581638 228392 581644 228404
rect 554096 228364 581644 228392
rect 554096 228352 554102 228364
rect 581638 228352 581644 228364
rect 581696 228352 581702 228404
rect 673276 228336 673328 228342
rect 673276 228278 673328 228284
rect 133598 228216 133604 228268
rect 133656 228256 133662 228268
rect 200390 228256 200396 228268
rect 133656 228228 200396 228256
rect 133656 228216 133662 228228
rect 200390 228216 200396 228228
rect 200448 228216 200454 228268
rect 210878 228216 210884 228268
rect 210936 228256 210942 228268
rect 260282 228256 260288 228268
rect 210936 228228 260288 228256
rect 210936 228216 210942 228228
rect 260282 228216 260288 228228
rect 260340 228216 260346 228268
rect 398742 228216 398748 228268
rect 398800 228256 398806 228268
rect 409046 228256 409052 228268
rect 398800 228228 409052 228256
rect 398800 228216 398806 228228
rect 409046 228216 409052 228228
rect 409104 228216 409110 228268
rect 672920 228228 673190 228256
rect 139302 228080 139308 228132
rect 139360 228120 139366 228132
rect 205542 228120 205548 228132
rect 139360 228092 205548 228120
rect 139360 228080 139366 228092
rect 205542 228080 205548 228092
rect 205600 228080 205606 228132
rect 222010 228080 222016 228132
rect 222068 228120 222074 228132
rect 269942 228120 269948 228132
rect 222068 228092 269948 228120
rect 222068 228080 222074 228092
rect 269942 228080 269948 228092
rect 270000 228080 270006 228132
rect 672920 228120 672948 228228
rect 672828 228092 672948 228120
rect 140498 227944 140504 227996
rect 140556 227984 140562 227996
rect 146202 227984 146208 227996
rect 140556 227956 146208 227984
rect 140556 227944 140562 227956
rect 146202 227944 146208 227956
rect 146260 227944 146266 227996
rect 152918 227944 152924 227996
rect 152976 227984 152982 227996
rect 215846 227984 215852 227996
rect 152976 227956 215852 227984
rect 152976 227944 152982 227956
rect 215846 227944 215852 227956
rect 215904 227944 215910 227996
rect 252278 227944 252284 227996
rect 252336 227984 252342 227996
rect 293126 227984 293132 227996
rect 252336 227956 293132 227984
rect 252336 227944 252342 227956
rect 293126 227944 293132 227956
rect 293184 227944 293190 227996
rect 671154 227944 671160 227996
rect 671212 227984 671218 227996
rect 672828 227984 672856 228092
rect 673040 228080 673046 228132
rect 673098 228080 673104 228132
rect 671212 227956 672856 227984
rect 671212 227944 671218 227956
rect 393958 227876 393964 227928
rect 394016 227916 394022 227928
rect 401318 227916 401324 227928
rect 394016 227888 401324 227916
rect 394016 227876 394022 227888
rect 401318 227876 401324 227888
rect 401376 227876 401382 227928
rect 402238 227876 402244 227928
rect 402296 227916 402302 227928
rect 402296 227888 402974 227916
rect 402296 227876 402302 227888
rect 143166 227808 143172 227860
rect 143224 227848 143230 227860
rect 148686 227848 148692 227860
rect 143224 227820 148692 227848
rect 143224 227808 143230 227820
rect 148686 227808 148692 227820
rect 148744 227808 148750 227860
rect 169478 227808 169484 227860
rect 169536 227848 169542 227860
rect 169938 227848 169944 227860
rect 169536 227820 169944 227848
rect 169536 227808 169542 227820
rect 169938 227808 169944 227820
rect 169996 227808 170002 227860
rect 200666 227808 200672 227860
rect 200724 227848 200730 227860
rect 230658 227848 230664 227860
rect 200724 227820 230664 227848
rect 200724 227808 200730 227820
rect 230658 227808 230664 227820
rect 230716 227808 230722 227860
rect 280798 227808 280804 227860
rect 280856 227848 280862 227860
rect 284754 227848 284760 227860
rect 280856 227820 284760 227848
rect 280856 227808 280862 227820
rect 284754 227808 284760 227820
rect 284812 227808 284818 227860
rect 297358 227808 297364 227860
rect 297416 227848 297422 227860
rect 305362 227848 305368 227860
rect 297416 227820 305368 227848
rect 297416 227808 297422 227820
rect 305362 227808 305368 227820
rect 305420 227808 305426 227860
rect 396718 227740 396724 227792
rect 396776 227780 396782 227792
rect 397454 227780 397460 227792
rect 396776 227752 397460 227780
rect 396776 227740 396782 227752
rect 397454 227740 397460 227752
rect 397512 227740 397518 227792
rect 400858 227740 400864 227792
rect 400916 227780 400922 227792
rect 402606 227780 402612 227792
rect 400916 227752 402612 227780
rect 400916 227740 400922 227752
rect 402606 227740 402612 227752
rect 402664 227740 402670 227792
rect 402946 227780 402974 227888
rect 403250 227780 403256 227792
rect 402946 227752 403256 227780
rect 403250 227740 403256 227752
rect 403308 227740 403314 227792
rect 409138 227740 409144 227792
rect 409196 227780 409202 227792
rect 410334 227780 410340 227792
rect 409196 227752 410340 227780
rect 409196 227740 409202 227752
rect 410334 227740 410340 227752
rect 410392 227740 410398 227792
rect 411898 227740 411904 227792
rect 411956 227780 411962 227792
rect 413554 227780 413560 227792
rect 411956 227752 413560 227780
rect 411956 227740 411962 227752
rect 413554 227740 413560 227752
rect 413612 227740 413618 227792
rect 416682 227740 416688 227792
rect 416740 227780 416746 227792
rect 420638 227780 420644 227792
rect 416740 227752 420644 227780
rect 416740 227740 416746 227752
rect 420638 227740 420644 227752
rect 420696 227740 420702 227792
rect 474734 227740 474740 227792
rect 474792 227780 474798 227792
rect 482738 227780 482744 227792
rect 474792 227752 482744 227780
rect 474792 227740 474798 227752
rect 482738 227740 482744 227752
rect 482796 227740 482802 227792
rect 659562 227740 659568 227792
rect 659620 227780 659626 227792
rect 665266 227780 665272 227792
rect 659620 227752 665272 227780
rect 659620 227740 659626 227752
rect 665266 227740 665272 227752
rect 665324 227740 665330 227792
rect 672954 227724 673006 227730
rect 117038 227672 117044 227724
rect 117096 227712 117102 227724
rect 187510 227712 187516 227724
rect 117096 227684 187516 227712
rect 117096 227672 117102 227684
rect 187510 227672 187516 227684
rect 187568 227672 187574 227724
rect 200022 227672 200028 227724
rect 200080 227712 200086 227724
rect 252002 227712 252008 227724
rect 200080 227684 252008 227712
rect 200080 227672 200086 227684
rect 252002 227672 252008 227684
rect 252060 227672 252066 227724
rect 263410 227672 263416 227724
rect 263468 227712 263474 227724
rect 301498 227712 301504 227724
rect 263468 227684 301504 227712
rect 263468 227672 263474 227684
rect 301498 227672 301504 227684
rect 301556 227672 301562 227724
rect 516594 227672 516600 227724
rect 516652 227712 516658 227724
rect 538858 227712 538864 227724
rect 516652 227684 538864 227712
rect 516652 227672 516658 227684
rect 538858 227672 538864 227684
rect 538916 227672 538922 227724
rect 672954 227666 673006 227672
rect 671614 227604 671620 227656
rect 671672 227644 671678 227656
rect 671672 227616 672842 227644
rect 671672 227604 671678 227616
rect 109862 227536 109868 227588
rect 109920 227576 109926 227588
rect 182358 227576 182364 227588
rect 109920 227548 182364 227576
rect 109920 227536 109926 227548
rect 182358 227536 182364 227548
rect 182416 227536 182422 227588
rect 182818 227536 182824 227588
rect 182876 227576 182882 227588
rect 236454 227576 236460 227588
rect 182876 227548 236460 227576
rect 182876 227536 182882 227548
rect 236454 227536 236460 227548
rect 236512 227536 236518 227588
rect 242710 227536 242716 227588
rect 242768 227576 242774 227588
rect 285398 227576 285404 227588
rect 242768 227548 285404 227576
rect 242768 227536 242774 227548
rect 285398 227536 285404 227548
rect 285456 227536 285462 227588
rect 293678 227536 293684 227588
rect 293736 227576 293742 227588
rect 325326 227576 325332 227588
rect 293736 227548 325332 227576
rect 293736 227536 293742 227548
rect 325326 227536 325332 227548
rect 325384 227536 325390 227588
rect 512086 227536 512092 227588
rect 512144 227576 512150 227588
rect 533154 227576 533160 227588
rect 512144 227548 533160 227576
rect 512144 227536 512150 227548
rect 533154 227536 533160 227548
rect 533212 227536 533218 227588
rect 103238 227400 103244 227452
rect 103296 227440 103302 227452
rect 177206 227440 177212 227452
rect 103296 227412 177212 227440
rect 103296 227400 103302 227412
rect 177206 227400 177212 227412
rect 177264 227400 177270 227452
rect 185394 227400 185400 227452
rect 185452 227440 185458 227452
rect 192662 227440 192668 227452
rect 185452 227412 192668 227440
rect 185452 227400 185458 227412
rect 192662 227400 192668 227412
rect 192720 227400 192726 227452
rect 198458 227400 198464 227452
rect 198516 227440 198522 227452
rect 253198 227440 253204 227452
rect 198516 227412 253204 227440
rect 198516 227400 198522 227412
rect 253198 227400 253204 227412
rect 253256 227400 253262 227452
rect 259362 227400 259368 227452
rect 259420 227440 259426 227452
rect 298278 227440 298284 227452
rect 259420 227412 298284 227440
rect 259420 227400 259426 227412
rect 298278 227400 298284 227412
rect 298336 227400 298342 227452
rect 301958 227400 301964 227452
rect 302016 227440 302022 227452
rect 331122 227440 331128 227452
rect 302016 227412 331128 227440
rect 302016 227400 302022 227412
rect 331122 227400 331128 227412
rect 331180 227400 331186 227452
rect 333882 227400 333888 227452
rect 333940 227440 333946 227452
rect 356238 227440 356244 227452
rect 333940 227412 356244 227440
rect 333940 227400 333946 227412
rect 356238 227400 356244 227412
rect 356296 227400 356302 227452
rect 493962 227400 493968 227452
rect 494020 227440 494026 227452
rect 505646 227440 505652 227452
rect 494020 227412 505652 227440
rect 494020 227400 494026 227412
rect 505646 227400 505652 227412
rect 505704 227400 505710 227452
rect 521102 227400 521108 227452
rect 521160 227440 521166 227452
rect 544562 227440 544568 227452
rect 521160 227412 544568 227440
rect 521160 227400 521166 227412
rect 544562 227400 544568 227412
rect 544620 227400 544626 227452
rect 672166 227400 672172 227452
rect 672224 227440 672230 227452
rect 672224 227412 672750 227440
rect 672224 227400 672230 227412
rect 81342 227264 81348 227316
rect 81400 227304 81406 227316
rect 95234 227304 95240 227316
rect 81400 227276 95240 227304
rect 81400 227264 81406 227276
rect 95234 227264 95240 227276
rect 95292 227264 95298 227316
rect 96522 227264 96528 227316
rect 96580 227304 96586 227316
rect 172054 227304 172060 227316
rect 96580 227276 172060 227304
rect 96580 227264 96586 227276
rect 172054 227264 172060 227276
rect 172112 227264 172118 227316
rect 173158 227264 173164 227316
rect 173216 227304 173222 227316
rect 185578 227304 185584 227316
rect 173216 227276 185584 227304
rect 173216 227264 173222 227276
rect 185578 227264 185584 227276
rect 185636 227264 185642 227316
rect 188982 227264 188988 227316
rect 189040 227304 189046 227316
rect 244182 227304 244188 227316
rect 189040 227276 244188 227304
rect 189040 227264 189046 227276
rect 244182 227264 244188 227276
rect 244240 227264 244246 227316
rect 251082 227264 251088 227316
rect 251140 227304 251146 227316
rect 294414 227304 294420 227316
rect 251140 227276 294420 227304
rect 251140 227264 251146 227276
rect 294414 227264 294420 227276
rect 294472 227264 294478 227316
rect 308858 227264 308864 227316
rect 308916 227304 308922 227316
rect 339494 227304 339500 227316
rect 308916 227276 339500 227304
rect 308916 227264 308922 227276
rect 339494 227264 339500 227276
rect 339552 227264 339558 227316
rect 351178 227264 351184 227316
rect 351236 227304 351242 227316
rect 363322 227304 363328 227316
rect 351236 227276 363328 227304
rect 351236 227264 351242 227276
rect 363322 227264 363328 227276
rect 363380 227264 363386 227316
rect 363598 227264 363604 227316
rect 363656 227304 363662 227316
rect 368474 227304 368480 227316
rect 363656 227276 368480 227304
rect 363656 227264 363662 227276
rect 368474 227264 368480 227276
rect 368532 227264 368538 227316
rect 467650 227264 467656 227316
rect 467708 227304 467714 227316
rect 476574 227304 476580 227316
rect 467708 227276 476580 227304
rect 467708 227264 467714 227276
rect 476574 227264 476580 227276
rect 476632 227264 476638 227316
rect 481174 227264 481180 227316
rect 481232 227304 481238 227316
rect 492674 227304 492680 227316
rect 481232 227276 492680 227304
rect 481232 227264 481238 227276
rect 492674 227264 492680 227276
rect 492732 227264 492738 227316
rect 495342 227264 495348 227316
rect 495400 227304 495406 227316
rect 511442 227304 511448 227316
rect 495400 227276 511448 227304
rect 495400 227264 495406 227276
rect 511442 227264 511448 227276
rect 511500 227264 511506 227316
rect 528186 227264 528192 227316
rect 528244 227304 528250 227316
rect 553670 227304 553676 227316
rect 528244 227276 553676 227304
rect 528244 227264 528250 227276
rect 553670 227264 553676 227276
rect 553728 227264 553734 227316
rect 671798 227196 671804 227248
rect 671856 227236 671862 227248
rect 671856 227208 672630 227236
rect 671856 227196 671862 227208
rect 68186 227128 68192 227180
rect 68244 227168 68250 227180
rect 143718 227168 143724 227180
rect 68244 227140 143724 227168
rect 68244 227128 68250 227140
rect 143718 227128 143724 227140
rect 143776 227128 143782 227180
rect 156598 227128 156604 227180
rect 156656 227168 156662 227180
rect 213270 227168 213276 227180
rect 156656 227140 213276 227168
rect 156656 227128 156662 227140
rect 213270 227128 213276 227140
rect 213328 227128 213334 227180
rect 224770 227128 224776 227180
rect 224828 227168 224834 227180
rect 273806 227168 273812 227180
rect 224828 227140 273812 227168
rect 224828 227128 224834 227140
rect 273806 227128 273812 227140
rect 273864 227128 273870 227180
rect 274450 227128 274456 227180
rect 274508 227168 274514 227180
rect 312446 227168 312452 227180
rect 274508 227140 312452 227168
rect 274508 227128 274514 227140
rect 312446 227128 312452 227140
rect 312504 227128 312510 227180
rect 319806 227128 319812 227180
rect 319864 227168 319870 227180
rect 345842 227168 345848 227180
rect 319864 227140 345848 227168
rect 319864 227128 319870 227140
rect 345842 227128 345848 227140
rect 345900 227128 345906 227180
rect 346026 227128 346032 227180
rect 346084 227168 346090 227180
rect 366542 227168 366548 227180
rect 346084 227140 366548 227168
rect 346084 227128 346090 227140
rect 366542 227128 366548 227140
rect 366600 227128 366606 227180
rect 369762 227128 369768 227180
rect 369820 227168 369826 227180
rect 384574 227168 384580 227180
rect 369820 227140 384580 227168
rect 369820 227128 369826 227140
rect 384574 227128 384580 227140
rect 384632 227128 384638 227180
rect 391382 227128 391388 227180
rect 391440 227168 391446 227180
rect 400674 227168 400680 227180
rect 391440 227140 400680 227168
rect 391440 227128 391446 227140
rect 400674 227128 400680 227140
rect 400732 227128 400738 227180
rect 401318 227128 401324 227180
rect 401376 227168 401382 227180
rect 408402 227168 408408 227180
rect 401376 227140 408408 227168
rect 401376 227128 401382 227140
rect 408402 227128 408408 227140
rect 408460 227128 408466 227180
rect 474090 227128 474096 227180
rect 474148 227168 474154 227180
rect 484854 227168 484860 227180
rect 474148 227140 484860 227168
rect 474148 227128 474154 227140
rect 484854 227128 484860 227140
rect 484912 227128 484918 227180
rect 488902 227128 488908 227180
rect 488960 227168 488966 227180
rect 503254 227168 503260 227180
rect 488960 227140 503260 227168
rect 488960 227128 488966 227140
rect 503254 227128 503260 227140
rect 503312 227128 503318 227180
rect 506290 227128 506296 227180
rect 506348 227168 506354 227180
rect 526438 227168 526444 227180
rect 506348 227140 526444 227168
rect 506348 227128 506354 227140
rect 526438 227128 526444 227140
rect 526496 227128 526502 227180
rect 533338 227128 533344 227180
rect 533396 227168 533402 227180
rect 561306 227168 561312 227180
rect 533396 227140 561312 227168
rect 533396 227128 533402 227140
rect 561306 227128 561312 227140
rect 561364 227128 561370 227180
rect 56502 226992 56508 227044
rect 56560 227032 56566 227044
rect 142430 227032 142436 227044
rect 56560 227004 142436 227032
rect 56560 226992 56566 227004
rect 142430 226992 142436 227004
rect 142488 226992 142494 227044
rect 143350 226992 143356 227044
rect 143408 227032 143414 227044
rect 208118 227032 208124 227044
rect 143408 227004 208124 227032
rect 143408 226992 143414 227004
rect 208118 226992 208124 227004
rect 208176 226992 208182 227044
rect 226150 227032 226156 227044
rect 209746 227004 226156 227032
rect 122742 226856 122748 226908
rect 122800 226896 122806 226908
rect 185394 226896 185400 226908
rect 122800 226868 185400 226896
rect 122800 226856 122806 226868
rect 185394 226856 185400 226868
rect 185452 226856 185458 226908
rect 185578 226856 185584 226908
rect 185636 226896 185642 226908
rect 209746 226896 209774 227004
rect 226150 226992 226156 227004
rect 226208 226992 226214 227044
rect 228726 226992 228732 227044
rect 228784 227032 228790 227044
rect 275094 227032 275100 227044
rect 228784 227004 275100 227032
rect 228784 226992 228790 227004
rect 275094 226992 275100 227004
rect 275152 226992 275158 227044
rect 284938 226992 284944 227044
rect 284996 227032 285002 227044
rect 320174 227032 320180 227044
rect 284996 227004 320180 227032
rect 284996 226992 285002 227004
rect 320174 226992 320180 227004
rect 320232 226992 320238 227044
rect 325510 226992 325516 227044
rect 325568 227032 325574 227044
rect 349154 227032 349160 227044
rect 325568 227004 349160 227032
rect 325568 226992 325574 227004
rect 349154 226992 349160 227004
rect 349212 226992 349218 227044
rect 357250 226992 357256 227044
rect 357308 227032 357314 227044
rect 374270 227032 374276 227044
rect 357308 227004 374276 227032
rect 357308 226992 357314 227004
rect 374270 226992 374276 227004
rect 374328 226992 374334 227044
rect 376478 226992 376484 227044
rect 376536 227032 376542 227044
rect 389726 227032 389732 227044
rect 376536 227004 389732 227032
rect 376536 226992 376542 227004
rect 389726 226992 389732 227004
rect 389784 226992 389790 227044
rect 395706 226992 395712 227044
rect 395764 227032 395770 227044
rect 406470 227032 406476 227044
rect 395764 227004 406476 227032
rect 395764 226992 395770 227004
rect 406470 226992 406476 227004
rect 406528 226992 406534 227044
rect 412542 226992 412548 227044
rect 412600 227032 412606 227044
rect 419350 227032 419356 227044
rect 412600 227004 419356 227032
rect 412600 226992 412606 227004
rect 419350 226992 419356 227004
rect 419408 226992 419414 227044
rect 477310 226992 477316 227044
rect 477368 227032 477374 227044
rect 488994 227032 489000 227044
rect 477368 227004 489000 227032
rect 477368 226992 477374 227004
rect 488994 226992 489000 227004
rect 489052 226992 489058 227044
rect 499206 226992 499212 227044
rect 499264 227032 499270 227044
rect 516410 227032 516416 227044
rect 499264 227004 516416 227032
rect 499264 226992 499270 227004
rect 516410 226992 516416 227004
rect 516468 226992 516474 227044
rect 523678 226992 523684 227044
rect 523736 227032 523742 227044
rect 548518 227032 548524 227044
rect 523736 227004 548524 227032
rect 523736 226992 523742 227004
rect 548518 226992 548524 227004
rect 548576 226992 548582 227044
rect 555418 226992 555424 227044
rect 555476 227032 555482 227044
rect 633710 227032 633716 227044
rect 555476 227004 633716 227032
rect 555476 226992 555482 227004
rect 633710 226992 633716 227004
rect 633768 226992 633774 227044
rect 672258 226992 672264 227044
rect 672316 227032 672322 227044
rect 672316 227004 672520 227032
rect 672316 226992 672322 227004
rect 185636 226868 209774 226896
rect 185636 226856 185642 226868
rect 212350 226856 212356 226908
rect 212408 226896 212414 226908
rect 262214 226896 262220 226908
rect 212408 226868 262220 226896
rect 212408 226856 212414 226868
rect 262214 226856 262220 226868
rect 262272 226856 262278 226908
rect 275462 226856 275468 226908
rect 275520 226896 275526 226908
rect 311158 226896 311164 226908
rect 275520 226868 311164 226896
rect 275520 226856 275526 226868
rect 311158 226856 311164 226868
rect 311216 226856 311222 226908
rect 384758 226856 384764 226908
rect 384816 226896 384822 226908
rect 395522 226896 395528 226908
rect 384816 226868 395528 226896
rect 384816 226856 384822 226868
rect 395522 226856 395528 226868
rect 395580 226856 395586 226908
rect 419442 226856 419448 226908
rect 419500 226896 419506 226908
rect 424502 226896 424508 226908
rect 419500 226868 424508 226896
rect 419500 226856 419506 226868
rect 424502 226856 424508 226868
rect 424560 226856 424566 226908
rect 672258 226856 672264 226908
rect 672316 226896 672322 226908
rect 672316 226868 672406 226896
rect 672316 226856 672322 226868
rect 129458 226720 129464 226772
rect 129516 226760 129522 226772
rect 197814 226760 197820 226772
rect 129516 226732 197820 226760
rect 129516 226720 129522 226732
rect 197814 226720 197820 226732
rect 197872 226720 197878 226772
rect 224586 226720 224592 226772
rect 224644 226760 224650 226772
rect 270586 226760 270592 226772
rect 224644 226732 270592 226760
rect 224644 226720 224650 226732
rect 270586 226720 270592 226732
rect 270644 226720 270650 226772
rect 150066 226584 150072 226636
rect 150124 226624 150130 226636
rect 156598 226624 156604 226636
rect 150124 226596 156604 226624
rect 150124 226584 150130 226596
rect 156598 226584 156604 226596
rect 156656 226584 156662 226636
rect 160002 226584 160008 226636
rect 160060 226624 160066 226636
rect 220998 226624 221004 226636
rect 160060 226596 221004 226624
rect 160060 226584 160066 226596
rect 220998 226584 221004 226596
rect 221056 226584 221062 226636
rect 671798 226584 671804 226636
rect 671856 226624 671862 226636
rect 671856 226596 672290 226624
rect 671856 226584 671862 226596
rect 177298 226448 177304 226500
rect 177356 226488 177362 226500
rect 231302 226488 231308 226500
rect 177356 226460 231308 226488
rect 177356 226448 177362 226460
rect 231302 226448 231308 226460
rect 231360 226448 231366 226500
rect 670694 226448 670700 226500
rect 670752 226488 670758 226500
rect 670752 226460 672182 226488
rect 670752 226448 670758 226460
rect 385678 226312 385684 226364
rect 385736 226352 385742 226364
rect 391658 226352 391664 226364
rect 385736 226324 391664 226352
rect 385736 226312 385742 226324
rect 391658 226312 391664 226324
rect 391716 226312 391722 226364
rect 407758 226312 407764 226364
rect 407816 226352 407822 226364
rect 411622 226352 411628 226364
rect 407816 226324 411628 226352
rect 407816 226312 407822 226324
rect 411622 226312 411628 226324
rect 411680 226312 411686 226364
rect 63402 226244 63408 226296
rect 63460 226284 63466 226296
rect 133966 226284 133972 226296
rect 63460 226256 133972 226284
rect 63460 226244 63466 226256
rect 133966 226244 133972 226256
rect 134024 226244 134030 226296
rect 135162 226244 135168 226296
rect 135220 226284 135226 226296
rect 204254 226284 204260 226296
rect 135220 226256 204260 226284
rect 135220 226244 135226 226256
rect 204254 226244 204260 226256
rect 204312 226244 204318 226296
rect 219158 226244 219164 226296
rect 219216 226284 219222 226296
rect 267366 226284 267372 226296
rect 219216 226256 267372 226284
rect 219216 226244 219222 226256
rect 267366 226244 267372 226256
rect 267424 226244 267430 226296
rect 286962 226244 286968 226296
rect 287020 226284 287026 226296
rect 319530 226284 319536 226296
rect 287020 226256 319536 226284
rect 287020 226244 287026 226256
rect 319530 226244 319536 226256
rect 319588 226244 319594 226296
rect 518894 226244 518900 226296
rect 518952 226284 518958 226296
rect 531958 226284 531964 226296
rect 518952 226256 531964 226284
rect 518952 226244 518958 226256
rect 531958 226244 531964 226256
rect 532016 226244 532022 226296
rect 539778 226284 539784 226296
rect 533356 226256 539784 226284
rect 99098 226108 99104 226160
rect 99156 226148 99162 226160
rect 175918 226148 175924 226160
rect 99156 226120 175924 226148
rect 99156 226108 99162 226120
rect 175918 226108 175924 226120
rect 175976 226108 175982 226160
rect 205450 226108 205456 226160
rect 205508 226148 205514 226160
rect 258350 226148 258356 226160
rect 205508 226120 258356 226148
rect 205508 226108 205514 226120
rect 258350 226108 258356 226120
rect 258408 226108 258414 226160
rect 296622 226108 296628 226160
rect 296680 226148 296686 226160
rect 329190 226148 329196 226160
rect 296680 226120 329196 226148
rect 296680 226108 296686 226120
rect 329190 226108 329196 226120
rect 329248 226108 329254 226160
rect 330478 226108 330484 226160
rect 330536 226148 330542 226160
rect 351914 226148 351920 226160
rect 330536 226120 351920 226148
rect 330536 226108 330542 226120
rect 351914 226108 351920 226120
rect 351972 226108 351978 226160
rect 352558 226108 352564 226160
rect 352616 226148 352622 226160
rect 358170 226148 358176 226160
rect 352616 226120 358176 226148
rect 352616 226108 352622 226120
rect 358170 226108 358176 226120
rect 358228 226108 358234 226160
rect 501138 226108 501144 226160
rect 501196 226148 501202 226160
rect 519262 226148 519268 226160
rect 501196 226120 519268 226148
rect 501196 226108 501202 226120
rect 519262 226108 519268 226120
rect 519320 226108 519326 226160
rect 525978 226108 525984 226160
rect 526036 226148 526042 226160
rect 533356 226148 533384 226256
rect 539778 226244 539784 226256
rect 539836 226244 539842 226296
rect 671706 226244 671712 226296
rect 671764 226284 671770 226296
rect 671764 226256 672060 226284
rect 671764 226244 671770 226256
rect 540606 226148 540612 226160
rect 526036 226120 533384 226148
rect 538186 226120 540612 226148
rect 526036 226108 526042 226120
rect 84102 225972 84108 226024
rect 84160 226012 84166 226024
rect 161750 226012 161756 226024
rect 84160 225984 161756 226012
rect 84160 225972 84166 225984
rect 161750 225972 161756 225984
rect 161808 225972 161814 226024
rect 186038 225972 186044 226024
rect 186096 226012 186102 226024
rect 241606 226012 241612 226024
rect 186096 225984 241612 226012
rect 186096 225972 186102 225984
rect 241606 225972 241612 225984
rect 241664 225972 241670 226024
rect 255130 225972 255136 226024
rect 255188 226012 255194 226024
rect 296990 226012 296996 226024
rect 255188 225984 296996 226012
rect 255188 225972 255194 225984
rect 296990 225972 296996 225984
rect 297048 225972 297054 226024
rect 303246 225972 303252 226024
rect 303304 226012 303310 226024
rect 333054 226012 333060 226024
rect 303304 225984 333060 226012
rect 303304 225972 303310 225984
rect 333054 225972 333060 225984
rect 333112 225972 333118 226024
rect 480714 225972 480720 226024
rect 480772 226012 480778 226024
rect 487798 226012 487804 226024
rect 480772 225984 487804 226012
rect 480772 225972 480778 225984
rect 487798 225972 487804 225984
rect 487856 225972 487862 226024
rect 517882 225972 517888 226024
rect 517940 226012 517946 226024
rect 538186 226012 538214 226120
rect 540606 226108 540612 226120
rect 540664 226108 540670 226160
rect 671798 226040 671804 226092
rect 671856 226080 671862 226092
rect 671856 226052 671968 226080
rect 671856 226040 671862 226052
rect 517940 225984 538214 226012
rect 517940 225972 517946 225984
rect 539594 225972 539600 226024
rect 539652 226012 539658 226024
rect 555326 226012 555332 226024
rect 539652 225984 555332 226012
rect 539652 225972 539658 225984
rect 555326 225972 555332 225984
rect 555384 225972 555390 226024
rect 350350 225904 350356 225956
rect 350408 225944 350414 225956
rect 354858 225944 354864 225956
rect 350408 225916 354864 225944
rect 350408 225904 350414 225916
rect 354858 225904 354864 225916
rect 354916 225904 354922 225956
rect 70118 225836 70124 225888
rect 70176 225876 70182 225888
rect 151446 225876 151452 225888
rect 70176 225848 151452 225876
rect 70176 225836 70182 225848
rect 151446 225836 151452 225848
rect 151504 225836 151510 225888
rect 155770 225836 155776 225888
rect 155828 225876 155834 225888
rect 219710 225876 219716 225888
rect 155828 225848 219716 225876
rect 155828 225836 155834 225848
rect 219710 225836 219716 225848
rect 219768 225836 219774 225888
rect 220630 225836 220636 225888
rect 220688 225876 220694 225888
rect 268010 225876 268016 225888
rect 220688 225848 268016 225876
rect 220688 225836 220694 225848
rect 268010 225836 268016 225848
rect 268068 225836 268074 225888
rect 268838 225836 268844 225888
rect 268896 225876 268902 225888
rect 306006 225876 306012 225888
rect 268896 225848 306012 225876
rect 268896 225836 268902 225848
rect 306006 225836 306012 225848
rect 306064 225836 306070 225888
rect 319990 225836 319996 225888
rect 320048 225876 320054 225888
rect 347222 225876 347228 225888
rect 320048 225848 347228 225876
rect 320048 225836 320054 225848
rect 347222 225836 347228 225848
rect 347280 225836 347286 225888
rect 355318 225836 355324 225888
rect 355376 225876 355382 225888
rect 372338 225876 372344 225888
rect 355376 225848 372344 225876
rect 355376 225836 355382 225848
rect 372338 225836 372344 225848
rect 372396 225836 372402 225888
rect 388438 225836 388444 225888
rect 388496 225876 388502 225888
rect 396534 225876 396540 225888
rect 388496 225848 396540 225876
rect 388496 225836 388502 225848
rect 396534 225836 396540 225848
rect 396592 225836 396598 225888
rect 486510 225836 486516 225888
rect 486568 225876 486574 225888
rect 494790 225876 494796 225888
rect 486568 225848 494796 225876
rect 486568 225836 486574 225848
rect 494790 225836 494796 225848
rect 494848 225836 494854 225888
rect 495986 225836 495992 225888
rect 496044 225876 496050 225888
rect 512270 225876 512276 225888
rect 496044 225848 512276 225876
rect 496044 225836 496050 225848
rect 512270 225836 512276 225848
rect 512328 225836 512334 225888
rect 525610 225836 525616 225888
rect 525668 225876 525674 225888
rect 551002 225876 551008 225888
rect 525668 225848 551008 225876
rect 525668 225836 525674 225848
rect 551002 225836 551008 225848
rect 551060 225836 551066 225888
rect 458634 225768 458640 225820
rect 458692 225808 458698 225820
rect 462590 225808 462596 225820
rect 458692 225780 462596 225808
rect 458692 225768 458698 225780
rect 462590 225768 462596 225780
rect 462648 225768 462654 225820
rect 671820 225752 671872 225758
rect 59998 225700 60004 225752
rect 60056 225740 60062 225752
rect 141786 225740 141792 225752
rect 60056 225712 141792 225740
rect 60056 225700 60062 225712
rect 141786 225700 141792 225712
rect 141844 225700 141850 225752
rect 142062 225700 142068 225752
rect 142120 225740 142126 225752
rect 209406 225740 209412 225752
rect 142120 225712 209412 225740
rect 142120 225700 142126 225712
rect 209406 225700 209412 225712
rect 209464 225700 209470 225752
rect 209590 225700 209596 225752
rect 209648 225740 209654 225752
rect 259638 225740 259644 225752
rect 209648 225712 259644 225740
rect 209648 225700 209654 225712
rect 259638 225700 259644 225712
rect 259696 225700 259702 225752
rect 264698 225700 264704 225752
rect 264756 225740 264762 225752
rect 304718 225740 304724 225752
rect 264756 225712 304724 225740
rect 264756 225700 264762 225712
rect 304718 225700 304724 225712
rect 304776 225700 304782 225752
rect 306098 225700 306104 225752
rect 306156 225740 306162 225752
rect 336918 225740 336924 225752
rect 306156 225712 336924 225740
rect 306156 225700 306162 225712
rect 336918 225700 336924 225712
rect 336976 225700 336982 225752
rect 340690 225700 340696 225752
rect 340748 225740 340754 225752
rect 361482 225740 361488 225752
rect 340748 225712 361488 225740
rect 340748 225700 340754 225712
rect 361482 225700 361488 225712
rect 361540 225700 361546 225752
rect 365530 225700 365536 225752
rect 365588 225740 365594 225752
rect 380066 225740 380072 225752
rect 365588 225712 380072 225740
rect 365588 225700 365594 225712
rect 380066 225700 380072 225712
rect 380124 225700 380130 225752
rect 380250 225700 380256 225752
rect 380308 225740 380314 225752
rect 391014 225740 391020 225752
rect 380308 225712 391020 225740
rect 380308 225700 380314 225712
rect 391014 225700 391020 225712
rect 391072 225700 391078 225752
rect 472158 225700 472164 225752
rect 472216 225740 472222 225752
rect 480806 225740 480812 225752
rect 472216 225712 480812 225740
rect 472216 225700 472222 225712
rect 480806 225700 480812 225712
rect 480864 225700 480870 225752
rect 487982 225700 487988 225752
rect 488040 225740 488046 225752
rect 501506 225740 501512 225752
rect 488040 225712 501512 225740
rect 488040 225700 488046 225712
rect 501506 225700 501512 225712
rect 501564 225700 501570 225752
rect 505002 225700 505008 225752
rect 505060 225740 505066 225752
rect 524138 225740 524144 225752
rect 505060 225712 524144 225740
rect 505060 225700 505066 225712
rect 524138 225700 524144 225712
rect 524196 225700 524202 225752
rect 537846 225700 537852 225752
rect 537904 225740 537910 225752
rect 566090 225740 566096 225752
rect 537904 225712 566096 225740
rect 537904 225700 537910 225712
rect 566090 225700 566096 225712
rect 566148 225700 566154 225752
rect 671820 225694 671872 225700
rect 667934 225632 667940 225684
rect 667992 225672 667998 225684
rect 667992 225644 671738 225672
rect 667992 225632 667998 225644
rect 61838 225564 61844 225616
rect 61896 225604 61902 225616
rect 144362 225604 144368 225616
rect 61896 225576 144368 225604
rect 61896 225564 61902 225576
rect 144362 225564 144368 225576
rect 144420 225564 144426 225616
rect 158438 225564 158444 225616
rect 158496 225604 158502 225616
rect 222286 225604 222292 225616
rect 158496 225576 222292 225604
rect 158496 225564 158502 225576
rect 222286 225564 222292 225576
rect 222344 225564 222350 225616
rect 239398 225564 239404 225616
rect 239456 225604 239462 225616
rect 284110 225604 284116 225616
rect 239456 225576 284116 225604
rect 239456 225564 239462 225576
rect 284110 225564 284116 225576
rect 284168 225564 284174 225616
rect 288158 225564 288164 225616
rect 288216 225604 288222 225616
rect 321462 225604 321468 225616
rect 288216 225576 321468 225604
rect 288216 225564 288222 225576
rect 321462 225564 321468 225576
rect 321520 225564 321526 225616
rect 324038 225564 324044 225616
rect 324096 225604 324102 225616
rect 348510 225604 348516 225616
rect 324096 225576 348516 225604
rect 324096 225564 324102 225576
rect 348510 225564 348516 225576
rect 348568 225564 348574 225616
rect 349062 225564 349068 225616
rect 349120 225604 349126 225616
rect 367186 225604 367192 225616
rect 349120 225576 367192 225604
rect 349120 225564 349126 225576
rect 367186 225564 367192 225576
rect 367244 225564 367250 225616
rect 375282 225564 375288 225616
rect 375340 225604 375346 225616
rect 387794 225604 387800 225616
rect 375340 225576 387800 225604
rect 375340 225564 375346 225576
rect 387794 225564 387800 225576
rect 387852 225564 387858 225616
rect 391750 225564 391756 225616
rect 391808 225604 391814 225616
rect 403526 225604 403532 225616
rect 391808 225576 403532 225604
rect 391808 225564 391814 225576
rect 403526 225564 403532 225576
rect 403584 225564 403590 225616
rect 469398 225564 469404 225616
rect 469456 225604 469462 225616
rect 473538 225604 473544 225616
rect 469456 225576 473544 225604
rect 469456 225564 469462 225576
rect 473538 225564 473544 225576
rect 473596 225564 473602 225616
rect 478598 225564 478604 225616
rect 478656 225604 478662 225616
rect 485866 225604 485872 225616
rect 478656 225576 485872 225604
rect 478656 225564 478662 225576
rect 485866 225564 485872 225576
rect 485924 225564 485930 225616
rect 491294 225564 491300 225616
rect 491352 225604 491358 225616
rect 505922 225604 505928 225616
rect 491352 225576 505928 225604
rect 491352 225564 491358 225576
rect 505922 225564 505928 225576
rect 505980 225564 505986 225616
rect 508222 225564 508228 225616
rect 508280 225604 508286 225616
rect 527358 225604 527364 225616
rect 508280 225576 527364 225604
rect 508280 225564 508286 225576
rect 527358 225564 527364 225576
rect 527416 225564 527422 225616
rect 535270 225564 535276 225616
rect 535328 225604 535334 225616
rect 563514 225604 563520 225616
rect 535328 225576 563520 225604
rect 535328 225564 535334 225576
rect 563514 225564 563520 225576
rect 563572 225564 563578 225616
rect 132218 225428 132224 225480
rect 132276 225468 132282 225480
rect 201678 225468 201684 225480
rect 132276 225440 201684 225468
rect 132276 225428 132282 225440
rect 201678 225428 201684 225440
rect 201736 225428 201742 225480
rect 202598 225428 202604 225480
rect 202656 225468 202662 225480
rect 254486 225468 254492 225480
rect 202656 225440 254492 225468
rect 202656 225428 202662 225440
rect 254486 225428 254492 225440
rect 254544 225428 254550 225480
rect 254946 225428 254952 225480
rect 255004 225468 255010 225480
rect 295702 225468 295708 225480
rect 255004 225440 295708 225468
rect 255004 225428 255010 225440
rect 295702 225428 295708 225440
rect 295760 225428 295766 225480
rect 670694 225428 670700 225480
rect 670752 225468 670758 225480
rect 670752 225440 671622 225468
rect 670752 225428 670758 225440
rect 506106 225360 506112 225412
rect 506164 225400 506170 225412
rect 510338 225400 510344 225412
rect 506164 225372 510344 225400
rect 506164 225360 506170 225372
rect 510338 225360 510344 225372
rect 510396 225360 510402 225412
rect 138842 225292 138848 225344
rect 138900 225332 138906 225344
rect 206370 225332 206376 225344
rect 138900 225304 206376 225332
rect 138900 225292 138906 225304
rect 206370 225292 206376 225304
rect 206428 225292 206434 225344
rect 206554 225292 206560 225344
rect 206612 225332 206618 225344
rect 228082 225332 228088 225344
rect 206612 225304 228088 225332
rect 206612 225292 206618 225304
rect 228082 225292 228088 225304
rect 228140 225292 228146 225344
rect 245562 225292 245568 225344
rect 245620 225332 245626 225344
rect 287974 225332 287980 225344
rect 245620 225304 287980 225332
rect 245620 225292 245626 225304
rect 287974 225292 287980 225304
rect 288032 225292 288038 225344
rect 463142 225224 463148 225276
rect 463200 225264 463206 225276
rect 467098 225264 467104 225276
rect 463200 225236 467104 225264
rect 463200 225224 463206 225236
rect 467098 225224 467104 225236
rect 467156 225224 467162 225276
rect 671154 225224 671160 225276
rect 671212 225264 671218 225276
rect 671212 225236 671508 225264
rect 671212 225224 671218 225236
rect 155586 225156 155592 225208
rect 155644 225196 155650 225208
rect 218422 225196 218428 225208
rect 155644 225168 218428 225196
rect 155644 225156 155650 225168
rect 218422 225156 218428 225168
rect 218480 225156 218486 225208
rect 225506 225156 225512 225208
rect 225564 225196 225570 225208
rect 246114 225196 246120 225208
rect 225564 225168 246120 225196
rect 225564 225156 225570 225168
rect 246114 225156 246120 225168
rect 246172 225156 246178 225208
rect 166074 225020 166080 225072
rect 166132 225060 166138 225072
rect 186866 225060 186872 225072
rect 166132 225032 186872 225060
rect 166132 225020 166138 225032
rect 186866 225020 186872 225032
rect 186924 225020 186930 225072
rect 195882 225020 195888 225072
rect 195940 225060 195946 225072
rect 249334 225060 249340 225072
rect 195940 225032 249340 225060
rect 195940 225020 195946 225032
rect 249334 225020 249340 225032
rect 249392 225020 249398 225072
rect 670694 225020 670700 225072
rect 670752 225060 670758 225072
rect 670752 225032 671398 225060
rect 670752 225020 670758 225032
rect 260098 224952 260104 225004
rect 260156 224992 260162 225004
rect 264146 224992 264152 225004
rect 260156 224964 264152 224992
rect 260156 224952 260162 224964
rect 264146 224952 264152 224964
rect 264204 224952 264210 225004
rect 367738 224952 367744 225004
rect 367796 224992 367802 225004
rect 373626 224992 373632 225004
rect 367796 224964 373632 224992
rect 367796 224952 367802 224964
rect 373626 224952 373632 224964
rect 373684 224952 373690 225004
rect 404170 224952 404176 225004
rect 404228 224992 404234 225004
rect 412266 224992 412272 225004
rect 404228 224964 412272 224992
rect 404228 224952 404234 224964
rect 412266 224952 412272 224964
rect 412324 224952 412330 225004
rect 529842 224952 529848 225004
rect 529900 224992 529906 225004
rect 619634 224992 619640 225004
rect 529900 224964 619640 224992
rect 529900 224952 529906 224964
rect 619634 224952 619640 224964
rect 619692 224952 619698 225004
rect 118602 224884 118608 224936
rect 118660 224924 118666 224936
rect 185578 224924 185584 224936
rect 118660 224896 185584 224924
rect 118660 224884 118666 224896
rect 185578 224884 185584 224896
rect 185636 224884 185642 224936
rect 191466 224884 191472 224936
rect 191524 224924 191530 224936
rect 248046 224924 248052 224936
rect 191524 224896 248052 224924
rect 191524 224884 191530 224896
rect 248046 224884 248052 224896
rect 248104 224884 248110 224936
rect 266262 224884 266268 224936
rect 266320 224924 266326 224936
rect 303430 224924 303436 224936
rect 266320 224896 303436 224924
rect 266320 224884 266326 224896
rect 303430 224884 303436 224896
rect 303488 224884 303494 224936
rect 321462 224884 321468 224936
rect 321520 224924 321526 224936
rect 346578 224924 346584 224936
rect 321520 224896 346584 224924
rect 321520 224884 321526 224896
rect 346578 224884 346584 224896
rect 346636 224884 346642 224936
rect 426434 224884 426440 224936
rect 426492 224924 426498 224936
rect 426986 224924 426992 224936
rect 426492 224896 426992 224924
rect 426492 224884 426498 224896
rect 426986 224884 426992 224896
rect 427044 224884 427050 224936
rect 466362 224816 466368 224868
rect 466420 224856 466426 224868
rect 471238 224856 471244 224868
rect 466420 224828 471244 224856
rect 466420 224816 466426 224828
rect 471238 224816 471244 224828
rect 471296 224816 471302 224868
rect 669038 224816 669044 224868
rect 669096 224856 669102 224868
rect 669096 224828 671278 224856
rect 669096 224816 669102 224828
rect 112898 224748 112904 224800
rect 112956 224788 112962 224800
rect 185854 224788 185860 224800
rect 112956 224760 185860 224788
rect 112956 224748 112962 224760
rect 185854 224748 185860 224760
rect 185912 224748 185918 224800
rect 242894 224788 242900 224800
rect 186148 224760 242900 224788
rect 105722 224612 105728 224664
rect 105780 224652 105786 224664
rect 181070 224652 181076 224664
rect 105780 224624 181076 224652
rect 105780 224612 105786 224624
rect 181070 224612 181076 224624
rect 181128 224612 181134 224664
rect 185762 224612 185768 224664
rect 185820 224652 185826 224664
rect 186148 224652 186176 224760
rect 242894 224748 242900 224760
rect 242952 224748 242958 224800
rect 271322 224748 271328 224800
rect 271380 224788 271386 224800
rect 309870 224788 309876 224800
rect 271380 224760 309876 224788
rect 271380 224748 271386 224760
rect 309870 224748 309876 224760
rect 309928 224748 309934 224800
rect 313090 224748 313096 224800
rect 313148 224788 313154 224800
rect 342070 224788 342076 224800
rect 313148 224760 342076 224788
rect 313148 224748 313154 224760
rect 342070 224748 342076 224760
rect 342128 224748 342134 224800
rect 365898 224788 365904 224800
rect 354646 224760 365904 224788
rect 185820 224624 186176 224652
rect 185820 224612 185826 224624
rect 186314 224612 186320 224664
rect 186372 224652 186378 224664
rect 240318 224652 240324 224664
rect 186372 224624 240324 224652
rect 186372 224612 186378 224624
rect 240318 224612 240324 224624
rect 240376 224612 240382 224664
rect 249610 224612 249616 224664
rect 249668 224652 249674 224664
rect 290550 224652 290556 224664
rect 249668 224624 290556 224652
rect 249668 224612 249674 224624
rect 290550 224612 290556 224624
rect 290608 224612 290614 224664
rect 295150 224612 295156 224664
rect 295208 224652 295214 224664
rect 325970 224652 325976 224664
rect 295208 224624 325976 224652
rect 295208 224612 295214 224624
rect 325970 224612 325976 224624
rect 326028 224612 326034 224664
rect 347038 224612 347044 224664
rect 347096 224652 347102 224664
rect 354646 224652 354674 224760
rect 365898 224748 365904 224760
rect 365956 224748 365962 224800
rect 534626 224748 534632 224800
rect 534684 224788 534690 224800
rect 547414 224788 547420 224800
rect 534684 224760 547420 224788
rect 534684 224748 534690 224760
rect 547414 224748 547420 224760
rect 547472 224748 547478 224800
rect 551830 224748 551836 224800
rect 551888 224788 551894 224800
rect 558178 224788 558184 224800
rect 551888 224760 558184 224788
rect 551888 224748 551894 224760
rect 558178 224748 558184 224760
rect 558236 224748 558242 224800
rect 558362 224748 558368 224800
rect 558420 224788 558426 224800
rect 562042 224788 562048 224800
rect 558420 224760 562048 224788
rect 558420 224748 558426 224760
rect 562042 224748 562048 224760
rect 562100 224748 562106 224800
rect 363966 224652 363972 224664
rect 347096 224624 354674 224652
rect 359292 224624 363972 224652
rect 347096 224612 347102 224624
rect 85482 224476 85488 224528
rect 85540 224516 85546 224528
rect 165614 224516 165620 224528
rect 85540 224488 165620 224516
rect 85540 224476 85546 224488
rect 165614 224476 165620 224488
rect 165672 224476 165678 224528
rect 172330 224476 172336 224528
rect 172388 224516 172394 224528
rect 232590 224516 232596 224528
rect 172388 224488 232596 224516
rect 172388 224476 172394 224488
rect 232590 224476 232596 224488
rect 232648 224476 232654 224528
rect 233142 224476 233148 224528
rect 233200 224516 233206 224528
rect 277670 224516 277676 224528
rect 233200 224488 277676 224516
rect 233200 224476 233206 224488
rect 277670 224476 277676 224488
rect 277728 224476 277734 224528
rect 282546 224476 282552 224528
rect 282604 224516 282610 224528
rect 316310 224516 316316 224528
rect 282604 224488 316316 224516
rect 282604 224476 282610 224488
rect 316310 224476 316316 224488
rect 316368 224476 316374 224528
rect 316862 224476 316868 224528
rect 316920 224516 316926 224528
rect 342990 224516 342996 224528
rect 316920 224488 342996 224516
rect 316920 224476 316926 224488
rect 342990 224476 342996 224488
rect 343048 224476 343054 224528
rect 343358 224476 343364 224528
rect 343416 224516 343422 224528
rect 359292 224516 359320 224624
rect 363966 224612 363972 224624
rect 364024 224612 364030 224664
rect 493042 224612 493048 224664
rect 493100 224652 493106 224664
rect 508590 224652 508596 224664
rect 493100 224624 508596 224652
rect 493100 224612 493106 224624
rect 508590 224612 508596 224624
rect 508648 224652 508654 224664
rect 598382 224652 598388 224664
rect 508648 224624 598388 224652
rect 508648 224612 508654 224624
rect 598382 224612 598388 224624
rect 598440 224612 598446 224664
rect 670878 224612 670884 224664
rect 670936 224652 670942 224664
rect 670936 224624 671186 224652
rect 670936 224612 670942 224624
rect 343416 224488 359320 224516
rect 343416 224476 343422 224488
rect 363782 224476 363788 224528
rect 363840 224516 363846 224528
rect 378134 224516 378140 224528
rect 363840 224488 378140 224516
rect 363840 224476 363846 224488
rect 378134 224476 378140 224488
rect 378192 224476 378198 224528
rect 394510 224476 394516 224528
rect 394568 224516 394574 224528
rect 404538 224516 404544 224528
rect 394568 224488 404544 224516
rect 394568 224476 394574 224488
rect 404538 224476 404544 224488
rect 404596 224476 404602 224528
rect 506934 224476 506940 224528
rect 506992 224516 506998 224528
rect 525794 224516 525800 224528
rect 506992 224488 525800 224516
rect 506992 224476 506998 224488
rect 525794 224476 525800 224488
rect 525852 224476 525858 224528
rect 526254 224476 526260 224528
rect 526312 224516 526318 224528
rect 551278 224516 551284 224528
rect 526312 224488 551284 224516
rect 526312 224476 526318 224488
rect 551278 224476 551284 224488
rect 551336 224476 551342 224528
rect 552750 224476 552756 224528
rect 552808 224516 552814 224528
rect 557994 224516 558000 224528
rect 552808 224488 558000 224516
rect 552808 224476 552814 224488
rect 557994 224476 558000 224488
rect 558052 224476 558058 224528
rect 558178 224476 558184 224528
rect 558236 224516 558242 224528
rect 625246 224516 625252 224528
rect 558236 224488 625252 224516
rect 558236 224476 558242 224488
rect 625246 224476 625252 224488
rect 625304 224476 625310 224528
rect 670804 224420 671048 224448
rect 76558 224340 76564 224392
rect 76616 224380 76622 224392
rect 157794 224380 157800 224392
rect 76616 224352 157800 224380
rect 76616 224340 76622 224352
rect 157794 224340 157800 224352
rect 157852 224340 157858 224392
rect 165338 224340 165344 224392
rect 165396 224380 165402 224392
rect 227438 224380 227444 224392
rect 165396 224352 227444 224380
rect 165396 224340 165402 224352
rect 227438 224340 227444 224352
rect 227496 224340 227502 224392
rect 241238 224340 241244 224392
rect 241296 224380 241302 224392
rect 286686 224380 286692 224392
rect 241296 224352 286692 224380
rect 241296 224340 241302 224352
rect 286686 224340 286692 224352
rect 286744 224340 286750 224392
rect 291102 224340 291108 224392
rect 291160 224380 291166 224392
rect 323854 224380 323860 224392
rect 291160 224352 323860 224380
rect 291160 224340 291166 224352
rect 323854 224340 323860 224352
rect 323912 224340 323918 224392
rect 341886 224340 341892 224392
rect 341944 224380 341950 224392
rect 365254 224380 365260 224392
rect 341944 224352 365260 224380
rect 341944 224340 341950 224352
rect 365254 224340 365260 224352
rect 365312 224340 365318 224392
rect 368198 224340 368204 224392
rect 368256 224380 368262 224392
rect 382550 224380 382556 224392
rect 368256 224352 382556 224380
rect 368256 224340 368262 224352
rect 382550 224340 382556 224352
rect 382608 224340 382614 224392
rect 382918 224340 382924 224392
rect 382976 224380 382982 224392
rect 396166 224380 396172 224392
rect 382976 224352 396172 224380
rect 382976 224340 382982 224352
rect 396166 224340 396172 224352
rect 396224 224340 396230 224392
rect 436370 224340 436376 224392
rect 436428 224380 436434 224392
rect 436830 224380 436836 224392
rect 436428 224352 436836 224380
rect 436428 224340 436434 224352
rect 436830 224340 436836 224352
rect 436888 224340 436894 224392
rect 480530 224340 480536 224392
rect 480588 224380 480594 224392
rect 492858 224380 492864 224392
rect 480588 224352 492864 224380
rect 480588 224340 480594 224352
rect 492858 224340 492864 224352
rect 492916 224340 492922 224392
rect 497274 224340 497280 224392
rect 497332 224380 497338 224392
rect 514018 224380 514024 224392
rect 497332 224352 514024 224380
rect 497332 224340 497338 224352
rect 514018 224340 514024 224352
rect 514076 224340 514082 224392
rect 519814 224340 519820 224392
rect 519872 224380 519878 224392
rect 542538 224380 542544 224392
rect 519872 224352 542544 224380
rect 519872 224340 519878 224352
rect 542538 224340 542544 224352
rect 542596 224340 542602 224392
rect 549530 224340 549536 224392
rect 549588 224380 549594 224392
rect 625430 224380 625436 224392
rect 549588 224352 625436 224380
rect 549588 224340 549594 224352
rect 625430 224340 625436 224352
rect 625488 224340 625494 224392
rect 63218 224204 63224 224256
rect 63276 224244 63282 224256
rect 147582 224244 147588 224256
rect 63276 224216 147588 224244
rect 63276 224204 63282 224216
rect 147582 224204 147588 224216
rect 147640 224204 147646 224256
rect 151722 224204 151728 224256
rect 151780 224244 151786 224256
rect 217134 224244 217140 224256
rect 151780 224216 217140 224244
rect 151780 224204 151786 224216
rect 217134 224204 217140 224216
rect 217192 224204 217198 224256
rect 223298 224204 223304 224256
rect 223356 224244 223362 224256
rect 224954 224244 224960 224256
rect 223356 224216 224960 224244
rect 223356 224204 223362 224216
rect 224954 224204 224960 224216
rect 225012 224204 225018 224256
rect 231578 224204 231584 224256
rect 231636 224244 231642 224256
rect 278958 224244 278964 224256
rect 231636 224216 278964 224244
rect 231636 224204 231642 224216
rect 278958 224204 278964 224216
rect 279016 224204 279022 224256
rect 281258 224204 281264 224256
rect 281316 224244 281322 224256
rect 317598 224244 317604 224256
rect 281316 224216 317604 224244
rect 281316 224204 281322 224216
rect 317598 224204 317604 224216
rect 317656 224204 317662 224256
rect 322566 224204 322572 224256
rect 322624 224244 322630 224256
rect 349798 224244 349804 224256
rect 322624 224216 349804 224244
rect 322624 224204 322630 224216
rect 349798 224204 349804 224216
rect 349856 224204 349862 224256
rect 351638 224204 351644 224256
rect 351696 224244 351702 224256
rect 369578 224244 369584 224256
rect 351696 224216 369584 224244
rect 351696 224204 351702 224216
rect 369578 224204 369584 224216
rect 369636 224204 369642 224256
rect 372338 224204 372344 224256
rect 372396 224244 372402 224256
rect 387426 224244 387432 224256
rect 372396 224216 387432 224244
rect 372396 224204 372402 224216
rect 387426 224204 387432 224216
rect 387484 224204 387490 224256
rect 387702 224204 387708 224256
rect 387760 224244 387766 224256
rect 398098 224244 398104 224256
rect 387760 224216 398104 224244
rect 387760 224204 387766 224216
rect 398098 224204 398104 224216
rect 398156 224204 398162 224256
rect 405458 224204 405464 224256
rect 405516 224244 405522 224256
rect 414198 224244 414204 224256
rect 405516 224216 414204 224244
rect 405516 224204 405522 224216
rect 414198 224204 414204 224216
rect 414256 224204 414262 224256
rect 420822 224204 420828 224256
rect 420880 224244 420886 224256
rect 425146 224244 425152 224256
rect 420880 224216 425152 224244
rect 420880 224204 420886 224216
rect 425146 224204 425152 224216
rect 425204 224204 425210 224256
rect 427814 224204 427820 224256
rect 427872 224244 427878 224256
rect 428734 224244 428740 224256
rect 427872 224216 428740 224244
rect 427872 224204 427878 224216
rect 428734 224204 428740 224216
rect 428792 224204 428798 224256
rect 436278 224204 436284 224256
rect 436336 224244 436342 224256
rect 437014 224244 437020 224256
rect 436336 224216 437020 224244
rect 436336 224204 436342 224216
rect 437014 224204 437020 224216
rect 437072 224204 437078 224256
rect 438946 224204 438952 224256
rect 439004 224244 439010 224256
rect 439590 224244 439596 224256
rect 439004 224216 439596 224244
rect 439004 224204 439010 224216
rect 439590 224204 439596 224216
rect 439648 224204 439654 224256
rect 451366 224204 451372 224256
rect 451424 224244 451430 224256
rect 452010 224244 452016 224256
rect 451424 224216 452016 224244
rect 451424 224204 451430 224216
rect 452010 224204 452016 224216
rect 452068 224204 452074 224256
rect 456150 224204 456156 224256
rect 456208 224244 456214 224256
rect 459738 224244 459744 224256
rect 456208 224216 459744 224244
rect 456208 224204 456214 224216
rect 459738 224204 459744 224216
rect 459796 224204 459802 224256
rect 462406 224204 462412 224256
rect 462464 224244 462470 224256
rect 469674 224244 469680 224256
rect 462464 224216 469680 224244
rect 462464 224204 462470 224216
rect 469674 224204 469680 224216
rect 469732 224204 469738 224256
rect 470870 224204 470876 224256
rect 470928 224244 470934 224256
rect 477494 224244 477500 224256
rect 470928 224216 477500 224244
rect 470928 224204 470934 224216
rect 477494 224204 477500 224216
rect 477552 224204 477558 224256
rect 489546 224204 489552 224256
rect 489604 224244 489610 224256
rect 504082 224244 504088 224256
rect 489604 224216 504088 224244
rect 489604 224204 489610 224216
rect 504082 224204 504088 224216
rect 504140 224204 504146 224256
rect 504634 224204 504640 224256
rect 504692 224244 504698 224256
rect 523034 224244 523040 224256
rect 504692 224216 523040 224244
rect 504692 224204 504698 224216
rect 523034 224204 523040 224216
rect 523092 224204 523098 224256
rect 527542 224204 527548 224256
rect 527600 224244 527606 224256
rect 552014 224244 552020 224256
rect 527600 224216 552020 224244
rect 527600 224204 527606 224216
rect 552014 224204 552020 224216
rect 552072 224204 552078 224256
rect 556798 224204 556804 224256
rect 556856 224244 556862 224256
rect 570322 224244 570328 224256
rect 556856 224216 570328 224244
rect 556856 224204 556862 224216
rect 570322 224204 570328 224216
rect 570380 224204 570386 224256
rect 115658 224068 115664 224120
rect 115716 224108 115722 224120
rect 188798 224108 188804 224120
rect 115716 224080 188804 224108
rect 115716 224068 115722 224080
rect 188798 224068 188804 224080
rect 188856 224068 188862 224120
rect 189902 224068 189908 224120
rect 189960 224108 189966 224120
rect 212626 224108 212632 224120
rect 189960 224080 212632 224108
rect 189960 224068 189966 224080
rect 212626 224068 212632 224080
rect 212684 224068 212690 224120
rect 216582 224068 216588 224120
rect 216640 224108 216646 224120
rect 264422 224108 264428 224120
rect 216640 224080 264428 224108
rect 216640 224068 216646 224080
rect 264422 224068 264428 224080
rect 264480 224068 264486 224120
rect 275830 224068 275836 224120
rect 275888 224108 275894 224120
rect 288710 224108 288716 224120
rect 275888 224080 288716 224108
rect 275888 224068 275894 224080
rect 288710 224068 288716 224080
rect 288768 224068 288774 224120
rect 510338 224000 510344 224052
rect 510396 224040 510402 224052
rect 615494 224040 615500 224052
rect 510396 224012 615500 224040
rect 510396 224000 510402 224012
rect 615494 224000 615500 224012
rect 615552 224000 615558 224052
rect 122282 223932 122288 223984
rect 122340 223972 122346 223984
rect 193950 223972 193956 223984
rect 122340 223944 193956 223972
rect 122340 223932 122346 223944
rect 193950 223932 193956 223944
rect 194008 223932 194014 223984
rect 196802 223932 196808 223984
rect 196860 223972 196866 223984
rect 222930 223972 222936 223984
rect 196860 223944 222936 223972
rect 196860 223932 196866 223944
rect 222930 223932 222936 223944
rect 222988 223932 222994 223984
rect 226150 223932 226156 223984
rect 226208 223972 226214 223984
rect 272518 223972 272524 223984
rect 226208 223944 272524 223972
rect 226208 223932 226214 223944
rect 272518 223932 272524 223944
rect 272576 223932 272582 223984
rect 289078 223864 289084 223916
rect 289136 223904 289142 223916
rect 294782 223904 294788 223916
rect 289136 223876 294788 223904
rect 289136 223864 289142 223876
rect 294782 223864 294788 223876
rect 294840 223864 294846 223916
rect 514846 223864 514852 223916
rect 514904 223904 514910 223916
rect 515214 223904 515220 223916
rect 514904 223876 515220 223904
rect 514904 223864 514910 223876
rect 515214 223864 515220 223876
rect 515272 223904 515278 223916
rect 616874 223904 616880 223916
rect 515272 223876 616880 223904
rect 515272 223864 515278 223876
rect 616874 223864 616880 223876
rect 616932 223864 616938 223916
rect 140038 223796 140044 223848
rect 140096 223836 140102 223848
rect 171410 223836 171416 223848
rect 140096 223808 171416 223836
rect 140096 223796 140102 223808
rect 171410 223796 171416 223808
rect 171468 223796 171474 223848
rect 175182 223796 175188 223848
rect 175240 223836 175246 223848
rect 235166 223836 235172 223848
rect 175240 223808 235172 223836
rect 175240 223796 175246 223808
rect 235166 223796 235172 223808
rect 235224 223796 235230 223848
rect 514662 223728 514668 223780
rect 514720 223768 514726 223780
rect 536374 223768 536380 223780
rect 514720 223740 536380 223768
rect 514720 223728 514726 223740
rect 536374 223728 536380 223740
rect 536432 223728 536438 223780
rect 539778 223728 539784 223780
rect 539836 223768 539842 223780
rect 622394 223768 622400 223780
rect 539836 223740 622400 223768
rect 539836 223728 539842 223740
rect 622394 223728 622400 223740
rect 622452 223728 622458 223780
rect 181898 223660 181904 223712
rect 181956 223700 181962 223712
rect 181956 223672 185440 223700
rect 181956 223660 181962 223672
rect 102042 223524 102048 223576
rect 102100 223564 102106 223576
rect 178494 223564 178500 223576
rect 102100 223536 178500 223564
rect 102100 223524 102106 223536
rect 178494 223524 178500 223536
rect 178552 223524 178558 223576
rect 185412 223564 185440 223672
rect 185578 223660 185584 223712
rect 185636 223700 185642 223712
rect 191006 223700 191012 223712
rect 185636 223672 191012 223700
rect 185636 223660 185642 223672
rect 191006 223660 191012 223672
rect 191064 223660 191070 223712
rect 227438 223660 227444 223712
rect 227496 223700 227502 223712
rect 273162 223700 273168 223712
rect 227496 223672 273168 223700
rect 227496 223660 227502 223672
rect 273162 223660 273168 223672
rect 273220 223660 273226 223712
rect 415302 223660 415308 223712
rect 415360 223700 415366 223712
rect 419626 223700 419632 223712
rect 415360 223672 419632 223700
rect 415360 223660 415366 223672
rect 419626 223660 419632 223672
rect 419684 223660 419690 223712
rect 460566 223660 460572 223712
rect 460624 223700 460630 223712
rect 462958 223700 462964 223712
rect 460624 223672 462964 223700
rect 460624 223660 460630 223672
rect 462958 223660 462964 223672
rect 463016 223660 463022 223712
rect 670510 223660 670516 223712
rect 670568 223700 670574 223712
rect 670804 223700 670832 224420
rect 670930 224120 670982 224126
rect 670930 224062 670982 224068
rect 670568 223672 670832 223700
rect 670568 223660 670574 223672
rect 543642 223592 543648 223644
rect 543700 223632 543706 223644
rect 557442 223632 557448 223644
rect 543700 223604 557448 223632
rect 543700 223592 543706 223604
rect 557442 223592 557448 223604
rect 557500 223632 557506 223644
rect 626534 223632 626540 223644
rect 557500 223604 626540 223632
rect 557500 223592 557506 223604
rect 626534 223592 626540 223604
rect 626592 223592 626598 223644
rect 654962 223592 654968 223644
rect 655020 223632 655026 223644
rect 656710 223632 656716 223644
rect 655020 223604 656716 223632
rect 655020 223592 655026 223604
rect 656710 223592 656716 223604
rect 656768 223592 656774 223644
rect 186314 223564 186320 223576
rect 185412 223536 186320 223564
rect 186314 223524 186320 223536
rect 186372 223524 186378 223576
rect 194318 223524 194324 223576
rect 194376 223564 194382 223576
rect 247402 223564 247408 223576
rect 194376 223536 247408 223564
rect 194376 223524 194382 223536
rect 247402 223524 247408 223536
rect 247460 223524 247466 223576
rect 253750 223524 253756 223576
rect 253808 223564 253814 223576
rect 293494 223564 293500 223576
rect 253808 223536 293500 223564
rect 253808 223524 253814 223536
rect 293494 223524 293500 223536
rect 293552 223524 293558 223576
rect 307018 223524 307024 223576
rect 307076 223564 307082 223576
rect 315390 223564 315396 223576
rect 307076 223536 315396 223564
rect 307076 223524 307082 223536
rect 315390 223524 315396 223536
rect 315448 223524 315454 223576
rect 454770 223524 454776 223576
rect 454828 223564 454834 223576
rect 460106 223564 460112 223576
rect 454828 223536 460112 223564
rect 454828 223524 454834 223536
rect 460106 223524 460112 223536
rect 460164 223524 460170 223576
rect 473722 223524 473728 223576
rect 473780 223564 473786 223576
rect 480990 223564 480996 223576
rect 473780 223536 480996 223564
rect 473780 223524 473786 223536
rect 480990 223524 480996 223536
rect 481048 223524 481054 223576
rect 670326 223524 670332 223576
rect 670384 223564 670390 223576
rect 670384 223536 670648 223564
rect 670384 223524 670390 223536
rect 88242 223388 88248 223440
rect 88300 223428 88306 223440
rect 164970 223428 164976 223440
rect 88300 223400 164976 223428
rect 88300 223388 88306 223400
rect 164970 223388 164976 223400
rect 165028 223388 165034 223440
rect 166442 223388 166448 223440
rect 166500 223428 166506 223440
rect 192018 223428 192024 223440
rect 166500 223400 192024 223428
rect 166500 223388 166506 223400
rect 192018 223388 192024 223400
rect 192076 223388 192082 223440
rect 197262 223388 197268 223440
rect 197320 223428 197326 223440
rect 249978 223428 249984 223440
rect 197320 223400 249984 223428
rect 197320 223388 197326 223400
rect 249978 223388 249984 223400
rect 250036 223388 250042 223440
rect 267366 223388 267372 223440
rect 267424 223428 267430 223440
rect 307294 223428 307300 223440
rect 267424 223400 307300 223428
rect 267424 223388 267430 223400
rect 307294 223388 307300 223400
rect 307352 223388 307358 223440
rect 322842 223388 322848 223440
rect 322900 223428 322906 223440
rect 332410 223428 332416 223440
rect 322900 223400 332416 223428
rect 322900 223388 322906 223400
rect 332410 223388 332416 223400
rect 332468 223388 332474 223440
rect 498562 223388 498568 223440
rect 498620 223428 498626 223440
rect 515766 223428 515772 223440
rect 498620 223400 515772 223428
rect 498620 223388 498626 223400
rect 515766 223388 515772 223400
rect 515824 223388 515830 223440
rect 516778 223388 516784 223440
rect 516836 223428 516842 223440
rect 527174 223428 527180 223440
rect 516836 223400 527180 223428
rect 516836 223388 516842 223400
rect 527174 223388 527180 223400
rect 527232 223388 527238 223440
rect 528554 223388 528560 223440
rect 528612 223428 528618 223440
rect 542354 223428 542360 223440
rect 528612 223400 542360 223428
rect 528612 223388 528618 223400
rect 542354 223388 542360 223400
rect 542412 223388 542418 223440
rect 670620 223304 670648 223536
rect 78398 223252 78404 223304
rect 78456 223292 78462 223304
rect 78456 223264 154528 223292
rect 78456 223252 78462 223264
rect 81158 223116 81164 223168
rect 81216 223156 81222 223168
rect 154298 223156 154304 223168
rect 81216 223128 154304 223156
rect 81216 223116 81222 223128
rect 154298 223116 154304 223128
rect 154356 223116 154362 223168
rect 154500 223156 154528 223264
rect 157058 223252 157064 223304
rect 157116 223292 157122 223304
rect 160186 223292 160192 223304
rect 157116 223264 160192 223292
rect 157116 223252 157122 223264
rect 160186 223252 160192 223264
rect 160244 223252 160250 223304
rect 181714 223292 181720 223304
rect 161446 223264 181720 223292
rect 157242 223156 157248 223168
rect 154500 223128 157248 223156
rect 157242 223116 157248 223128
rect 157300 223116 157306 223168
rect 159266 223116 159272 223168
rect 159324 223156 159330 223168
rect 161446 223156 161474 223264
rect 181714 223252 181720 223264
rect 181772 223252 181778 223304
rect 191650 223252 191656 223304
rect 191708 223292 191714 223304
rect 244826 223292 244832 223304
rect 191708 223264 244832 223292
rect 191708 223252 191714 223264
rect 244826 223252 244832 223264
rect 244884 223252 244890 223304
rect 262122 223252 262128 223304
rect 262180 223292 262186 223304
rect 300854 223292 300860 223304
rect 262180 223264 300860 223292
rect 262180 223252 262186 223264
rect 300854 223252 300860 223264
rect 300912 223252 300918 223304
rect 315666 223252 315672 223304
rect 315724 223292 315730 223304
rect 341426 223292 341432 223304
rect 315724 223264 341432 223292
rect 315724 223252 315730 223264
rect 341426 223252 341432 223264
rect 341484 223252 341490 223304
rect 342070 223252 342076 223304
rect 342128 223292 342134 223304
rect 362034 223292 362040 223304
rect 342128 223264 362040 223292
rect 342128 223252 342134 223264
rect 362034 223252 362040 223264
rect 362092 223252 362098 223304
rect 366910 223252 366916 223304
rect 366968 223292 366974 223304
rect 381998 223292 382004 223304
rect 366968 223264 382004 223292
rect 366968 223252 366974 223264
rect 381998 223252 382004 223264
rect 382056 223252 382062 223304
rect 407022 223252 407028 223304
rect 407080 223292 407086 223304
rect 414842 223292 414848 223304
rect 407080 223264 414848 223292
rect 407080 223252 407086 223264
rect 414842 223252 414848 223264
rect 414900 223252 414906 223304
rect 503438 223252 503444 223304
rect 503496 223292 503502 223304
rect 521746 223292 521752 223304
rect 503496 223264 521752 223292
rect 503496 223252 503502 223264
rect 521746 223252 521752 223264
rect 521804 223252 521810 223304
rect 522482 223252 522488 223304
rect 522540 223292 522546 223304
rect 534902 223292 534908 223304
rect 522540 223264 534908 223292
rect 522540 223252 522546 223264
rect 534902 223252 534908 223264
rect 534960 223252 534966 223304
rect 536742 223252 536748 223304
rect 536800 223292 536806 223304
rect 559926 223292 559932 223304
rect 536800 223264 559932 223292
rect 536800 223252 536806 223264
rect 559926 223252 559932 223264
rect 559984 223292 559990 223304
rect 567746 223292 567752 223304
rect 559984 223264 567752 223292
rect 559984 223252 559990 223264
rect 567746 223252 567752 223264
rect 567804 223252 567810 223304
rect 670602 223252 670608 223304
rect 670660 223252 670666 223304
rect 159324 223128 161474 223156
rect 159324 223116 159330 223128
rect 168282 223116 168288 223168
rect 168340 223156 168346 223168
rect 226794 223156 226800 223168
rect 168340 223128 226800 223156
rect 168340 223116 168346 223128
rect 226794 223116 226800 223128
rect 226852 223116 226858 223168
rect 248138 223116 248144 223168
rect 248196 223156 248202 223168
rect 291838 223156 291844 223168
rect 248196 223128 291844 223156
rect 248196 223116 248202 223128
rect 291838 223116 291844 223128
rect 291896 223116 291902 223168
rect 300762 223116 300768 223168
rect 300820 223156 300826 223168
rect 330110 223156 330116 223168
rect 300820 223128 330116 223156
rect 300820 223116 300826 223128
rect 330110 223116 330116 223128
rect 330168 223116 330174 223168
rect 336458 223116 336464 223168
rect 336516 223156 336522 223168
rect 359734 223156 359740 223168
rect 336516 223128 359740 223156
rect 336516 223116 336522 223128
rect 359734 223116 359740 223128
rect 359792 223116 359798 223168
rect 366726 223116 366732 223168
rect 366784 223156 366790 223168
rect 383930 223156 383936 223168
rect 366784 223128 383936 223156
rect 366784 223116 366790 223128
rect 383930 223116 383936 223128
rect 383988 223116 383994 223168
rect 483106 223116 483112 223168
rect 483164 223156 483170 223168
rect 495802 223156 495808 223168
rect 483164 223128 495808 223156
rect 483164 223116 483170 223128
rect 495802 223116 495808 223128
rect 495860 223116 495866 223168
rect 515950 223116 515956 223168
rect 516008 223156 516014 223168
rect 538306 223156 538312 223168
rect 516008 223128 538312 223156
rect 516008 223116 516014 223128
rect 538306 223116 538312 223128
rect 538364 223156 538370 223168
rect 539042 223156 539048 223168
rect 538364 223128 539048 223156
rect 538364 223116 538370 223128
rect 539042 223116 539048 223128
rect 539100 223116 539106 223168
rect 75822 222980 75828 223032
rect 75880 223020 75886 223032
rect 154666 223020 154672 223032
rect 75880 222992 154672 223020
rect 75880 222980 75886 222992
rect 154666 222980 154672 222992
rect 154724 222980 154730 223032
rect 164050 222980 164056 223032
rect 164108 223020 164114 223032
rect 224218 223020 224224 223032
rect 164108 222992 224224 223020
rect 164108 222980 164114 222992
rect 224218 222980 224224 222992
rect 224276 222980 224282 223032
rect 238662 222980 238668 223032
rect 238720 223020 238726 223032
rect 282822 223020 282828 223032
rect 238720 222992 282828 223020
rect 238720 222980 238726 222992
rect 282822 222980 282828 222992
rect 282880 222980 282886 223032
rect 292482 222980 292488 223032
rect 292540 223020 292546 223032
rect 326614 223020 326620 223032
rect 292540 222992 326620 223020
rect 292540 222980 292546 222992
rect 326614 222980 326620 222992
rect 326672 222980 326678 223032
rect 329742 222980 329748 223032
rect 329800 223020 329806 223032
rect 353662 223020 353668 223032
rect 329800 222992 353668 223020
rect 329800 222980 329806 222992
rect 353662 222980 353668 222992
rect 353720 222980 353726 223032
rect 355778 222980 355784 223032
rect 355836 223020 355842 223032
rect 375558 223020 375564 223032
rect 355836 222992 375564 223020
rect 355836 222980 355842 222992
rect 375558 222980 375564 222992
rect 375616 222980 375622 223032
rect 382090 222980 382096 223032
rect 382148 223020 382154 223032
rect 392946 223020 392952 223032
rect 382148 222992 392952 223020
rect 382148 222980 382154 222992
rect 392946 222980 392952 222992
rect 393004 222980 393010 223032
rect 479886 222980 479892 223032
rect 479944 223020 479950 223032
rect 491938 223020 491944 223032
rect 479944 222992 491944 223020
rect 479944 222980 479950 222992
rect 491938 222980 491944 222992
rect 491996 222980 492002 223032
rect 500494 222980 500500 223032
rect 500552 223020 500558 223032
rect 518434 223020 518440 223032
rect 500552 222992 518440 223020
rect 500552 222980 500558 222992
rect 518434 222980 518440 222992
rect 518492 222980 518498 223032
rect 518802 222980 518808 223032
rect 518860 223020 518866 223032
rect 618254 223020 618260 223032
rect 518860 222992 618260 223020
rect 518860 222980 518866 222992
rect 618254 222980 618260 222992
rect 618312 222980 618318 223032
rect 68922 222844 68928 222896
rect 68980 222884 68986 222896
rect 149514 222884 149520 222896
rect 68980 222856 149520 222884
rect 68980 222844 68986 222856
rect 149514 222844 149520 222856
rect 149572 222844 149578 222896
rect 154482 222844 154488 222896
rect 154540 222884 154546 222896
rect 216214 222884 216220 222896
rect 154540 222856 216220 222884
rect 154540 222844 154546 222856
rect 216214 222844 216220 222856
rect 216272 222844 216278 222896
rect 217778 222844 217784 222896
rect 217836 222884 217842 222896
rect 268654 222884 268660 222896
rect 217836 222856 268660 222884
rect 217836 222844 217842 222856
rect 268654 222844 268660 222856
rect 268712 222844 268718 222896
rect 278406 222844 278412 222896
rect 278464 222884 278470 222896
rect 313734 222884 313740 222896
rect 278464 222856 313740 222884
rect 278464 222844 278470 222856
rect 313734 222844 313740 222856
rect 313792 222844 313798 222896
rect 315850 222844 315856 222896
rect 315908 222884 315914 222896
rect 344646 222884 344652 222896
rect 315908 222856 344652 222884
rect 315908 222844 315914 222856
rect 344646 222844 344652 222856
rect 344704 222844 344710 222896
rect 346210 222844 346216 222896
rect 346268 222884 346274 222896
rect 367462 222884 367468 222896
rect 346268 222856 367468 222884
rect 346268 222844 346274 222856
rect 367462 222844 367468 222856
rect 367520 222844 367526 222896
rect 386322 222844 386328 222896
rect 386380 222884 386386 222896
rect 398374 222884 398380 222896
rect 386380 222856 398380 222884
rect 386380 222844 386386 222856
rect 398374 222844 398380 222856
rect 398432 222844 398438 222896
rect 398558 222844 398564 222896
rect 398616 222884 398622 222896
rect 405826 222884 405832 222896
rect 398616 222856 405832 222884
rect 398616 222844 398622 222856
rect 405826 222844 405832 222856
rect 405884 222844 405890 222896
rect 459922 222844 459928 222896
rect 459980 222884 459986 222896
rect 466730 222884 466736 222896
rect 459980 222856 466736 222884
rect 459980 222844 459986 222856
rect 466730 222844 466736 222856
rect 466788 222844 466794 222896
rect 467282 222844 467288 222896
rect 467340 222884 467346 222896
rect 475010 222884 475016 222896
rect 467340 222856 475016 222884
rect 467340 222844 467346 222856
rect 475010 222844 475016 222856
rect 475068 222844 475074 222896
rect 486326 222844 486332 222896
rect 486384 222884 486390 222896
rect 499850 222884 499856 222896
rect 486384 222856 499856 222884
rect 486384 222844 486390 222856
rect 499850 222844 499856 222856
rect 499908 222844 499914 222896
rect 508866 222844 508872 222896
rect 508924 222884 508930 222896
rect 528922 222884 528928 222896
rect 508924 222856 528928 222884
rect 508924 222844 508930 222856
rect 528922 222844 528928 222856
rect 528980 222844 528986 222896
rect 537202 222844 537208 222896
rect 537260 222884 537266 222896
rect 565630 222884 565636 222896
rect 537260 222856 565636 222884
rect 537260 222844 537266 222856
rect 565630 222844 565636 222856
rect 565688 222884 565694 222896
rect 571610 222884 571616 222896
rect 565688 222856 571616 222884
rect 565688 222844 565694 222856
rect 571610 222844 571616 222856
rect 571668 222844 571674 222896
rect 131022 222708 131028 222760
rect 131080 222748 131086 222760
rect 196066 222748 196072 222760
rect 131080 222720 196072 222748
rect 131080 222708 131086 222720
rect 196066 222708 196072 222720
rect 196124 222708 196130 222760
rect 208118 222708 208124 222760
rect 208176 222748 208182 222760
rect 260926 222748 260932 222760
rect 208176 222720 260932 222748
rect 208176 222708 208182 222720
rect 260926 222708 260932 222720
rect 260984 222708 260990 222760
rect 290918 222708 290924 222760
rect 290976 222748 290982 222760
rect 321830 222748 321836 222760
rect 290976 222720 321836 222748
rect 290976 222708 290982 222720
rect 321830 222708 321836 222720
rect 321888 222708 321894 222760
rect 525150 222708 525156 222760
rect 525208 222748 525214 222760
rect 537570 222748 537576 222760
rect 525208 222720 537576 222748
rect 525208 222708 525214 222720
rect 537570 222708 537576 222720
rect 537628 222748 537634 222760
rect 537628 222720 538536 222748
rect 537628 222708 537634 222720
rect 146018 222572 146024 222624
rect 146076 222612 146082 222624
rect 211982 222612 211988 222624
rect 146076 222584 211988 222612
rect 146076 222572 146082 222584
rect 211982 222572 211988 222584
rect 212040 222572 212046 222624
rect 213822 222572 213828 222624
rect 213880 222612 213886 222624
rect 262858 222612 262864 222624
rect 213880 222584 262864 222612
rect 213880 222572 213886 222584
rect 262858 222572 262864 222584
rect 262916 222572 262922 222624
rect 538508 222612 538536 222720
rect 542354 222708 542360 222760
rect 542412 222748 542418 222760
rect 622578 222748 622584 222760
rect 542412 222720 622584 222748
rect 542412 222708 542418 222720
rect 622578 222708 622584 222720
rect 622636 222708 622642 222760
rect 622762 222612 622768 222624
rect 538508 222584 622768 222612
rect 622762 222572 622768 222584
rect 622820 222572 622826 222624
rect 528526 222516 538444 222544
rect 134702 222436 134708 222488
rect 134760 222476 134766 222488
rect 197446 222476 197452 222488
rect 134760 222448 197452 222476
rect 134760 222436 134766 222448
rect 197446 222436 197452 222448
rect 197504 222436 197510 222488
rect 204162 222436 204168 222488
rect 204220 222476 204226 222488
rect 254762 222476 254768 222488
rect 204220 222448 254768 222476
rect 204220 222436 204226 222448
rect 254762 222436 254768 222448
rect 254820 222436 254826 222488
rect 527174 222436 527180 222488
rect 527232 222476 527238 222488
rect 528526 222476 528554 222516
rect 527232 222448 528554 222476
rect 538416 222476 538444 222516
rect 620002 222476 620008 222488
rect 538416 222448 620008 222476
rect 527232 222436 527238 222448
rect 620002 222436 620008 222448
rect 620060 222436 620066 222488
rect 416498 222368 416504 222420
rect 416556 222408 416562 222420
rect 422202 222408 422208 222420
rect 416556 222380 422208 222408
rect 416556 222368 416562 222380
rect 422202 222368 422208 222380
rect 422260 222368 422266 222420
rect 533356 222380 534074 222408
rect 154298 222300 154304 222352
rect 154356 222340 154362 222352
rect 159818 222340 159824 222352
rect 154356 222312 159824 222340
rect 154356 222300 154362 222312
rect 159818 222300 159824 222312
rect 159876 222300 159882 222352
rect 178678 222300 178684 222352
rect 178736 222340 178742 222352
rect 204898 222340 204904 222352
rect 178736 222312 204904 222340
rect 178736 222300 178742 222312
rect 204898 222300 204904 222312
rect 204956 222300 204962 222352
rect 243998 222300 244004 222352
rect 244056 222340 244062 222352
rect 286042 222340 286048 222352
rect 244056 222312 286048 222340
rect 244056 222300 244062 222312
rect 286042 222300 286048 222312
rect 286100 222300 286106 222352
rect 524782 222300 524788 222352
rect 524840 222340 524846 222352
rect 533356 222340 533384 222380
rect 524840 222312 533384 222340
rect 534046 222340 534074 222380
rect 619818 222340 619824 222352
rect 534046 222312 619824 222340
rect 524840 222300 524846 222312
rect 619818 222300 619824 222312
rect 619876 222300 619882 222352
rect 529474 222164 529480 222216
rect 529532 222204 529538 222216
rect 555694 222204 555700 222216
rect 529532 222176 555700 222204
rect 529532 222164 529538 222176
rect 555694 222164 555700 222176
rect 555752 222164 555758 222216
rect 567746 222164 567752 222216
rect 567804 222204 567810 222216
rect 627086 222204 627092 222216
rect 567804 222176 627092 222204
rect 567804 222164 567810 222176
rect 627086 222164 627092 222176
rect 627144 222164 627150 222216
rect 670326 222164 670332 222216
rect 670384 222204 670390 222216
rect 670786 222204 670792 222216
rect 670384 222176 670792 222204
rect 670384 222164 670390 222176
rect 670786 222164 670792 222176
rect 670844 222164 670850 222216
rect 111426 222096 111432 222148
rect 111484 222136 111490 222148
rect 182542 222136 182548 222148
rect 111484 222108 182548 222136
rect 111484 222096 111490 222108
rect 182542 222096 182548 222108
rect 182600 222096 182606 222148
rect 184014 222096 184020 222148
rect 184072 222136 184078 222148
rect 239214 222136 239220 222148
rect 184072 222108 239220 222136
rect 184072 222096 184078 222108
rect 239214 222096 239220 222108
rect 239272 222096 239278 222148
rect 267090 222096 267096 222148
rect 267148 222136 267154 222148
rect 303798 222136 303804 222148
rect 267148 222108 303804 222136
rect 267148 222096 267154 222108
rect 303798 222096 303804 222108
rect 303856 222096 303862 222148
rect 330846 222096 330852 222148
rect 330904 222136 330910 222148
rect 345658 222136 345664 222148
rect 330904 222108 345664 222136
rect 330904 222096 330910 222108
rect 345658 222096 345664 222108
rect 345716 222096 345722 222148
rect 424962 222096 424968 222148
rect 425020 222136 425026 222148
rect 429286 222136 429292 222148
rect 425020 222108 429292 222136
rect 425020 222096 425026 222108
rect 429286 222096 429292 222108
rect 429344 222096 429350 222148
rect 462130 222096 462136 222148
rect 462188 222136 462194 222148
rect 468478 222136 468484 222148
rect 462188 222108 468484 222136
rect 462188 222096 462194 222108
rect 468478 222096 468484 222108
rect 468536 222096 468542 222148
rect 471882 222096 471888 222148
rect 471940 222136 471946 222148
rect 479242 222136 479248 222148
rect 471940 222108 479248 222136
rect 471940 222096 471946 222108
rect 479242 222096 479248 222108
rect 479300 222096 479306 222148
rect 509878 222096 509884 222148
rect 509936 222136 509942 222148
rect 518802 222136 518808 222148
rect 509936 222108 518808 222136
rect 509936 222096 509942 222108
rect 518802 222096 518808 222108
rect 518860 222136 518866 222148
rect 519814 222136 519820 222148
rect 518860 222108 519820 222136
rect 518860 222096 518866 222108
rect 519814 222096 519820 222108
rect 519872 222096 519878 222148
rect 533338 222028 533344 222080
rect 533396 222068 533402 222080
rect 538674 222068 538680 222080
rect 533396 222040 538680 222068
rect 533396 222028 533402 222040
rect 538674 222028 538680 222040
rect 538732 222028 538738 222080
rect 104618 221960 104624 222012
rect 104676 222000 104682 222012
rect 177482 222000 177488 222012
rect 104676 221972 177488 222000
rect 104676 221960 104682 221972
rect 177482 221960 177488 221972
rect 177540 221960 177546 222012
rect 195146 221960 195152 222012
rect 195204 222000 195210 222012
rect 250162 222000 250168 222012
rect 195204 221972 250168 222000
rect 195204 221960 195210 221972
rect 250162 221960 250168 221972
rect 250220 221960 250226 222012
rect 269942 221960 269948 222012
rect 270000 222000 270006 222012
rect 306558 222000 306564 222012
rect 270000 221972 306564 222000
rect 270000 221960 270006 221972
rect 306558 221960 306564 221972
rect 306616 221960 306622 222012
rect 306834 221960 306840 222012
rect 306892 222000 306898 222012
rect 335446 222000 335452 222012
rect 306892 221972 335452 222000
rect 306892 221960 306898 221972
rect 335446 221960 335452 221972
rect 335504 221960 335510 222012
rect 513742 221960 513748 222012
rect 513800 222000 513806 222012
rect 524782 222000 524788 222012
rect 513800 221972 524788 222000
rect 513800 221960 513806 221972
rect 524782 221960 524788 221972
rect 524840 221960 524846 222012
rect 539042 221960 539048 222012
rect 539100 222000 539106 222012
rect 604454 222000 604460 222012
rect 539100 221972 604460 222000
rect 539100 221960 539106 221972
rect 604454 221960 604460 221972
rect 604512 221960 604518 222012
rect 101490 221824 101496 221876
rect 101548 221864 101554 221876
rect 175458 221864 175464 221876
rect 101548 221836 175464 221864
rect 101548 221824 101554 221836
rect 175458 221824 175464 221836
rect 175516 221824 175522 221876
rect 189442 221824 189448 221876
rect 189500 221864 189506 221876
rect 245102 221864 245108 221876
rect 189500 221836 245108 221864
rect 189500 221824 189506 221836
rect 245102 221824 245108 221836
rect 245160 221824 245166 221876
rect 258074 221824 258080 221876
rect 258132 221864 258138 221876
rect 269206 221864 269212 221876
rect 258132 221836 269212 221864
rect 258132 221824 258138 221836
rect 269206 221824 269212 221836
rect 269264 221824 269270 221876
rect 277854 221824 277860 221876
rect 277912 221864 277918 221876
rect 314838 221864 314844 221876
rect 277912 221836 314844 221864
rect 277912 221824 277918 221836
rect 314838 221824 314844 221836
rect 314896 221824 314902 221876
rect 344922 221824 344928 221876
rect 344980 221864 344986 221876
rect 364518 221864 364524 221876
rect 344980 221836 364524 221864
rect 344980 221824 344986 221836
rect 364518 221824 364524 221836
rect 364576 221824 364582 221876
rect 484302 221824 484308 221876
rect 484360 221864 484366 221876
rect 496906 221864 496912 221876
rect 484360 221836 496912 221864
rect 484360 221824 484366 221836
rect 496906 221824 496912 221836
rect 496964 221824 496970 221876
rect 523954 221824 523960 221876
rect 524012 221864 524018 221876
rect 548978 221864 548984 221876
rect 524012 221836 548984 221864
rect 524012 221824 524018 221836
rect 548978 221824 548984 221836
rect 549036 221824 549042 221876
rect 560754 221824 560760 221876
rect 560812 221864 560818 221876
rect 561306 221864 561312 221876
rect 560812 221836 561312 221864
rect 560812 221824 560818 221836
rect 561306 221824 561312 221836
rect 561364 221824 561370 221876
rect 565078 221824 565084 221876
rect 565136 221864 565142 221876
rect 567286 221864 567292 221876
rect 565136 221836 567292 221864
rect 565136 221824 565142 221836
rect 567286 221824 567292 221836
rect 567344 221824 567350 221876
rect 60642 221688 60648 221740
rect 60700 221728 60706 221740
rect 94498 221728 94504 221740
rect 60700 221700 94504 221728
rect 60700 221688 60706 221700
rect 94498 221688 94504 221700
rect 94556 221688 94562 221740
rect 94866 221688 94872 221740
rect 94924 221728 94930 221740
rect 161474 221728 161480 221740
rect 94924 221700 161480 221728
rect 94924 221688 94930 221700
rect 161474 221688 161480 221700
rect 161532 221688 161538 221740
rect 167270 221728 167276 221740
rect 161676 221700 167276 221728
rect 74166 221552 74172 221604
rect 74224 221592 74230 221604
rect 86218 221592 86224 221604
rect 74224 221564 86224 221592
rect 74224 221552 74230 221564
rect 86218 221552 86224 221564
rect 86276 221552 86282 221604
rect 91554 221552 91560 221604
rect 91612 221592 91618 221604
rect 161676 221592 161704 221700
rect 167270 221688 167276 221700
rect 167328 221688 167334 221740
rect 177666 221688 177672 221740
rect 177724 221728 177730 221740
rect 234154 221728 234160 221740
rect 177724 221700 234160 221728
rect 177724 221688 177730 221700
rect 234154 221688 234160 221700
rect 234212 221688 234218 221740
rect 247126 221688 247132 221740
rect 247184 221728 247190 221740
rect 253382 221728 253388 221740
rect 247184 221700 253388 221728
rect 247184 221688 247190 221700
rect 253382 221688 253388 221700
rect 253440 221688 253446 221740
rect 253566 221688 253572 221740
rect 253624 221728 253630 221740
rect 258626 221728 258632 221740
rect 253624 221700 258632 221728
rect 253624 221688 253630 221700
rect 258626 221688 258632 221700
rect 258684 221688 258690 221740
rect 260466 221688 260472 221740
rect 260524 221728 260530 221740
rect 298370 221728 298376 221740
rect 260524 221700 298376 221728
rect 260524 221688 260530 221700
rect 298370 221688 298376 221700
rect 298428 221688 298434 221740
rect 298554 221688 298560 221740
rect 298612 221728 298618 221740
rect 328546 221728 328552 221740
rect 298612 221700 328552 221728
rect 298612 221688 298618 221700
rect 328546 221688 328552 221700
rect 328604 221688 328610 221740
rect 331674 221688 331680 221740
rect 331732 221728 331738 221740
rect 353938 221728 353944 221740
rect 331732 221700 353944 221728
rect 331732 221688 331738 221700
rect 353938 221688 353944 221700
rect 353996 221688 354002 221740
rect 362310 221688 362316 221740
rect 362368 221728 362374 221740
rect 376018 221728 376024 221740
rect 362368 221700 376024 221728
rect 362368 221688 362374 221700
rect 376018 221688 376024 221700
rect 376076 221688 376082 221740
rect 382734 221728 382740 221740
rect 378428 221700 382740 221728
rect 162026 221592 162032 221604
rect 91612 221564 161704 221592
rect 161768 221564 162032 221592
rect 91612 221552 91618 221564
rect 84930 221416 84936 221468
rect 84988 221456 84994 221468
rect 161768 221456 161796 221564
rect 162026 221552 162032 221564
rect 162084 221552 162090 221604
rect 178494 221552 178500 221604
rect 178552 221592 178558 221604
rect 237374 221592 237380 221604
rect 178552 221564 237380 221592
rect 178552 221552 178558 221564
rect 237374 221552 237380 221564
rect 237432 221552 237438 221604
rect 238846 221552 238852 221604
rect 238904 221592 238910 221604
rect 248598 221592 248604 221604
rect 238904 221564 248604 221592
rect 238904 221552 238910 221564
rect 248598 221552 248604 221564
rect 248656 221552 248662 221604
rect 250530 221552 250536 221604
rect 250588 221592 250594 221604
rect 291378 221592 291384 221604
rect 250588 221564 291384 221592
rect 250588 221552 250594 221564
rect 291378 221552 291384 221564
rect 291436 221552 291442 221604
rect 296438 221552 296444 221604
rect 296496 221592 296502 221604
rect 327534 221592 327540 221604
rect 296496 221564 327540 221592
rect 296496 221552 296502 221564
rect 327534 221552 327540 221564
rect 327592 221552 327598 221604
rect 328362 221552 328368 221604
rect 328420 221592 328426 221604
rect 351362 221592 351368 221604
rect 328420 221564 351368 221592
rect 328420 221552 328426 221564
rect 351362 221552 351368 221564
rect 351420 221552 351426 221604
rect 353386 221552 353392 221604
rect 353444 221592 353450 221604
rect 369946 221592 369952 221604
rect 353444 221564 369952 221592
rect 353444 221552 353450 221564
rect 369946 221552 369952 221564
rect 370004 221552 370010 221604
rect 370498 221552 370504 221604
rect 370556 221592 370562 221604
rect 378428 221592 378456 221700
rect 382734 221688 382740 221700
rect 382792 221688 382798 221740
rect 494330 221688 494336 221740
rect 494388 221728 494394 221740
rect 510706 221728 510712 221740
rect 494388 221700 510712 221728
rect 494388 221688 494394 221700
rect 510706 221688 510712 221700
rect 510764 221688 510770 221740
rect 522850 221688 522856 221740
rect 522908 221728 522914 221740
rect 546494 221728 546500 221740
rect 522908 221700 546500 221728
rect 522908 221688 522914 221700
rect 546494 221688 546500 221700
rect 546552 221688 546558 221740
rect 548518 221688 548524 221740
rect 548576 221728 548582 221740
rect 607214 221728 607220 221740
rect 548576 221700 607220 221728
rect 548576 221688 548582 221700
rect 607214 221688 607220 221700
rect 607272 221688 607278 221740
rect 370556 221564 378456 221592
rect 370556 221552 370562 221564
rect 382734 221552 382740 221604
rect 382792 221592 382798 221604
rect 394878 221592 394884 221604
rect 382792 221564 394884 221592
rect 382792 221552 382798 221564
rect 394878 221552 394884 221564
rect 394936 221552 394942 221604
rect 397086 221552 397092 221604
rect 397144 221592 397150 221604
rect 407298 221592 407304 221604
rect 397144 221564 407304 221592
rect 397144 221552 397150 221564
rect 407298 221552 407304 221564
rect 407356 221552 407362 221604
rect 456702 221552 456708 221604
rect 456760 221592 456766 221604
rect 461762 221592 461768 221604
rect 456760 221564 461768 221592
rect 456760 221552 456766 221564
rect 461762 221552 461768 221564
rect 461820 221552 461826 221604
rect 468754 221552 468760 221604
rect 468812 221592 468818 221604
rect 474274 221592 474280 221604
rect 468812 221564 474280 221592
rect 468812 221552 468818 221564
rect 474274 221552 474280 221564
rect 474332 221552 474338 221604
rect 478782 221552 478788 221604
rect 478840 221592 478846 221604
rect 489178 221592 489184 221604
rect 478840 221564 489184 221592
rect 478840 221552 478846 221564
rect 489178 221552 489184 221564
rect 489236 221552 489242 221604
rect 496170 221552 496176 221604
rect 496228 221592 496234 221604
rect 513466 221592 513472 221604
rect 496228 221564 513472 221592
rect 496228 221552 496234 221564
rect 513466 221552 513472 221564
rect 513524 221552 513530 221604
rect 533706 221552 533712 221604
rect 533764 221592 533770 221604
rect 533764 221564 535132 221592
rect 533764 221552 533770 221564
rect 535104 221524 535132 221564
rect 535454 221552 535460 221604
rect 535512 221592 535518 221604
rect 538490 221592 538496 221604
rect 535512 221564 538496 221592
rect 535512 221552 535518 221564
rect 538490 221552 538496 221564
rect 538548 221552 538554 221604
rect 538674 221552 538680 221604
rect 538732 221592 538738 221604
rect 603074 221592 603080 221604
rect 538732 221564 603080 221592
rect 538732 221552 538738 221564
rect 603074 221552 603080 221564
rect 603132 221552 603138 221604
rect 535104 221496 535316 221524
rect 84988 221428 161796 221456
rect 84988 221416 84994 221428
rect 161934 221416 161940 221468
rect 161992 221456 161998 221468
rect 224402 221456 224408 221468
rect 161992 221428 224408 221456
rect 161992 221416 161998 221428
rect 224402 221416 224408 221428
rect 224460 221416 224466 221468
rect 234338 221416 234344 221468
rect 234396 221456 234402 221468
rect 281718 221456 281724 221468
rect 234396 221428 281724 221456
rect 234396 221416 234402 221428
rect 281718 221416 281724 221428
rect 281776 221416 281782 221468
rect 284018 221416 284024 221468
rect 284076 221456 284082 221468
rect 289906 221456 289912 221468
rect 284076 221428 289912 221456
rect 284076 221416 284082 221428
rect 289906 221416 289912 221428
rect 289964 221416 289970 221468
rect 292298 221416 292304 221468
rect 292356 221456 292362 221468
rect 299750 221456 299756 221468
rect 292356 221428 299756 221456
rect 292356 221416 292362 221428
rect 299750 221416 299756 221428
rect 299808 221416 299814 221468
rect 302694 221416 302700 221468
rect 302752 221456 302758 221468
rect 334066 221456 334072 221468
rect 302752 221428 334072 221456
rect 302752 221416 302758 221428
rect 334066 221416 334072 221428
rect 334124 221416 334130 221468
rect 335262 221416 335268 221468
rect 335320 221456 335326 221468
rect 357526 221456 357532 221468
rect 335320 221428 357532 221456
rect 335320 221416 335326 221428
rect 357526 221416 357532 221428
rect 357584 221416 357590 221468
rect 358170 221416 358176 221468
rect 358228 221456 358234 221468
rect 374546 221456 374552 221468
rect 358228 221428 374552 221456
rect 358228 221416 358234 221428
rect 374546 221416 374552 221428
rect 374604 221416 374610 221468
rect 375466 221416 375472 221468
rect 375524 221456 375530 221468
rect 386506 221456 386512 221468
rect 375524 221428 386512 221456
rect 375524 221416 375530 221428
rect 386506 221416 386512 221428
rect 386564 221416 386570 221468
rect 390462 221416 390468 221468
rect 390520 221456 390526 221468
rect 401686 221456 401692 221468
rect 390520 221428 401692 221456
rect 390520 221416 390526 221428
rect 401686 221416 401692 221428
rect 401744 221416 401750 221468
rect 408402 221416 408408 221468
rect 408460 221456 408466 221468
rect 416866 221456 416872 221468
rect 408460 221428 416872 221456
rect 408460 221416 408466 221428
rect 416866 221416 416872 221428
rect 416924 221416 416930 221468
rect 452562 221416 452568 221468
rect 452620 221456 452626 221468
rect 456702 221456 456708 221468
rect 452620 221428 456708 221456
rect 452620 221416 452626 221428
rect 456702 221416 456708 221428
rect 456760 221416 456766 221468
rect 484026 221416 484032 221468
rect 484084 221456 484090 221468
rect 534626 221456 534632 221468
rect 484084 221428 534632 221456
rect 484084 221416 484090 221428
rect 534626 221416 534632 221428
rect 534684 221416 534690 221468
rect 535288 221456 535316 221496
rect 560754 221456 560760 221468
rect 535288 221428 560760 221456
rect 560754 221416 560760 221428
rect 560812 221416 560818 221468
rect 560938 221348 560944 221400
rect 560996 221388 561002 221400
rect 568666 221388 568672 221400
rect 560996 221360 568672 221388
rect 560996 221348 561002 221360
rect 568666 221348 568672 221360
rect 568724 221348 568730 221400
rect 121362 221280 121368 221332
rect 121420 221320 121426 221332
rect 190638 221320 190644 221332
rect 121420 221292 190644 221320
rect 121420 221280 121426 221292
rect 190638 221280 190644 221292
rect 190696 221280 190702 221332
rect 201402 221280 201408 221332
rect 201460 221320 201466 221332
rect 255406 221320 255412 221332
rect 201460 221292 255412 221320
rect 201460 221280 201466 221292
rect 255406 221280 255412 221292
rect 255464 221280 255470 221332
rect 282822 221280 282828 221332
rect 282880 221320 282886 221332
rect 283558 221320 283564 221332
rect 282880 221292 283564 221320
rect 282880 221280 282886 221292
rect 283558 221280 283564 221292
rect 283616 221280 283622 221332
rect 530946 221212 530952 221264
rect 531004 221252 531010 221264
rect 603350 221252 603356 221264
rect 531004 221224 603356 221252
rect 531004 221212 531010 221224
rect 603350 221212 603356 221224
rect 603408 221212 603414 221264
rect 667934 221212 667940 221264
rect 667992 221252 667998 221264
rect 670786 221252 670792 221264
rect 667992 221224 670792 221252
rect 667992 221212 667998 221224
rect 670786 221212 670792 221224
rect 670844 221212 670850 221264
rect 148686 221144 148692 221196
rect 148744 221184 148750 221196
rect 214098 221184 214104 221196
rect 148744 221156 214104 221184
rect 148744 221144 148750 221156
rect 214098 221144 214104 221156
rect 214156 221144 214162 221196
rect 215202 221144 215208 221196
rect 215260 221184 215266 221196
rect 263134 221184 263140 221196
rect 215260 221156 263140 221184
rect 215260 221144 215266 221156
rect 263134 221144 263140 221156
rect 263192 221144 263198 221196
rect 373994 221144 374000 221196
rect 374052 221184 374058 221196
rect 381078 221184 381084 221196
rect 374052 221156 381084 221184
rect 374052 221144 374058 221156
rect 381078 221144 381084 221156
rect 381136 221144 381142 221196
rect 527358 221076 527364 221128
rect 527416 221116 527422 221128
rect 528002 221116 528008 221128
rect 527416 221088 528008 221116
rect 527416 221076 527422 221088
rect 528002 221076 528008 221088
rect 528060 221116 528066 221128
rect 603534 221116 603540 221128
rect 528060 221088 603540 221116
rect 528060 221076 528066 221088
rect 603534 221076 603540 221088
rect 603592 221076 603598 221128
rect 141234 221008 141240 221060
rect 141292 221048 141298 221060
rect 205818 221048 205824 221060
rect 141292 221020 205824 221048
rect 141292 221008 141298 221020
rect 205818 221008 205824 221020
rect 205876 221008 205882 221060
rect 222562 221008 222568 221060
rect 222620 221048 222626 221060
rect 270862 221048 270868 221060
rect 222620 221020 270868 221048
rect 222620 221008 222626 221020
rect 270862 221008 270868 221020
rect 270920 221008 270926 221060
rect 387150 220940 387156 220992
rect 387208 220980 387214 220992
rect 389910 220980 389916 220992
rect 387208 220952 389916 220980
rect 387208 220940 387214 220952
rect 389910 220940 389916 220952
rect 389968 220940 389974 220992
rect 526438 220940 526444 220992
rect 526496 220980 526502 220992
rect 601786 220980 601792 220992
rect 526496 220952 601792 220980
rect 526496 220940 526502 220952
rect 601786 220940 601792 220952
rect 601844 220940 601850 220992
rect 161474 220872 161480 220924
rect 161532 220912 161538 220924
rect 169754 220912 169760 220924
rect 161532 220884 169760 220912
rect 161532 220872 161538 220884
rect 169754 220872 169760 220884
rect 169812 220872 169818 220924
rect 172514 220872 172520 220924
rect 172572 220912 172578 220924
rect 194962 220912 194968 220924
rect 172572 220884 194968 220912
rect 172572 220872 172578 220884
rect 194962 220872 194968 220884
rect 195020 220872 195026 220924
rect 228174 220872 228180 220924
rect 228232 220912 228238 220924
rect 276106 220912 276112 220924
rect 228232 220884 276112 220912
rect 228232 220872 228238 220884
rect 276106 220872 276112 220884
rect 276164 220872 276170 220924
rect 420638 220804 420644 220856
rect 420696 220844 420702 220856
rect 423858 220844 423864 220856
rect 420696 220816 423864 220844
rect 420696 220804 420702 220816
rect 423858 220804 423864 220816
rect 423916 220804 423922 220856
rect 521286 220804 521292 220856
rect 521344 220844 521350 220856
rect 600406 220844 600412 220856
rect 521344 220816 600412 220844
rect 521344 220804 521350 220816
rect 600406 220804 600412 220816
rect 600464 220804 600470 220856
rect 108114 220736 108120 220788
rect 108172 220776 108178 220788
rect 179966 220776 179972 220788
rect 108172 220748 179972 220776
rect 108172 220736 108178 220748
rect 179966 220736 179972 220748
rect 180024 220736 180030 220788
rect 187602 220736 187608 220788
rect 187660 220776 187666 220788
rect 241790 220776 241796 220788
rect 187660 220748 241796 220776
rect 187660 220736 187666 220748
rect 241790 220736 241796 220748
rect 241848 220736 241854 220788
rect 261294 220736 261300 220788
rect 261352 220776 261358 220788
rect 301774 220776 301780 220788
rect 261352 220748 301780 220776
rect 261352 220736 261358 220748
rect 301774 220736 301780 220748
rect 301832 220736 301838 220788
rect 313918 220736 313924 220788
rect 313976 220776 313982 220788
rect 320358 220776 320364 220788
rect 313976 220748 320364 220776
rect 313976 220736 313982 220748
rect 320358 220736 320364 220748
rect 320416 220736 320422 220788
rect 338942 220736 338948 220788
rect 339000 220776 339006 220788
rect 342438 220776 342444 220788
rect 339000 220748 342444 220776
rect 339000 220736 339006 220748
rect 342438 220736 342444 220748
rect 342496 220736 342502 220788
rect 455322 220736 455328 220788
rect 455380 220776 455386 220788
rect 458542 220776 458548 220788
rect 455380 220748 458548 220776
rect 455380 220736 455386 220748
rect 458542 220736 458548 220748
rect 458600 220736 458606 220788
rect 465718 220736 465724 220788
rect 465776 220776 465782 220788
rect 469306 220776 469312 220788
rect 465776 220748 469312 220776
rect 465776 220736 465782 220748
rect 469306 220736 469312 220748
rect 469364 220736 469370 220788
rect 476758 220736 476764 220788
rect 476816 220776 476822 220788
rect 478414 220776 478420 220788
rect 476816 220748 478420 220776
rect 476816 220736 476822 220748
rect 478414 220736 478420 220748
rect 478472 220736 478478 220788
rect 518158 220668 518164 220720
rect 518216 220708 518222 220720
rect 529842 220708 529848 220720
rect 518216 220680 529848 220708
rect 518216 220668 518222 220680
rect 529842 220668 529848 220680
rect 529900 220668 529906 220720
rect 534626 220668 534632 220720
rect 534684 220708 534690 220720
rect 534684 220680 534856 220708
rect 534684 220668 534690 220680
rect 66714 220600 66720 220652
rect 66772 220640 66778 220652
rect 144178 220640 144184 220652
rect 66772 220612 144184 220640
rect 66772 220600 66778 220612
rect 144178 220600 144184 220612
rect 144236 220600 144242 220652
rect 144546 220600 144552 220652
rect 144604 220640 144610 220652
rect 208578 220640 208584 220652
rect 144604 220612 208584 220640
rect 144604 220600 144610 220612
rect 208578 220600 208584 220612
rect 208636 220600 208642 220652
rect 216398 220600 216404 220652
rect 216456 220640 216462 220652
rect 217318 220640 217324 220652
rect 216456 220612 217324 220640
rect 216456 220600 216462 220612
rect 217318 220600 217324 220612
rect 217376 220600 217382 220652
rect 217502 220600 217508 220652
rect 217560 220640 217566 220652
rect 265066 220640 265072 220652
rect 217560 220612 265072 220640
rect 217560 220600 217566 220612
rect 265066 220600 265072 220612
rect 265124 220600 265130 220652
rect 277026 220600 277032 220652
rect 277084 220640 277090 220652
rect 311434 220640 311440 220652
rect 277084 220612 311440 220640
rect 277084 220600 277090 220612
rect 311434 220600 311440 220612
rect 311492 220600 311498 220652
rect 311618 220600 311624 220652
rect 311676 220640 311682 220652
rect 338574 220640 338580 220652
rect 311676 220612 338580 220640
rect 311676 220600 311682 220612
rect 338574 220600 338580 220612
rect 338632 220600 338638 220652
rect 534828 220572 534856 220680
rect 535086 220668 535092 220720
rect 535144 220708 535150 220720
rect 543734 220708 543740 220720
rect 535144 220680 543740 220708
rect 535144 220668 535150 220680
rect 543734 220668 543740 220680
rect 543792 220668 543798 220720
rect 544470 220668 544476 220720
rect 544528 220708 544534 220720
rect 551830 220708 551836 220720
rect 544528 220680 551836 220708
rect 544528 220668 544534 220680
rect 551830 220668 551836 220680
rect 551888 220668 551894 220720
rect 557994 220668 558000 220720
rect 558052 220708 558058 220720
rect 558546 220708 558552 220720
rect 558052 220680 558552 220708
rect 558052 220668 558058 220680
rect 558546 220668 558552 220680
rect 558604 220668 558610 220720
rect 559742 220668 559748 220720
rect 559800 220708 559806 220720
rect 563514 220708 563520 220720
rect 559800 220680 563520 220708
rect 559800 220668 559806 220680
rect 563514 220668 563520 220680
rect 563572 220668 563578 220720
rect 563698 220600 563704 220652
rect 563756 220640 563762 220652
rect 563756 220612 571518 220640
rect 563756 220600 563762 220612
rect 535454 220572 535460 220584
rect 534828 220544 535460 220572
rect 535454 220532 535460 220544
rect 535512 220532 535518 220584
rect 535730 220532 535736 220584
rect 535788 220572 535794 220584
rect 553302 220572 553308 220584
rect 535788 220544 553308 220572
rect 535788 220532 535794 220544
rect 553302 220532 553308 220544
rect 553360 220532 553366 220584
rect 553486 220532 553492 220584
rect 553544 220572 553550 220584
rect 558914 220572 558920 220584
rect 553544 220544 558920 220572
rect 553544 220532 553550 220544
rect 558914 220532 558920 220544
rect 558972 220532 558978 220584
rect 86586 220464 86592 220516
rect 86644 220504 86650 220516
rect 164326 220504 164332 220516
rect 86644 220476 164332 220504
rect 86644 220464 86650 220476
rect 164326 220464 164332 220476
rect 164384 220464 164390 220516
rect 180702 220464 180708 220516
rect 180760 220504 180766 220516
rect 180760 220476 231716 220504
rect 180760 220464 180766 220476
rect 79778 220328 79784 220380
rect 79836 220368 79842 220380
rect 158898 220368 158904 220380
rect 79836 220340 158904 220368
rect 79836 220328 79842 220340
rect 158898 220328 158904 220340
rect 158956 220328 158962 220380
rect 171042 220328 171048 220380
rect 171100 220368 171106 220380
rect 229094 220368 229100 220380
rect 171100 220340 229100 220368
rect 171100 220328 171106 220340
rect 229094 220328 229100 220340
rect 229152 220328 229158 220380
rect 231688 220368 231716 220476
rect 231854 220464 231860 220516
rect 231912 220504 231918 220516
rect 238018 220504 238024 220516
rect 231912 220476 238024 220504
rect 231912 220464 231918 220476
rect 238018 220464 238024 220476
rect 238076 220464 238082 220516
rect 246942 220464 246948 220516
rect 247000 220504 247006 220516
rect 288526 220504 288532 220516
rect 247000 220476 288532 220504
rect 247000 220464 247006 220476
rect 288526 220464 288532 220476
rect 288584 220464 288590 220516
rect 310146 220464 310152 220516
rect 310204 220504 310210 220516
rect 338206 220504 338212 220516
rect 310204 220476 338212 220504
rect 310204 220464 310210 220476
rect 338206 220464 338212 220476
rect 338264 220464 338270 220516
rect 342714 220464 342720 220516
rect 342772 220504 342778 220516
rect 352374 220504 352380 220516
rect 342772 220476 352380 220504
rect 342772 220464 342778 220476
rect 352374 220464 352380 220476
rect 352432 220464 352438 220516
rect 353202 220464 353208 220516
rect 353260 220504 353266 220516
rect 371418 220504 371424 220516
rect 353260 220476 371424 220504
rect 353260 220464 353266 220476
rect 371418 220464 371424 220476
rect 371476 220464 371482 220516
rect 432230 220464 432236 220516
rect 432288 220504 432294 220516
rect 434806 220504 434812 220516
rect 432288 220476 434812 220504
rect 432288 220464 432294 220476
rect 434806 220464 434812 220476
rect 434864 220464 434870 220516
rect 482922 220464 482928 220516
rect 482980 220504 482986 220516
rect 495342 220504 495348 220516
rect 482980 220476 495348 220504
rect 482980 220464 482986 220476
rect 495342 220464 495348 220476
rect 495400 220464 495406 220516
rect 500218 220464 500224 220516
rect 500276 220504 500282 220516
rect 509234 220504 509240 220516
rect 500276 220476 509240 220504
rect 500276 220464 500282 220476
rect 509234 220464 509240 220476
rect 509292 220464 509298 220516
rect 513282 220464 513288 220516
rect 513340 220504 513346 220516
rect 534626 220504 534632 220516
rect 513340 220476 534632 220504
rect 513340 220464 513346 220476
rect 534626 220464 534632 220476
rect 534684 220464 534690 220516
rect 562502 220464 562508 220516
rect 562560 220504 562566 220516
rect 571334 220504 571340 220516
rect 562560 220476 571340 220504
rect 562560 220464 562566 220476
rect 571334 220464 571340 220476
rect 571392 220464 571398 220516
rect 571490 220504 571518 220612
rect 571610 220600 571616 220652
rect 571668 220640 571674 220652
rect 611354 220640 611360 220652
rect 571668 220612 611360 220640
rect 571668 220600 571674 220612
rect 611354 220600 611360 220612
rect 611412 220600 611418 220652
rect 610526 220504 610532 220516
rect 571490 220476 610532 220504
rect 610526 220464 610532 220476
rect 610584 220464 610590 220516
rect 543734 220436 543740 220448
rect 543706 220396 543740 220436
rect 543792 220396 543798 220448
rect 552014 220396 552020 220448
rect 552072 220436 552078 220448
rect 552750 220436 552756 220448
rect 552072 220408 552756 220436
rect 552072 220396 552078 220408
rect 552750 220396 552756 220408
rect 552808 220436 552814 220448
rect 552808 220408 558132 220436
rect 552808 220396 552814 220408
rect 236638 220368 236644 220380
rect 231688 220340 236644 220368
rect 236638 220328 236644 220340
rect 236696 220328 236702 220380
rect 240594 220328 240600 220380
rect 240652 220368 240658 220380
rect 283098 220368 283104 220380
rect 240652 220340 283104 220368
rect 240652 220328 240658 220340
rect 283098 220328 283104 220340
rect 283156 220328 283162 220380
rect 299198 220328 299204 220380
rect 299256 220368 299262 220380
rect 331398 220368 331404 220380
rect 299256 220340 331404 220368
rect 299256 220328 299262 220340
rect 331398 220328 331404 220340
rect 331456 220328 331462 220380
rect 338022 220328 338028 220380
rect 338080 220368 338086 220380
rect 358998 220368 359004 220380
rect 338080 220340 359004 220368
rect 338080 220328 338086 220340
rect 358998 220328 359004 220340
rect 359056 220328 359062 220380
rect 372522 220328 372528 220380
rect 372580 220368 372586 220380
rect 385402 220368 385408 220380
rect 372580 220340 385408 220368
rect 372580 220328 372586 220340
rect 385402 220328 385408 220340
rect 385460 220328 385466 220380
rect 469122 220328 469128 220380
rect 469180 220368 469186 220380
rect 476114 220368 476120 220380
rect 469180 220340 476120 220368
rect 469180 220328 469186 220340
rect 476114 220328 476120 220340
rect 476172 220328 476178 220380
rect 485682 220328 485688 220380
rect 485740 220368 485746 220380
rect 499114 220368 499120 220380
rect 485740 220340 499120 220368
rect 485740 220328 485746 220340
rect 499114 220328 499120 220340
rect 499172 220328 499178 220380
rect 504358 220328 504364 220380
rect 504416 220368 504422 220380
rect 517698 220368 517704 220380
rect 504416 220340 517704 220368
rect 504416 220328 504422 220340
rect 517698 220328 517704 220340
rect 517756 220368 517762 220380
rect 518802 220368 518808 220380
rect 517756 220340 518808 220368
rect 517756 220328 517762 220340
rect 518802 220328 518808 220340
rect 518860 220328 518866 220380
rect 521562 220328 521568 220380
rect 521620 220368 521626 220380
rect 543706 220368 543734 220396
rect 521620 220340 543734 220368
rect 558104 220368 558132 220408
rect 608686 220368 608692 220380
rect 558104 220340 608692 220368
rect 521620 220328 521626 220340
rect 608686 220328 608692 220340
rect 608744 220328 608750 220380
rect 556246 220300 556252 220312
rect 548536 220272 556252 220300
rect 76374 220192 76380 220244
rect 76432 220232 76438 220244
rect 156138 220232 156144 220244
rect 76432 220204 156144 220232
rect 76432 220192 76438 220204
rect 156138 220192 156144 220204
rect 156196 220192 156202 220244
rect 161474 220192 161480 220244
rect 161532 220232 161538 220244
rect 161532 220204 219434 220232
rect 161532 220192 161538 220204
rect 73062 220056 73068 220108
rect 73120 220096 73126 220108
rect 153746 220096 153752 220108
rect 73120 220068 153752 220096
rect 73120 220056 73126 220068
rect 153746 220056 153752 220068
rect 153804 220056 153810 220108
rect 157794 220056 157800 220108
rect 157852 220096 157858 220108
rect 218606 220096 218612 220108
rect 157852 220068 218612 220096
rect 157852 220056 157858 220068
rect 218606 220056 218612 220068
rect 218664 220056 218670 220108
rect 219406 220096 219434 220204
rect 220814 220192 220820 220244
rect 220872 220232 220878 220244
rect 233418 220232 233424 220244
rect 220872 220204 233424 220232
rect 220872 220192 220878 220204
rect 233418 220192 233424 220204
rect 233476 220192 233482 220244
rect 237282 220192 237288 220244
rect 237340 220232 237346 220244
rect 280522 220232 280528 220244
rect 237340 220204 280528 220232
rect 237340 220192 237346 220204
rect 280522 220192 280528 220204
rect 280580 220192 280586 220244
rect 283650 220192 283656 220244
rect 283708 220232 283714 220244
rect 316586 220232 316592 220244
rect 283708 220204 316592 220232
rect 283708 220192 283714 220204
rect 316586 220192 316592 220204
rect 316644 220192 316650 220244
rect 329190 220192 329196 220244
rect 329248 220232 329254 220244
rect 354674 220232 354680 220244
rect 329248 220204 354680 220232
rect 329248 220192 329254 220204
rect 354674 220192 354680 220204
rect 354732 220192 354738 220244
rect 361482 220192 361488 220244
rect 361540 220232 361546 220244
rect 376846 220232 376852 220244
rect 361540 220204 376852 220232
rect 361540 220192 361546 220204
rect 376846 220192 376852 220204
rect 376904 220192 376910 220244
rect 377030 220192 377036 220244
rect 377088 220232 377094 220244
rect 388622 220232 388628 220244
rect 377088 220204 388628 220232
rect 377088 220192 377094 220204
rect 388622 220192 388628 220204
rect 388680 220192 388686 220244
rect 459462 220192 459468 220244
rect 459520 220232 459526 220244
rect 465166 220232 465172 220244
rect 459520 220204 465172 220232
rect 459520 220192 459526 220204
rect 465166 220192 465172 220204
rect 465224 220192 465230 220244
rect 473262 220192 473268 220244
rect 473320 220232 473326 220244
rect 481726 220232 481732 220244
rect 473320 220204 481732 220232
rect 473320 220192 473326 220204
rect 481726 220192 481732 220204
rect 481784 220192 481790 220244
rect 488166 220192 488172 220244
rect 488224 220232 488230 220244
rect 502426 220232 502432 220244
rect 488224 220204 502432 220232
rect 488224 220192 488230 220204
rect 502426 220192 502432 220204
rect 502484 220192 502490 220244
rect 507118 220192 507124 220244
rect 507176 220232 507182 220244
rect 521930 220232 521936 220244
rect 507176 220204 521936 220232
rect 507176 220192 507182 220204
rect 521930 220192 521936 220204
rect 521988 220192 521994 220244
rect 531222 220192 531228 220244
rect 531280 220232 531286 220244
rect 548536 220232 548564 220272
rect 556246 220260 556252 220272
rect 556304 220260 556310 220312
rect 531280 220204 548564 220232
rect 531280 220192 531286 220204
rect 558546 220192 558552 220244
rect 558604 220232 558610 220244
rect 609422 220232 609428 220244
rect 558604 220204 609428 220232
rect 558604 220192 558610 220204
rect 609422 220192 609428 220204
rect 609480 220192 609486 220244
rect 548702 220124 548708 220176
rect 548760 220164 548766 220176
rect 548760 220136 553900 220164
rect 548760 220124 548766 220136
rect 221274 220096 221280 220108
rect 219406 220068 221280 220096
rect 221274 220056 221280 220068
rect 221332 220056 221338 220108
rect 230198 220056 230204 220108
rect 230256 220096 230262 220108
rect 275278 220096 275284 220108
rect 230256 220068 275284 220096
rect 230256 220056 230262 220068
rect 275278 220056 275284 220068
rect 275336 220056 275342 220108
rect 280062 220056 280068 220108
rect 280120 220096 280126 220108
rect 313734 220096 313740 220108
rect 280120 220068 313740 220096
rect 280120 220056 280126 220068
rect 313734 220056 313740 220068
rect 313792 220056 313798 220108
rect 318426 220056 318432 220108
rect 318484 220096 318490 220108
rect 318484 220068 335354 220096
rect 318484 220056 318490 220068
rect 114462 219920 114468 219972
rect 114520 219960 114526 219972
rect 185118 219960 185124 219972
rect 114520 219932 185124 219960
rect 114520 219920 114526 219932
rect 185118 219920 185124 219932
rect 185176 219920 185182 219972
rect 200850 219920 200856 219972
rect 200908 219960 200914 219972
rect 252738 219960 252744 219972
rect 200908 219932 252744 219960
rect 200908 219920 200914 219932
rect 252738 219920 252744 219932
rect 252796 219920 252802 219972
rect 257154 219920 257160 219972
rect 257212 219960 257218 219972
rect 295978 219960 295984 219972
rect 257212 219932 295984 219960
rect 257212 219920 257218 219932
rect 295978 219920 295984 219932
rect 296036 219920 296042 219972
rect 335326 219960 335354 220068
rect 343634 220056 343640 220108
rect 343692 220096 343698 220108
rect 347866 220096 347872 220108
rect 343692 220068 347872 220096
rect 343692 220056 343698 220068
rect 347866 220056 347872 220068
rect 347924 220056 347930 220108
rect 354306 220056 354312 220108
rect 354364 220096 354370 220108
rect 372798 220096 372804 220108
rect 354364 220068 372804 220096
rect 354364 220056 354370 220068
rect 372798 220056 372804 220068
rect 372856 220056 372862 220108
rect 379422 220056 379428 220108
rect 379480 220096 379486 220108
rect 392118 220096 392124 220108
rect 379480 220068 392124 220096
rect 379480 220056 379486 220068
rect 392118 220056 392124 220068
rect 392176 220056 392182 220108
rect 395982 220056 395988 220108
rect 396040 220096 396046 220108
rect 404722 220096 404728 220108
rect 396040 220068 404728 220096
rect 396040 220056 396046 220068
rect 404722 220056 404728 220068
rect 404780 220056 404786 220108
rect 421926 220056 421932 220108
rect 421984 220096 421990 220108
rect 426802 220096 426808 220108
rect 421984 220068 426808 220096
rect 421984 220056 421990 220068
rect 426802 220056 426808 220068
rect 426860 220056 426866 220108
rect 475930 220056 475936 220108
rect 475988 220096 475994 220108
rect 485866 220096 485872 220108
rect 475988 220068 485872 220096
rect 475988 220056 475994 220068
rect 485866 220056 485872 220068
rect 485924 220056 485930 220108
rect 491662 220056 491668 220108
rect 491720 220096 491726 220108
rect 507762 220096 507768 220108
rect 491720 220068 507768 220096
rect 491720 220056 491726 220068
rect 507762 220056 507768 220068
rect 507820 220056 507826 220108
rect 511810 220056 511816 220108
rect 511868 220096 511874 220108
rect 531498 220096 531504 220108
rect 511868 220068 531504 220096
rect 511868 220056 511874 220068
rect 531498 220056 531504 220068
rect 531556 220056 531562 220108
rect 532510 220056 532516 220108
rect 532568 220096 532574 220108
rect 553872 220096 553900 220136
rect 532568 220068 543734 220096
rect 553872 220068 582374 220096
rect 532568 220056 532574 220068
rect 414474 219988 414480 220040
rect 414532 220028 414538 220040
rect 418338 220028 418344 220040
rect 414532 220000 418344 220028
rect 414532 219988 414538 220000
rect 418338 219988 418344 220000
rect 418396 219988 418402 220040
rect 543706 220028 543734 220068
rect 553486 220028 553492 220040
rect 543706 220000 553492 220028
rect 553486 219988 553492 220000
rect 553544 219988 553550 220040
rect 582346 220028 582374 220068
rect 592678 220056 592684 220108
rect 592736 220096 592742 220108
rect 633434 220096 633440 220108
rect 592736 220068 633440 220096
rect 592736 220056 592742 220068
rect 633434 220056 633440 220068
rect 633492 220056 633498 220108
rect 636470 220056 636476 220108
rect 636528 220096 636534 220108
rect 653398 220096 653404 220108
rect 636528 220068 653404 220096
rect 636528 220056 636534 220068
rect 653398 220056 653404 220068
rect 653456 220056 653462 220108
rect 675846 220056 675852 220108
rect 675904 220096 675910 220108
rect 676490 220096 676496 220108
rect 675904 220068 676496 220096
rect 675904 220056 675910 220068
rect 676490 220056 676496 220068
rect 676548 220056 676554 220108
rect 582558 220028 582564 220040
rect 582346 220000 582564 220028
rect 582558 219988 582564 220000
rect 582616 219988 582622 220040
rect 343818 219960 343824 219972
rect 335326 219932 343824 219960
rect 343818 219920 343824 219932
rect 343876 219920 343882 219972
rect 528554 219920 528560 219972
rect 528612 219960 528618 219972
rect 534258 219960 534264 219972
rect 528612 219932 534264 219960
rect 528612 219920 528618 219932
rect 534258 219920 534264 219932
rect 534316 219920 534322 219972
rect 542538 219852 542544 219904
rect 542596 219892 542602 219904
rect 543090 219892 543096 219904
rect 542596 219864 543096 219892
rect 542596 219852 542602 219864
rect 543090 219852 543096 219864
rect 543148 219892 543154 219904
rect 605834 219892 605840 219904
rect 543148 219864 605840 219892
rect 543148 219852 543154 219864
rect 605834 219852 605840 219864
rect 605892 219852 605898 219904
rect 127986 219784 127992 219836
rect 128044 219824 128050 219836
rect 195606 219824 195612 219836
rect 128044 219796 195612 219824
rect 128044 219784 128050 219796
rect 195606 219784 195612 219796
rect 195664 219784 195670 219836
rect 207474 219784 207480 219836
rect 207532 219824 207538 219836
rect 257338 219824 257344 219836
rect 207532 219796 257344 219824
rect 207532 219784 207538 219796
rect 257338 219784 257344 219796
rect 257396 219784 257402 219836
rect 288526 219784 288532 219836
rect 288584 219824 288590 219836
rect 310514 219824 310520 219836
rect 288584 219796 310520 219824
rect 288584 219784 288590 219796
rect 310514 219784 310520 219796
rect 310572 219784 310578 219836
rect 543734 219716 543740 219768
rect 543792 219756 543798 219768
rect 548702 219756 548708 219768
rect 543792 219728 548708 219756
rect 543792 219716 543798 219728
rect 548702 219716 548708 219728
rect 548760 219716 548766 219768
rect 551002 219716 551008 219768
rect 551060 219756 551066 219768
rect 607766 219756 607772 219768
rect 551060 219728 607772 219756
rect 551060 219716 551066 219728
rect 607766 219716 607772 219728
rect 607824 219716 607830 219768
rect 137922 219648 137928 219700
rect 137980 219688 137986 219700
rect 203150 219688 203156 219700
rect 137980 219660 203156 219688
rect 137980 219648 137986 219660
rect 203150 219648 203156 219660
rect 203208 219648 203214 219700
rect 236454 219648 236460 219700
rect 236512 219688 236518 219700
rect 261478 219688 261484 219700
rect 236512 219660 261484 219688
rect 236512 219648 236518 219660
rect 261478 219648 261484 219660
rect 261536 219648 261542 219700
rect 464982 219580 464988 219632
rect 465040 219620 465046 219632
rect 471974 219620 471980 219632
rect 465040 219592 471980 219620
rect 465040 219580 465046 219592
rect 471974 219580 471980 219592
rect 472032 219580 472038 219632
rect 545758 219580 545764 219632
rect 545816 219620 545822 219632
rect 606662 219620 606668 219632
rect 545816 219592 606668 219620
rect 545816 219580 545822 219592
rect 606662 219580 606668 219592
rect 606720 219580 606726 219632
rect 179506 219512 179512 219564
rect 179564 219552 179570 219564
rect 232038 219552 232044 219564
rect 179564 219524 232044 219552
rect 179564 219512 179570 219524
rect 232038 219512 232044 219524
rect 232096 219512 232102 219564
rect 235902 219512 235908 219564
rect 235960 219552 235966 219564
rect 243078 219552 243084 219564
rect 235960 219524 243084 219552
rect 235960 219512 235966 219524
rect 243078 219512 243084 219524
rect 243136 219512 243142 219564
rect 273070 219512 273076 219564
rect 273128 219552 273134 219564
rect 279234 219552 279240 219564
rect 273128 219524 279240 219552
rect 273128 219512 273134 219524
rect 279234 219512 279240 219524
rect 279292 219512 279298 219564
rect 406194 219512 406200 219564
rect 406252 219552 406258 219564
rect 412726 219552 412732 219564
rect 406252 219524 412732 219552
rect 406252 219512 406258 219524
rect 412726 219512 412732 219524
rect 412784 219512 412790 219564
rect 432046 219552 432052 219564
rect 429212 219524 432052 219552
rect 421006 219484 421012 219496
rect 418172 219456 421012 219484
rect 108298 219376 108304 219428
rect 108356 219416 108362 219428
rect 146846 219416 146852 219428
rect 108356 219388 146852 219416
rect 108356 219376 108362 219388
rect 146846 219376 146852 219388
rect 146904 219376 146910 219428
rect 153654 219376 153660 219428
rect 153712 219416 153718 219428
rect 160738 219416 160744 219428
rect 153712 219388 160744 219416
rect 153712 219376 153718 219388
rect 160738 219376 160744 219388
rect 160796 219376 160802 219428
rect 163590 219376 163596 219428
rect 163648 219416 163654 219428
rect 184198 219416 184204 219428
rect 163648 219388 184204 219416
rect 163648 219376 163654 219388
rect 184198 219376 184204 219388
rect 184256 219376 184262 219428
rect 192938 219376 192944 219428
rect 192996 219416 193002 219428
rect 233878 219416 233884 219428
rect 192996 219388 233884 219416
rect 192996 219376 193002 219388
rect 233878 219376 233884 219388
rect 233936 219376 233942 219428
rect 253014 219376 253020 219428
rect 253072 219416 253078 219428
rect 253072 219388 258074 219416
rect 253072 219376 253078 219388
rect 140038 219280 140044 219292
rect 103486 219252 140044 219280
rect 93578 219104 93584 219156
rect 93636 219144 93642 219156
rect 103486 219144 103514 219252
rect 140038 219240 140044 219252
rect 140096 219240 140102 219292
rect 147030 219240 147036 219292
rect 147088 219280 147094 219292
rect 189902 219280 189908 219292
rect 147088 219252 189908 219280
rect 147088 219240 147094 219252
rect 189902 219240 189908 219252
rect 189960 219240 189966 219292
rect 209682 219240 209688 219292
rect 209740 219280 209746 219292
rect 210418 219280 210424 219292
rect 209740 219252 210424 219280
rect 209740 219240 209746 219252
rect 210418 219240 210424 219252
rect 210476 219240 210482 219292
rect 214374 219240 214380 219292
rect 214432 219280 214438 219292
rect 253566 219280 253572 219292
rect 214432 219252 253572 219280
rect 214432 219240 214438 219252
rect 253566 219240 253572 219252
rect 253624 219240 253630 219292
rect 93636 219116 103514 219144
rect 93636 219104 93642 219116
rect 123846 219104 123852 219156
rect 123904 219144 123910 219156
rect 123904 219116 166304 219144
rect 123904 219104 123910 219116
rect 87414 218968 87420 219020
rect 87472 219008 87478 219020
rect 106918 219008 106924 219020
rect 87472 218980 106924 219008
rect 87472 218968 87478 218980
rect 106918 218968 106924 218980
rect 106976 218968 106982 219020
rect 107286 218968 107292 219020
rect 107344 219008 107350 219020
rect 107344 218980 113174 219008
rect 107344 218968 107350 218980
rect 100478 218832 100484 218884
rect 100536 218872 100542 218884
rect 108298 218872 108304 218884
rect 100536 218844 108304 218872
rect 100536 218832 100542 218844
rect 108298 218832 108304 218844
rect 108356 218832 108362 218884
rect 113146 218872 113174 218980
rect 113910 218968 113916 219020
rect 113968 219008 113974 219020
rect 166074 219008 166080 219020
rect 113968 218980 166080 219008
rect 113968 218968 113974 218980
rect 166074 218968 166080 218980
rect 166132 218968 166138 219020
rect 159266 218872 159272 218884
rect 113146 218844 159272 218872
rect 159266 218832 159272 218844
rect 159324 218832 159330 218884
rect 166276 218872 166304 219116
rect 183094 219104 183100 219156
rect 183152 219144 183158 219156
rect 189718 219144 189724 219156
rect 183152 219116 189724 219144
rect 183152 219104 183158 219116
rect 189718 219104 189724 219116
rect 189776 219104 189782 219156
rect 199838 219104 199844 219156
rect 199896 219144 199902 219156
rect 247126 219144 247132 219156
rect 199896 219116 247132 219144
rect 199896 219104 199902 219116
rect 247126 219104 247132 219116
rect 247184 219104 247190 219156
rect 258046 219144 258074 219388
rect 272518 219376 272524 219428
rect 272576 219416 272582 219428
rect 297358 219416 297364 219428
rect 272576 219388 297364 219416
rect 272576 219376 272582 219388
rect 297358 219376 297364 219388
rect 297416 219376 297422 219428
rect 323394 219376 323400 219428
rect 323452 219416 323458 219428
rect 324038 219416 324044 219428
rect 323452 219388 324044 219416
rect 323452 219376 323458 219388
rect 324038 219376 324044 219388
rect 324096 219376 324102 219428
rect 324222 219376 324228 219428
rect 324280 219416 324286 219428
rect 324866 219416 324872 219428
rect 324280 219388 324872 219416
rect 324280 219376 324286 219388
rect 324866 219376 324872 219388
rect 324924 219376 324930 219428
rect 325050 219376 325056 219428
rect 325108 219416 325114 219428
rect 325510 219416 325516 219428
rect 325108 219388 325516 219416
rect 325108 219376 325114 219388
rect 325510 219376 325516 219388
rect 325568 219376 325574 219428
rect 327718 219416 327724 219428
rect 325712 219388 327724 219416
rect 259178 219240 259184 219292
rect 259236 219280 259242 219292
rect 292298 219280 292304 219292
rect 259236 219252 292304 219280
rect 259236 219240 259242 219252
rect 292298 219240 292304 219252
rect 292356 219240 292362 219292
rect 307662 219240 307668 219292
rect 307720 219280 307726 219292
rect 325712 219280 325740 219388
rect 327718 219376 327724 219388
rect 327776 219376 327782 219428
rect 373626 219376 373632 219428
rect 373684 219416 373690 219428
rect 377030 219416 377036 219428
rect 373684 219388 377036 219416
rect 373684 219376 373690 219388
rect 377030 219376 377036 219388
rect 377088 219376 377094 219428
rect 417786 219376 417792 219428
rect 417844 219416 417850 219428
rect 418172 219416 418200 219456
rect 421006 219444 421012 219456
rect 421064 219444 421070 219496
rect 417844 219388 418200 219416
rect 417844 219376 417850 219388
rect 428274 219376 428280 219428
rect 428332 219416 428338 219428
rect 429212 219416 429240 219524
rect 432046 219512 432052 219524
rect 432104 219512 432110 219564
rect 528738 219552 528744 219564
rect 528526 219524 528744 219552
rect 521930 219444 521936 219496
rect 521988 219484 521994 219496
rect 522574 219484 522580 219496
rect 521988 219456 522580 219484
rect 521988 219444 521994 219456
rect 522574 219444 522580 219456
rect 522632 219484 522638 219496
rect 528526 219484 528554 219524
rect 528738 219512 528744 219524
rect 528796 219512 528802 219564
rect 522632 219456 528554 219484
rect 522632 219444 522638 219456
rect 540606 219444 540612 219496
rect 540664 219484 540670 219496
rect 606018 219484 606024 219496
rect 540664 219456 606024 219484
rect 540664 219444 540670 219456
rect 606018 219444 606024 219456
rect 606076 219444 606082 219496
rect 428332 219388 429240 219416
rect 428332 219376 428338 219388
rect 430206 219376 430212 219428
rect 430264 219416 430270 219428
rect 432690 219416 432696 219428
rect 430264 219388 432696 219416
rect 430264 219376 430270 219388
rect 432690 219376 432696 219388
rect 432748 219376 432754 219428
rect 676214 219376 676220 219428
rect 676272 219416 676278 219428
rect 678606 219416 678612 219428
rect 676272 219388 678612 219416
rect 676272 219376 676278 219388
rect 678606 219376 678612 219388
rect 678664 219376 678670 219428
rect 504542 219308 504548 219360
rect 504600 219348 504606 219360
rect 504600 219320 514616 219348
rect 504600 219308 504606 219320
rect 307720 219252 325740 219280
rect 307720 219240 307726 219252
rect 327534 219240 327540 219292
rect 327592 219280 327598 219292
rect 342714 219280 342720 219292
rect 327592 219252 342720 219280
rect 327592 219240 327598 219252
rect 342714 219240 342720 219252
rect 342772 219240 342778 219292
rect 354582 219240 354588 219292
rect 354640 219280 354646 219292
rect 355318 219280 355324 219292
rect 354640 219252 355324 219280
rect 354640 219240 354646 219252
rect 355318 219240 355324 219252
rect 355376 219240 355382 219292
rect 457990 219240 457996 219292
rect 458048 219280 458054 219292
rect 461118 219280 461124 219292
rect 458048 219252 461124 219280
rect 458048 219240 458054 219252
rect 461118 219240 461124 219252
rect 461176 219240 461182 219292
rect 258046 219116 287054 219144
rect 166626 218968 166632 219020
rect 166684 219008 166690 219020
rect 173158 219008 173164 219020
rect 166684 218980 173164 219008
rect 166684 218968 166690 218980
rect 173158 218968 173164 218980
rect 173216 218968 173222 219020
rect 173526 218968 173532 219020
rect 173584 219008 173590 219020
rect 173584 218980 178908 219008
rect 173584 218968 173590 218980
rect 172514 218872 172520 218884
rect 166276 218844 172520 218872
rect 172514 218832 172520 218844
rect 172572 218832 172578 218884
rect 174906 218832 174912 218884
rect 174964 218872 174970 218884
rect 178678 218872 178684 218884
rect 174964 218844 178684 218872
rect 174964 218832 174970 218844
rect 178678 218832 178684 218844
rect 178736 218832 178742 218884
rect 178880 218872 178908 218980
rect 179322 218968 179328 219020
rect 179380 219008 179386 219020
rect 182818 219008 182824 219020
rect 179380 218980 182824 219008
rect 179380 218968 179386 218980
rect 182818 218968 182824 218980
rect 182876 218968 182882 219020
rect 186774 218968 186780 219020
rect 186832 219008 186838 219020
rect 235902 219008 235908 219020
rect 186832 218980 235908 219008
rect 186832 218968 186838 218980
rect 235902 218968 235908 218980
rect 235960 218968 235966 219020
rect 238110 218968 238116 219020
rect 238168 219008 238174 219020
rect 239398 219008 239404 219020
rect 238168 218980 239404 219008
rect 238168 218968 238174 218980
rect 239398 218968 239404 218980
rect 239456 218968 239462 219020
rect 239766 218968 239772 219020
rect 239824 219008 239830 219020
rect 246482 219008 246488 219020
rect 239824 218980 246488 219008
rect 239824 218968 239830 218980
rect 246482 218968 246488 218980
rect 246540 218968 246546 219020
rect 249242 218968 249248 219020
rect 249300 219008 249306 219020
rect 284018 219008 284024 219020
rect 249300 218980 284024 219008
rect 249300 218968 249306 218980
rect 284018 218968 284024 218980
rect 284076 218968 284082 219020
rect 287026 219008 287054 219116
rect 300578 219104 300584 219156
rect 300636 219144 300642 219156
rect 322842 219144 322848 219156
rect 300636 219116 322848 219144
rect 300636 219104 300642 219116
rect 322842 219104 322848 219116
rect 322900 219104 322906 219156
rect 325602 219104 325608 219156
rect 325660 219144 325666 219156
rect 330478 219144 330484 219156
rect 325660 219116 330484 219144
rect 325660 219104 325666 219116
rect 330478 219104 330484 219116
rect 330536 219104 330542 219156
rect 363966 219104 363972 219156
rect 364024 219144 364030 219156
rect 373994 219144 374000 219156
rect 364024 219116 374000 219144
rect 364024 219104 364030 219116
rect 373994 219104 374000 219116
rect 374052 219104 374058 219156
rect 388806 219104 388812 219156
rect 388864 219144 388870 219156
rect 393958 219144 393964 219156
rect 388864 219116 393964 219144
rect 388864 219104 388870 219116
rect 393958 219104 393964 219116
rect 394016 219104 394022 219156
rect 419258 219104 419264 219156
rect 419316 219144 419322 219156
rect 422662 219144 422668 219156
rect 419316 219116 422668 219144
rect 419316 219104 419322 219116
rect 422662 219104 422668 219116
rect 422720 219104 422726 219156
rect 496906 219104 496912 219156
rect 496964 219144 496970 219156
rect 504726 219144 504732 219156
rect 496964 219116 504732 219144
rect 496964 219104 496970 219116
rect 504726 219104 504732 219116
rect 504784 219104 504790 219156
rect 289078 219008 289084 219020
rect 287026 218980 289084 219008
rect 289078 218968 289084 218980
rect 289136 218968 289142 219020
rect 294414 218968 294420 219020
rect 294472 219008 294478 219020
rect 309778 219008 309784 219020
rect 294472 218980 309784 219008
rect 294472 218968 294478 218980
rect 309778 218968 309784 218980
rect 309836 218968 309842 219020
rect 314286 218968 314292 219020
rect 314344 219008 314350 219020
rect 338942 219008 338948 219020
rect 314344 218980 338948 219008
rect 314344 218968 314350 218980
rect 338942 218968 338948 218980
rect 339000 218968 339006 219020
rect 340506 218968 340512 219020
rect 340564 219008 340570 219020
rect 351178 219008 351184 219020
rect 340564 218980 351184 219008
rect 340564 218968 340570 218980
rect 351178 218968 351184 218980
rect 351236 218968 351242 219020
rect 383562 218968 383568 219020
rect 383620 219008 383626 219020
rect 388438 219008 388444 219020
rect 383620 218980 388444 219008
rect 383620 218968 383626 218980
rect 388438 218968 388444 218980
rect 388496 218968 388502 219020
rect 407574 218968 407580 219020
rect 407632 219008 407638 219020
rect 411898 219008 411904 219020
rect 407632 218980 411904 219008
rect 407632 218968 407638 218980
rect 411898 218968 411904 218980
rect 411956 218968 411962 219020
rect 499850 218900 499856 218952
rect 499908 218940 499914 218952
rect 499908 218912 506796 218940
rect 499908 218900 499914 218912
rect 214558 218872 214564 218884
rect 178880 218844 214564 218872
rect 214558 218832 214564 218844
rect 214616 218832 214622 218884
rect 232958 218832 232964 218884
rect 233016 218872 233022 218884
rect 273070 218872 273076 218884
rect 233016 218844 273076 218872
rect 233016 218832 233022 218844
rect 273070 218832 273076 218844
rect 273128 218832 273134 218884
rect 286134 218832 286140 218884
rect 286192 218872 286198 218884
rect 313918 218872 313924 218884
rect 286192 218844 313924 218872
rect 286192 218832 286198 218844
rect 313918 218832 313924 218844
rect 313976 218832 313982 218884
rect 343634 218872 343640 218884
rect 331186 218844 343640 218872
rect 59814 218696 59820 218748
rect 59872 218736 59878 218748
rect 68186 218736 68192 218748
rect 59872 218708 68192 218736
rect 59872 218696 59878 218708
rect 68186 218696 68192 218708
rect 68244 218696 68250 218748
rect 83918 218696 83924 218748
rect 83976 218736 83982 218748
rect 160186 218736 160192 218748
rect 83976 218708 160192 218736
rect 83976 218696 83982 218708
rect 160186 218696 160192 218708
rect 160244 218696 160250 218748
rect 162762 218696 162768 218748
rect 162820 218736 162826 218748
rect 169018 218736 169024 218748
rect 162820 218708 169024 218736
rect 162820 218696 162826 218708
rect 169018 218696 169024 218708
rect 169076 218696 169082 218748
rect 174354 218696 174360 218748
rect 174412 218736 174418 218748
rect 179506 218736 179512 218748
rect 174412 218708 179512 218736
rect 174412 218696 174418 218708
rect 179506 218696 179512 218708
rect 179564 218696 179570 218748
rect 180150 218696 180156 218748
rect 180208 218736 180214 218748
rect 231854 218736 231860 218748
rect 180208 218708 231860 218736
rect 180208 218696 180214 218708
rect 231854 218696 231860 218708
rect 231912 218696 231918 218748
rect 233878 218696 233884 218748
rect 233936 218736 233942 218748
rect 238846 218736 238852 218748
rect 233936 218708 238852 218736
rect 233936 218696 233942 218708
rect 238846 218696 238852 218708
rect 238904 218696 238910 218748
rect 244734 218696 244740 218748
rect 244792 218736 244798 218748
rect 246298 218736 246304 218748
rect 244792 218708 246304 218736
rect 244792 218696 244798 218708
rect 246298 218696 246304 218708
rect 246356 218696 246362 218748
rect 246482 218696 246488 218748
rect 246540 218736 246546 218748
rect 280798 218736 280804 218748
rect 246540 218708 280804 218736
rect 246540 218696 246546 218708
rect 280798 218696 280804 218708
rect 280856 218696 280862 218748
rect 291930 218696 291936 218748
rect 291988 218736 291994 218748
rect 323578 218736 323584 218748
rect 291988 218708 323584 218736
rect 291988 218696 291994 218708
rect 323578 218696 323584 218708
rect 323636 218696 323642 218748
rect 120534 218560 120540 218612
rect 120592 218600 120598 218612
rect 166442 218600 166448 218612
rect 120592 218572 166448 218600
rect 120592 218560 120598 218572
rect 166442 218560 166448 218572
rect 166500 218560 166506 218612
rect 170214 218560 170220 218612
rect 170272 218600 170278 218612
rect 200666 218600 200672 218612
rect 170272 218572 200672 218600
rect 170272 218560 170278 218572
rect 200666 218560 200672 218572
rect 200724 218560 200730 218612
rect 206646 218560 206652 218612
rect 206704 218600 206710 218612
rect 214374 218600 214380 218612
rect 206704 218572 214380 218600
rect 206704 218560 206710 218572
rect 214374 218560 214380 218572
rect 214432 218560 214438 218612
rect 214742 218560 214748 218612
rect 214800 218600 214806 218612
rect 260098 218600 260104 218612
rect 214800 218572 260104 218600
rect 214800 218560 214806 218572
rect 260098 218560 260104 218572
rect 260156 218560 260162 218612
rect 262950 218560 262956 218612
rect 263008 218600 263014 218612
rect 276658 218600 276664 218612
rect 263008 218572 276664 218600
rect 263008 218560 263014 218572
rect 276658 218560 276664 218572
rect 276716 218560 276722 218612
rect 279510 218560 279516 218612
rect 279568 218600 279574 218612
rect 279568 218572 296714 218600
rect 279568 218560 279574 218572
rect 137094 218424 137100 218476
rect 137152 218464 137158 218476
rect 174906 218464 174912 218476
rect 137152 218436 174912 218464
rect 137152 218424 137158 218436
rect 174906 218424 174912 218436
rect 174964 218424 174970 218476
rect 176286 218424 176292 218476
rect 176344 218464 176350 218476
rect 183094 218464 183100 218476
rect 176344 218436 183100 218464
rect 176344 218424 176350 218436
rect 183094 218424 183100 218436
rect 183152 218424 183158 218476
rect 183278 218424 183284 218476
rect 183336 218464 183342 218476
rect 202138 218464 202144 218476
rect 183336 218436 202144 218464
rect 183336 218424 183342 218436
rect 202138 218424 202144 218436
rect 202196 218424 202202 218476
rect 203334 218424 203340 218476
rect 203392 218464 203398 218476
rect 213086 218464 213092 218476
rect 203392 218436 213092 218464
rect 203392 218424 203398 218436
rect 213086 218424 213092 218436
rect 213144 218424 213150 218476
rect 214558 218424 214564 218476
rect 214616 218464 214622 218476
rect 220814 218464 220820 218476
rect 214616 218436 220820 218464
rect 214616 218424 214622 218436
rect 220814 218424 220820 218436
rect 220872 218424 220878 218476
rect 225966 218424 225972 218476
rect 226024 218464 226030 218476
rect 265618 218464 265624 218476
rect 226024 218436 265624 218464
rect 226024 218424 226030 218436
rect 265618 218424 265624 218436
rect 265676 218424 265682 218476
rect 266078 218424 266084 218476
rect 266136 218464 266142 218476
rect 272518 218464 272524 218476
rect 266136 218436 272524 218464
rect 266136 218424 266142 218436
rect 272518 218424 272524 218436
rect 272576 218424 272582 218476
rect 272886 218424 272892 218476
rect 272944 218464 272950 218476
rect 288526 218464 288532 218476
rect 272944 218436 288532 218464
rect 272944 218424 272950 218436
rect 288526 218424 288532 218436
rect 288584 218424 288590 218476
rect 296686 218464 296714 218572
rect 320910 218560 320916 218612
rect 320968 218600 320974 218612
rect 331186 218600 331214 218844
rect 343634 218832 343640 218844
rect 343692 218832 343698 218884
rect 347406 218832 347412 218884
rect 347464 218872 347470 218884
rect 363598 218872 363604 218884
rect 347464 218844 363604 218872
rect 347464 218832 347470 218844
rect 363598 218832 363604 218844
rect 363656 218832 363662 218884
rect 402054 218832 402060 218884
rect 402112 218872 402118 218884
rect 407758 218872 407764 218884
rect 402112 218844 407764 218872
rect 402112 218832 402118 218844
rect 407758 218832 407764 218844
rect 407816 218832 407822 218884
rect 411990 218832 411996 218884
rect 412048 218872 412054 218884
rect 412542 218872 412548 218884
rect 412048 218844 412548 218872
rect 412048 218832 412054 218844
rect 412542 218832 412548 218844
rect 412600 218832 412606 218884
rect 333698 218696 333704 218748
rect 333756 218736 333762 218748
rect 352558 218736 352564 218748
rect 333756 218708 352564 218736
rect 333756 218696 333762 218708
rect 352558 218696 352564 218708
rect 352616 218696 352622 218748
rect 354030 218696 354036 218748
rect 354088 218736 354094 218748
rect 367738 218736 367744 218748
rect 354088 218708 367744 218736
rect 354088 218696 354094 218708
rect 367738 218696 367744 218708
rect 367796 218696 367802 218748
rect 386138 218696 386144 218748
rect 386196 218736 386202 218748
rect 396718 218736 396724 218748
rect 386196 218708 396724 218736
rect 386196 218696 386202 218708
rect 396718 218696 396724 218708
rect 396776 218696 396782 218748
rect 402698 218696 402704 218748
rect 402756 218736 402762 218748
rect 409138 218736 409144 218748
rect 402756 218708 409144 218736
rect 402756 218696 402762 218708
rect 409138 218696 409144 218708
rect 409196 218696 409202 218748
rect 412542 218696 412548 218748
rect 412600 218736 412606 218748
rect 417142 218736 417148 218748
rect 412600 218708 417148 218736
rect 412600 218696 412606 218708
rect 417142 218696 417148 218708
rect 417200 218696 417206 218748
rect 484854 218696 484860 218748
rect 484912 218736 484918 218748
rect 506290 218736 506296 218748
rect 484912 218708 506296 218736
rect 484912 218696 484918 218708
rect 506290 218696 506296 218708
rect 506348 218696 506354 218748
rect 320968 218572 331214 218600
rect 320968 218560 320974 218572
rect 392946 218560 392952 218612
rect 393004 218600 393010 218612
rect 400858 218600 400864 218612
rect 393004 218572 400864 218600
rect 393004 218560 393010 218572
rect 400858 218560 400864 218572
rect 400916 218560 400922 218612
rect 504726 218560 504732 218612
rect 504784 218600 504790 218612
rect 505278 218600 505284 218612
rect 504784 218572 505284 218600
rect 504784 218560 504790 218572
rect 505278 218560 505284 218572
rect 505336 218560 505342 218612
rect 506768 218600 506796 218912
rect 514588 218804 514616 219320
rect 534074 219308 534080 219360
rect 534132 219348 534138 219360
rect 543918 219348 543924 219360
rect 534132 219320 543924 219348
rect 534132 219308 534138 219320
rect 543918 219308 543924 219320
rect 543976 219308 543982 219360
rect 553118 219308 553124 219360
rect 553176 219348 553182 219360
rect 553176 219320 572714 219348
rect 553176 219308 553182 219320
rect 572686 219280 572714 219320
rect 582466 219308 582472 219360
rect 582524 219348 582530 219360
rect 596818 219348 596824 219360
rect 582524 219320 596824 219348
rect 582524 219308 582530 219320
rect 596818 219308 596824 219320
rect 596876 219308 596882 219360
rect 579430 219280 579436 219292
rect 572686 219252 579436 219280
rect 579430 219240 579436 219252
rect 579488 219240 579494 219292
rect 579706 219240 579712 219292
rect 579764 219280 579770 219292
rect 579764 219252 582374 219280
rect 579764 219240 579770 219252
rect 524046 219172 524052 219224
rect 524104 219212 524110 219224
rect 528462 219212 528468 219224
rect 524104 219184 528468 219212
rect 524104 219172 524110 219184
rect 528462 219172 528468 219184
rect 528520 219172 528526 219224
rect 544654 219172 544660 219224
rect 544712 219212 544718 219224
rect 558362 219212 558368 219224
rect 544712 219184 558368 219212
rect 544712 219172 544718 219184
rect 558362 219172 558368 219184
rect 558420 219172 558426 219224
rect 563238 219172 563244 219224
rect 563296 219212 563302 219224
rect 563698 219212 563704 219224
rect 563296 219184 563704 219212
rect 563296 219172 563302 219184
rect 563698 219172 563704 219184
rect 563756 219172 563762 219224
rect 564434 219172 564440 219224
rect 564492 219212 564498 219224
rect 565170 219212 565176 219224
rect 564492 219184 565176 219212
rect 564492 219172 564498 219184
rect 565170 219172 565176 219184
rect 565228 219172 565234 219224
rect 582346 219212 582374 219252
rect 583110 219212 583116 219224
rect 582346 219184 583116 219212
rect 583110 219172 583116 219184
rect 583168 219172 583174 219224
rect 534258 219104 534264 219156
rect 534316 219144 534322 219156
rect 544286 219144 544292 219156
rect 534316 219116 544292 219144
rect 534316 219104 534322 219116
rect 544286 219104 544292 219116
rect 544344 219104 544350 219156
rect 562778 219104 562784 219156
rect 562836 219144 562842 219156
rect 563054 219144 563060 219156
rect 562836 219116 563060 219144
rect 562836 219104 562842 219116
rect 563054 219104 563060 219116
rect 563112 219104 563118 219156
rect 567010 219104 567016 219156
rect 567068 219144 567074 219156
rect 577498 219144 577504 219156
rect 567068 219116 577504 219144
rect 567068 219104 567074 219116
rect 577498 219104 577504 219116
rect 577556 219104 577562 219156
rect 547414 219036 547420 219088
rect 547472 219076 547478 219088
rect 558178 219076 558184 219088
rect 547472 219048 558184 219076
rect 547472 219036 547478 219048
rect 558178 219036 558184 219048
rect 558236 219036 558242 219088
rect 558380 219048 558500 219076
rect 514754 218900 514760 218952
rect 514812 218940 514818 218952
rect 524046 218940 524052 218952
rect 514812 218912 524052 218940
rect 514812 218900 514818 218912
rect 524046 218900 524052 218912
rect 524104 218900 524110 218952
rect 534074 218900 534080 218952
rect 534132 218940 534138 218952
rect 543642 218940 543648 218952
rect 534132 218912 543648 218940
rect 534132 218900 534138 218912
rect 543642 218900 543648 218912
rect 543700 218900 543706 218952
rect 543918 218900 543924 218952
rect 543976 218940 543982 218952
rect 543976 218912 544148 218940
rect 543976 218900 543982 218912
rect 528278 218832 528284 218884
rect 528336 218872 528342 218884
rect 529014 218872 529020 218884
rect 528336 218844 529020 218872
rect 528336 218832 528342 218844
rect 529014 218832 529020 218844
rect 529072 218832 529078 218884
rect 514588 218776 514754 218804
rect 514726 218736 514754 218776
rect 543458 218764 543464 218816
rect 543516 218804 543522 218816
rect 543918 218804 543924 218816
rect 543516 218776 543924 218804
rect 543516 218764 543522 218776
rect 543918 218764 543924 218776
rect 543976 218764 543982 218816
rect 544120 218804 544148 218912
rect 552566 218900 552572 218952
rect 552624 218940 552630 218952
rect 553854 218940 553860 218952
rect 552624 218912 553860 218940
rect 552624 218900 552630 218912
rect 553854 218900 553860 218912
rect 553912 218900 553918 218952
rect 555326 218900 555332 218952
rect 555384 218940 555390 218952
rect 558380 218940 558408 219048
rect 558472 219008 558500 219048
rect 567470 219008 567476 219020
rect 558472 218980 567476 219008
rect 567470 218968 567476 218980
rect 567528 218968 567534 219020
rect 567654 218968 567660 219020
rect 567712 219008 567718 219020
rect 572162 219008 572168 219020
rect 567712 218980 572168 219008
rect 567712 218968 567718 218980
rect 572162 218968 572168 218980
rect 572220 218968 572226 219020
rect 572318 218980 576440 219008
rect 555384 218912 558408 218940
rect 555384 218900 555390 218912
rect 558730 218832 558736 218884
rect 558788 218872 558794 218884
rect 568114 218872 568120 218884
rect 558788 218844 568120 218872
rect 558788 218832 558794 218844
rect 568114 218832 568120 218844
rect 568172 218832 568178 218884
rect 568298 218832 568304 218884
rect 568356 218872 568362 218884
rect 572318 218872 572346 218980
rect 568356 218844 572346 218872
rect 568356 218832 568362 218844
rect 572438 218832 572444 218884
rect 572496 218872 572502 218884
rect 576210 218872 576216 218884
rect 572496 218844 576216 218872
rect 572496 218832 572502 218844
rect 576210 218832 576216 218844
rect 576268 218832 576274 218884
rect 553302 218804 553308 218816
rect 544120 218776 553308 218804
rect 553302 218764 553308 218776
rect 553360 218764 553366 218816
rect 523954 218736 523960 218748
rect 514726 218708 523960 218736
rect 523954 218696 523960 218708
rect 524012 218696 524018 218748
rect 531958 218696 531964 218748
rect 532016 218736 532022 218748
rect 532602 218736 532608 218748
rect 532016 218708 532608 218736
rect 532016 218696 532022 218708
rect 532602 218696 532608 218708
rect 532660 218736 532666 218748
rect 532660 218708 538904 218736
rect 532660 218696 532666 218708
rect 528278 218628 528284 218680
rect 528336 218668 528342 218680
rect 528336 218640 528554 218668
rect 528336 218628 528342 218640
rect 514938 218600 514944 218612
rect 506768 218572 514944 218600
rect 514938 218560 514944 218572
rect 514996 218560 515002 218612
rect 528526 218600 528554 218640
rect 534258 218600 534264 218612
rect 528526 218572 534264 218600
rect 534258 218560 534264 218572
rect 534316 218560 534322 218612
rect 469858 218492 469864 218544
rect 469916 218532 469922 218544
rect 470962 218532 470968 218544
rect 469916 218504 470968 218532
rect 469916 218492 469922 218504
rect 470962 218492 470968 218504
rect 471020 218492 471026 218544
rect 307018 218464 307024 218476
rect 296686 218436 307024 218464
rect 307018 218424 307024 218436
rect 307076 218424 307082 218476
rect 365346 218424 365352 218476
rect 365404 218464 365410 218476
rect 370498 218464 370504 218476
rect 365404 218436 370504 218464
rect 365404 218424 365410 218436
rect 370498 218424 370504 218436
rect 370556 218424 370562 218476
rect 523770 218424 523776 218476
rect 523828 218464 523834 218476
rect 528462 218464 528468 218476
rect 523828 218436 528468 218464
rect 523828 218424 523834 218436
rect 528462 218424 528468 218436
rect 528520 218424 528526 218476
rect 528646 218424 528652 218476
rect 528704 218464 528710 218476
rect 534442 218464 534448 218476
rect 528704 218436 534448 218464
rect 528704 218424 528710 218436
rect 534442 218424 534448 218436
rect 534500 218424 534506 218476
rect 538876 218464 538904 218708
rect 553486 218696 553492 218748
rect 553544 218736 553550 218748
rect 563054 218736 563060 218748
rect 553544 218708 563060 218736
rect 553544 218696 553550 218708
rect 563054 218696 563060 218708
rect 563112 218696 563118 218748
rect 576210 218736 576216 218748
rect 567580 218708 576216 218736
rect 543458 218560 543464 218612
rect 543516 218600 543522 218612
rect 544102 218600 544108 218612
rect 543516 218572 544108 218600
rect 543516 218560 543522 218572
rect 544102 218560 544108 218572
rect 544160 218560 544166 218612
rect 544286 218560 544292 218612
rect 544344 218600 544350 218612
rect 552934 218600 552940 218612
rect 544344 218572 552940 218600
rect 544344 218560 544350 218572
rect 552934 218560 552940 218572
rect 552992 218560 552998 218612
rect 553118 218560 553124 218612
rect 553176 218600 553182 218612
rect 553854 218600 553860 218612
rect 553176 218572 553860 218600
rect 553176 218560 553182 218572
rect 553854 218560 553860 218572
rect 553912 218560 553918 218612
rect 558178 218560 558184 218612
rect 558236 218600 558242 218612
rect 567580 218600 567608 218708
rect 576210 218696 576216 218708
rect 576268 218696 576274 218748
rect 576412 218736 576440 218980
rect 576578 218968 576584 219020
rect 576636 219008 576642 219020
rect 577682 219008 577688 219020
rect 576636 218980 577688 219008
rect 576636 218968 576642 218980
rect 577682 218968 577688 218980
rect 577740 218968 577746 219020
rect 576578 218832 576584 218884
rect 576636 218872 576642 218884
rect 582374 218872 582380 218884
rect 576636 218844 582380 218872
rect 576636 218832 576642 218844
rect 582374 218832 582380 218844
rect 582432 218832 582438 218884
rect 595898 218832 595904 218884
rect 595956 218872 595962 218884
rect 597554 218872 597560 218884
rect 595956 218844 597560 218872
rect 595956 218832 595962 218844
rect 597554 218832 597560 218844
rect 597612 218832 597618 218884
rect 611814 218736 611820 218748
rect 576412 218708 611820 218736
rect 611814 218696 611820 218708
rect 611872 218696 611878 218748
rect 558236 218572 567608 218600
rect 558236 218560 558242 218572
rect 567746 218560 567752 218612
rect 567804 218600 567810 218612
rect 577866 218600 577872 218612
rect 567804 218572 577872 218600
rect 567804 218560 567810 218572
rect 577866 218560 577872 218572
rect 577924 218560 577930 218612
rect 578050 218464 578056 218476
rect 538876 218436 578056 218464
rect 578050 218424 578056 218436
rect 578108 218424 578114 218476
rect 582374 218424 582380 218476
rect 582432 218464 582438 218476
rect 596082 218464 596088 218476
rect 582432 218436 596088 218464
rect 582432 218424 582438 218436
rect 596082 218424 596088 218436
rect 596140 218424 596146 218476
rect 450538 218356 450544 218408
rect 450596 218396 450602 218408
rect 453574 218396 453580 218408
rect 450596 218368 453580 218396
rect 450596 218356 450602 218368
rect 453574 218356 453580 218368
rect 453632 218356 453638 218408
rect 57606 218288 57612 218340
rect 57664 218328 57670 218340
rect 64138 218328 64144 218340
rect 57664 218300 64144 218328
rect 57664 218288 57670 218300
rect 64138 218288 64144 218300
rect 64196 218288 64202 218340
rect 68738 218288 68744 218340
rect 68796 218328 68802 218340
rect 72418 218328 72424 218340
rect 68796 218300 72424 218328
rect 68796 218288 68802 218300
rect 72418 218288 72424 218300
rect 72476 218288 72482 218340
rect 159818 218288 159824 218340
rect 159876 218328 159882 218340
rect 196802 218328 196808 218340
rect 159876 218300 196808 218328
rect 159876 218288 159882 218300
rect 196802 218288 196808 218300
rect 196860 218288 196866 218340
rect 199194 218288 199200 218340
rect 199252 218328 199258 218340
rect 200022 218328 200028 218340
rect 199252 218300 200028 218328
rect 199252 218288 199258 218300
rect 200022 218288 200028 218300
rect 200080 218288 200086 218340
rect 203886 218288 203892 218340
rect 203944 218328 203950 218340
rect 207658 218328 207664 218340
rect 203944 218300 207664 218328
rect 203944 218288 203950 218300
rect 207658 218288 207664 218300
rect 207716 218288 207722 218340
rect 213270 218288 213276 218340
rect 213328 218328 213334 218340
rect 214742 218328 214748 218340
rect 213328 218300 214748 218328
rect 213328 218288 213334 218300
rect 214742 218288 214748 218300
rect 214800 218288 214806 218340
rect 219894 218288 219900 218340
rect 219952 218328 219958 218340
rect 258074 218328 258080 218340
rect 219952 218300 258080 218328
rect 219952 218288 219958 218300
rect 258074 218288 258080 218300
rect 258132 218288 258138 218340
rect 344094 218288 344100 218340
rect 344152 218328 344158 218340
rect 347038 218328 347044 218340
rect 344152 218300 347044 218328
rect 344152 218288 344158 218300
rect 347038 218288 347044 218300
rect 347096 218288 347102 218340
rect 370590 218288 370596 218340
rect 370648 218328 370654 218340
rect 375466 218328 375472 218340
rect 370648 218300 375472 218328
rect 370648 218288 370654 218300
rect 375466 218288 375472 218300
rect 375524 218288 375530 218340
rect 377214 218288 377220 218340
rect 377272 218328 377278 218340
rect 385678 218328 385684 218340
rect 377272 218300 385684 218328
rect 377272 218288 377278 218300
rect 385678 218288 385684 218300
rect 385736 218288 385742 218340
rect 426802 218288 426808 218340
rect 426860 218328 426866 218340
rect 429562 218328 429568 218340
rect 426860 218300 429568 218328
rect 426860 218288 426866 218300
rect 429562 218288 429568 218300
rect 429620 218288 429626 218340
rect 479518 218288 479524 218340
rect 479576 218328 479582 218340
rect 480346 218328 480352 218340
rect 479576 218300 480352 218328
rect 479576 218288 479582 218300
rect 480346 218288 480352 218300
rect 480404 218288 480410 218340
rect 534902 218288 534908 218340
rect 534960 218328 534966 218340
rect 567746 218328 567752 218340
rect 534960 218300 567752 218328
rect 534960 218288 534966 218300
rect 567746 218288 567752 218300
rect 567804 218288 567810 218340
rect 568114 218288 568120 218340
rect 568172 218328 568178 218340
rect 568172 218300 596174 218328
rect 568172 218288 568178 218300
rect 55950 218152 55956 218204
rect 56008 218192 56014 218204
rect 56502 218192 56508 218204
rect 56008 218164 56508 218192
rect 56008 218152 56014 218164
rect 56502 218152 56508 218164
rect 56560 218152 56566 218204
rect 64230 218152 64236 218204
rect 64288 218192 64294 218204
rect 65518 218192 65524 218204
rect 64288 218164 65524 218192
rect 64288 218152 64294 218164
rect 65518 218152 65524 218164
rect 65576 218152 65582 218204
rect 67542 218152 67548 218204
rect 67600 218192 67606 218204
rect 71038 218192 71044 218204
rect 67600 218164 71044 218192
rect 67600 218152 67606 218164
rect 71038 218152 71044 218164
rect 71096 218152 71102 218204
rect 75638 218152 75644 218204
rect 75696 218192 75702 218204
rect 76558 218192 76564 218204
rect 75696 218164 76564 218192
rect 75696 218152 75702 218164
rect 76558 218152 76564 218164
rect 76616 218152 76622 218204
rect 130470 218152 130476 218204
rect 130528 218192 130534 218204
rect 167546 218192 167552 218204
rect 130528 218164 167552 218192
rect 130528 218152 130534 218164
rect 167546 218152 167552 218164
rect 167604 218152 167610 218204
rect 168098 218152 168104 218204
rect 168156 218192 168162 218204
rect 170582 218192 170588 218204
rect 168156 218164 170588 218192
rect 168156 218152 168162 218164
rect 170582 218152 170588 218164
rect 170640 218152 170646 218204
rect 172146 218152 172152 218204
rect 172204 218192 172210 218204
rect 177298 218192 177304 218204
rect 172204 218164 177304 218192
rect 172204 218152 172210 218164
rect 177298 218152 177304 218164
rect 177356 218152 177362 218204
rect 190086 218152 190092 218204
rect 190144 218192 190150 218204
rect 225506 218192 225512 218204
rect 190144 218164 225512 218192
rect 190144 218152 190150 218164
rect 225506 218152 225512 218164
rect 225564 218152 225570 218204
rect 246390 218152 246396 218204
rect 246448 218192 246454 218204
rect 249242 218192 249248 218204
rect 246448 218164 249248 218192
rect 246448 218152 246454 218164
rect 249242 218152 249248 218164
rect 249300 218152 249306 218204
rect 249426 218152 249432 218204
rect 249484 218192 249490 218204
rect 251818 218192 251824 218204
rect 249484 218164 251824 218192
rect 249484 218152 249490 218164
rect 251818 218152 251824 218164
rect 251876 218152 251882 218204
rect 289446 218152 289452 218204
rect 289504 218192 289510 218204
rect 294598 218192 294604 218204
rect 289504 218164 294604 218192
rect 289504 218152 289510 218164
rect 294598 218152 294604 218164
rect 294656 218152 294662 218204
rect 332502 218152 332508 218204
rect 332560 218192 332566 218204
rect 335262 218192 335268 218204
rect 332560 218164 335268 218192
rect 332560 218152 332566 218164
rect 335262 218152 335268 218164
rect 335320 218152 335326 218204
rect 339126 218152 339132 218204
rect 339184 218192 339190 218204
rect 340138 218192 340144 218204
rect 339184 218164 340144 218192
rect 339184 218152 339190 218164
rect 340138 218152 340144 218164
rect 340196 218152 340202 218204
rect 348878 218152 348884 218204
rect 348936 218192 348942 218204
rect 353386 218192 353392 218204
rect 348936 218164 353392 218192
rect 348936 218152 348942 218164
rect 353386 218152 353392 218164
rect 353444 218152 353450 218204
rect 358722 218152 358728 218204
rect 358780 218192 358786 218204
rect 363782 218192 363788 218204
rect 358780 218164 363788 218192
rect 358780 218152 358786 218164
rect 363782 218152 363788 218164
rect 363840 218152 363846 218204
rect 375098 218152 375104 218204
rect 375156 218192 375162 218204
rect 380158 218192 380164 218204
rect 375156 218164 380164 218192
rect 375156 218152 375162 218164
rect 380158 218152 380164 218164
rect 380216 218152 380222 218204
rect 381906 218152 381912 218204
rect 381964 218192 381970 218204
rect 382918 218192 382924 218204
rect 381964 218164 382924 218192
rect 381964 218152 381970 218164
rect 382918 218152 382924 218164
rect 382976 218152 382982 218204
rect 394326 218152 394332 218204
rect 394384 218192 394390 218204
rect 402238 218192 402244 218204
rect 394384 218164 402244 218192
rect 394384 218152 394390 218164
rect 402238 218152 402244 218164
rect 402296 218152 402302 218204
rect 424410 218152 424416 218204
rect 424468 218192 424474 218204
rect 426986 218192 426992 218204
rect 424468 218164 426992 218192
rect 424468 218152 424474 218164
rect 426986 218152 426992 218164
rect 427044 218152 427050 218204
rect 433242 218152 433248 218204
rect 433300 218192 433306 218204
rect 435266 218192 435272 218204
rect 433300 218164 435272 218192
rect 433300 218152 433306 218164
rect 435266 218152 435272 218164
rect 435324 218152 435330 218204
rect 436002 218152 436008 218204
rect 436060 218192 436066 218204
rect 436830 218192 436836 218204
rect 436060 218164 436836 218192
rect 436060 218152 436066 218164
rect 436830 218152 436836 218164
rect 436888 218152 436894 218204
rect 461946 218152 461952 218204
rect 462004 218192 462010 218204
rect 465994 218192 466000 218204
rect 462004 218164 466000 218192
rect 462004 218152 462010 218164
rect 465994 218152 466000 218164
rect 466052 218152 466058 218204
rect 505646 218152 505652 218204
rect 505704 218192 505710 218204
rect 558178 218192 558184 218204
rect 505704 218164 558184 218192
rect 505704 218152 505710 218164
rect 558178 218152 558184 218164
rect 558236 218152 558242 218204
rect 558362 218152 558368 218204
rect 558420 218192 558426 218204
rect 567010 218192 567016 218204
rect 558420 218164 567016 218192
rect 558420 218152 558426 218164
rect 567010 218152 567016 218164
rect 567068 218152 567074 218204
rect 567470 218152 567476 218204
rect 567528 218192 567534 218204
rect 594978 218192 594984 218204
rect 567528 218164 594984 218192
rect 567528 218152 567534 218164
rect 594978 218152 594984 218164
rect 595036 218152 595042 218204
rect 596146 218192 596174 218300
rect 613010 218192 613016 218204
rect 596146 218164 613016 218192
rect 613010 218152 613016 218164
rect 613068 218152 613074 218204
rect 56502 218016 56508 218068
rect 56560 218056 56566 218068
rect 57238 218056 57244 218068
rect 56560 218028 57244 218056
rect 56560 218016 56566 218028
rect 57238 218016 57244 218028
rect 57296 218016 57302 218068
rect 58434 218016 58440 218068
rect 58492 218056 58498 218068
rect 59998 218056 60004 218068
rect 58492 218028 60004 218056
rect 58492 218016 58498 218028
rect 59998 218016 60004 218028
rect 60056 218016 60062 218068
rect 62574 218016 62580 218068
rect 62632 218056 62638 218068
rect 63218 218056 63224 218068
rect 62632 218028 63224 218056
rect 62632 218016 62638 218028
rect 63218 218016 63224 218028
rect 63276 218016 63282 218068
rect 65886 218016 65892 218068
rect 65944 218056 65950 218068
rect 66898 218056 66904 218068
rect 65944 218028 66904 218056
rect 65944 218016 65950 218028
rect 66898 218016 66904 218028
rect 66956 218016 66962 218068
rect 68370 218016 68376 218068
rect 68428 218056 68434 218068
rect 68922 218056 68928 218068
rect 68428 218028 68928 218056
rect 68428 218016 68434 218028
rect 68922 218016 68928 218028
rect 68980 218016 68986 218068
rect 72510 218016 72516 218068
rect 72568 218056 72574 218068
rect 73798 218056 73804 218068
rect 72568 218028 73804 218056
rect 72568 218016 72574 218028
rect 73798 218016 73804 218028
rect 73856 218016 73862 218068
rect 74994 218016 75000 218068
rect 75052 218056 75058 218068
rect 75822 218056 75828 218068
rect 75052 218028 75828 218056
rect 75052 218016 75058 218028
rect 75822 218016 75828 218028
rect 75880 218016 75886 218068
rect 79042 218016 79048 218068
rect 79100 218056 79106 218068
rect 79962 218056 79968 218068
rect 79100 218028 79968 218056
rect 79100 218016 79106 218028
rect 79962 218016 79968 218028
rect 80020 218016 80026 218068
rect 80790 218016 80796 218068
rect 80848 218056 80854 218068
rect 81342 218056 81348 218068
rect 80848 218028 81348 218056
rect 80848 218016 80854 218028
rect 81342 218016 81348 218028
rect 81400 218016 81406 218068
rect 83274 218016 83280 218068
rect 83332 218056 83338 218068
rect 84102 218056 84108 218068
rect 83332 218028 84108 218056
rect 83332 218016 83338 218028
rect 84102 218016 84108 218028
rect 84160 218016 84166 218068
rect 93210 218016 93216 218068
rect 93268 218056 93274 218068
rect 93762 218056 93768 218068
rect 93268 218028 93768 218056
rect 93268 218016 93274 218028
rect 93762 218016 93768 218028
rect 93820 218016 93826 218068
rect 97350 218016 97356 218068
rect 97408 218056 97414 218068
rect 97902 218056 97908 218068
rect 97408 218028 97908 218056
rect 97408 218016 97414 218028
rect 97902 218016 97908 218028
rect 97960 218016 97966 218068
rect 99834 218016 99840 218068
rect 99892 218056 99898 218068
rect 100662 218056 100668 218068
rect 99892 218028 100668 218056
rect 99892 218016 99898 218028
rect 100662 218016 100668 218028
rect 100720 218016 100726 218068
rect 103974 218016 103980 218068
rect 104032 218056 104038 218068
rect 104802 218056 104808 218068
rect 104032 218028 104808 218056
rect 104032 218016 104038 218028
rect 104802 218016 104808 218028
rect 104860 218016 104866 218068
rect 112254 218016 112260 218068
rect 112312 218056 112318 218068
rect 112898 218056 112904 218068
rect 112312 218028 112904 218056
rect 112312 218016 112318 218028
rect 112898 218016 112904 218028
rect 112956 218016 112962 218068
rect 116394 218016 116400 218068
rect 116452 218056 116458 218068
rect 117038 218056 117044 218068
rect 116452 218028 117044 218056
rect 116452 218016 116458 218028
rect 117038 218016 117044 218028
rect 117096 218016 117102 218068
rect 128630 218016 128636 218068
rect 128688 218056 128694 218068
rect 129642 218056 129648 218068
rect 128688 218028 129648 218056
rect 128688 218016 128694 218028
rect 129642 218016 129648 218028
rect 129700 218016 129706 218068
rect 132954 218016 132960 218068
rect 133012 218056 133018 218068
rect 133598 218056 133604 218068
rect 133012 218028 133604 218056
rect 133012 218016 133018 218028
rect 133598 218016 133604 218028
rect 133656 218016 133662 218068
rect 142890 218016 142896 218068
rect 142948 218056 142954 218068
rect 143350 218056 143356 218068
rect 142948 218028 143356 218056
rect 142948 218016 142954 218028
rect 143350 218016 143356 218028
rect 143408 218016 143414 218068
rect 145374 218016 145380 218068
rect 145432 218056 145438 218068
rect 146018 218056 146024 218068
rect 145432 218028 146024 218056
rect 145432 218016 145438 218028
rect 146018 218016 146024 218028
rect 146076 218016 146082 218068
rect 149514 218016 149520 218068
rect 149572 218056 149578 218068
rect 150066 218056 150072 218068
rect 149572 218028 150072 218056
rect 149572 218016 149578 218028
rect 150066 218016 150072 218028
rect 150124 218016 150130 218068
rect 155310 218016 155316 218068
rect 155368 218056 155374 218068
rect 155770 218056 155776 218068
rect 155368 218028 155776 218056
rect 155368 218016 155374 218028
rect 155770 218016 155776 218028
rect 155828 218016 155834 218068
rect 159450 218016 159456 218068
rect 159508 218056 159514 218068
rect 160002 218056 160008 218068
rect 159508 218028 160008 218056
rect 159508 218016 159514 218028
rect 160002 218016 160008 218028
rect 160060 218016 160066 218068
rect 160186 218016 160192 218068
rect 160244 218056 160250 218068
rect 163222 218056 163228 218068
rect 160244 218028 163228 218056
rect 160244 218016 160250 218028
rect 163222 218016 163228 218028
rect 163280 218016 163286 218068
rect 166074 218016 166080 218068
rect 166132 218056 166138 218068
rect 166626 218056 166632 218068
rect 166132 218028 166632 218056
rect 166132 218016 166138 218028
rect 166626 218016 166632 218028
rect 166684 218016 166690 218068
rect 167730 218016 167736 218068
rect 167788 218056 167794 218068
rect 168282 218056 168288 218068
rect 167788 218028 168288 218056
rect 167788 218016 167794 218028
rect 168282 218016 168288 218028
rect 168340 218016 168346 218068
rect 171870 218016 171876 218068
rect 171928 218056 171934 218068
rect 172330 218056 172336 218068
rect 171928 218028 172336 218056
rect 171928 218016 171934 218028
rect 172330 218016 172336 218028
rect 172388 218016 172394 218068
rect 176010 218016 176016 218068
rect 176068 218056 176074 218068
rect 176470 218056 176476 218068
rect 176068 218028 176476 218056
rect 176068 218016 176074 218028
rect 176470 218016 176476 218028
rect 176528 218016 176534 218068
rect 182634 218016 182640 218068
rect 182692 218056 182698 218068
rect 183462 218056 183468 218068
rect 182692 218028 183468 218056
rect 182692 218016 182698 218028
rect 183462 218016 183468 218028
rect 183520 218016 183526 218068
rect 184842 218016 184848 218068
rect 184900 218056 184906 218068
rect 185578 218056 185584 218068
rect 184900 218028 185584 218056
rect 184900 218016 184906 218028
rect 185578 218016 185584 218028
rect 185636 218016 185642 218068
rect 188430 218016 188436 218068
rect 188488 218056 188494 218068
rect 189442 218056 189448 218068
rect 188488 218028 189448 218056
rect 188488 218016 188494 218028
rect 189442 218016 189448 218028
rect 189500 218016 189506 218068
rect 190914 218016 190920 218068
rect 190972 218056 190978 218068
rect 191650 218056 191656 218068
rect 190972 218028 191656 218056
rect 190972 218016 190978 218028
rect 191650 218016 191656 218028
rect 191708 218016 191714 218068
rect 192570 218016 192576 218068
rect 192628 218056 192634 218068
rect 193122 218056 193128 218068
rect 192628 218028 193128 218056
rect 192628 218016 192634 218028
rect 193122 218016 193128 218028
rect 193180 218016 193186 218068
rect 196710 218016 196716 218068
rect 196768 218056 196774 218068
rect 203886 218056 203892 218068
rect 196768 218028 203892 218056
rect 196768 218016 196774 218028
rect 203886 218016 203892 218028
rect 203944 218016 203950 218068
rect 204990 218016 204996 218068
rect 205048 218056 205054 218068
rect 205450 218056 205456 218068
rect 205048 218028 205456 218056
rect 205048 218016 205054 218028
rect 205450 218016 205456 218028
rect 205508 218016 205514 218068
rect 211614 218016 211620 218068
rect 211672 218056 211678 218068
rect 215202 218056 215208 218068
rect 211672 218028 215208 218056
rect 211672 218016 211678 218028
rect 215202 218016 215208 218028
rect 215260 218016 215266 218068
rect 215754 218016 215760 218068
rect 215812 218056 215818 218068
rect 216582 218056 216588 218068
rect 215812 218028 216588 218056
rect 215812 218016 215818 218028
rect 216582 218016 216588 218028
rect 216640 218016 216646 218068
rect 221550 218016 221556 218068
rect 221608 218056 221614 218068
rect 222562 218056 222568 218068
rect 221608 218028 222568 218056
rect 221608 218016 221614 218028
rect 222562 218016 222568 218028
rect 222620 218016 222626 218068
rect 224034 218016 224040 218068
rect 224092 218056 224098 218068
rect 224586 218056 224592 218068
rect 224092 218028 224592 218056
rect 224092 218016 224098 218028
rect 224586 218016 224592 218028
rect 224644 218016 224650 218068
rect 225690 218016 225696 218068
rect 225748 218056 225754 218068
rect 226150 218056 226156 218068
rect 225748 218028 226156 218056
rect 225748 218016 225754 218028
rect 226150 218016 226156 218028
rect 226208 218016 226214 218068
rect 229830 218016 229836 218068
rect 229888 218056 229894 218068
rect 230382 218056 230388 218068
rect 229888 218028 230388 218056
rect 229888 218016 229894 218028
rect 230382 218016 230388 218028
rect 230440 218016 230446 218068
rect 232314 218016 232320 218068
rect 232372 218056 232378 218068
rect 233142 218056 233148 218068
rect 232372 218028 233148 218056
rect 232372 218016 232378 218028
rect 233142 218016 233148 218028
rect 233200 218016 233206 218068
rect 233970 218016 233976 218068
rect 234028 218056 234034 218068
rect 234522 218056 234528 218068
rect 234028 218028 234528 218056
rect 234028 218016 234034 218028
rect 234522 218016 234528 218028
rect 234580 218016 234586 218068
rect 242250 218016 242256 218068
rect 242308 218056 242314 218068
rect 242710 218056 242716 218068
rect 242308 218028 242716 218056
rect 242308 218016 242314 218028
rect 242710 218016 242716 218028
rect 242768 218016 242774 218068
rect 248874 218016 248880 218068
rect 248932 218056 248938 218068
rect 249610 218056 249616 218068
rect 248932 218028 249616 218056
rect 248932 218016 248938 218028
rect 249610 218016 249616 218028
rect 249668 218016 249674 218068
rect 254670 218016 254676 218068
rect 254728 218056 254734 218068
rect 255130 218056 255136 218068
rect 254728 218028 255136 218056
rect 254728 218016 254734 218028
rect 255130 218016 255136 218028
rect 255188 218016 255194 218068
rect 258810 218016 258816 218068
rect 258868 218056 258874 218068
rect 259362 218056 259368 218068
rect 258868 218028 259368 218056
rect 258868 218016 258874 218028
rect 259362 218016 259368 218028
rect 259420 218016 259426 218068
rect 265434 218016 265440 218068
rect 265492 218056 265498 218068
rect 266262 218056 266268 218068
rect 265492 218028 266268 218056
rect 265492 218016 265498 218028
rect 266262 218016 266268 218028
rect 266320 218016 266326 218068
rect 269574 218016 269580 218068
rect 269632 218056 269638 218068
rect 270126 218056 270132 218068
rect 269632 218028 270132 218056
rect 269632 218016 269638 218028
rect 270126 218016 270132 218028
rect 270184 218016 270190 218068
rect 273714 218016 273720 218068
rect 273772 218056 273778 218068
rect 274266 218056 274272 218068
rect 273772 218028 274272 218056
rect 273772 218016 273778 218028
rect 274266 218016 274272 218028
rect 274324 218016 274330 218068
rect 281994 218016 282000 218068
rect 282052 218056 282058 218068
rect 282546 218056 282552 218068
rect 282052 218028 282552 218056
rect 282052 218016 282058 218028
rect 282546 218016 282552 218028
rect 282604 218016 282610 218068
rect 284202 218016 284208 218068
rect 284260 218056 284266 218068
rect 284938 218056 284944 218068
rect 284260 218028 284944 218056
rect 284260 218016 284266 218028
rect 284938 218016 284944 218028
rect 284996 218016 285002 218068
rect 287790 218016 287796 218068
rect 287848 218056 287854 218068
rect 288342 218056 288348 218068
rect 287848 218028 288348 218056
rect 287848 218016 287854 218028
rect 288342 218016 288348 218028
rect 288400 218016 288406 218068
rect 290274 218016 290280 218068
rect 290332 218056 290338 218068
rect 290918 218056 290924 218068
rect 290332 218028 290924 218056
rect 290332 218016 290338 218028
rect 290918 218016 290924 218028
rect 290976 218016 290982 218068
rect 296070 218016 296076 218068
rect 296128 218056 296134 218068
rect 296622 218056 296628 218068
rect 296128 218028 296628 218056
rect 296128 218016 296134 218028
rect 296622 218016 296628 218028
rect 296680 218016 296686 218068
rect 297726 218016 297732 218068
rect 297784 218056 297790 218068
rect 300026 218056 300032 218068
rect 297784 218028 300032 218056
rect 297784 218016 297790 218028
rect 300026 218016 300032 218028
rect 300084 218016 300090 218068
rect 300210 218016 300216 218068
rect 300268 218056 300274 218068
rect 300762 218056 300768 218068
rect 300268 218028 300768 218056
rect 300268 218016 300274 218028
rect 300762 218016 300768 218028
rect 300820 218016 300826 218068
rect 304350 218016 304356 218068
rect 304408 218056 304414 218068
rect 305638 218056 305644 218068
rect 304408 218028 305644 218056
rect 304408 218016 304414 218028
rect 305638 218016 305644 218028
rect 305696 218016 305702 218068
rect 308490 218016 308496 218068
rect 308548 218056 308554 218068
rect 309042 218056 309048 218068
rect 308548 218028 309048 218056
rect 308548 218016 308554 218028
rect 309042 218016 309048 218028
rect 309100 218016 309106 218068
rect 310974 218016 310980 218068
rect 311032 218056 311038 218068
rect 311802 218056 311808 218068
rect 311032 218028 311808 218056
rect 311032 218016 311038 218028
rect 311802 218016 311808 218028
rect 311860 218016 311866 218068
rect 312630 218016 312636 218068
rect 312688 218056 312694 218068
rect 313090 218056 313096 218068
rect 312688 218028 313096 218056
rect 312688 218016 312694 218028
rect 313090 218016 313096 218028
rect 313148 218016 313154 218068
rect 315114 218016 315120 218068
rect 315172 218056 315178 218068
rect 315666 218056 315672 218068
rect 315172 218028 315672 218056
rect 315172 218016 315178 218028
rect 315666 218016 315672 218028
rect 315724 218016 315730 218068
rect 317322 218016 317328 218068
rect 317380 218056 317386 218068
rect 318058 218056 318064 218068
rect 317380 218028 318064 218056
rect 317380 218016 317386 218028
rect 318058 218016 318064 218028
rect 318116 218016 318122 218068
rect 319254 218016 319260 218068
rect 319312 218056 319318 218068
rect 319990 218056 319996 218068
rect 319312 218028 319996 218056
rect 319312 218016 319318 218028
rect 319990 218016 319996 218028
rect 320048 218016 320054 218068
rect 333330 218016 333336 218068
rect 333388 218056 333394 218068
rect 333882 218056 333888 218068
rect 333388 218028 333888 218056
rect 333388 218016 333394 218028
rect 333882 218016 333888 218028
rect 333940 218016 333946 218068
rect 335814 218016 335820 218068
rect 335872 218056 335878 218068
rect 336458 218056 336464 218068
rect 335872 218028 336464 218056
rect 335872 218016 335878 218028
rect 336458 218016 336464 218028
rect 336516 218016 336522 218068
rect 339954 218016 339960 218068
rect 340012 218056 340018 218068
rect 340690 218056 340696 218068
rect 340012 218028 340696 218056
rect 340012 218016 340018 218028
rect 340690 218016 340696 218028
rect 340748 218016 340754 218068
rect 341610 218016 341616 218068
rect 341668 218056 341674 218068
rect 342070 218056 342076 218068
rect 341668 218028 342076 218056
rect 341668 218016 341674 218028
rect 342070 218016 342076 218028
rect 342128 218016 342134 218068
rect 345750 218016 345756 218068
rect 345808 218056 345814 218068
rect 346210 218056 346216 218068
rect 345808 218028 346216 218056
rect 345808 218016 345814 218028
rect 346210 218016 346216 218028
rect 346268 218016 346274 218068
rect 348234 218016 348240 218068
rect 348292 218056 348298 218068
rect 349062 218056 349068 218068
rect 348292 218028 349068 218056
rect 348292 218016 348298 218028
rect 349062 218016 349068 218028
rect 349120 218016 349126 218068
rect 352374 218016 352380 218068
rect 352432 218056 352438 218068
rect 354306 218056 354312 218068
rect 352432 218028 354312 218056
rect 352432 218016 352438 218028
rect 354306 218016 354312 218028
rect 354364 218016 354370 218068
rect 356514 218016 356520 218068
rect 356572 218056 356578 218068
rect 357250 218056 357256 218068
rect 356572 218028 357256 218056
rect 356572 218016 356578 218028
rect 357250 218016 357256 218028
rect 357308 218016 357314 218068
rect 360654 218016 360660 218068
rect 360712 218056 360718 218068
rect 361298 218056 361304 218068
rect 360712 218028 361304 218056
rect 360712 218016 360718 218028
rect 361298 218016 361304 218028
rect 361356 218016 361362 218068
rect 364794 218016 364800 218068
rect 364852 218056 364858 218068
rect 365530 218056 365536 218068
rect 364852 218028 365536 218056
rect 364852 218016 364858 218028
rect 365530 218016 365536 218028
rect 365588 218016 365594 218068
rect 366450 218016 366456 218068
rect 366508 218056 366514 218068
rect 366910 218056 366916 218068
rect 366508 218028 366916 218056
rect 366508 218016 366514 218028
rect 366910 218016 366916 218028
rect 366968 218016 366974 218068
rect 368934 218016 368940 218068
rect 368992 218056 368998 218068
rect 372522 218056 372528 218068
rect 368992 218028 372528 218056
rect 368992 218016 368998 218028
rect 372522 218016 372528 218028
rect 372580 218016 372586 218068
rect 372982 218016 372988 218068
rect 373040 218056 373046 218068
rect 373810 218056 373816 218068
rect 373040 218028 373816 218056
rect 373040 218016 373046 218028
rect 373810 218016 373816 218028
rect 373868 218016 373874 218068
rect 374730 218016 374736 218068
rect 374788 218056 374794 218068
rect 375282 218056 375288 218068
rect 374788 218028 375288 218056
rect 374788 218016 374794 218028
rect 375282 218016 375288 218028
rect 375340 218016 375346 218068
rect 381354 218016 381360 218068
rect 381412 218056 381418 218068
rect 382090 218056 382096 218068
rect 381412 218028 382096 218056
rect 381412 218016 381418 218028
rect 382090 218016 382096 218028
rect 382148 218016 382154 218068
rect 385494 218016 385500 218068
rect 385552 218056 385558 218068
rect 386322 218056 386328 218068
rect 385552 218028 386328 218056
rect 385552 218016 385558 218028
rect 386322 218016 386328 218028
rect 386380 218016 386386 218068
rect 389634 218016 389640 218068
rect 389692 218056 389698 218068
rect 390186 218056 390192 218068
rect 389692 218028 390192 218056
rect 389692 218016 389698 218028
rect 390186 218016 390192 218028
rect 390244 218016 390250 218068
rect 393774 218016 393780 218068
rect 393832 218056 393838 218068
rect 394510 218056 394516 218068
rect 393832 218028 394516 218056
rect 393832 218016 393838 218028
rect 394510 218016 394516 218028
rect 394568 218016 394574 218068
rect 397914 218016 397920 218068
rect 397972 218056 397978 218068
rect 398558 218056 398564 218068
rect 397972 218028 398564 218056
rect 397972 218016 397978 218028
rect 398558 218016 398564 218028
rect 398616 218016 398622 218068
rect 399570 218016 399576 218068
rect 399628 218056 399634 218068
rect 400030 218056 400036 218068
rect 399628 218028 400036 218056
rect 399628 218016 399634 218028
rect 400030 218016 400036 218028
rect 400088 218016 400094 218068
rect 403710 218016 403716 218068
rect 403768 218056 403774 218068
rect 404170 218056 404176 218068
rect 403768 218028 404176 218056
rect 403768 218016 403774 218028
rect 404170 218016 404176 218028
rect 404228 218016 404234 218068
rect 410334 218016 410340 218068
rect 410392 218056 410398 218068
rect 410886 218056 410892 218068
rect 410392 218028 410892 218056
rect 410392 218016 410398 218028
rect 410886 218016 410892 218028
rect 410944 218016 410950 218068
rect 416130 218016 416136 218068
rect 416188 218056 416194 218068
rect 416682 218056 416688 218068
rect 416188 218028 416688 218056
rect 416188 218016 416194 218028
rect 416682 218016 416688 218028
rect 416740 218016 416746 218068
rect 418614 218016 418620 218068
rect 418672 218056 418678 218068
rect 419442 218056 419448 218068
rect 418672 218028 419448 218056
rect 418672 218016 418678 218028
rect 419442 218016 419448 218028
rect 419500 218016 419506 218068
rect 420270 218016 420276 218068
rect 420328 218056 420334 218068
rect 420822 218056 420828 218068
rect 420328 218028 420828 218056
rect 420328 218016 420334 218028
rect 420822 218016 420828 218028
rect 420880 218016 420886 218068
rect 422754 218016 422760 218068
rect 422812 218056 422818 218068
rect 425422 218056 425428 218068
rect 422812 218028 425428 218056
rect 422812 218016 422818 218028
rect 425422 218016 425428 218028
rect 425480 218016 425486 218068
rect 426066 218016 426072 218068
rect 426124 218056 426130 218068
rect 428458 218056 428464 218068
rect 426124 218028 428464 218056
rect 426124 218016 426130 218028
rect 428458 218016 428464 218028
rect 428516 218016 428522 218068
rect 429102 218016 429108 218068
rect 429160 218056 429166 218068
rect 430666 218056 430672 218068
rect 429160 218028 430672 218056
rect 429160 218016 429166 218028
rect 430666 218016 430672 218028
rect 430724 218016 430730 218068
rect 432690 218016 432696 218068
rect 432748 218056 432754 218068
rect 433794 218056 433800 218068
rect 432748 218028 433800 218056
rect 432748 218016 432754 218028
rect 433794 218016 433800 218028
rect 433852 218016 433858 218068
rect 434990 218016 434996 218068
rect 435048 218056 435054 218068
rect 436278 218056 436284 218068
rect 435048 218028 436284 218056
rect 435048 218016 435054 218028
rect 436278 218016 436284 218028
rect 436336 218016 436342 218068
rect 436462 218016 436468 218068
rect 436520 218056 436526 218068
rect 437474 218056 437480 218068
rect 436520 218028 437480 218056
rect 436520 218016 436526 218028
rect 437474 218016 437480 218028
rect 437532 218016 437538 218068
rect 438486 218016 438492 218068
rect 438544 218056 438550 218068
rect 438946 218056 438952 218068
rect 438544 218028 438952 218056
rect 438544 218016 438550 218028
rect 438946 218016 438952 218028
rect 439004 218016 439010 218068
rect 440142 218016 440148 218068
rect 440200 218056 440206 218068
rect 440694 218056 440700 218068
rect 440200 218028 440700 218056
rect 440200 218016 440206 218028
rect 440694 218016 440700 218028
rect 440752 218016 440758 218068
rect 453298 218016 453304 218068
rect 453356 218056 453362 218068
rect 455414 218056 455420 218068
rect 453356 218028 455420 218056
rect 453356 218016 453362 218028
rect 455414 218016 455420 218028
rect 455472 218016 455478 218068
rect 462958 218016 462964 218068
rect 463016 218056 463022 218068
rect 464338 218056 464344 218068
rect 463016 218028 464344 218056
rect 463016 218016 463022 218028
rect 464338 218016 464344 218028
rect 464396 218016 464402 218068
rect 467098 218016 467104 218068
rect 467156 218056 467162 218068
rect 467834 218056 467840 218068
rect 467156 218028 467840 218056
rect 467156 218016 467162 218028
rect 467834 218016 467840 218028
rect 467892 218016 467898 218068
rect 471238 218016 471244 218068
rect 471296 218056 471302 218068
rect 472618 218056 472624 218068
rect 471296 218028 472624 218056
rect 471296 218016 471302 218028
rect 472618 218016 472624 218028
rect 472676 218016 472682 218068
rect 480990 218016 480996 218068
rect 481048 218056 481054 218068
rect 482554 218056 482560 218068
rect 481048 218028 482560 218056
rect 481048 218016 481054 218028
rect 482554 218016 482560 218028
rect 482612 218016 482618 218068
rect 482738 218016 482744 218068
rect 482796 218056 482802 218068
rect 485038 218056 485044 218068
rect 482796 218028 485044 218056
rect 482796 218016 482802 218028
rect 485038 218016 485044 218028
rect 485096 218016 485102 218068
rect 495342 218016 495348 218068
rect 495400 218056 495406 218068
rect 500218 218056 500224 218068
rect 495400 218028 500224 218056
rect 495400 218016 495406 218028
rect 500218 218016 500224 218028
rect 500276 218016 500282 218068
rect 502426 218016 502432 218068
rect 502484 218056 502490 218068
rect 502484 218028 608640 218056
rect 502484 218016 502490 218028
rect 608612 217988 608640 218028
rect 648246 218016 648252 218068
rect 648304 218056 648310 218068
rect 654778 218056 654784 218068
rect 648304 218028 654784 218056
rect 648304 218016 648310 218028
rect 654778 218016 654784 218028
rect 654836 218016 654842 218068
rect 614482 217988 614488 218000
rect 608612 217960 614488 217988
rect 614482 217948 614488 217960
rect 614540 217948 614546 218000
rect 565170 217880 565176 217932
rect 565228 217920 565234 217932
rect 568298 217920 568304 217932
rect 565228 217892 568304 217920
rect 565228 217880 565234 217892
rect 568298 217880 568304 217892
rect 568356 217880 568362 217932
rect 572162 217880 572168 217932
rect 572220 217920 572226 217932
rect 576026 217920 576032 217932
rect 572220 217892 576032 217920
rect 572220 217880 572226 217892
rect 576026 217880 576032 217892
rect 576084 217880 576090 217932
rect 576210 217880 576216 217932
rect 576268 217920 576274 217932
rect 576268 217892 576854 217920
rect 576268 217880 576274 217892
rect 447134 217812 447140 217864
rect 447192 217852 447198 217864
rect 447778 217852 447784 217864
rect 447192 217824 447784 217852
rect 447192 217812 447198 217824
rect 447778 217812 447784 217824
rect 447836 217812 447842 217864
rect 525794 217812 525800 217864
rect 525852 217852 525858 217864
rect 526438 217852 526444 217864
rect 525852 217824 526444 217852
rect 525852 217812 525858 217824
rect 526438 217812 526444 217824
rect 526496 217812 526502 217864
rect 555694 217812 555700 217864
rect 555752 217852 555758 217864
rect 562870 217852 562876 217864
rect 555752 217824 562876 217852
rect 555752 217812 555758 217824
rect 562870 217812 562876 217824
rect 562928 217812 562934 217864
rect 572346 217744 572352 217796
rect 572404 217784 572410 217796
rect 576578 217784 576584 217796
rect 572404 217756 576584 217784
rect 572404 217744 572410 217756
rect 576578 217744 576584 217756
rect 576636 217744 576642 217796
rect 576826 217784 576854 217892
rect 578234 217784 578240 217796
rect 576826 217756 578240 217784
rect 578234 217744 578240 217756
rect 578292 217744 578298 217796
rect 561122 217676 561128 217728
rect 561180 217716 561186 217728
rect 563238 217716 563244 217728
rect 561180 217688 563244 217716
rect 561180 217676 561186 217688
rect 563238 217676 563244 217688
rect 563296 217676 563302 217728
rect 605098 217676 605104 217728
rect 605156 217716 605162 217728
rect 614114 217716 614120 217728
rect 605156 217688 614120 217716
rect 605156 217676 605162 217688
rect 614114 217676 614120 217688
rect 614172 217676 614178 217728
rect 577314 217648 577320 217660
rect 572686 217620 577320 217648
rect 553210 217540 553216 217592
rect 553268 217580 553274 217592
rect 554222 217580 554228 217592
rect 553268 217552 554228 217580
rect 553268 217540 553274 217552
rect 554222 217540 554228 217552
rect 554280 217540 554286 217592
rect 563054 217540 563060 217592
rect 563112 217580 563118 217592
rect 572686 217580 572714 217620
rect 577314 217608 577320 217620
rect 577372 217608 577378 217660
rect 563112 217552 572714 217580
rect 563112 217540 563118 217552
rect 597554 217540 597560 217592
rect 597612 217580 597618 217592
rect 613378 217580 613384 217592
rect 597612 217552 613384 217580
rect 597612 217540 597618 217552
rect 613378 217540 613384 217552
rect 613436 217540 613442 217592
rect 576578 217472 576584 217524
rect 576636 217512 576642 217524
rect 576946 217512 576952 217524
rect 576636 217484 576952 217512
rect 576636 217472 576642 217484
rect 576946 217472 576952 217484
rect 577004 217472 577010 217524
rect 591574 217472 591580 217524
rect 591632 217512 591638 217524
rect 595714 217512 595720 217524
rect 591632 217484 595720 217512
rect 591632 217472 591638 217484
rect 595714 217472 595720 217484
rect 595772 217472 595778 217524
rect 611814 217404 611820 217456
rect 611872 217444 611878 217456
rect 628282 217444 628288 217456
rect 611872 217416 628288 217444
rect 611872 217404 611878 217416
rect 628282 217404 628288 217416
rect 628340 217404 628346 217456
rect 571702 217336 571708 217388
rect 571760 217376 571766 217388
rect 577130 217376 577136 217388
rect 571760 217348 577136 217376
rect 571760 217336 571766 217348
rect 577130 217336 577136 217348
rect 577188 217336 577194 217388
rect 594978 217268 594984 217320
rect 595036 217308 595042 217320
rect 626074 217308 626080 217320
rect 595036 217280 626080 217308
rect 595036 217268 595042 217280
rect 626074 217268 626080 217280
rect 626132 217268 626138 217320
rect 563054 217200 563060 217252
rect 563112 217240 563118 217252
rect 563112 217212 572714 217240
rect 563112 217200 563118 217212
rect 562686 217064 562692 217116
rect 562744 217104 562750 217116
rect 572530 217104 572536 217116
rect 562744 217076 572536 217104
rect 562744 217064 562750 217076
rect 572530 217064 572536 217076
rect 572588 217064 572594 217116
rect 572686 217104 572714 217212
rect 582374 217200 582380 217252
rect 582432 217240 582438 217252
rect 591942 217240 591948 217252
rect 582432 217212 591948 217240
rect 582432 217200 582438 217212
rect 591942 217200 591948 217212
rect 592000 217200 592006 217252
rect 572686 217076 576854 217104
rect 576826 216832 576854 217076
rect 591758 217064 591764 217116
rect 591816 217104 591822 217116
rect 595162 217104 595168 217116
rect 591816 217076 595168 217104
rect 591816 217064 591822 217076
rect 595162 217064 595168 217076
rect 595220 217064 595226 217116
rect 576826 216804 582374 216832
rect 582346 216764 582374 216804
rect 582558 216764 582564 216776
rect 582346 216736 582564 216764
rect 582558 216724 582564 216736
rect 582616 216724 582622 216776
rect 663242 216112 663248 216164
rect 663300 216152 663306 216164
rect 664438 216152 664444 216164
rect 663300 216124 664444 216152
rect 663300 216112 663306 216124
rect 664438 216112 664444 216124
rect 664496 216112 664502 216164
rect 622946 216044 622952 216096
rect 623004 216084 623010 216096
rect 629938 216084 629944 216096
rect 623004 216056 629944 216084
rect 623004 216044 623010 216056
rect 629938 216044 629944 216056
rect 629996 216044 630002 216096
rect 577682 215908 577688 215960
rect 577740 215948 577746 215960
rect 628834 215948 628840 215960
rect 577740 215920 628840 215948
rect 577740 215908 577746 215920
rect 628834 215908 628840 215920
rect 628892 215908 628898 215960
rect 655422 215296 655428 215348
rect 655480 215336 655486 215348
rect 656158 215336 656164 215348
rect 655480 215308 656164 215336
rect 655480 215296 655486 215308
rect 656158 215296 656164 215308
rect 656216 215296 656222 215348
rect 577314 215092 577320 215144
rect 577372 215132 577378 215144
rect 612274 215132 612280 215144
rect 577372 215104 612280 215132
rect 577372 215092 577378 215104
rect 612274 215092 612280 215104
rect 612332 215092 612338 215144
rect 675846 215092 675852 215144
rect 675904 215132 675910 215144
rect 676858 215132 676864 215144
rect 675904 215104 676864 215132
rect 675904 215092 675910 215104
rect 676858 215092 676864 215104
rect 676916 215092 676922 215144
rect 577866 214956 577872 215008
rect 577924 214996 577930 215008
rect 621842 214996 621848 215008
rect 577924 214968 621848 214996
rect 577924 214956 577930 214968
rect 621842 214956 621848 214968
rect 621900 214956 621906 215008
rect 578050 214820 578056 214872
rect 578108 214860 578114 214872
rect 621106 214860 621112 214872
rect 578108 214832 621112 214860
rect 578108 214820 578114 214832
rect 621106 214820 621112 214832
rect 621164 214820 621170 214872
rect 621658 214820 621664 214872
rect 621716 214860 621722 214872
rect 632882 214860 632888 214872
rect 621716 214832 632888 214860
rect 621716 214820 621722 214832
rect 632882 214820 632888 214832
rect 632940 214820 632946 214872
rect 578234 214684 578240 214736
rect 578292 214724 578298 214736
rect 624418 214724 624424 214736
rect 578292 214696 624424 214724
rect 578292 214684 578298 214696
rect 624418 214684 624424 214696
rect 624476 214684 624482 214736
rect 648430 214684 648436 214736
rect 648488 214724 648494 214736
rect 658918 214724 658924 214736
rect 648488 214696 658924 214724
rect 648488 214684 648494 214696
rect 658918 214684 658924 214696
rect 658976 214684 658982 214736
rect 577498 214548 577504 214600
rect 577556 214588 577562 214600
rect 577556 214560 616736 214588
rect 577556 214548 577562 214560
rect 599026 214412 599032 214464
rect 599084 214452 599090 214464
rect 599578 214452 599584 214464
rect 599084 214424 599584 214452
rect 599084 214412 599090 214424
rect 599578 214412 599584 214424
rect 599636 214412 599642 214464
rect 600406 214412 600412 214464
rect 600464 214452 600470 214464
rect 601234 214452 601240 214464
rect 600464 214424 601240 214452
rect 600464 214412 600470 214424
rect 601234 214412 601240 214424
rect 601292 214412 601298 214464
rect 615494 214412 615500 214464
rect 615552 214452 615558 214464
rect 616138 214452 616144 214464
rect 615552 214424 616144 214452
rect 615552 214412 615558 214424
rect 616138 214412 616144 214424
rect 616196 214412 616202 214464
rect 616708 214452 616736 214560
rect 616874 214548 616880 214600
rect 616932 214588 616938 214600
rect 617334 214588 617340 214600
rect 616932 214560 617340 214588
rect 616932 214548 616938 214560
rect 617334 214548 617340 214560
rect 617392 214548 617398 214600
rect 619634 214548 619640 214600
rect 619692 214588 619698 214600
rect 620554 214588 620560 214600
rect 619692 214560 620560 214588
rect 619692 214548 619698 214560
rect 620554 214548 620560 214560
rect 620612 214548 620618 214600
rect 622578 214548 622584 214600
rect 622636 214588 622642 214600
rect 623314 214588 623320 214600
rect 622636 214560 623320 214588
rect 622636 214548 622642 214560
rect 623314 214548 623320 214560
rect 623372 214548 623378 214600
rect 623774 214548 623780 214600
rect 623832 214588 623838 214600
rect 623832 214560 625154 214588
rect 623832 214548 623838 214560
rect 623866 214452 623872 214464
rect 616708 214424 623872 214452
rect 623866 214412 623872 214424
rect 623924 214412 623930 214464
rect 625126 214452 625154 214560
rect 625246 214548 625252 214600
rect 625304 214588 625310 214600
rect 625614 214588 625620 214600
rect 625304 214560 625620 214588
rect 625304 214548 625310 214560
rect 625614 214548 625620 214560
rect 625672 214548 625678 214600
rect 636286 214548 636292 214600
rect 636344 214588 636350 214600
rect 639598 214588 639604 214600
rect 636344 214560 639604 214588
rect 636344 214548 636350 214560
rect 639598 214548 639604 214560
rect 639656 214548 639662 214600
rect 652754 214548 652760 214600
rect 652812 214588 652818 214600
rect 665818 214588 665824 214600
rect 652812 214560 665824 214588
rect 652812 214548 652818 214560
rect 665818 214548 665824 214560
rect 665876 214548 665882 214600
rect 631594 214452 631600 214464
rect 625126 214424 631600 214452
rect 631594 214412 631600 214424
rect 631652 214412 631658 214464
rect 675846 214412 675852 214464
rect 675904 214452 675910 214464
rect 677410 214452 677416 214464
rect 675904 214424 677416 214452
rect 675904 214412 675910 214424
rect 677410 214412 677416 214424
rect 677468 214412 677474 214464
rect 600498 214276 600504 214328
rect 600556 214316 600562 214328
rect 600866 214316 600872 214328
rect 600556 214288 600872 214316
rect 600556 214276 600562 214288
rect 600866 214276 600872 214288
rect 600924 214276 600930 214328
rect 41322 213936 41328 213988
rect 41380 213976 41386 213988
rect 41690 213976 41696 213988
rect 41380 213948 41696 213976
rect 41380 213936 41386 213948
rect 41690 213936 41696 213948
rect 41748 213936 41754 213988
rect 638310 213868 638316 213920
rect 638368 213908 638374 213920
rect 640610 213908 640616 213920
rect 638368 213880 640616 213908
rect 638368 213868 638374 213880
rect 640610 213868 640616 213880
rect 640668 213868 640674 213920
rect 648614 213868 648620 213920
rect 648672 213908 648678 213920
rect 649258 213908 649264 213920
rect 648672 213880 649264 213908
rect 648672 213868 648678 213880
rect 649258 213868 649264 213880
rect 649316 213868 649322 213920
rect 650454 213868 650460 213920
rect 650512 213908 650518 213920
rect 653122 213908 653128 213920
rect 650512 213880 653128 213908
rect 650512 213868 650518 213880
rect 653122 213868 653128 213880
rect 653180 213868 653186 213920
rect 660390 213868 660396 213920
rect 660448 213908 660454 213920
rect 660942 213908 660948 213920
rect 660448 213880 660948 213908
rect 660448 213868 660454 213880
rect 660942 213868 660948 213880
rect 661000 213868 661006 213920
rect 641622 213732 641628 213784
rect 641680 213772 641686 213784
rect 650638 213772 650644 213784
rect 641680 213744 650644 213772
rect 641680 213732 641686 213744
rect 650638 213732 650644 213744
rect 650696 213732 650702 213784
rect 660942 213732 660948 213784
rect 661000 213772 661006 213784
rect 662966 213772 662972 213784
rect 661000 213744 662972 213772
rect 661000 213732 661006 213744
rect 662966 213732 662972 213744
rect 663024 213732 663030 213784
rect 640242 213596 640248 213648
rect 640300 213636 640306 213648
rect 649718 213636 649724 213648
rect 640300 213608 649724 213636
rect 640300 213596 640306 213608
rect 649718 213596 649724 213608
rect 649776 213596 649782 213648
rect 651834 213596 651840 213648
rect 651892 213636 651898 213648
rect 657538 213636 657544 213648
rect 651892 213608 657544 213636
rect 651892 213596 651898 213608
rect 657538 213596 657544 213608
rect 657596 213596 657602 213648
rect 676030 213528 676036 213580
rect 676088 213568 676094 213580
rect 677042 213568 677048 213580
rect 676088 213540 677048 213568
rect 676088 213528 676094 213540
rect 677042 213528 677048 213540
rect 677100 213528 677106 213580
rect 635550 213460 635556 213512
rect 635608 213500 635614 213512
rect 652386 213500 652392 213512
rect 635608 213472 652392 213500
rect 635608 213460 635614 213472
rect 652386 213460 652392 213472
rect 652444 213460 652450 213512
rect 638862 213324 638868 213376
rect 638920 213364 638926 213376
rect 660206 213364 660212 213376
rect 638920 213336 660212 213364
rect 638920 213324 638926 213336
rect 660206 213324 660212 213336
rect 660264 213324 660270 213376
rect 642174 213188 642180 213240
rect 642232 213228 642238 213240
rect 642232 213200 644474 213228
rect 642232 213188 642238 213200
rect 644446 213024 644474 213200
rect 661494 213120 661500 213172
rect 661552 213160 661558 213172
rect 666278 213160 666284 213172
rect 661552 213132 666284 213160
rect 661552 213120 661558 213132
rect 666278 213120 666284 213132
rect 666336 213120 666342 213172
rect 644446 212996 663794 213024
rect 613010 212848 613016 212900
rect 613068 212888 613074 212900
rect 615034 212888 615040 212900
rect 613068 212860 615040 212888
rect 613068 212848 613074 212860
rect 615034 212848 615040 212860
rect 615092 212848 615098 212900
rect 663766 212888 663794 212996
rect 664254 212984 664260 213036
rect 664312 213024 664318 213036
rect 665082 213024 665088 213036
rect 664312 212996 665088 213024
rect 664312 212984 664318 212996
rect 665082 212984 665088 212996
rect 665140 212984 665146 213036
rect 665450 212888 665456 212900
rect 663766 212860 665456 212888
rect 665450 212848 665456 212860
rect 665508 212848 665514 212900
rect 632698 212712 632704 212764
rect 632756 212752 632762 212764
rect 634354 212752 634360 212764
rect 632756 212724 634360 212752
rect 632756 212712 632762 212724
rect 634354 212712 634360 212724
rect 634412 212712 634418 212764
rect 658734 212712 658740 212764
rect 658792 212752 658798 212764
rect 659562 212752 659568 212764
rect 658792 212724 659568 212752
rect 658792 212712 658798 212724
rect 659562 212712 659568 212724
rect 659620 212712 659626 212764
rect 601786 212372 601792 212424
rect 601844 212412 601850 212424
rect 602338 212412 602344 212424
rect 601844 212384 602344 212412
rect 601844 212372 601850 212384
rect 602338 212372 602344 212384
rect 602396 212372 602402 212424
rect 603074 212372 603080 212424
rect 603132 212412 603138 212424
rect 603994 212412 604000 212424
rect 603132 212384 604000 212412
rect 603132 212372 603138 212384
rect 603994 212372 604000 212384
rect 604052 212372 604058 212424
rect 604454 212372 604460 212424
rect 604512 212412 604518 212424
rect 605098 212412 605104 212424
rect 604512 212384 605104 212412
rect 604512 212372 604518 212384
rect 605098 212372 605104 212384
rect 605156 212372 605162 212424
rect 41322 211284 41328 211336
rect 41380 211324 41386 211336
rect 41690 211324 41696 211336
rect 41380 211296 41696 211324
rect 41380 211284 41386 211296
rect 41690 211284 41696 211296
rect 41748 211284 41754 211336
rect 41138 211148 41144 211200
rect 41196 211188 41202 211200
rect 41506 211188 41512 211200
rect 41196 211160 41512 211188
rect 41196 211148 41202 211160
rect 41506 211148 41512 211160
rect 41564 211148 41570 211200
rect 578510 211148 578516 211200
rect 578568 211188 578574 211200
rect 580902 211188 580908 211200
rect 578568 211160 580908 211188
rect 578568 211148 578574 211160
rect 580902 211148 580908 211160
rect 580960 211148 580966 211200
rect 603258 211012 603264 211064
rect 603316 211052 603322 211064
rect 603626 211052 603632 211064
rect 603316 211024 603632 211052
rect 603316 211012 603322 211024
rect 603626 211012 603632 211024
rect 603684 211012 603690 211064
rect 605834 210060 605840 210112
rect 605892 210100 605898 210112
rect 606202 210100 606208 210112
rect 605892 210072 606208 210100
rect 605892 210060 605898 210072
rect 606202 210060 606208 210072
rect 606260 210060 606266 210112
rect 622394 210060 622400 210112
rect 622452 210100 622458 210112
rect 622762 210100 622768 210112
rect 622452 210072 622768 210100
rect 622452 210060 622458 210072
rect 622762 210060 622768 210072
rect 622820 210060 622826 210112
rect 578418 209788 578424 209840
rect 578476 209828 578482 209840
rect 580074 209828 580080 209840
rect 578476 209800 580080 209828
rect 578476 209788 578482 209800
rect 580074 209788 580080 209800
rect 580132 209788 580138 209840
rect 652202 209692 652208 209704
rect 651852 209664 652208 209692
rect 632146 209556 632152 209568
rect 625126 209528 632152 209556
rect 580258 208564 580264 208616
rect 580316 208604 580322 208616
rect 625126 208604 625154 209528
rect 632146 209516 632152 209528
rect 632204 209516 632210 209568
rect 651852 209420 651880 209664
rect 652202 209652 652208 209664
rect 652260 209652 652266 209704
rect 652018 209516 652024 209568
rect 652076 209556 652082 209568
rect 652076 209528 654134 209556
rect 652076 209516 652082 209528
rect 651852 209392 651972 209420
rect 651944 209080 651972 209392
rect 654106 209216 654134 209528
rect 666830 209216 666836 209228
rect 654106 209188 666836 209216
rect 666830 209176 666836 209188
rect 666888 209176 666894 209228
rect 667014 209080 667020 209092
rect 651944 209052 667020 209080
rect 667014 209040 667020 209052
rect 667072 209040 667078 209092
rect 580316 208576 625154 208604
rect 580316 208564 580322 208576
rect 578878 208292 578884 208344
rect 578936 208332 578942 208344
rect 589458 208332 589464 208344
rect 578936 208304 589464 208332
rect 578936 208292 578942 208304
rect 589458 208292 589464 208304
rect 589516 208292 589522 208344
rect 580074 207612 580080 207664
rect 580132 207652 580138 207664
rect 589642 207652 589648 207664
rect 580132 207624 589648 207652
rect 580132 207612 580138 207624
rect 589642 207612 589648 207624
rect 589700 207612 589706 207664
rect 580902 206864 580908 206916
rect 580960 206904 580966 206916
rect 589458 206904 589464 206916
rect 580960 206876 589464 206904
rect 580960 206864 580966 206876
rect 589458 206864 589464 206876
rect 589516 206864 589522 206916
rect 579522 205776 579528 205828
rect 579580 205816 579586 205828
rect 582374 205816 582380 205828
rect 579580 205788 582380 205816
rect 579580 205776 579586 205788
rect 582374 205776 582380 205788
rect 582432 205776 582438 205828
rect 579706 204212 579712 204264
rect 579764 204252 579770 204264
rect 589458 204252 589464 204264
rect 579764 204224 589464 204252
rect 579764 204212 579770 204224
rect 589458 204212 589464 204224
rect 589516 204212 589522 204264
rect 578510 202920 578516 202972
rect 578568 202960 578574 202972
rect 580442 202960 580448 202972
rect 578568 202932 580448 202960
rect 578568 202920 578574 202932
rect 580442 202920 580448 202932
rect 580500 202920 580506 202972
rect 582374 202784 582380 202836
rect 582432 202824 582438 202836
rect 589458 202824 589464 202836
rect 582432 202796 589464 202824
rect 582432 202784 582438 202796
rect 589458 202784 589464 202796
rect 589516 202784 589522 202836
rect 578786 200132 578792 200184
rect 578844 200172 578850 200184
rect 590378 200172 590384 200184
rect 578844 200144 590384 200172
rect 578844 200132 578850 200144
rect 590378 200132 590384 200144
rect 590436 200132 590442 200184
rect 580442 199996 580448 200048
rect 580500 200036 580506 200048
rect 589458 200036 589464 200048
rect 580500 200008 589464 200036
rect 580500 199996 580506 200008
rect 589458 199996 589464 200008
rect 589516 199996 589522 200048
rect 579522 198704 579528 198756
rect 579580 198744 579586 198756
rect 589458 198744 589464 198756
rect 579580 198716 589464 198744
rect 579580 198704 579586 198716
rect 589458 198704 589464 198716
rect 589516 198704 589522 198756
rect 578510 195984 578516 196036
rect 578568 196024 578574 196036
rect 589274 196024 589280 196036
rect 578568 195996 589280 196024
rect 578568 195984 578574 195996
rect 589274 195984 589280 195996
rect 589332 195984 589338 196036
rect 579522 194556 579528 194608
rect 579580 194596 579586 194608
rect 589458 194596 589464 194608
rect 579580 194568 589464 194596
rect 579580 194556 579586 194568
rect 589458 194556 589464 194568
rect 589516 194556 589522 194608
rect 668026 192448 668032 192500
rect 668084 192488 668090 192500
rect 669314 192488 669320 192500
rect 668084 192460 669320 192488
rect 668084 192448 668090 192460
rect 669314 192448 669320 192460
rect 669372 192448 669378 192500
rect 579522 191836 579528 191888
rect 579580 191876 579586 191888
rect 589458 191876 589464 191888
rect 579580 191848 589464 191876
rect 579580 191836 579586 191848
rect 589458 191836 589464 191848
rect 589516 191836 589522 191888
rect 579522 190476 579528 190528
rect 579580 190516 579586 190528
rect 590562 190516 590568 190528
rect 579580 190488 590568 190516
rect 579580 190476 579586 190488
rect 590562 190476 590568 190488
rect 590620 190476 590626 190528
rect 669130 188436 669136 188488
rect 669188 188436 669194 188488
rect 669148 188204 669176 188436
rect 669314 188204 669320 188216
rect 669148 188176 669320 188204
rect 669314 188164 669320 188176
rect 669372 188164 669378 188216
rect 579522 187688 579528 187740
rect 579580 187728 579586 187740
rect 589458 187728 589464 187740
rect 579580 187700 589464 187728
rect 579580 187688 579586 187700
rect 589458 187688 589464 187700
rect 589516 187688 589522 187740
rect 579522 186260 579528 186312
rect 579580 186300 579586 186312
rect 589642 186300 589648 186312
rect 579580 186272 589648 186300
rect 579580 186260 579586 186272
rect 589642 186260 589648 186272
rect 589700 186260 589706 186312
rect 579522 184832 579528 184884
rect 579580 184872 579586 184884
rect 589458 184872 589464 184884
rect 579580 184844 589464 184872
rect 579580 184832 579586 184844
rect 589458 184832 589464 184844
rect 589516 184832 589522 184884
rect 667934 184492 667940 184544
rect 667992 184532 667998 184544
rect 669590 184532 669596 184544
rect 667992 184504 669596 184532
rect 667992 184492 667998 184504
rect 669590 184492 669596 184504
rect 669648 184492 669654 184544
rect 579522 182112 579528 182164
rect 579580 182152 579586 182164
rect 589458 182152 589464 182164
rect 579580 182124 589464 182152
rect 579580 182112 579586 182124
rect 589458 182112 589464 182124
rect 589516 182112 589522 182164
rect 578786 180752 578792 180804
rect 578844 180792 578850 180804
rect 590562 180792 590568 180804
rect 578844 180764 590568 180792
rect 578844 180752 578850 180764
rect 590562 180752 590568 180764
rect 590620 180752 590626 180804
rect 578786 178032 578792 178084
rect 578844 178072 578850 178084
rect 589458 178072 589464 178084
rect 578844 178044 589464 178072
rect 578844 178032 578850 178044
rect 589458 178032 589464 178044
rect 589516 178032 589522 178084
rect 579522 177896 579528 177948
rect 579580 177936 579586 177948
rect 589642 177936 589648 177948
rect 579580 177908 589648 177936
rect 579580 177896 579586 177908
rect 589642 177896 589648 177908
rect 589700 177896 589706 177948
rect 589458 175352 589464 175364
rect 586486 175324 589464 175352
rect 582374 175244 582380 175296
rect 582432 175284 582438 175296
rect 586486 175284 586514 175324
rect 589458 175312 589464 175324
rect 589516 175312 589522 175364
rect 582432 175256 586514 175284
rect 582432 175244 582438 175256
rect 667934 174836 667940 174888
rect 667992 174876 667998 174888
rect 669774 174876 669780 174888
rect 667992 174848 669780 174876
rect 667992 174836 667998 174848
rect 669774 174836 669780 174848
rect 669832 174836 669838 174888
rect 578418 174496 578424 174548
rect 578476 174536 578482 174548
rect 589642 174536 589648 174548
rect 578476 174508 589648 174536
rect 578476 174496 578482 174508
rect 589642 174496 589648 174508
rect 589700 174496 589706 174548
rect 578234 173204 578240 173256
rect 578292 173244 578298 173256
rect 582374 173244 582380 173256
rect 578292 173216 582380 173244
rect 578292 173204 578298 173216
rect 582374 173204 582380 173216
rect 582432 173204 582438 173256
rect 589458 172564 589464 172576
rect 582392 172536 589464 172564
rect 578418 172456 578424 172508
rect 578476 172496 578482 172508
rect 582392 172496 582420 172536
rect 589458 172524 589464 172536
rect 589516 172524 589522 172576
rect 578476 172468 582420 172496
rect 578476 172456 578482 172468
rect 579798 171096 579804 171148
rect 579856 171136 579862 171148
rect 589458 171136 589464 171148
rect 579856 171108 589464 171136
rect 579856 171096 579862 171108
rect 589458 171096 589464 171108
rect 589516 171096 589522 171148
rect 668026 169668 668032 169720
rect 668084 169708 668090 169720
rect 670326 169708 670332 169720
rect 668084 169680 670332 169708
rect 668084 169668 668090 169680
rect 670326 169668 670332 169680
rect 670384 169668 670390 169720
rect 582374 167016 582380 167068
rect 582432 167056 582438 167068
rect 589458 167056 589464 167068
rect 582432 167028 589464 167056
rect 582432 167016 582438 167028
rect 589458 167016 589464 167028
rect 589516 167016 589522 167068
rect 579522 166268 579528 166320
rect 579580 166308 579586 166320
rect 589182 166308 589188 166320
rect 579580 166280 589188 166308
rect 579580 166268 579586 166280
rect 589182 166268 589188 166280
rect 589240 166268 589246 166320
rect 667934 165180 667940 165232
rect 667992 165220 667998 165232
rect 670142 165220 670148 165232
rect 667992 165192 670148 165220
rect 667992 165180 667998 165192
rect 670142 165180 670148 165192
rect 670200 165180 670206 165232
rect 579338 164840 579344 164892
rect 579396 164880 579402 164892
rect 589826 164880 589832 164892
rect 579396 164852 589832 164880
rect 579396 164840 579402 164852
rect 589826 164840 589832 164852
rect 589884 164840 589890 164892
rect 580902 162868 580908 162920
rect 580960 162908 580966 162920
rect 589458 162908 589464 162920
rect 580960 162880 589464 162908
rect 580960 162868 580966 162880
rect 589458 162868 589464 162880
rect 589516 162868 589522 162920
rect 578234 162528 578240 162580
rect 578292 162568 578298 162580
rect 582374 162568 582380 162580
rect 578292 162540 582380 162568
rect 578292 162528 578298 162540
rect 582374 162528 582380 162540
rect 582432 162528 582438 162580
rect 675846 162528 675852 162580
rect 675904 162568 675910 162580
rect 680998 162568 681004 162580
rect 675904 162540 681004 162568
rect 675904 162528 675910 162540
rect 680998 162528 681004 162540
rect 681056 162528 681062 162580
rect 578418 162120 578424 162172
rect 578476 162160 578482 162172
rect 589642 162160 589648 162172
rect 578476 162132 589648 162160
rect 578476 162120 578482 162132
rect 589642 162120 589648 162132
rect 589700 162120 589706 162172
rect 582374 160080 582380 160132
rect 582432 160120 582438 160132
rect 589458 160120 589464 160132
rect 582432 160092 589464 160120
rect 582432 160080 582438 160092
rect 589458 160080 589464 160092
rect 589516 160080 589522 160132
rect 667934 160012 667940 160064
rect 667992 160052 667998 160064
rect 669958 160052 669964 160064
rect 667992 160024 669964 160052
rect 667992 160012 667998 160024
rect 669958 160012 669964 160024
rect 670016 160012 670022 160064
rect 583754 159332 583760 159384
rect 583812 159372 583818 159384
rect 590562 159372 590568 159384
rect 583812 159344 590568 159372
rect 583812 159332 583818 159344
rect 590562 159332 590568 159344
rect 590620 159332 590626 159384
rect 578510 157564 578516 157616
rect 578568 157604 578574 157616
rect 580902 157604 580908 157616
rect 578568 157576 580908 157604
rect 578568 157564 578574 157576
rect 580902 157564 580908 157576
rect 580960 157564 580966 157616
rect 587158 157360 587164 157412
rect 587216 157400 587222 157412
rect 589274 157400 589280 157412
rect 587216 157372 589280 157400
rect 587216 157360 587222 157372
rect 589274 157360 589280 157372
rect 589332 157360 589338 157412
rect 585778 154572 585784 154624
rect 585836 154612 585842 154624
rect 589458 154612 589464 154624
rect 585836 154584 589464 154612
rect 585836 154572 585842 154584
rect 589458 154572 589464 154584
rect 589516 154572 589522 154624
rect 578694 154164 578700 154216
rect 578752 154204 578758 154216
rect 583754 154204 583760 154216
rect 578752 154176 583760 154204
rect 578752 154164 578758 154176
rect 583754 154164 583760 154176
rect 583812 154164 583818 154216
rect 584398 153212 584404 153264
rect 584456 153252 584462 153264
rect 589458 153252 589464 153264
rect 584456 153224 589464 153252
rect 584456 153212 584462 153224
rect 589458 153212 589464 153224
rect 589516 153212 589522 153264
rect 578234 152600 578240 152652
rect 578292 152640 578298 152652
rect 582374 152640 582380 152652
rect 578292 152612 582380 152640
rect 578292 152600 578298 152612
rect 582374 152600 582380 152612
rect 582432 152600 582438 152652
rect 583018 151784 583024 151836
rect 583076 151824 583082 151836
rect 589458 151824 589464 151836
rect 583076 151796 589464 151824
rect 583076 151784 583082 151796
rect 589458 151784 589464 151796
rect 589516 151784 589522 151836
rect 578326 151036 578332 151088
rect 578384 151076 578390 151088
rect 588538 151076 588544 151088
rect 578384 151048 588544 151076
rect 578384 151036 578390 151048
rect 588538 151036 588544 151048
rect 588596 151036 588602 151088
rect 668302 150220 668308 150272
rect 668360 150260 668366 150272
rect 670786 150260 670792 150272
rect 668360 150232 670792 150260
rect 668360 150220 668366 150232
rect 670786 150220 670792 150232
rect 670844 150220 670850 150272
rect 579522 148316 579528 148368
rect 579580 148356 579586 148368
rect 587158 148356 587164 148368
rect 579580 148328 587164 148356
rect 579580 148316 579586 148328
rect 587158 148316 587164 148328
rect 587216 148316 587222 148368
rect 585962 146276 585968 146328
rect 586020 146316 586026 146328
rect 589458 146316 589464 146328
rect 586020 146288 589464 146316
rect 586020 146276 586026 146288
rect 589458 146276 589464 146288
rect 589516 146276 589522 146328
rect 578878 145528 578884 145580
rect 578936 145568 578942 145580
rect 589182 145568 589188 145580
rect 578936 145540 589188 145568
rect 578936 145528 578942 145540
rect 589182 145528 589188 145540
rect 589240 145528 589246 145580
rect 579430 144644 579436 144696
rect 579488 144684 579494 144696
rect 585778 144684 585784 144696
rect 579488 144656 585784 144684
rect 579488 144644 579494 144656
rect 585778 144644 585784 144656
rect 585836 144644 585842 144696
rect 587158 143556 587164 143608
rect 587216 143596 587222 143608
rect 589458 143596 589464 143608
rect 587216 143568 589464 143596
rect 587216 143556 587222 143568
rect 589458 143556 589464 143568
rect 589516 143556 589522 143608
rect 579522 143420 579528 143472
rect 579580 143460 579586 143472
rect 584398 143460 584404 143472
rect 579580 143432 584404 143460
rect 579580 143420 579586 143432
rect 584398 143420 584404 143432
rect 584456 143420 584462 143472
rect 583202 140768 583208 140820
rect 583260 140808 583266 140820
rect 589458 140808 589464 140820
rect 583260 140780 589464 140808
rect 583260 140768 583266 140780
rect 589458 140768 589464 140780
rect 589516 140768 589522 140820
rect 579522 140564 579528 140616
rect 579580 140604 579586 140616
rect 583018 140604 583024 140616
rect 579580 140576 583024 140604
rect 579580 140564 579586 140576
rect 583018 140564 583024 140576
rect 583076 140564 583082 140616
rect 584398 139408 584404 139460
rect 584456 139448 584462 139460
rect 589458 139448 589464 139460
rect 584456 139420 589464 139448
rect 584456 139408 584462 139420
rect 589458 139408 589464 139420
rect 589516 139408 589522 139460
rect 578602 139272 578608 139324
rect 578660 139312 578666 139324
rect 589918 139312 589924 139324
rect 578660 139284 589924 139312
rect 578660 139272 578666 139284
rect 589918 139272 589924 139284
rect 589976 139272 589982 139324
rect 579522 138116 579528 138168
rect 579580 138156 579586 138168
rect 585962 138156 585968 138168
rect 579580 138128 585968 138156
rect 579580 138116 579586 138128
rect 585962 138116 585968 138128
rect 586020 138116 586026 138168
rect 580442 137368 580448 137420
rect 580500 137408 580506 137420
rect 589642 137408 589648 137420
rect 580500 137380 589648 137408
rect 580500 137368 580506 137380
rect 589642 137368 589648 137380
rect 589700 137368 589706 137420
rect 579062 137232 579068 137284
rect 579120 137272 579126 137284
rect 588722 137272 588728 137284
rect 579120 137244 588728 137272
rect 579120 137232 579126 137244
rect 588722 137232 588728 137244
rect 588780 137232 588786 137284
rect 585962 135260 585968 135312
rect 586020 135300 586026 135312
rect 589458 135300 589464 135312
rect 586020 135272 589464 135300
rect 586020 135260 586026 135272
rect 589458 135260 589464 135272
rect 589516 135260 589522 135312
rect 581822 131860 581828 131912
rect 581880 131900 581886 131912
rect 590286 131900 590292 131912
rect 581880 131872 590292 131900
rect 581880 131860 581886 131872
rect 590286 131860 590292 131872
rect 590344 131860 590350 131912
rect 578694 131724 578700 131776
rect 578752 131764 578758 131776
rect 587158 131764 587164 131776
rect 578752 131736 587164 131764
rect 578752 131724 578758 131736
rect 587158 131724 587164 131736
rect 587216 131724 587222 131776
rect 587526 131112 587532 131164
rect 587584 131152 587590 131164
rect 590102 131152 590108 131164
rect 587584 131124 590108 131152
rect 587584 131112 587590 131124
rect 590102 131112 590108 131124
rect 590160 131112 590166 131164
rect 578510 127984 578516 128036
rect 578568 128024 578574 128036
rect 580442 128024 580448 128036
rect 578568 127996 580448 128024
rect 578568 127984 578574 127996
rect 580442 127984 580448 127996
rect 580500 127984 580506 128036
rect 579062 126964 579068 127016
rect 579120 127004 579126 127016
rect 589458 127004 589464 127016
rect 579120 126976 589464 127004
rect 579120 126964 579126 126976
rect 589458 126964 589464 126976
rect 589516 126964 589522 127016
rect 580626 125604 580632 125656
rect 580684 125644 580690 125656
rect 589458 125644 589464 125656
rect 580684 125616 589464 125644
rect 580684 125604 580690 125616
rect 589458 125604 589464 125616
rect 589516 125604 589522 125656
rect 579522 125332 579528 125384
rect 579580 125372 579586 125384
rect 583202 125372 583208 125384
rect 579580 125344 583208 125372
rect 579580 125332 579586 125344
rect 583202 125332 583208 125344
rect 583260 125332 583266 125384
rect 583018 124856 583024 124908
rect 583076 124896 583082 124908
rect 589274 124896 589280 124908
rect 583076 124868 589280 124896
rect 583076 124856 583082 124868
rect 589274 124856 589280 124868
rect 589332 124856 589338 124908
rect 579246 124108 579252 124160
rect 579304 124148 579310 124160
rect 584398 124148 584404 124160
rect 579304 124120 584404 124148
rect 579304 124108 579310 124120
rect 584398 124108 584404 124120
rect 584456 124108 584462 124160
rect 584582 122816 584588 122868
rect 584640 122856 584646 122868
rect 589458 122856 589464 122868
rect 584640 122828 589464 122856
rect 584640 122816 584646 122828
rect 589458 122816 589464 122828
rect 589516 122816 589522 122868
rect 578878 122204 578884 122256
rect 578936 122244 578942 122256
rect 587526 122244 587532 122256
rect 578936 122216 587532 122244
rect 578936 122204 578942 122216
rect 587526 122204 587532 122216
rect 587584 122204 587590 122256
rect 580442 122068 580448 122120
rect 580500 122108 580506 122120
rect 589734 122108 589740 122120
rect 580500 122080 589740 122108
rect 580500 122068 580506 122080
rect 589734 122068 589740 122080
rect 589792 122068 589798 122120
rect 587342 121456 587348 121508
rect 587400 121496 587406 121508
rect 589274 121496 589280 121508
rect 587400 121468 589280 121496
rect 587400 121456 587406 121468
rect 589274 121456 589280 121468
rect 589332 121456 589338 121508
rect 578510 121320 578516 121372
rect 578568 121360 578574 121372
rect 588538 121360 588544 121372
rect 578568 121332 588544 121360
rect 578568 121320 578574 121332
rect 588538 121320 588544 121332
rect 588596 121320 588602 121372
rect 667934 120708 667940 120760
rect 667992 120748 667998 120760
rect 669774 120748 669780 120760
rect 667992 120720 669780 120748
rect 667992 120708 667998 120720
rect 669774 120708 669780 120720
rect 669832 120708 669838 120760
rect 579522 118396 579528 118448
rect 579580 118436 579586 118448
rect 585962 118436 585968 118448
rect 579580 118408 585968 118436
rect 579580 118396 579586 118408
rect 585962 118396 585968 118408
rect 586020 118396 586026 118448
rect 667934 118056 667940 118108
rect 667992 118096 667998 118108
rect 670142 118096 670148 118108
rect 667992 118068 670148 118096
rect 667992 118056 667998 118068
rect 670142 118056 670148 118068
rect 670200 118056 670206 118108
rect 585778 117308 585784 117360
rect 585836 117348 585842 117360
rect 589458 117348 589464 117360
rect 585836 117320 589464 117348
rect 585836 117308 585842 117320
rect 589458 117308 589464 117320
rect 589516 117308 589522 117360
rect 675846 117240 675852 117292
rect 675904 117280 675910 117292
rect 679618 117280 679624 117292
rect 675904 117252 679624 117280
rect 675904 117240 675910 117252
rect 679618 117240 679624 117252
rect 679676 117240 679682 117292
rect 579338 117172 579344 117224
rect 579396 117212 579402 117224
rect 581822 117212 581828 117224
rect 579396 117184 581828 117212
rect 579396 117172 579402 117184
rect 581822 117172 581828 117184
rect 581880 117172 581886 117224
rect 585962 115948 585968 116000
rect 586020 115988 586026 116000
rect 589458 115988 589464 116000
rect 586020 115960 589464 115988
rect 586020 115948 586026 115960
rect 589458 115948 589464 115960
rect 589516 115948 589522 116000
rect 578510 114452 578516 114504
rect 578568 114492 578574 114504
rect 580258 114492 580264 114504
rect 578568 114464 580264 114492
rect 578568 114452 578574 114464
rect 580258 114452 580264 114464
rect 580316 114452 580322 114504
rect 588538 113704 588544 113756
rect 588596 113744 588602 113756
rect 589550 113744 589556 113756
rect 588596 113716 589556 113744
rect 588596 113704 588602 113716
rect 589550 113704 589556 113716
rect 589608 113704 589614 113756
rect 579522 113092 579528 113144
rect 579580 113132 579586 113144
rect 589918 113132 589924 113144
rect 579580 113104 589924 113132
rect 579580 113092 579586 113104
rect 589918 113092 589924 113104
rect 589976 113092 589982 113144
rect 667934 111392 667940 111444
rect 667992 111432 667998 111444
rect 669958 111432 669964 111444
rect 667992 111404 669964 111432
rect 667992 111392 667998 111404
rect 669958 111392 669964 111404
rect 670016 111392 670022 111444
rect 583202 111052 583208 111104
rect 583260 111092 583266 111104
rect 590286 111092 590292 111104
rect 583260 111064 590292 111092
rect 583260 111052 583266 111064
rect 590286 111052 590292 111064
rect 590344 111052 590350 111104
rect 581822 109692 581828 109744
rect 581880 109732 581886 109744
rect 589366 109732 589372 109744
rect 581880 109704 589372 109732
rect 581880 109692 581886 109704
rect 589366 109692 589372 109704
rect 589424 109692 589430 109744
rect 578326 108672 578332 108724
rect 578384 108712 578390 108724
rect 580626 108712 580632 108724
rect 578384 108684 580632 108712
rect 578384 108672 578390 108684
rect 580626 108672 580632 108684
rect 580684 108672 580690 108724
rect 583754 107652 583760 107704
rect 583812 107692 583818 107704
rect 589458 107692 589464 107704
rect 583812 107664 589464 107692
rect 583812 107652 583818 107664
rect 589458 107652 589464 107664
rect 589516 107652 589522 107704
rect 580258 106292 580264 106344
rect 580316 106332 580322 106344
rect 589458 106332 589464 106344
rect 580316 106304 589464 106332
rect 580316 106292 580322 106304
rect 589458 106292 589464 106304
rect 589516 106292 589522 106344
rect 668394 106156 668400 106208
rect 668452 106196 668458 106208
rect 670786 106196 670792 106208
rect 668452 106168 670792 106196
rect 668452 106156 668458 106168
rect 670786 106156 670792 106168
rect 670844 106156 670850 106208
rect 579430 105136 579436 105188
rect 579488 105176 579494 105188
rect 583754 105176 583760 105188
rect 579488 105148 583760 105176
rect 579488 105136 579494 105148
rect 583754 105136 583760 105148
rect 583812 105136 583818 105188
rect 587158 104864 587164 104916
rect 587216 104904 587222 104916
rect 589826 104904 589832 104916
rect 587216 104876 589832 104904
rect 587216 104864 587222 104876
rect 589826 104864 589832 104876
rect 589884 104864 589890 104916
rect 579246 103300 579252 103352
rect 579304 103340 579310 103352
rect 583018 103340 583024 103352
rect 579304 103312 583024 103340
rect 579304 103300 579310 103312
rect 583018 103300 583024 103312
rect 583076 103300 583082 103352
rect 578326 101668 578332 101720
rect 578384 101708 578390 101720
rect 584582 101708 584588 101720
rect 578384 101680 584588 101708
rect 578384 101668 578390 101680
rect 584582 101668 584588 101680
rect 584640 101668 584646 101720
rect 584398 101396 584404 101448
rect 584456 101436 584462 101448
rect 590286 101436 590292 101448
rect 584456 101408 590292 101436
rect 584456 101396 584462 101408
rect 590286 101396 590292 101408
rect 590344 101396 590350 101448
rect 624786 100104 624792 100156
rect 624844 100144 624850 100156
rect 667934 100144 667940 100156
rect 624844 100116 667940 100144
rect 624844 100104 624850 100116
rect 667934 100104 667940 100116
rect 667992 100104 667998 100156
rect 668118 100008 668124 100020
rect 615466 99980 668124 100008
rect 614850 99900 614856 99952
rect 614908 99940 614914 99952
rect 615466 99940 615494 99980
rect 668118 99968 668124 99980
rect 668176 99968 668182 100020
rect 614908 99912 615494 99940
rect 614908 99900 614914 99912
rect 578602 99288 578608 99340
rect 578660 99328 578666 99340
rect 580442 99328 580448 99340
rect 578660 99300 580448 99328
rect 578660 99288 578666 99300
rect 580442 99288 580448 99300
rect 580500 99288 580506 99340
rect 622302 99288 622308 99340
rect 622360 99328 622366 99340
rect 630766 99328 630772 99340
rect 622360 99300 630772 99328
rect 622360 99288 622366 99300
rect 630766 99288 630772 99300
rect 630824 99288 630830 99340
rect 623682 99152 623688 99204
rect 623740 99192 623746 99204
rect 633526 99192 633532 99204
rect 623740 99164 633532 99192
rect 623740 99152 623746 99164
rect 633526 99152 633532 99164
rect 633584 99152 633590 99204
rect 625062 99016 625068 99068
rect 625120 99056 625126 99068
rect 636286 99056 636292 99068
rect 625120 99028 636292 99056
rect 625120 99016 625126 99028
rect 636286 99016 636292 99028
rect 636344 99016 636350 99068
rect 627546 98880 627552 98932
rect 627604 98920 627610 98932
rect 640702 98920 640708 98932
rect 627604 98892 640708 98920
rect 627604 98880 627610 98892
rect 640702 98880 640708 98892
rect 640760 98880 640766 98932
rect 579246 98744 579252 98796
rect 579304 98784 579310 98796
rect 587342 98784 587348 98796
rect 579304 98756 587348 98784
rect 579304 98744 579310 98756
rect 587342 98744 587348 98756
rect 587400 98744 587406 98796
rect 629018 98744 629024 98796
rect 629076 98784 629082 98796
rect 643646 98784 643652 98796
rect 629076 98756 643652 98784
rect 629076 98744 629082 98756
rect 643646 98744 643652 98756
rect 643704 98744 643710 98796
rect 580626 98608 580632 98660
rect 580684 98648 580690 98660
rect 590102 98648 590108 98660
rect 580684 98620 590108 98648
rect 580684 98608 580690 98620
rect 590102 98608 590108 98620
rect 590160 98608 590166 98660
rect 647142 98608 647148 98660
rect 647200 98648 647206 98660
rect 661954 98648 661960 98660
rect 647200 98620 661960 98648
rect 647200 98608 647206 98620
rect 661954 98608 661960 98620
rect 662012 98608 662018 98660
rect 630490 98472 630496 98524
rect 630548 98512 630554 98524
rect 646590 98512 646596 98524
rect 630548 98484 646596 98512
rect 630548 98472 630554 98484
rect 646590 98472 646596 98484
rect 646648 98472 646654 98524
rect 631410 98200 631416 98252
rect 631468 98240 631474 98252
rect 642174 98240 642180 98252
rect 631468 98212 642180 98240
rect 631468 98200 631474 98212
rect 642174 98200 642180 98212
rect 642232 98200 642238 98252
rect 595254 98104 595260 98116
rect 592512 98076 595260 98104
rect 581638 97928 581644 97980
rect 581696 97968 581702 97980
rect 592512 97968 592540 98076
rect 595254 98064 595260 98076
rect 595312 98064 595318 98116
rect 631980 98076 634814 98104
rect 581696 97940 592540 97968
rect 581696 97928 581702 97940
rect 592678 97928 592684 97980
rect 592736 97968 592742 97980
rect 597554 97968 597560 97980
rect 592736 97940 597560 97968
rect 592736 97928 592742 97940
rect 597554 97928 597560 97940
rect 597612 97928 597618 97980
rect 618714 97928 618720 97980
rect 618772 97968 618778 97980
rect 625798 97968 625804 97980
rect 618772 97940 625804 97968
rect 618772 97928 618778 97940
rect 625798 97928 625804 97940
rect 625856 97928 625862 97980
rect 629754 97928 629760 97980
rect 629812 97968 629818 97980
rect 631980 97968 632008 98076
rect 634786 98036 634814 98076
rect 645302 98036 645308 98048
rect 634786 98008 645308 98036
rect 645302 97996 645308 98008
rect 645360 97996 645366 98048
rect 629812 97940 632008 97968
rect 629812 97928 629818 97940
rect 592862 97792 592868 97844
rect 592920 97832 592926 97844
rect 598198 97832 598204 97844
rect 592920 97804 598204 97832
rect 592920 97792 592926 97804
rect 598198 97792 598204 97804
rect 598256 97792 598262 97844
rect 628282 97792 628288 97844
rect 628340 97832 628346 97844
rect 631410 97832 631416 97844
rect 628340 97804 631416 97832
rect 628340 97792 628346 97804
rect 631410 97792 631416 97804
rect 631468 97792 631474 97844
rect 633342 97792 633348 97844
rect 633400 97832 633406 97844
rect 650546 97832 650552 97844
rect 633400 97804 650552 97832
rect 633400 97792 633406 97804
rect 650546 97792 650552 97804
rect 650604 97792 650610 97844
rect 653950 97792 653956 97844
rect 654008 97832 654014 97844
rect 655054 97832 655060 97844
rect 654008 97804 655060 97832
rect 654008 97792 654014 97804
rect 655054 97792 655060 97804
rect 655112 97792 655118 97844
rect 659194 97792 659200 97844
rect 659252 97832 659258 97844
rect 663886 97832 663892 97844
rect 659252 97804 663892 97832
rect 659252 97792 659258 97804
rect 663886 97792 663892 97804
rect 663944 97792 663950 97844
rect 590102 97656 590108 97708
rect 590160 97696 590166 97708
rect 600406 97696 600412 97708
rect 590160 97668 600412 97696
rect 590160 97656 590166 97668
rect 600406 97656 600412 97668
rect 600464 97656 600470 97708
rect 626074 97656 626080 97708
rect 626132 97696 626138 97708
rect 637758 97696 637764 97708
rect 626132 97668 637764 97696
rect 626132 97656 626138 97668
rect 637758 97656 637764 97668
rect 637816 97656 637822 97708
rect 643002 97656 643008 97708
rect 643060 97696 643066 97708
rect 659746 97696 659752 97708
rect 643060 97668 659752 97696
rect 643060 97656 643066 97668
rect 659746 97656 659752 97668
rect 659804 97656 659810 97708
rect 659930 97656 659936 97708
rect 659988 97696 659994 97708
rect 665358 97696 665364 97708
rect 659988 97668 665364 97696
rect 659988 97656 659994 97668
rect 665358 97656 665364 97668
rect 665416 97656 665422 97708
rect 583018 97520 583024 97572
rect 583076 97560 583082 97572
rect 596174 97560 596180 97572
rect 583076 97532 596180 97560
rect 583076 97520 583082 97532
rect 596174 97520 596180 97532
rect 596232 97520 596238 97572
rect 623130 97520 623136 97572
rect 623188 97560 623194 97572
rect 632054 97560 632060 97572
rect 623188 97532 632060 97560
rect 623188 97520 623194 97532
rect 632054 97520 632060 97532
rect 632112 97520 632118 97572
rect 634722 97520 634728 97572
rect 634780 97560 634786 97572
rect 649074 97560 649080 97572
rect 634780 97532 649080 97560
rect 634780 97520 634786 97532
rect 649074 97520 649080 97532
rect 649132 97520 649138 97572
rect 651834 97520 651840 97572
rect 651892 97560 651898 97572
rect 659562 97560 659568 97572
rect 651892 97532 659568 97560
rect 651892 97520 651898 97532
rect 659562 97520 659568 97532
rect 659620 97520 659626 97572
rect 577682 97384 577688 97436
rect 577740 97424 577746 97436
rect 596726 97424 596732 97436
rect 577740 97396 596732 97424
rect 577740 97384 577746 97396
rect 596726 97384 596732 97396
rect 596784 97384 596790 97436
rect 605466 97384 605472 97436
rect 605524 97424 605530 97436
rect 613378 97424 613384 97436
rect 605524 97396 613384 97424
rect 605524 97384 605530 97396
rect 613378 97384 613384 97396
rect 613436 97384 613442 97436
rect 620186 97384 620192 97436
rect 620244 97424 620250 97436
rect 625982 97424 625988 97436
rect 620244 97396 625988 97424
rect 620244 97384 620250 97396
rect 625982 97384 625988 97396
rect 626040 97384 626046 97436
rect 632698 97384 632704 97436
rect 632756 97424 632762 97436
rect 650178 97424 650184 97436
rect 632756 97396 650184 97424
rect 632756 97384 632762 97396
rect 650178 97384 650184 97396
rect 650236 97384 650242 97436
rect 658182 97384 658188 97436
rect 658240 97424 658246 97436
rect 663058 97424 663064 97436
rect 658240 97396 663064 97424
rect 658240 97384 658246 97396
rect 663058 97384 663064 97396
rect 663116 97384 663122 97436
rect 577498 97248 577504 97300
rect 577556 97288 577562 97300
rect 601878 97288 601884 97300
rect 577556 97260 601884 97288
rect 577556 97248 577562 97260
rect 601878 97248 601884 97260
rect 601936 97248 601942 97300
rect 612642 97248 612648 97300
rect 612700 97288 612706 97300
rect 620278 97288 620284 97300
rect 612700 97260 620284 97288
rect 612700 97248 612706 97260
rect 620278 97248 620284 97260
rect 620336 97248 620342 97300
rect 621658 97248 621664 97300
rect 621716 97288 621722 97300
rect 629294 97288 629300 97300
rect 621716 97260 629300 97288
rect 621716 97248 621722 97260
rect 629294 97248 629300 97260
rect 629352 97248 629358 97300
rect 631870 97248 631876 97300
rect 631928 97288 631934 97300
rect 648614 97288 648620 97300
rect 631928 97260 648620 97288
rect 631928 97248 631934 97260
rect 648614 97248 648620 97260
rect 648672 97248 648678 97300
rect 650362 97248 650368 97300
rect 650420 97288 650426 97300
rect 658274 97288 658280 97300
rect 650420 97260 658280 97288
rect 650420 97248 650426 97260
rect 658274 97248 658280 97260
rect 658332 97248 658338 97300
rect 634170 97112 634176 97164
rect 634228 97152 634234 97164
rect 647602 97152 647608 97164
rect 634228 97124 647608 97152
rect 634228 97112 634234 97124
rect 647602 97112 647608 97124
rect 647660 97112 647666 97164
rect 656802 97112 656808 97164
rect 656860 97152 656866 97164
rect 661402 97152 661408 97164
rect 656860 97124 661408 97152
rect 656860 97112 656866 97124
rect 661402 97112 661408 97124
rect 661460 97112 661466 97164
rect 615034 96976 615040 97028
rect 615092 97016 615098 97028
rect 616138 97016 616144 97028
rect 615092 96988 616144 97016
rect 615092 96976 615098 96988
rect 616138 96976 616144 96988
rect 616196 96976 616202 97028
rect 626810 96976 626816 97028
rect 626868 97016 626874 97028
rect 639230 97016 639236 97028
rect 626868 96988 639236 97016
rect 626868 96976 626874 96988
rect 639230 96976 639236 96988
rect 639288 96976 639294 97028
rect 644290 96976 644296 97028
rect 644348 97016 644354 97028
rect 658826 97016 658832 97028
rect 644348 96988 658832 97016
rect 644348 96976 644354 96988
rect 658826 96976 658832 96988
rect 658884 96976 658890 97028
rect 612090 96908 612096 96960
rect 612148 96948 612154 96960
rect 612642 96948 612648 96960
rect 612148 96920 612648 96948
rect 612148 96908 612154 96920
rect 612642 96908 612648 96920
rect 612700 96908 612706 96960
rect 617242 96908 617248 96960
rect 617300 96948 617306 96960
rect 618162 96948 618168 96960
rect 617300 96920 618168 96948
rect 617300 96908 617306 96920
rect 618162 96908 618168 96920
rect 618220 96908 618226 96960
rect 613562 96840 613568 96892
rect 613620 96880 613626 96892
rect 615034 96880 615040 96892
rect 613620 96852 615040 96880
rect 613620 96840 613626 96852
rect 615034 96840 615040 96852
rect 615092 96840 615098 96892
rect 624602 96840 624608 96892
rect 624660 96880 624666 96892
rect 634998 96880 635004 96892
rect 624660 96852 635004 96880
rect 624660 96840 624666 96852
rect 634998 96840 635004 96852
rect 635056 96840 635062 96892
rect 654778 96840 654784 96892
rect 654836 96880 654842 96892
rect 655422 96880 655428 96892
rect 654836 96852 655428 96880
rect 654836 96840 654842 96852
rect 655422 96840 655428 96852
rect 655480 96840 655486 96892
rect 660666 96840 660672 96892
rect 660724 96880 660730 96892
rect 663242 96880 663248 96892
rect 660724 96852 663248 96880
rect 660724 96840 660730 96852
rect 663242 96840 663248 96852
rect 663300 96840 663306 96892
rect 615770 96772 615776 96824
rect 615828 96812 615834 96824
rect 618898 96812 618904 96824
rect 615828 96784 618904 96812
rect 615828 96772 615834 96784
rect 618898 96772 618904 96784
rect 618956 96772 618962 96824
rect 606202 96704 606208 96756
rect 606260 96744 606266 96756
rect 607122 96744 607128 96756
rect 606260 96716 607128 96744
rect 606260 96704 606266 96716
rect 607122 96704 607128 96716
rect 607180 96704 607186 96756
rect 610618 96704 610624 96756
rect 610676 96744 610682 96756
rect 611170 96744 611176 96756
rect 610676 96716 611176 96744
rect 610676 96704 610682 96716
rect 611170 96704 611176 96716
rect 611228 96704 611234 96756
rect 638586 96704 638592 96756
rect 638644 96744 638650 96756
rect 647234 96744 647240 96756
rect 638644 96716 647240 96744
rect 638644 96704 638650 96716
rect 647234 96704 647240 96716
rect 647292 96704 647298 96756
rect 655238 96704 655244 96756
rect 655296 96744 655302 96756
rect 662506 96744 662512 96756
rect 655296 96716 662512 96744
rect 655296 96704 655302 96716
rect 662506 96704 662512 96716
rect 662564 96704 662570 96756
rect 639046 96568 639052 96620
rect 639104 96608 639110 96620
rect 649258 96608 649264 96620
rect 639104 96580 649264 96608
rect 639104 96568 639110 96580
rect 649258 96568 649264 96580
rect 649316 96568 649322 96620
rect 653306 96568 653312 96620
rect 653364 96608 653370 96620
rect 665174 96608 665180 96620
rect 653364 96580 665180 96608
rect 653364 96568 653370 96580
rect 665174 96568 665180 96580
rect 665232 96568 665238 96620
rect 640058 96432 640064 96484
rect 640116 96472 640122 96484
rect 645118 96472 645124 96484
rect 640116 96444 645124 96472
rect 640116 96432 640122 96444
rect 645118 96432 645124 96444
rect 645176 96432 645182 96484
rect 645762 96432 645768 96484
rect 645820 96472 645826 96484
rect 652018 96472 652024 96484
rect 645820 96444 652024 96472
rect 645820 96432 645826 96444
rect 652018 96432 652024 96444
rect 652076 96432 652082 96484
rect 652570 96432 652576 96484
rect 652628 96472 652634 96484
rect 664162 96472 664168 96484
rect 652628 96444 664168 96472
rect 652628 96432 652634 96444
rect 664162 96432 664168 96444
rect 664220 96432 664226 96484
rect 640518 96296 640524 96348
rect 640576 96336 640582 96348
rect 648430 96336 648436 96348
rect 640576 96308 648436 96336
rect 640576 96296 640582 96308
rect 648430 96296 648436 96308
rect 648488 96296 648494 96348
rect 648890 96296 648896 96348
rect 648948 96336 648954 96348
rect 664346 96336 664352 96348
rect 648948 96308 664352 96336
rect 648948 96296 648954 96308
rect 664346 96296 664352 96308
rect 664404 96296 664410 96348
rect 637574 96160 637580 96212
rect 637632 96200 637638 96212
rect 660666 96200 660672 96212
rect 637632 96172 660672 96200
rect 637632 96160 637638 96172
rect 660666 96160 660672 96172
rect 660724 96160 660730 96212
rect 641530 96024 641536 96076
rect 641588 96064 641594 96076
rect 663702 96064 663708 96076
rect 641588 96036 663708 96064
rect 641588 96024 641594 96036
rect 663702 96024 663708 96036
rect 663760 96024 663766 96076
rect 609146 95888 609152 95940
rect 609204 95928 609210 95940
rect 621658 95928 621664 95940
rect 609204 95900 621664 95928
rect 609204 95888 609210 95900
rect 621658 95888 621664 95900
rect 621716 95888 621722 95940
rect 644934 95888 644940 95940
rect 644992 95928 644998 95940
rect 648062 95928 648068 95940
rect 644992 95900 648068 95928
rect 644992 95888 644998 95900
rect 648062 95888 648068 95900
rect 648120 95888 648126 95940
rect 648430 95888 648436 95940
rect 648488 95928 648494 95940
rect 664530 95928 664536 95940
rect 648488 95900 664536 95928
rect 648488 95888 648494 95900
rect 664530 95888 664536 95900
rect 664588 95888 664594 95940
rect 645118 95752 645124 95804
rect 645176 95792 645182 95804
rect 652202 95792 652208 95804
rect 645176 95764 652208 95792
rect 645176 95752 645182 95764
rect 652202 95752 652208 95764
rect 652260 95752 652266 95804
rect 656158 95792 656164 95804
rect 654106 95764 656164 95792
rect 646406 95616 646412 95668
rect 646464 95656 646470 95668
rect 653398 95656 653404 95668
rect 646464 95628 653404 95656
rect 646464 95616 646470 95628
rect 653398 95616 653404 95628
rect 653456 95616 653462 95668
rect 648062 95480 648068 95532
rect 648120 95520 648126 95532
rect 654106 95520 654134 95764
rect 656158 95752 656164 95764
rect 656216 95752 656222 95804
rect 648120 95492 654134 95520
rect 648120 95480 648126 95492
rect 631226 95412 631232 95464
rect 631284 95452 631290 95464
rect 631284 95424 634814 95452
rect 631284 95412 631290 95424
rect 634786 95248 634814 95424
rect 643462 95412 643468 95464
rect 643520 95452 643526 95464
rect 647878 95452 647884 95464
rect 643520 95424 647884 95452
rect 643520 95412 643526 95424
rect 647878 95412 647884 95424
rect 647936 95412 647942 95464
rect 647142 95248 647148 95260
rect 634786 95220 647148 95248
rect 647142 95208 647148 95220
rect 647200 95208 647206 95260
rect 579246 95140 579252 95192
rect 579304 95180 579310 95192
rect 588722 95180 588728 95192
rect 579304 95152 588728 95180
rect 579304 95140 579310 95152
rect 588722 95140 588728 95152
rect 588780 95140 588786 95192
rect 620922 95140 620928 95192
rect 620980 95180 620986 95192
rect 626442 95180 626448 95192
rect 620980 95152 626448 95180
rect 620980 95140 620986 95152
rect 626442 95140 626448 95152
rect 626500 95140 626506 95192
rect 647602 95140 647608 95192
rect 647660 95180 647666 95192
rect 649994 95180 650000 95192
rect 647660 95152 650000 95180
rect 647660 95140 647666 95152
rect 649994 95140 650000 95152
rect 650052 95140 650058 95192
rect 616506 95004 616512 95056
rect 616564 95044 616570 95056
rect 623222 95044 623228 95056
rect 616564 95016 623228 95044
rect 616564 95004 616570 95016
rect 623222 95004 623228 95016
rect 623280 95004 623286 95056
rect 648246 94732 648252 94784
rect 648304 94772 648310 94784
rect 654778 94772 654784 94784
rect 648304 94744 654784 94772
rect 648304 94732 648310 94744
rect 654778 94732 654784 94744
rect 654836 94732 654842 94784
rect 596818 94528 596824 94580
rect 596876 94568 596882 94580
rect 598934 94568 598940 94580
rect 596876 94540 598940 94568
rect 596876 94528 596882 94540
rect 598934 94528 598940 94540
rect 598992 94528 598998 94580
rect 607674 94460 607680 94512
rect 607732 94500 607738 94512
rect 620922 94500 620928 94512
rect 607732 94472 620928 94500
rect 607732 94460 607738 94472
rect 620922 94460 620928 94472
rect 620980 94460 620986 94512
rect 619542 93780 619548 93832
rect 619600 93820 619606 93832
rect 626442 93820 626448 93832
rect 619600 93792 626448 93820
rect 619600 93780 619606 93792
rect 626442 93780 626448 93792
rect 626500 93780 626506 93832
rect 651282 93508 651288 93560
rect 651340 93548 651346 93560
rect 655422 93548 655428 93560
rect 651340 93520 655428 93548
rect 651340 93508 651346 93520
rect 655422 93508 655428 93520
rect 655480 93508 655486 93560
rect 579338 93100 579344 93152
rect 579396 93140 579402 93152
rect 585778 93140 585784 93152
rect 579396 93112 585784 93140
rect 579396 93100 579402 93112
rect 585778 93100 585784 93112
rect 585836 93100 585842 93152
rect 611170 93100 611176 93152
rect 611228 93140 611234 93152
rect 622394 93140 622400 93152
rect 611228 93112 622400 93140
rect 611228 93100 611234 93112
rect 622394 93100 622400 93112
rect 622452 93100 622458 93152
rect 617978 92420 617984 92472
rect 618036 92460 618042 92472
rect 626442 92460 626448 92472
rect 618036 92432 626448 92460
rect 618036 92420 618042 92432
rect 626442 92420 626448 92432
rect 626500 92420 626506 92472
rect 578234 91808 578240 91860
rect 578292 91848 578298 91860
rect 585962 91848 585968 91860
rect 578292 91820 585968 91848
rect 578292 91808 578298 91820
rect 585962 91808 585968 91820
rect 586020 91808 586026 91860
rect 606938 91740 606944 91792
rect 606996 91780 607002 91792
rect 626258 91780 626264 91792
rect 606996 91752 626264 91780
rect 606996 91740 607002 91752
rect 626258 91740 626264 91752
rect 626316 91740 626322 91792
rect 647234 91672 647240 91724
rect 647292 91712 647298 91724
rect 654686 91712 654692 91724
rect 647292 91684 654692 91712
rect 647292 91672 647298 91684
rect 654686 91672 654692 91684
rect 654744 91672 654750 91724
rect 610986 90992 610992 91044
rect 611044 91032 611050 91044
rect 617518 91032 617524 91044
rect 611044 91004 617524 91032
rect 611044 90992 611050 91004
rect 617518 90992 617524 91004
rect 617576 90992 617582 91044
rect 618162 90992 618168 91044
rect 618220 91032 618226 91044
rect 626442 91032 626448 91044
rect 618220 91004 626448 91032
rect 618220 90992 618226 91004
rect 626442 90992 626448 91004
rect 626500 90992 626506 91044
rect 649258 90652 649264 90704
rect 649316 90692 649322 90704
rect 655422 90692 655428 90704
rect 649316 90664 655428 90692
rect 649316 90652 649322 90664
rect 655422 90652 655428 90664
rect 655480 90652 655486 90704
rect 584582 90312 584588 90364
rect 584640 90352 584646 90364
rect 590102 90352 590108 90364
rect 584640 90324 590108 90352
rect 584640 90312 584646 90324
rect 590102 90312 590108 90324
rect 590160 90312 590166 90364
rect 620922 89632 620928 89684
rect 620980 89672 620986 89684
rect 625430 89672 625436 89684
rect 620980 89644 625436 89672
rect 620980 89632 620986 89644
rect 625430 89632 625436 89644
rect 625488 89632 625494 89684
rect 623222 89496 623228 89548
rect 623280 89536 623286 89548
rect 626442 89536 626448 89548
rect 623280 89508 626448 89536
rect 623280 89496 623286 89508
rect 626442 89496 626448 89508
rect 626500 89496 626506 89548
rect 649718 88748 649724 88800
rect 649776 88788 649782 88800
rect 658550 88788 658556 88800
rect 649776 88760 658556 88788
rect 649776 88748 649782 88760
rect 658550 88748 658556 88760
rect 658608 88748 658614 88800
rect 662322 88748 662328 88800
rect 662380 88788 662386 88800
rect 663886 88788 663892 88800
rect 662380 88760 663892 88788
rect 662380 88748 662386 88760
rect 663886 88748 663892 88760
rect 663944 88748 663950 88800
rect 579338 88272 579344 88324
rect 579396 88312 579402 88324
rect 588538 88312 588544 88324
rect 579396 88284 588544 88312
rect 579396 88272 579402 88284
rect 588538 88272 588544 88284
rect 588596 88272 588602 88324
rect 617518 88272 617524 88324
rect 617576 88312 617582 88324
rect 626442 88312 626448 88324
rect 617576 88284 626448 88312
rect 617576 88272 617582 88284
rect 626442 88272 626448 88284
rect 626500 88272 626506 88324
rect 655238 88272 655244 88324
rect 655296 88312 655302 88324
rect 658458 88312 658464 88324
rect 655296 88284 658464 88312
rect 655296 88272 655302 88284
rect 658458 88272 658464 88284
rect 658516 88272 658522 88324
rect 659562 86912 659568 86964
rect 659620 86952 659626 86964
rect 663242 86952 663248 86964
rect 659620 86924 663248 86952
rect 659620 86912 659626 86924
rect 663242 86912 663248 86924
rect 663300 86912 663306 86964
rect 653398 86844 653404 86896
rect 653456 86884 653462 86896
rect 657170 86884 657176 86896
rect 653456 86856 657176 86884
rect 653456 86844 653462 86856
rect 657170 86844 657176 86856
rect 657228 86844 657234 86896
rect 647878 86708 647884 86760
rect 647936 86748 647942 86760
rect 661402 86748 661408 86760
rect 647936 86720 661408 86748
rect 647936 86708 647942 86720
rect 661402 86708 661408 86720
rect 661460 86708 661466 86760
rect 656158 86572 656164 86624
rect 656216 86612 656222 86624
rect 660666 86612 660672 86624
rect 656216 86584 660672 86612
rect 656216 86572 656222 86584
rect 660666 86572 660672 86584
rect 660724 86572 660730 86624
rect 578786 86436 578792 86488
rect 578844 86476 578850 86488
rect 580626 86476 580632 86488
rect 578844 86448 580632 86476
rect 578844 86436 578850 86448
rect 580626 86436 580632 86448
rect 580684 86436 580690 86488
rect 652202 86436 652208 86488
rect 652260 86476 652266 86488
rect 660114 86476 660120 86488
rect 652260 86448 660120 86476
rect 652260 86436 652266 86448
rect 660114 86436 660120 86448
rect 660172 86436 660178 86488
rect 622394 86300 622400 86352
rect 622452 86340 622458 86352
rect 626442 86340 626448 86352
rect 622452 86312 626448 86340
rect 622452 86300 622458 86312
rect 626442 86300 626448 86312
rect 626500 86300 626506 86352
rect 654870 86300 654876 86352
rect 654928 86340 654934 86352
rect 662506 86340 662512 86352
rect 654928 86312 662512 86340
rect 654928 86300 654934 86312
rect 662506 86300 662512 86312
rect 662564 86300 662570 86352
rect 652018 86164 652024 86216
rect 652076 86204 652082 86216
rect 657722 86204 657728 86216
rect 652076 86176 657728 86204
rect 652076 86164 652082 86176
rect 657722 86164 657728 86176
rect 657780 86164 657786 86216
rect 609882 85484 609888 85536
rect 609940 85524 609946 85536
rect 626442 85524 626448 85536
rect 609940 85496 626448 85524
rect 609940 85484 609946 85496
rect 626442 85484 626448 85496
rect 626500 85484 626506 85536
rect 621658 85348 621664 85400
rect 621716 85388 621722 85400
rect 625246 85388 625252 85400
rect 621716 85360 625252 85388
rect 621716 85348 621722 85360
rect 625246 85348 625252 85360
rect 625304 85348 625310 85400
rect 608502 84124 608508 84176
rect 608560 84164 608566 84176
rect 625798 84164 625804 84176
rect 608560 84136 625804 84164
rect 608560 84124 608566 84136
rect 625798 84124 625804 84136
rect 625856 84124 625862 84176
rect 579338 83988 579344 84040
rect 579396 84028 579402 84040
rect 581822 84028 581828 84040
rect 579396 84000 581828 84028
rect 579396 83988 579402 84000
rect 581822 83988 581828 84000
rect 581880 83988 581886 84040
rect 581638 83444 581644 83496
rect 581696 83484 581702 83496
rect 589918 83484 589924 83496
rect 581696 83456 589924 83484
rect 581696 83444 581702 83456
rect 589918 83444 589924 83456
rect 589976 83444 589982 83496
rect 578694 82764 578700 82816
rect 578752 82804 578758 82816
rect 583202 82804 583208 82816
rect 578752 82776 583208 82804
rect 578752 82764 578758 82776
rect 583202 82764 583208 82776
rect 583260 82764 583266 82816
rect 578878 82084 578884 82136
rect 578936 82124 578942 82136
rect 587158 82124 587164 82136
rect 578936 82096 587164 82124
rect 578936 82084 578942 82096
rect 587158 82084 587164 82096
rect 587216 82084 587222 82136
rect 628742 80928 628748 80980
rect 628800 80968 628806 80980
rect 642450 80968 642456 80980
rect 628800 80940 642456 80968
rect 628800 80928 628806 80940
rect 642450 80928 642456 80940
rect 642508 80928 642514 80980
rect 618898 80792 618904 80844
rect 618956 80832 618962 80844
rect 648982 80832 648988 80844
rect 618956 80804 648988 80832
rect 618956 80792 618962 80804
rect 648982 80792 648988 80804
rect 649040 80792 649046 80844
rect 595438 80656 595444 80708
rect 595496 80696 595502 80708
rect 636746 80696 636752 80708
rect 595496 80668 636752 80696
rect 595496 80656 595502 80668
rect 636746 80656 636752 80668
rect 636804 80656 636810 80708
rect 629202 79976 629208 80028
rect 629260 80016 629266 80028
rect 633434 80016 633440 80028
rect 629260 79988 633440 80016
rect 629260 79976 629266 79988
rect 633434 79976 633440 79988
rect 633492 79976 633498 80028
rect 614022 79432 614028 79484
rect 614080 79472 614086 79484
rect 646038 79472 646044 79484
rect 614080 79444 646044 79472
rect 614080 79432 614086 79444
rect 646038 79432 646044 79444
rect 646096 79432 646102 79484
rect 588538 79296 588544 79348
rect 588596 79336 588602 79348
rect 592862 79336 592868 79348
rect 588596 79308 592868 79336
rect 588596 79296 588602 79308
rect 592862 79296 592868 79308
rect 592920 79296 592926 79348
rect 612642 79296 612648 79348
rect 612700 79336 612706 79348
rect 646314 79336 646320 79348
rect 612700 79308 646320 79336
rect 612700 79296 612706 79308
rect 646314 79296 646320 79308
rect 646372 79296 646378 79348
rect 578602 78208 578608 78260
rect 578660 78248 578666 78260
rect 580258 78248 580264 78260
rect 578660 78220 580264 78248
rect 578660 78208 578666 78220
rect 580258 78208 580264 78220
rect 580316 78208 580322 78260
rect 633434 78208 633440 78260
rect 633492 78248 633498 78260
rect 645302 78248 645308 78260
rect 633492 78220 645308 78248
rect 633492 78208 633498 78220
rect 645302 78208 645308 78220
rect 645360 78208 645366 78260
rect 631042 78072 631048 78124
rect 631100 78112 631106 78124
rect 643094 78112 643100 78124
rect 631100 78084 643100 78112
rect 631100 78072 631106 78084
rect 643094 78072 643100 78084
rect 643152 78072 643158 78124
rect 615034 77936 615040 77988
rect 615092 77976 615098 77988
rect 649166 77976 649172 77988
rect 615092 77948 649172 77976
rect 615092 77936 615098 77948
rect 649166 77936 649172 77948
rect 649224 77936 649230 77988
rect 631042 77432 631048 77444
rect 625126 77404 631048 77432
rect 622026 77256 622032 77308
rect 622084 77296 622090 77308
rect 625126 77296 625154 77404
rect 631042 77392 631048 77404
rect 631100 77392 631106 77444
rect 622084 77268 625154 77296
rect 622084 77256 622090 77268
rect 628466 77256 628472 77308
rect 628524 77296 628530 77308
rect 632790 77296 632796 77308
rect 628524 77268 632796 77296
rect 628524 77256 628530 77268
rect 632790 77256 632796 77268
rect 632848 77256 632854 77308
rect 578694 77188 578700 77240
rect 578752 77228 578758 77240
rect 584582 77228 584588 77240
rect 578752 77200 584588 77228
rect 578752 77188 578758 77200
rect 584582 77188 584588 77200
rect 584640 77188 584646 77240
rect 616138 76644 616144 76696
rect 616196 76684 616202 76696
rect 646866 76684 646872 76696
rect 616196 76656 646872 76684
rect 616196 76644 616202 76656
rect 646866 76644 646872 76656
rect 646924 76644 646930 76696
rect 579062 76508 579068 76560
rect 579120 76548 579126 76560
rect 666554 76548 666560 76560
rect 579120 76520 666560 76548
rect 579120 76508 579126 76520
rect 666554 76508 666560 76520
rect 666612 76508 666618 76560
rect 621658 75896 621664 75948
rect 621716 75936 621722 75948
rect 628466 75936 628472 75948
rect 621716 75908 628472 75936
rect 621716 75896 621722 75908
rect 628466 75896 628472 75908
rect 628524 75896 628530 75948
rect 618898 75624 618904 75676
rect 618956 75664 618962 75676
rect 622026 75664 622032 75676
rect 618956 75636 622032 75664
rect 618956 75624 618962 75636
rect 622026 75624 622032 75636
rect 622084 75624 622090 75676
rect 620278 75420 620284 75472
rect 620336 75460 620342 75472
rect 648798 75460 648804 75472
rect 620336 75432 648804 75460
rect 620336 75420 620342 75432
rect 648798 75420 648804 75432
rect 648856 75420 648862 75472
rect 607122 75284 607128 75336
rect 607180 75324 607186 75336
rect 646498 75324 646504 75336
rect 607180 75296 646504 75324
rect 607180 75284 607186 75296
rect 646498 75284 646504 75296
rect 646556 75284 646562 75336
rect 613378 75148 613384 75200
rect 613436 75188 613442 75200
rect 662598 75188 662604 75200
rect 613436 75160 662604 75188
rect 613436 75148 613442 75160
rect 662598 75148 662604 75160
rect 662656 75148 662662 75200
rect 579522 73108 579528 73160
rect 579580 73148 579586 73160
rect 584398 73148 584404 73160
rect 579580 73120 584404 73148
rect 579580 73108 579586 73120
rect 584398 73108 584404 73120
rect 584456 73108 584462 73160
rect 579246 71476 579252 71528
rect 579304 71516 579310 71528
rect 581638 71516 581644 71528
rect 579304 71488 581644 71516
rect 579304 71476 579310 71488
rect 581638 71476 581644 71488
rect 581696 71476 581702 71528
rect 579522 66240 579528 66292
rect 579580 66280 579586 66292
rect 623038 66280 623044 66292
rect 579580 66252 623044 66280
rect 579580 66240 579586 66252
rect 623038 66240 623044 66252
rect 623096 66240 623102 66292
rect 578510 62024 578516 62076
rect 578568 62064 578574 62076
rect 611998 62064 612004 62076
rect 578568 62036 612004 62064
rect 578568 62024 578574 62036
rect 611998 62024 612004 62036
rect 612056 62024 612062 62076
rect 579522 60664 579528 60716
rect 579580 60704 579586 60716
rect 624418 60704 624424 60716
rect 579580 60676 624424 60704
rect 579580 60664 579586 60676
rect 624418 60664 624424 60676
rect 624476 60664 624482 60716
rect 579522 57876 579528 57928
rect 579580 57916 579586 57928
rect 614850 57916 614856 57928
rect 579580 57888 614856 57916
rect 579580 57876 579586 57888
rect 614850 57876 614856 57888
rect 614908 57876 614914 57928
rect 579522 56516 579528 56568
rect 579580 56556 579586 56568
rect 621658 56556 621664 56568
rect 579580 56528 621664 56556
rect 579580 56516 579586 56528
rect 621658 56516 621664 56528
rect 621716 56516 621722 56568
rect 576118 53048 576124 53100
rect 576176 53088 576182 53100
rect 617518 53088 617524 53100
rect 576176 53060 617524 53088
rect 576176 53048 576182 53060
rect 617518 53048 617524 53060
rect 617576 53048 617582 53100
rect 464982 52776 464988 52828
rect 465040 52816 465046 52828
rect 467006 52816 467012 52828
rect 465040 52788 467012 52816
rect 465040 52776 465046 52788
rect 467006 52776 467012 52788
rect 467064 52776 467070 52828
rect 463602 52640 463608 52692
rect 463660 52680 463666 52692
rect 466822 52680 466828 52692
rect 463660 52652 466828 52680
rect 463660 52640 463666 52652
rect 466822 52640 466828 52652
rect 466880 52640 466886 52692
rect 464062 52504 464068 52556
rect 464120 52544 464126 52556
rect 466454 52544 466460 52556
rect 464120 52516 466460 52544
rect 464120 52504 464126 52516
rect 466454 52504 466460 52516
rect 466512 52504 466518 52556
rect 459462 52368 459468 52420
rect 459520 52408 459526 52420
rect 464982 52408 464988 52420
rect 459520 52380 464988 52408
rect 459520 52368 459526 52380
rect 464982 52368 464988 52380
rect 465040 52368 465046 52420
rect 465442 52368 465448 52420
rect 465500 52408 465506 52420
rect 475378 52408 475384 52420
rect 465500 52380 475384 52408
rect 465500 52368 465506 52380
rect 475378 52368 475384 52380
rect 475436 52368 475442 52420
rect 475562 52368 475568 52420
rect 475620 52408 475626 52420
rect 577682 52408 577688 52420
rect 475620 52380 577688 52408
rect 475620 52368 475626 52380
rect 577682 52368 577688 52380
rect 577740 52368 577746 52420
rect 457714 52232 457720 52284
rect 457772 52272 457778 52284
rect 459738 52272 459744 52284
rect 457772 52244 459744 52272
rect 457772 52232 457778 52244
rect 459738 52232 459744 52244
rect 459796 52232 459802 52284
rect 462222 52232 462228 52284
rect 462280 52272 462286 52284
rect 462280 52244 465764 52272
rect 462280 52232 462286 52244
rect 457898 52096 457904 52148
rect 457956 52136 457962 52148
rect 460842 52136 460848 52148
rect 457956 52108 460848 52136
rect 457956 52096 457962 52108
rect 460842 52096 460848 52108
rect 460900 52096 460906 52148
rect 463142 52096 463148 52148
rect 463200 52136 463206 52148
rect 465736 52136 465764 52244
rect 465902 52232 465908 52284
rect 465960 52272 465966 52284
rect 465960 52244 571932 52272
rect 465960 52232 465966 52244
rect 571904 52136 571932 52244
rect 572070 52232 572076 52284
rect 572128 52272 572134 52284
rect 625798 52272 625804 52284
rect 572128 52244 625804 52272
rect 572128 52232 572134 52244
rect 625798 52232 625804 52244
rect 625856 52232 625862 52284
rect 576118 52136 576124 52148
rect 463200 52108 464844 52136
rect 465736 52108 470594 52136
rect 571904 52108 576124 52136
rect 463200 52096 463206 52108
rect 50338 51960 50344 52012
rect 50396 52000 50402 52012
rect 130378 52000 130384 52012
rect 50396 51972 130384 52000
rect 50396 51960 50402 51972
rect 130378 51960 130384 51972
rect 130436 51960 130442 52012
rect 458082 51960 458088 52012
rect 458140 52000 458146 52012
rect 460198 52000 460204 52012
rect 458140 51972 460204 52000
rect 458140 51960 458146 51972
rect 460198 51960 460204 51972
rect 460256 51960 460262 52012
rect 464522 51960 464528 52012
rect 464580 51960 464586 52012
rect 49142 51824 49148 51876
rect 49200 51864 49206 51876
rect 129366 51864 129372 51876
rect 49200 51836 129372 51864
rect 49200 51824 49206 51836
rect 129366 51824 129372 51836
rect 129424 51824 129430 51876
rect 47578 51688 47584 51740
rect 47636 51728 47642 51740
rect 128998 51728 129004 51740
rect 47636 51700 129004 51728
rect 47636 51688 47642 51700
rect 128998 51688 129004 51700
rect 129056 51688 129062 51740
rect 145374 51688 145380 51740
rect 145432 51728 145438 51740
rect 306006 51728 306012 51740
rect 145432 51700 306012 51728
rect 145432 51688 145438 51700
rect 306006 51688 306012 51700
rect 306064 51688 306070 51740
rect 464540 51592 464568 51960
rect 464816 51796 464844 52108
rect 470566 52068 470594 52108
rect 576118 52096 576124 52108
rect 576176 52096 576182 52148
rect 576302 52096 576308 52148
rect 576360 52136 576366 52148
rect 583018 52136 583024 52148
rect 576360 52108 583024 52136
rect 576360 52096 576366 52108
rect 583018 52096 583024 52108
rect 583076 52096 583082 52148
rect 571702 52068 571708 52080
rect 470566 52040 571708 52068
rect 571702 52028 571708 52040
rect 571760 52028 571766 52080
rect 464982 51960 464988 52012
rect 465040 52000 465046 52012
rect 465040 51972 470456 52000
rect 465040 51960 465046 51972
rect 470428 51932 470456 51972
rect 475194 51932 475200 51944
rect 470428 51904 475200 51932
rect 475194 51892 475200 51904
rect 475252 51892 475258 51944
rect 475378 51892 475384 51944
rect 475436 51932 475442 51944
rect 572070 51932 572076 51944
rect 475436 51904 572076 51932
rect 475436 51892 475442 51904
rect 572070 51892 572076 51904
rect 572128 51892 572134 51944
rect 600314 51796 600320 51808
rect 464816 51768 600320 51796
rect 600314 51756 600320 51768
rect 600372 51756 600378 51808
rect 592678 51592 592684 51604
rect 464540 51564 592684 51592
rect 592678 51552 592684 51564
rect 592736 51552 592742 51604
rect 466454 51416 466460 51468
rect 466512 51456 466518 51468
rect 466512 51428 470594 51456
rect 466512 51416 466518 51428
rect 470566 51320 470594 51428
rect 475194 51416 475200 51468
rect 475252 51456 475258 51468
rect 475252 51428 567194 51456
rect 475252 51416 475258 51428
rect 475562 51320 475568 51332
rect 470566 51292 475568 51320
rect 475562 51280 475568 51292
rect 475620 51280 475626 51332
rect 567166 51320 567194 51428
rect 571702 51416 571708 51468
rect 571760 51456 571766 51468
rect 578878 51456 578884 51468
rect 571760 51428 578884 51456
rect 571760 51416 571766 51428
rect 578878 51416 578884 51428
rect 578936 51416 578942 51468
rect 576302 51320 576308 51332
rect 567166 51292 576308 51320
rect 576302 51280 576308 51292
rect 576360 51280 576366 51332
rect 467006 51008 467012 51060
rect 467064 51048 467070 51060
rect 596818 51048 596824 51060
rect 467064 51020 596824 51048
rect 467064 51008 467070 51020
rect 596818 51008 596824 51020
rect 596876 51008 596882 51060
rect 466822 50872 466828 50924
rect 466880 50912 466886 50924
rect 588538 50912 588544 50924
rect 466880 50884 588544 50912
rect 466880 50872 466886 50884
rect 588538 50872 588544 50884
rect 588596 50872 588602 50924
rect 50522 50600 50528 50652
rect 50580 50640 50586 50652
rect 128446 50640 128452 50652
rect 50580 50612 128452 50640
rect 50580 50600 50586 50612
rect 128446 50600 128452 50612
rect 128504 50600 128510 50652
rect 47762 50464 47768 50516
rect 47820 50504 47826 50516
rect 131022 50504 131028 50516
rect 47820 50476 131028 50504
rect 47820 50464 47826 50476
rect 131022 50464 131028 50476
rect 131080 50464 131086 50516
rect 318334 50464 318340 50516
rect 318392 50504 318398 50516
rect 458266 50504 458272 50516
rect 318392 50476 458272 50504
rect 318392 50464 318398 50476
rect 458266 50464 458272 50476
rect 458324 50464 458330 50516
rect 46198 50328 46204 50380
rect 46256 50368 46262 50380
rect 128630 50368 128636 50380
rect 46256 50340 128636 50368
rect 46256 50328 46262 50340
rect 128630 50328 128636 50340
rect 128688 50328 128694 50380
rect 314010 50328 314016 50380
rect 314068 50368 314074 50380
rect 458450 50368 458456 50380
rect 314068 50340 458456 50368
rect 314068 50328 314074 50340
rect 458450 50328 458456 50340
rect 458508 50328 458514 50380
rect 521102 50328 521108 50380
rect 521160 50368 521166 50380
rect 544010 50368 544016 50380
rect 521160 50340 544016 50368
rect 521160 50328 521166 50340
rect 544010 50328 544016 50340
rect 544068 50328 544074 50380
rect 467006 49376 467012 49428
rect 467064 49416 467070 49428
rect 577498 49416 577504 49428
rect 467064 49388 577504 49416
rect 467064 49376 467070 49388
rect 577498 49376 577504 49388
rect 577556 49376 577562 49428
rect 48958 49240 48964 49292
rect 49016 49280 49022 49292
rect 129550 49280 129556 49292
rect 49016 49252 129556 49280
rect 49016 49240 49022 49252
rect 129550 49240 129556 49252
rect 129608 49240 129614 49292
rect 466638 49240 466644 49292
rect 466696 49280 466702 49292
rect 599118 49280 599124 49292
rect 466696 49252 599124 49280
rect 466696 49240 466702 49252
rect 599118 49240 599124 49252
rect 599176 49240 599182 49292
rect 45462 49104 45468 49156
rect 45520 49144 45526 49156
rect 128814 49144 128820 49156
rect 45520 49116 128820 49144
rect 45520 49104 45526 49116
rect 128814 49104 128820 49116
rect 128872 49104 128878 49156
rect 466454 49104 466460 49156
rect 466512 49144 466518 49156
rect 601694 49144 601700 49156
rect 466512 49116 601700 49144
rect 466512 49104 466518 49116
rect 601694 49104 601700 49116
rect 601752 49104 601758 49156
rect 46382 48968 46388 49020
rect 46440 49008 46446 49020
rect 130470 49008 130476 49020
rect 46440 48980 130476 49008
rect 46440 48968 46446 48980
rect 130470 48968 130476 48980
rect 130528 48968 130534 49020
rect 466822 48968 466828 49020
rect 466880 49008 466886 49020
rect 618898 49008 618904 49020
rect 466880 48980 618904 49008
rect 466880 48968 466886 48980
rect 618898 48968 618904 48980
rect 618956 48968 618962 49020
rect 128446 48084 128452 48136
rect 128504 48124 128510 48136
rect 131942 48124 131948 48136
rect 128504 48096 131948 48124
rect 128504 48084 128510 48096
rect 131942 48084 131948 48096
rect 132000 48084 132006 48136
rect 128630 47812 128636 47864
rect 128688 47852 128694 47864
rect 131758 47852 131764 47864
rect 128688 47824 131764 47852
rect 128688 47812 128694 47824
rect 131758 47812 131764 47824
rect 131816 47812 131822 47864
rect 623038 46452 623044 46504
rect 623096 46492 623102 46504
rect 661586 46492 661592 46504
rect 623096 46464 661592 46492
rect 623096 46452 623102 46464
rect 661586 46452 661592 46464
rect 661644 46452 661650 46504
rect 129550 45024 129556 45076
rect 129608 45064 129614 45076
rect 129608 45036 131160 45064
rect 129608 45024 129614 45036
rect 131224 44964 131376 44992
rect 128998 44888 129004 44940
rect 129056 44928 129062 44940
rect 131224 44928 131252 44964
rect 129056 44900 131252 44928
rect 129056 44888 129062 44900
rect 129182 44752 129188 44804
rect 129240 44792 129246 44804
rect 131546 44792 131574 44894
rect 129240 44764 131574 44792
rect 131638 44796 131790 44824
rect 129240 44752 129246 44764
rect 129366 44616 129372 44668
rect 129424 44656 129430 44668
rect 131638 44656 131666 44796
rect 131758 44684 131764 44736
rect 131816 44724 131822 44736
rect 131960 44724 131988 44726
rect 131816 44696 131988 44724
rect 131816 44684 131822 44696
rect 129424 44628 131666 44656
rect 132052 44628 132158 44656
rect 129424 44616 129430 44628
rect 132052 44588 132080 44628
rect 131960 44584 132080 44588
rect 131942 44532 131948 44584
rect 132000 44560 132080 44584
rect 132000 44532 132006 44560
rect 132328 44316 132356 44558
rect 132604 44328 132632 44474
rect 132052 44288 132356 44316
rect 132052 44264 132080 44288
rect 132586 44276 132592 44328
rect 132644 44276 132650 44328
rect 128814 44208 128820 44260
rect 128872 44248 128878 44260
rect 131960 44248 132080 44264
rect 128872 44236 132080 44248
rect 128872 44220 131988 44236
rect 128872 44208 128878 44220
rect 132788 44180 132816 44362
rect 132052 44152 132816 44180
rect 130654 44072 130660 44124
rect 130712 44112 130718 44124
rect 132052 44112 132080 44152
rect 130712 44084 132080 44112
rect 130712 44072 130718 44084
rect 131022 43936 131028 43988
rect 131080 43976 131086 43988
rect 132972 43976 133000 44250
rect 131080 43948 133000 43976
rect 131080 43936 131086 43948
rect 43622 42780 43628 42832
rect 43680 42820 43686 42832
rect 133156 42820 133184 44138
rect 431218 43636 431224 43648
rect 412606 43608 431224 43636
rect 187326 43528 187332 43580
rect 187384 43568 187390 43580
rect 412606 43568 412634 43608
rect 431218 43596 431224 43608
rect 431276 43596 431282 43648
rect 439590 43596 439596 43648
rect 439648 43636 439654 43648
rect 441614 43636 441620 43648
rect 439648 43608 441620 43636
rect 439648 43596 439654 43608
rect 441614 43596 441620 43608
rect 441672 43596 441678 43648
rect 187384 43540 412634 43568
rect 187384 43528 187390 43540
rect 43680 42792 133184 42820
rect 43680 42780 43686 42792
rect 310422 42712 310428 42764
rect 310480 42752 310486 42764
rect 431218 42752 431224 42764
rect 310480 42724 431224 42752
rect 310480 42712 310486 42724
rect 431218 42712 431224 42724
rect 431276 42712 431282 42764
rect 456058 42712 456064 42764
rect 456116 42752 456122 42764
rect 463050 42752 463056 42764
rect 456116 42724 463056 42752
rect 456116 42712 456122 42724
rect 463050 42712 463056 42724
rect 463108 42712 463114 42764
rect 404446 42304 404452 42356
rect 404504 42344 404510 42356
rect 405550 42344 405556 42356
rect 404504 42316 405556 42344
rect 404504 42304 404510 42316
rect 405550 42304 405556 42316
rect 405608 42304 405614 42356
rect 420730 42304 420736 42356
rect 420788 42344 420794 42356
rect 427078 42344 427084 42356
rect 420788 42316 427084 42344
rect 420788 42304 420794 42316
rect 427078 42304 427084 42316
rect 427136 42304 427142 42356
rect 662414 42173 662420 42225
rect 662472 42173 662478 42225
rect 431218 42032 431224 42084
rect 431276 42072 431282 42084
rect 456058 42072 456064 42084
rect 431276 42044 456064 42072
rect 431276 42032 431282 42044
rect 456058 42032 456064 42044
rect 456116 42032 456122 42084
rect 404446 41420 404452 41472
rect 404504 41460 404510 41472
rect 420730 41460 420736 41472
rect 404504 41432 420736 41460
rect 404504 41420 404510 41432
rect 420730 41420 420736 41432
rect 420788 41420 420794 41472
rect 427078 41420 427084 41472
rect 427136 41460 427142 41472
rect 459186 41460 459192 41472
rect 427136 41432 459192 41460
rect 427136 41420 427142 41432
rect 459186 41420 459192 41432
rect 459244 41420 459250 41472
<< via1 >>
rect 366180 1027828 366232 1027880
rect 366548 1027828 366600 1027880
rect 366180 1024360 366232 1024412
rect 366548 1024360 366600 1024412
rect 200028 1007360 200080 1007412
rect 202696 1007360 202748 1007412
rect 505376 1007088 505428 1007140
rect 513840 1007088 513892 1007140
rect 428004 1006884 428056 1006936
rect 357716 1006816 357768 1006868
rect 369860 1006816 369912 1006868
rect 430856 1006748 430908 1006800
rect 434628 1006748 434680 1006800
rect 360200 1006680 360252 1006732
rect 373264 1006680 373316 1006732
rect 145748 1006544 145800 1006596
rect 153752 1006544 153804 1006596
rect 430028 1006476 430080 1006528
rect 433984 1006476 434036 1006528
rect 93308 1006408 93360 1006460
rect 102324 1006408 102376 1006460
rect 145564 1006408 145616 1006460
rect 152096 1006408 152148 1006460
rect 157432 1006408 157484 1006460
rect 166264 1006408 166316 1006460
rect 93124 1006000 93176 1006052
rect 101956 1006272 102008 1006324
rect 144184 1006272 144236 1006324
rect 151728 1006272 151780 1006324
rect 158260 1006272 158312 1006324
rect 171784 1006408 171836 1006460
rect 206192 1006408 206244 1006460
rect 210056 1006408 210108 1006460
rect 300308 1006408 300360 1006460
rect 306932 1006408 306984 1006460
rect 505376 1006884 505428 1006936
rect 518164 1006884 518216 1006936
rect 554780 1006884 554832 1006936
rect 569224 1006884 569276 1006936
rect 506204 1006748 506256 1006800
rect 555976 1006748 556028 1006800
rect 565820 1006748 565872 1006800
rect 520924 1006680 520976 1006732
rect 447784 1006408 447836 1006460
rect 508228 1006408 508280 1006460
rect 210424 1006272 210476 1006324
rect 228364 1006272 228416 1006324
rect 249248 1006272 249300 1006324
rect 256148 1006272 256200 1006324
rect 298928 1006272 298980 1006324
rect 311808 1006272 311860 1006324
rect 361396 1006272 361448 1006324
rect 375012 1006272 375064 1006324
rect 402244 1006272 402296 1006324
rect 429200 1006272 429252 1006324
rect 434628 1006272 434680 1006324
rect 469864 1006272 469916 1006324
rect 556988 1006408 557040 1006460
rect 559656 1006408 559708 1006460
rect 522304 1006272 522356 1006324
rect 431684 1006204 431736 1006256
rect 101404 1006136 101456 1006188
rect 103980 1006136 104032 1006188
rect 107660 1006136 107712 1006188
rect 124864 1006136 124916 1006188
rect 144736 1006136 144788 1006188
rect 150900 1006136 150952 1006188
rect 160284 1006136 160336 1006188
rect 164884 1006136 164936 1006188
rect 166264 1006136 166316 1006188
rect 175924 1006136 175976 1006188
rect 208400 1006136 208452 1006188
rect 94504 1006000 94556 1006052
rect 98276 1006000 98328 1006052
rect 102784 1006000 102836 1006052
rect 104808 1006000 104860 1006052
rect 108488 1006000 108540 1006052
rect 126244 1006000 126296 1006052
rect 147588 1006000 147640 1006052
rect 150072 1006000 150124 1006052
rect 159456 1006000 159508 1006052
rect 177304 1006000 177356 1006052
rect 196808 1006000 196860 1006052
rect 201040 1006000 201092 1006052
rect 209228 1006000 209280 1006052
rect 211804 1006000 211856 1006052
rect 249064 1006136 249116 1006188
rect 255320 1006136 255372 1006188
rect 261852 1006136 261904 1006188
rect 279424 1006136 279476 1006188
rect 300124 1006136 300176 1006188
rect 306104 1006136 306156 1006188
rect 357348 1006136 357400 1006188
rect 362224 1006136 362276 1006188
rect 229744 1006000 229796 1006052
rect 247040 1006000 247092 1006052
rect 252468 1006000 252520 1006052
rect 260196 1006000 260248 1006052
rect 280804 1006000 280856 1006052
rect 298744 1006000 298796 1006052
rect 303252 1006000 303304 1006052
rect 304080 1006000 304132 1006052
rect 314660 1006000 314712 1006052
rect 319444 1006000 319496 1006052
rect 356888 1006000 356940 1006052
rect 360844 1006000 360896 1006052
rect 363420 1006000 363472 1006052
rect 382924 1006000 382976 1006052
rect 400864 1006000 400916 1006052
rect 431500 1006136 431552 1006188
rect 428372 1006000 428424 1006052
rect 438124 1006000 438176 1006052
rect 507032 1006136 507084 1006188
rect 471244 1006000 471296 1006052
rect 496728 1006000 496780 1006052
rect 498844 1006000 498896 1006052
rect 502524 1006000 502576 1006052
rect 505744 1006000 505796 1006052
rect 509056 1006000 509108 1006052
rect 556804 1006136 556856 1006188
rect 567844 1006136 567896 1006188
rect 523684 1006000 523736 1006052
rect 555148 1006000 555200 1006052
rect 556436 1006000 556488 1006052
rect 557172 1006000 557224 1006052
rect 571984 1006000 572036 1006052
rect 514024 1005932 514076 1005984
rect 304080 1005796 304132 1005848
rect 425520 1005660 425572 1005712
rect 452568 1005660 452620 1005712
rect 505008 1005660 505060 1005712
rect 515404 1005660 515456 1005712
rect 360568 1005524 360620 1005576
rect 378784 1005524 378836 1005576
rect 427176 1005524 427228 1005576
rect 458824 1005524 458876 1005576
rect 556436 1005524 556488 1005576
rect 573364 1005524 573416 1005576
rect 358544 1005388 358596 1005440
rect 371884 1005388 371936 1005440
rect 428372 1005388 428424 1005440
rect 465724 1005388 465776 1005440
rect 502156 1005388 502208 1005440
rect 519544 1005388 519596 1005440
rect 553124 1005388 553176 1005440
rect 570604 1005388 570656 1005440
rect 149704 1005320 149756 1005372
rect 152924 1005320 152976 1005372
rect 357716 1005252 357768 1005304
rect 376760 1005252 376812 1005304
rect 423496 1005252 423548 1005304
rect 467104 1005252 467156 1005304
rect 499672 1005252 499724 1005304
rect 516784 1005252 516836 1005304
rect 551468 1005252 551520 1005304
rect 574744 1005252 574796 1005304
rect 208400 1005116 208452 1005168
rect 209872 1005116 209924 1005168
rect 149888 1005048 149940 1005100
rect 152924 1005048 152976 1005100
rect 500500 1005048 500552 1005100
rect 508504 1005048 508556 1005100
rect 207572 1004980 207624 1005032
rect 210056 1004980 210108 1005032
rect 151084 1004912 151136 1004964
rect 153752 1004912 153804 1004964
rect 158628 1004912 158680 1004964
rect 162124 1004912 162176 1004964
rect 263048 1004912 263100 1004964
rect 268384 1004912 268436 1004964
rect 313832 1004912 313884 1004964
rect 316040 1004912 316092 1004964
rect 361396 1004912 361448 1004964
rect 364892 1004912 364944 1004964
rect 431224 1004912 431276 1004964
rect 433524 1004912 433576 1004964
rect 160652 1004776 160704 1004828
rect 163136 1004776 163188 1004828
rect 209228 1004776 209280 1004828
rect 211160 1004776 211212 1004828
rect 314660 1004776 314712 1004828
rect 316684 1004776 316736 1004828
rect 353208 1004776 353260 1004828
rect 355692 1004776 355744 1004828
rect 362592 1004776 362644 1004828
rect 365260 1004776 365312 1004828
rect 420644 1004776 420696 1004828
rect 422668 1004776 422720 1004828
rect 432052 1004776 432104 1004828
rect 435548 1004776 435600 1004828
rect 498108 1004776 498160 1004828
rect 500500 1004776 500552 1004828
rect 507860 1004776 507912 1004828
rect 509700 1004776 509752 1004828
rect 555976 1004776 556028 1004828
rect 558184 1004776 558236 1004828
rect 151268 1004640 151320 1004692
rect 154120 1004640 154172 1004692
rect 161112 1004640 161164 1004692
rect 162952 1004640 163004 1004692
rect 212540 1004640 212592 1004692
rect 217324 1004640 217376 1004692
rect 315488 1004640 315540 1004692
rect 318064 1004640 318116 1004692
rect 354404 1004640 354456 1004692
rect 356520 1004640 356572 1004692
rect 364248 1004640 364300 1004692
rect 366364 1004640 366416 1004692
rect 430028 1004640 430080 1004692
rect 431960 1004640 432012 1004692
rect 499488 1004640 499540 1004692
rect 501328 1004640 501380 1004692
rect 507400 1004640 507452 1004692
rect 509240 1004640 509292 1004692
rect 557632 1004640 557684 1004692
rect 559564 1004640 559616 1004692
rect 560852 1004640 560904 1004692
rect 566464 1004640 566516 1004692
rect 424692 1004028 424744 1004080
rect 446036 1004028 446088 1004080
rect 551100 1004028 551152 1004080
rect 564440 1004028 564492 1004080
rect 360568 1003892 360620 1003944
rect 375380 1003892 375432 1003944
rect 426348 1003892 426400 1003944
rect 449900 1003892 449952 1003944
rect 452568 1003892 452620 1003944
rect 460940 1003892 460992 1003944
rect 504548 1003892 504600 1003944
rect 520280 1003892 520332 1003944
rect 552296 1003892 552348 1003944
rect 567384 1003892 567436 1003944
rect 565820 1003620 565872 1003672
rect 568580 1003620 568632 1003672
rect 513840 1003348 513892 1003400
rect 518900 1003348 518952 1003400
rect 355692 1003280 355744 1003332
rect 363604 1003280 363656 1003332
rect 375012 1003212 375064 1003264
rect 379428 1003212 379480 1003264
rect 421840 1002668 421892 1002720
rect 462964 1002668 463016 1002720
rect 97448 1002600 97500 1002652
rect 100300 1002600 100352 1002652
rect 106832 1002600 106884 1002652
rect 109500 1002600 109552 1002652
rect 253204 1002600 253256 1002652
rect 256148 1002600 256200 1002652
rect 558828 1002600 558880 1002652
rect 562508 1002600 562560 1002652
rect 358544 1002532 358596 1002584
rect 371148 1002532 371200 1002584
rect 423496 1002532 423548 1002584
rect 468484 1002532 468536 1002584
rect 92664 1002464 92716 1002516
rect 99472 1002464 99524 1002516
rect 100024 1002464 100076 1002516
rect 103152 1002464 103204 1002516
rect 108028 1002464 108080 1002516
rect 110696 1002464 110748 1002516
rect 153844 1002464 153896 1002516
rect 155776 1002464 155828 1002516
rect 211252 1002464 211304 1002516
rect 215944 1002464 215996 1002516
rect 251824 1002464 251876 1002516
rect 254492 1002464 254544 1002516
rect 560852 1002464 560904 1002516
rect 565084 1002464 565136 1002516
rect 97264 1002328 97316 1002380
rect 100300 1002328 100352 1002380
rect 106004 1002328 106056 1002380
rect 108304 1002328 108356 1002380
rect 156604 1002328 156656 1002380
rect 158720 1002328 158772 1002380
rect 261024 1002328 261076 1002380
rect 264244 1002328 264296 1002380
rect 500868 1002328 500920 1002380
rect 503352 1002328 503404 1002380
rect 558000 1002328 558052 1002380
rect 560944 1002328 560996 1002380
rect 365076 1002260 365128 1002312
rect 367928 1002260 367980 1002312
rect 98828 1002192 98880 1002244
rect 101128 1002192 101180 1002244
rect 105636 1002192 105688 1002244
rect 107936 1002192 107988 1002244
rect 108856 1002192 108908 1002244
rect 112076 1002192 112128 1002244
rect 148508 1002192 148560 1002244
rect 151728 1002192 151780 1002244
rect 155776 1002192 155828 1002244
rect 157340 1002192 157392 1002244
rect 211252 1002192 211304 1002244
rect 213184 1002192 213236 1002244
rect 262680 1002192 262732 1002244
rect 265808 1002192 265860 1002244
rect 357348 1002192 357400 1002244
rect 359372 1002192 359424 1002244
rect 502248 1002192 502300 1002244
rect 504180 1002192 504232 1002244
rect 553308 1002192 553360 1002244
rect 553952 1002192 554004 1002244
rect 560484 1002192 560536 1002244
rect 563060 1002192 563112 1002244
rect 365904 1002124 365956 1002176
rect 369124 1002124 369176 1002176
rect 95884 1002056 95936 1002108
rect 99104 1002056 99156 1002108
rect 96068 1001920 96120 1001972
rect 98276 1001920 98328 1001972
rect 98644 1001920 98696 1001972
rect 101956 1002056 102008 1002108
rect 106832 1002056 106884 1002108
rect 109040 1002056 109092 1002108
rect 109684 1002056 109736 1002108
rect 111892 1002056 111944 1002108
rect 144000 1002056 144052 1002108
rect 147588 1002056 147640 1002108
rect 148324 1002056 148376 1002108
rect 150900 1002056 150952 1002108
rect 155224 1002056 155276 1002108
rect 156604 1002056 156656 1002108
rect 203524 1002056 203576 1002108
rect 206376 1002056 206428 1002108
rect 210884 1002056 210936 1002108
rect 212540 1002056 212592 1002108
rect 252008 1002056 252060 1002108
rect 254124 1002056 254176 1002108
rect 263876 1002056 263928 1002108
rect 267004 1002056 267056 1002108
rect 301504 1002056 301556 1002108
rect 304908 1002056 304960 1002108
rect 310152 1002056 310204 1002108
rect 311900 1002056 311952 1002108
rect 424508 1002056 424560 1002108
rect 425520 1002056 425572 1002108
rect 427544 1002056 427596 1002108
rect 429844 1002056 429896 1002108
rect 433340 1002056 433392 1002108
rect 435364 1002056 435416 1002108
rect 502524 1002056 502576 1002108
rect 503720 1002056 503772 1002108
rect 509884 1002056 509936 1002108
rect 512828 1002056 512880 1002108
rect 560024 1002056 560076 1002108
rect 562324 1002056 562376 1002108
rect 365076 1001988 365128 1002040
rect 367744 1001988 367796 1002040
rect 369860 1001988 369912 1002040
rect 374644 1001988 374696 1002040
rect 423588 1001988 423640 1002040
rect 424324 1001988 424376 1002040
rect 100208 1001920 100260 1001972
rect 103152 1001920 103204 1001972
rect 106004 1001920 106056 1001972
rect 107752 1001920 107804 1001972
rect 108856 1001920 108908 1001972
rect 110512 1001920 110564 1001972
rect 146944 1001920 146996 1001972
rect 149244 1001920 149296 1001972
rect 152464 1001920 152516 1001972
rect 154580 1001920 154632 1001972
rect 154948 1001920 155000 1001972
rect 155960 1001920 156012 1001972
rect 157800 1001920 157852 1001972
rect 160100 1001920 160152 1001972
rect 204168 1001920 204220 1001972
rect 205548 1001920 205600 1001972
rect 206744 1001920 206796 1001972
rect 208400 1001920 208452 1001972
rect 212080 1001920 212132 1001972
rect 213920 1001920 213972 1001972
rect 253388 1001920 253440 1001972
rect 255320 1001920 255372 1001972
rect 263508 1001920 263560 1001972
rect 265624 1001920 265676 1001972
rect 310980 1001920 311032 1001972
rect 313280 1001920 313332 1001972
rect 351828 1001920 351880 1001972
rect 354036 1001920 354088 1001972
rect 358728 1001920 358780 1001972
rect 359372 1001920 359424 1001972
rect 419448 1001920 419500 1001972
rect 421472 1001920 421524 1001972
rect 429200 1001920 429252 1001972
rect 431224 1001920 431276 1001972
rect 432880 1001920 432932 1001972
rect 436744 1001920 436796 1001972
rect 496544 1001920 496596 1001972
rect 498476 1001920 498528 1001972
rect 501696 1001920 501748 1001972
rect 502984 1001920 503036 1001972
rect 503352 1001920 503404 1001972
rect 504364 1001920 504416 1001972
rect 510344 1001920 510396 1001972
rect 512644 1001920 512696 1001972
rect 558828 1001920 558880 1001972
rect 560300 1001920 560352 1001972
rect 561680 1001920 561732 1001972
rect 563704 1001920 563756 1001972
rect 354864 1001308 354916 1001360
rect 377956 1001308 378008 1001360
rect 499488 1001308 499540 1001360
rect 516968 1001308 517020 1001360
rect 353208 1001172 353260 1001224
rect 380900 1001172 380952 1001224
rect 429844 1001172 429896 1001224
rect 447140 1001172 447192 1001224
rect 496544 1001172 496596 1001224
rect 522764 1001172 522816 1001224
rect 550272 1001172 550324 1001224
rect 574100 1001172 574152 1001224
rect 449900 1001104 449952 1001156
rect 453764 1001104 453816 1001156
rect 447784 1000764 447836 1000816
rect 449900 1000764 449952 1000816
rect 98000 1000492 98052 1000544
rect 100208 1000492 100260 1000544
rect 447140 1000016 447192 1000068
rect 450084 1000016 450136 1000068
rect 95148 999132 95200 999184
rect 98828 999132 98880 999184
rect 376760 999132 376812 999184
rect 383384 999132 383436 999184
rect 618168 999132 618220 999184
rect 625528 999132 625580 999184
rect 564440 999064 564492 999116
rect 567936 999064 567988 999116
rect 196624 998792 196676 998844
rect 203892 998792 203944 998844
rect 449900 998792 449952 998844
rect 472624 998792 472676 998844
rect 515404 998792 515456 998844
rect 517152 998792 517204 998844
rect 198004 998656 198056 998708
rect 202696 998656 202748 998708
rect 427084 998656 427136 998708
rect 472440 998656 472492 998708
rect 201040 998520 201092 998572
rect 203892 998520 203944 998572
rect 303252 998520 303304 998572
rect 308956 998520 309008 998572
rect 371884 998520 371936 998572
rect 382740 998520 382792 998572
rect 424508 998520 424560 998572
rect 472256 998520 472308 998572
rect 502248 998520 502300 998572
rect 516508 998520 516560 998572
rect 92296 998384 92348 998436
rect 98000 998384 98052 998436
rect 143724 998384 143776 998436
rect 153844 998384 153896 998436
rect 195244 998384 195296 998436
rect 204168 998384 204220 998436
rect 304264 998384 304316 998436
rect 307300 998384 307352 998436
rect 351828 998384 351880 998436
rect 382280 998384 382332 998436
rect 423588 998384 423640 998436
rect 472072 998384 472124 998436
rect 503720 998384 503772 998436
rect 524052 998384 524104 998436
rect 552296 998384 552348 998436
rect 570788 998384 570840 998436
rect 247224 998248 247276 998300
rect 199384 998112 199436 998164
rect 201868 998112 201920 998164
rect 250444 998112 250496 998164
rect 253664 998112 253716 998164
rect 195796 997976 195848 998028
rect 200672 997976 200724 998028
rect 202328 997976 202380 998028
rect 205548 997976 205600 998028
rect 250628 997908 250680 997960
rect 253664 997908 253716 997960
rect 144184 997840 144236 997892
rect 151268 997840 151320 997892
rect 195428 997840 195480 997892
rect 200028 997840 200080 997892
rect 202144 997840 202196 997892
rect 204720 997840 204772 997892
rect 246580 997840 246632 997892
rect 247040 997840 247092 997892
rect 247684 997772 247736 997824
rect 252468 997772 252520 997824
rect 259368 998248 259420 998300
rect 260932 998248 260984 998300
rect 302884 998248 302936 998300
rect 306104 998248 306156 998300
rect 258172 998112 258224 998164
rect 259460 998112 259512 998164
rect 305644 998112 305696 998164
rect 308128 998112 308180 998164
rect 254768 998044 254820 998096
rect 257344 998044 257396 998096
rect 259828 998044 259880 998096
rect 262312 998044 262364 998096
rect 304448 997976 304500 998028
rect 306932 997976 306984 998028
rect 308404 997976 308456 998028
rect 310612 997976 310664 998028
rect 549168 997976 549220 998028
rect 551468 997976 551520 998028
rect 254584 997908 254636 997960
rect 256516 997908 256568 997960
rect 260196 997908 260248 997960
rect 262496 997908 262548 997960
rect 379428 997908 379480 997960
rect 383200 997908 383252 997960
rect 303068 997840 303120 997892
rect 305276 997840 305328 997892
rect 307024 997840 307076 997892
rect 308956 997840 309008 997892
rect 551560 997840 551612 997892
rect 553124 997840 553176 997892
rect 278136 997772 278188 997824
rect 378784 997772 378836 997824
rect 383568 997772 383620 997824
rect 520280 997772 520332 997824
rect 523868 997772 523920 997824
rect 108304 997704 108356 997756
rect 116308 997704 116360 997756
rect 143816 997704 143868 997756
rect 160100 997704 160152 997756
rect 162124 997704 162176 997756
rect 170312 997704 170364 997756
rect 195612 997704 195664 997756
rect 207020 997704 207072 997756
rect 298744 997704 298796 997756
rect 311900 997704 311952 997756
rect 371148 997704 371200 997756
rect 372528 997704 372580 997756
rect 375380 997704 375432 997756
rect 378600 997704 378652 997756
rect 399944 997704 399996 997756
rect 431960 997704 432012 997756
rect 438124 997704 438176 997756
rect 439872 997704 439924 997756
rect 489000 997704 489052 997756
rect 506480 997704 506532 997756
rect 509700 997704 509752 997756
rect 517336 997704 517388 997756
rect 540888 997704 540940 997756
rect 556988 997704 557040 997756
rect 246948 997636 247000 997688
rect 258080 997636 258132 997688
rect 571984 997636 572036 997688
rect 590568 997636 590620 997688
rect 92480 997568 92532 997620
rect 100024 997568 100076 997620
rect 109500 997568 109552 997620
rect 117228 997568 117280 997620
rect 144828 997568 144880 997620
rect 158720 997568 158772 997620
rect 299388 997568 299440 997620
rect 310520 997568 310572 997620
rect 365260 997568 365312 997620
rect 372344 997568 372396 997620
rect 431224 997568 431276 997620
rect 439688 997568 439740 997620
rect 498108 997568 498160 997620
rect 516876 997568 516928 997620
rect 246764 997500 246816 997552
rect 255964 997500 256016 997552
rect 553308 997500 553360 997552
rect 625712 997772 625764 997824
rect 504364 997432 504416 997484
rect 516692 997432 516744 997484
rect 568580 997364 568632 997416
rect 590384 997364 590436 997416
rect 551560 997296 551612 997348
rect 567568 997296 567620 997348
rect 591304 997296 591356 997348
rect 618168 997296 618220 997348
rect 200212 997228 200264 997280
rect 206192 997228 206244 997280
rect 303252 997228 303304 997280
rect 304448 997228 304500 997280
rect 446036 997228 446088 997280
rect 160744 997160 160796 997212
rect 162952 997160 163004 997212
rect 362224 997160 362276 997212
rect 372712 997160 372764 997212
rect 400128 997092 400180 997144
rect 446128 997092 446180 997144
rect 106924 997024 106976 997076
rect 111892 997024 111944 997076
rect 298376 997024 298428 997076
rect 307208 997024 307260 997076
rect 357348 997024 357400 997076
rect 372344 997024 372396 997076
rect 450084 997160 450136 997212
rect 471888 997160 471940 997212
rect 553492 997160 553544 997212
rect 570144 997160 570196 997212
rect 573364 997160 573416 997212
rect 622400 997160 622452 997212
rect 469220 997024 469272 997076
rect 500868 997024 500920 997076
rect 522948 997024 523000 997076
rect 567384 997024 567436 997076
rect 620284 997024 620336 997076
rect 92480 996956 92532 997008
rect 100760 996956 100812 997008
rect 569224 996888 569276 996940
rect 590568 996888 590620 996940
rect 143816 996684 143868 996736
rect 148508 996684 148560 996736
rect 200764 996684 200816 996736
rect 202512 996684 202564 996736
rect 251640 996684 251692 996736
rect 253388 996684 253440 996736
rect 199384 996344 199436 996396
rect 195612 996208 195664 996260
rect 246948 996208 247000 996260
rect 252008 996208 252060 996260
rect 144000 996072 144052 996124
rect 143816 995936 143868 995988
rect 136456 995800 136508 995852
rect 137744 995800 137796 995852
rect 144644 995800 144696 995852
rect 171784 996072 171836 996124
rect 211160 996072 211212 996124
rect 211804 996072 211856 996124
rect 262496 996072 262548 996124
rect 265808 996072 265860 996124
rect 316040 996072 316092 996124
rect 382924 996072 382976 996124
rect 433524 996072 433576 996124
rect 522304 996072 522356 996124
rect 563060 996072 563112 996124
rect 570604 996072 570656 996124
rect 169392 995936 169444 995988
rect 171508 995936 171560 995988
rect 175924 995936 175976 995988
rect 209872 995936 209924 995988
rect 213184 995936 213236 995988
rect 261116 995936 261168 995988
rect 280804 995936 280856 995988
rect 313280 995936 313332 995988
rect 366364 995936 366416 995988
rect 400864 995936 400916 995988
rect 152464 995800 152516 995852
rect 170680 995800 170732 995852
rect 171692 995800 171744 995852
rect 177304 995800 177356 995852
rect 212540 995800 212592 995852
rect 229744 995800 229796 995852
rect 262312 995800 262364 995852
rect 264244 995800 264296 995852
rect 298928 995800 298980 995852
rect 364892 995800 364944 995852
rect 402244 995800 402296 995852
rect 453764 995800 453816 995852
rect 558184 995936 558236 995988
rect 625896 995936 625948 995988
rect 488908 995868 488960 995920
rect 523684 995800 523736 995852
rect 560300 995800 560352 995852
rect 642088 995868 642140 995920
rect 143448 995528 143500 995580
rect 144184 995528 144236 995580
rect 171048 995528 171100 995580
rect 246212 995528 246264 995580
rect 257344 995528 257396 995580
rect 382740 995528 382792 995580
rect 384948 995528 385000 995580
rect 472624 995528 472676 995580
rect 473360 995528 473412 995580
rect 496820 995528 496872 995580
rect 520188 995528 520240 995580
rect 524052 995528 524104 995580
rect 525340 995528 525392 995580
rect 386696 995460 386748 995512
rect 388628 995460 388680 995512
rect 473820 995460 473872 995512
rect 478236 995460 478288 995512
rect 529572 995460 529624 995512
rect 530216 995460 530268 995512
rect 625896 995460 625948 995512
rect 629668 995460 629720 995512
rect 415400 995392 415452 995444
rect 171692 995277 171744 995329
rect 180708 995324 180760 995376
rect 182640 995324 182692 995376
rect 193128 995324 193180 995376
rect 195060 995324 195112 995376
rect 245568 995324 245620 995376
rect 246764 995324 246816 995376
rect 378140 995256 378192 995308
rect 397644 995256 397696 995308
rect 171508 995165 171560 995217
rect 180478 995188 180530 995240
rect 184664 995188 184716 995240
rect 190368 995188 190420 995240
rect 190552 995188 190604 995240
rect 192484 995188 192536 995240
rect 194140 995188 194192 995240
rect 194324 995188 194376 995240
rect 195244 995188 195296 995240
rect 234942 995188 234994 995240
rect 253204 995188 253256 995240
rect 292488 995188 292540 995240
rect 303068 995188 303120 995240
rect 416136 995235 416188 995287
rect 360844 995120 360896 995172
rect 389640 995120 389692 995172
rect 537760 995120 537812 995172
rect 538404 995120 538456 995172
rect 172428 995052 172480 995104
rect 181444 995052 181496 995104
rect 210056 995052 210108 995104
rect 234528 995052 234580 995104
rect 259460 995052 259512 995104
rect 283472 995052 283524 995104
rect 305644 995052 305696 995104
rect 425704 995052 425756 995104
rect 484124 995052 484176 995104
rect 505744 995052 505796 995104
rect 528744 995052 528796 995104
rect 567568 995052 567620 995104
rect 637028 995052 637080 995104
rect 358728 994984 358780 995036
rect 398840 994984 398892 995036
rect 180708 994916 180760 994968
rect 208400 994916 208452 994968
rect 232872 994916 232924 994968
rect 260932 994916 260984 994968
rect 284116 994916 284168 994968
rect 308404 994916 308456 994968
rect 419448 994916 419500 994968
rect 660580 994983 660632 995035
rect 80152 994780 80204 994832
rect 103520 994780 103572 994832
rect 128452 994780 128504 994832
rect 157340 994780 157392 994832
rect 170864 994829 170916 994881
rect 171232 994829 171284 994881
rect 372712 994848 372764 994900
rect 393320 994848 393372 994900
rect 287152 994780 287204 994832
rect 304264 994780 304316 994832
rect 433984 994780 434036 994832
rect 509240 994780 509292 994832
rect 523868 994780 523920 994832
rect 527916 994780 527968 994832
rect 529020 994780 529072 994832
rect 538220 994780 538272 994832
rect 567936 994780 567988 994832
rect 169392 994712 169444 994764
rect 247684 994712 247736 994764
rect 378600 994712 378652 994764
rect 397000 994712 397052 994764
rect 77668 994644 77720 994696
rect 93308 994644 93360 994696
rect 104900 994644 104952 994696
rect 110512 994644 110564 994696
rect 131580 994644 131632 994696
rect 155960 994644 156012 994696
rect 420644 994644 420696 994696
rect 590568 994644 590620 994696
rect 625712 994780 625764 994832
rect 630864 994780 630916 994832
rect 639512 994644 639564 994696
rect 171048 994576 171100 994628
rect 298560 994576 298612 994628
rect 363604 994576 363656 994628
rect 393964 994576 394016 994628
rect 660764 994576 660816 994628
rect 78312 994508 78364 994560
rect 102784 994508 102836 994560
rect 129740 994508 129792 994560
rect 155316 994508 155368 994560
rect 462964 994508 463016 994560
rect 474648 994508 474700 994560
rect 180156 994440 180208 994492
rect 207388 994440 207440 994492
rect 235908 994440 235960 994492
rect 243728 994440 243780 994492
rect 354404 994440 354456 994492
rect 392676 994440 392728 994492
rect 80704 994372 80756 994424
rect 93124 994372 93176 994424
rect 132132 994372 132184 994424
rect 145748 994372 145800 994424
rect 278136 994372 278188 994424
rect 316408 994372 316460 994424
rect 465724 994372 465776 994424
rect 485964 994508 486016 994560
rect 508504 994508 508556 994560
rect 534356 994508 534408 994560
rect 567752 994508 567804 994560
rect 639052 994508 639104 994560
rect 660948 994508 661000 994560
rect 184664 994304 184716 994356
rect 202328 994304 202380 994356
rect 231584 994304 231636 994356
rect 243360 994304 243412 994356
rect 243544 994304 243596 994356
rect 254584 994304 254636 994356
rect 88984 994236 89036 994288
rect 121736 994236 121788 994288
rect 294144 994236 294196 994288
rect 381176 994236 381228 994288
rect 474648 994236 474700 994288
rect 486608 994372 486660 994424
rect 502984 994372 503036 994424
rect 533712 994372 533764 994424
rect 570144 994372 570196 994424
rect 591304 994372 591356 994424
rect 625528 994372 625580 994424
rect 630220 994372 630272 994424
rect 494060 994236 494112 994288
rect 511080 994236 511132 994288
rect 518164 994236 518216 994288
rect 170680 994100 170732 994152
rect 301504 994100 301556 994152
rect 519544 994100 519596 994152
rect 529020 994100 529072 994152
rect 529388 994236 529440 994288
rect 539232 994236 539284 994288
rect 538404 994100 538456 994152
rect 574100 994032 574152 994084
rect 232228 993964 232280 994016
rect 243544 993964 243596 994016
rect 243728 993964 243780 994016
rect 249248 993964 249300 994016
rect 286508 993964 286560 994016
rect 298376 993964 298428 994016
rect 522948 993964 523000 994016
rect 529388 993964 529440 994016
rect 142068 993896 142120 993948
rect 142344 993896 142396 993948
rect 574744 993896 574796 993948
rect 243360 993828 243412 993880
rect 246212 993828 246264 993880
rect 171232 993760 171284 993812
rect 195796 993760 195848 993812
rect 522764 993760 522816 993812
rect 660764 993760 660816 993812
rect 142068 993692 142120 993744
rect 142252 993624 142304 993676
rect 170864 993624 170916 993676
rect 195612 993624 195664 993676
rect 516324 993624 516376 993676
rect 660948 993624 661000 993676
rect 549168 993488 549220 993540
rect 635832 993488 635884 993540
rect 554780 993352 554832 993404
rect 640708 993352 640760 993404
rect 51724 993148 51776 993200
rect 107936 993148 107988 993200
rect 50344 993012 50396 993064
rect 107752 993012 107804 993064
rect 563704 993012 563756 993064
rect 608600 993012 608652 993064
rect 55864 992876 55916 992928
rect 146944 992876 146996 992928
rect 147680 992876 147732 992928
rect 186504 992876 186556 992928
rect 202880 992876 202932 992928
rect 213920 992876 213972 992928
rect 316684 992876 316736 992928
rect 364984 992876 365036 992928
rect 367928 992876 367980 992928
rect 429936 992876 429988 992928
rect 435548 992876 435600 992928
rect 494704 992876 494756 992928
rect 512828 992876 512880 992928
rect 527272 992876 527324 992928
rect 562508 992876 562560 992928
rect 667204 992876 667256 992928
rect 638868 992264 638920 992316
rect 640800 992264 640852 992316
rect 47584 991720 47636 991772
rect 96068 991720 96120 991772
rect 48964 991584 49016 991636
rect 110696 991584 110748 991636
rect 138296 991584 138348 991636
rect 163136 991584 163188 991636
rect 54484 991448 54536 991500
rect 148324 991448 148376 991500
rect 267004 991448 267056 991500
rect 284300 991448 284352 991500
rect 318064 991448 318116 991500
rect 349160 991448 349212 991500
rect 367744 991448 367796 991500
rect 397828 991448 397880 991500
rect 435364 991448 435416 991500
rect 478972 991448 479024 991500
rect 512644 991448 512696 991500
rect 543832 991448 543884 991500
rect 559564 991448 559616 991500
rect 658924 991448 658976 991500
rect 164884 990836 164936 990888
rect 170772 990836 170824 990888
rect 265624 990836 265676 990888
rect 267648 990836 267700 990888
rect 73436 990224 73488 990276
rect 112076 990224 112128 990276
rect 562324 990224 562376 990276
rect 669964 990224 670016 990276
rect 44824 990088 44876 990140
rect 109040 990088 109092 990140
rect 319444 990088 319496 990140
rect 332968 990088 333020 990140
rect 369124 990088 369176 990140
rect 414112 990088 414164 990140
rect 560944 990088 560996 990140
rect 668584 990088 668636 990140
rect 53288 988728 53340 988780
rect 95884 988728 95936 988780
rect 104900 986620 104952 986672
rect 105820 986620 105872 986672
rect 217324 986620 217376 986672
rect 219440 986620 219492 986672
rect 566464 986076 566516 986128
rect 592500 986076 592552 986128
rect 89628 985940 89680 985992
rect 106924 985940 106976 985992
rect 215944 985940 215996 985992
rect 235632 985940 235684 985992
rect 268384 985940 268436 985992
rect 300492 985940 300544 985992
rect 436744 985940 436796 985992
rect 462780 985940 462832 985992
rect 514024 985940 514076 985992
rect 560116 985940 560168 985992
rect 565084 985940 565136 985992
rect 624976 985940 625028 985992
rect 154488 985668 154540 985720
rect 160744 985668 160796 985720
rect 43444 975672 43496 975724
rect 62120 975672 62172 975724
rect 651656 975672 651708 975724
rect 672724 975672 672776 975724
rect 43444 961868 43496 961920
rect 62120 961868 62172 961920
rect 651472 961868 651524 961920
rect 665824 961868 665876 961920
rect 36544 952416 36596 952468
rect 41696 952416 41748 952468
rect 37924 952212 37976 952264
rect 41696 952212 41748 952264
rect 675852 949424 675904 949476
rect 682384 949424 682436 949476
rect 652208 948064 652260 948116
rect 660304 948064 660356 948116
rect 45560 945956 45612 946008
rect 62120 945956 62172 946008
rect 41236 942556 41288 942608
rect 41696 942556 41748 942608
rect 41236 941196 41288 941248
rect 41696 941196 41748 941248
rect 40960 938612 41012 938664
rect 41420 938612 41472 938664
rect 41144 938408 41196 938460
rect 41512 938408 41564 938460
rect 651472 936980 651524 937032
rect 661684 936980 661736 937032
rect 675852 928752 675904 928804
rect 683120 928752 683172 928804
rect 53104 923244 53156 923296
rect 62120 923244 62172 923296
rect 651472 921816 651524 921868
rect 663064 921816 663116 921868
rect 50344 909440 50396 909492
rect 62120 909440 62172 909492
rect 652392 909440 652444 909492
rect 665824 909440 665876 909492
rect 47768 896996 47820 897048
rect 62120 896996 62172 897048
rect 651472 895636 651524 895688
rect 671344 895636 671396 895688
rect 44088 892712 44140 892764
rect 42938 892270 42990 892322
rect 43076 891896 43128 891948
rect 44088 891828 44140 891880
rect 651656 881832 651708 881884
rect 664444 881832 664496 881884
rect 46204 870816 46256 870868
rect 62120 870816 62172 870868
rect 651472 869388 651524 869440
rect 658924 869388 658976 869440
rect 51724 858372 51776 858424
rect 62120 858372 62172 858424
rect 651472 852116 651524 852168
rect 664444 852116 664496 852168
rect 54484 844568 54536 844620
rect 62120 844568 62172 844620
rect 651840 841780 651892 841832
rect 669964 841780 670016 841832
rect 651472 829404 651524 829456
rect 660304 829404 660356 829456
rect 47584 818320 47636 818372
rect 62120 818320 62172 818372
rect 41236 817028 41288 817080
rect 41696 817028 41748 817080
rect 41236 815600 41288 815652
rect 41604 815600 41656 815652
rect 651472 815600 651524 815652
rect 661684 815600 661736 815652
rect 40776 810704 40828 810756
rect 41696 810704 41748 810756
rect 41144 807372 41196 807424
rect 41604 807372 41656 807424
rect 50344 805944 50396 805996
rect 62120 805944 62172 805996
rect 651472 803224 651524 803276
rect 667204 803156 667256 803208
rect 33048 802408 33100 802460
rect 41696 802408 41748 802460
rect 39304 801728 39356 801780
rect 41604 801660 41656 801712
rect 55864 793568 55916 793620
rect 62120 793568 62172 793620
rect 651472 789352 651524 789404
rect 668584 789352 668636 789404
rect 652392 775548 652444 775600
rect 668768 775548 668820 775600
rect 35808 772828 35860 772880
rect 41696 772828 41748 772880
rect 35808 768952 35860 769004
rect 40040 768952 40092 769004
rect 35532 768816 35584 768868
rect 39304 768816 39356 768868
rect 35348 768680 35400 768732
rect 41696 768680 41748 768732
rect 35808 767456 35860 767508
rect 36544 767456 36596 767508
rect 35624 767320 35676 767372
rect 41328 767320 41380 767372
rect 48964 767320 49016 767372
rect 62120 767320 62172 767372
rect 40040 764736 40092 764788
rect 41696 764736 41748 764788
rect 35808 763240 35860 763292
rect 37924 763240 37976 763292
rect 651472 763240 651524 763292
rect 660304 763172 660356 763224
rect 31024 759636 31076 759688
rect 41696 759636 41748 759688
rect 35164 758276 35216 758328
rect 40316 758276 40368 758328
rect 37924 757732 37976 757784
rect 40316 757732 40368 757784
rect 676036 757120 676088 757172
rect 683396 757120 683448 757172
rect 51724 753516 51776 753568
rect 62120 753516 62172 753568
rect 651472 749368 651524 749420
rect 665824 749368 665876 749420
rect 668400 742704 668452 742756
rect 668768 742704 668820 742756
rect 54484 741072 54536 741124
rect 62120 741072 62172 741124
rect 651840 735564 651892 735616
rect 661868 735564 661920 735616
rect 35808 730056 35860 730108
rect 41696 730056 41748 730108
rect 674380 728560 674432 728612
rect 672172 728424 672224 728476
rect 672356 728288 672408 728340
rect 673184 728084 673236 728136
rect 41328 725908 41380 725960
rect 41696 725908 41748 725960
rect 41328 724752 41380 724804
rect 41696 724752 41748 724804
rect 677324 724208 677376 724260
rect 683212 724208 683264 724260
rect 651472 723120 651524 723172
rect 663064 723120 663116 723172
rect 34152 720264 34204 720316
rect 38660 720264 38712 720316
rect 36544 717340 36596 717392
rect 41696 717340 41748 717392
rect 39304 716184 39356 716236
rect 41512 716184 41564 716236
rect 34520 715504 34572 715556
rect 40316 715504 40368 715556
rect 50344 714824 50396 714876
rect 62120 714824 62172 714876
rect 652576 709316 652628 709368
rect 664444 709316 664496 709368
rect 55864 701020 55916 701072
rect 62120 701020 62172 701072
rect 652392 696940 652444 696992
rect 669964 696940 670016 696992
rect 53104 688644 53156 688696
rect 62120 688644 62172 688696
rect 35808 687216 35860 687268
rect 41420 687216 41472 687268
rect 35808 683136 35860 683188
rect 41696 683136 41748 683188
rect 651840 683136 651892 683188
rect 658924 683136 658976 683188
rect 35808 681980 35860 682032
rect 36544 681980 36596 682032
rect 35624 681844 35676 681896
rect 41696 681844 41748 681896
rect 35440 681708 35492 681760
rect 41604 681640 41656 681692
rect 51724 674840 51776 674892
rect 62120 674840 62172 674892
rect 32404 672732 32456 672784
rect 41604 672732 41656 672784
rect 36544 671644 36596 671696
rect 39672 671644 39724 671696
rect 35164 671304 35216 671356
rect 41328 671304 41380 671356
rect 652392 669332 652444 669384
rect 668400 669332 668452 669384
rect 671988 665660 672040 665712
rect 673000 665660 673052 665712
rect 47584 662396 47636 662448
rect 62120 662396 62172 662448
rect 651656 656888 651708 656940
rect 663064 656888 663116 656940
rect 54484 647844 54536 647896
rect 62120 647844 62172 647896
rect 651472 643084 651524 643136
rect 668584 643084 668636 643136
rect 35808 639072 35860 639124
rect 36544 639072 36596 639124
rect 35624 638936 35676 638988
rect 41512 638936 41564 638988
rect 35808 636828 35860 636880
rect 41696 636828 41748 636880
rect 51724 636216 51776 636268
rect 62120 636216 62172 636268
rect 675852 634176 675904 634228
rect 682384 634176 682436 634228
rect 32404 629892 32456 629944
rect 41696 629892 41748 629944
rect 651564 628532 651616 628584
rect 667204 628532 667256 628584
rect 48964 623772 49016 623824
rect 62120 623772 62172 623824
rect 675852 622820 675904 622872
rect 676680 622820 676732 622872
rect 651472 616836 651524 616888
rect 660304 616836 660356 616888
rect 43260 612892 43312 612944
rect 46940 612688 46992 612740
rect 43720 612484 43772 612536
rect 43582 612280 43634 612332
rect 43904 612076 43956 612128
rect 45560 611872 45612 611924
rect 43931 611668 43983 611720
rect 44916 611464 44968 611516
rect 44155 611328 44207 611380
rect 44732 611056 44784 611108
rect 45744 610852 45796 610904
rect 44502 610716 44554 610768
rect 56048 608608 56100 608660
rect 62120 608608 62172 608660
rect 651472 603100 651524 603152
rect 661684 603100 661736 603152
rect 673460 598612 673512 598664
rect 673828 598612 673880 598664
rect 48964 597524 49016 597576
rect 62120 597524 62172 597576
rect 40868 592832 40920 592884
rect 41604 592832 41656 592884
rect 673828 592424 673880 592476
rect 40316 592288 40368 592340
rect 41420 592288 41472 592340
rect 673552 592152 673604 592204
rect 675852 591336 675904 591388
rect 682384 591336 682436 591388
rect 652392 590656 652444 590708
rect 665824 590656 665876 590708
rect 33048 587120 33100 587172
rect 40408 587120 40460 587172
rect 39948 586100 40000 586152
rect 41696 586100 41748 586152
rect 35164 585896 35216 585948
rect 41696 585896 41748 585948
rect 31024 585760 31076 585812
rect 41696 585692 41748 585744
rect 40868 584536 40920 584588
rect 41604 584536 41656 584588
rect 50344 583720 50396 583772
rect 62120 583720 62172 583772
rect 672172 579028 672224 579080
rect 673184 579028 673236 579080
rect 651472 576852 651524 576904
rect 664444 576852 664496 576904
rect 651656 563048 651708 563100
rect 658924 563048 658976 563100
rect 55864 558084 55916 558136
rect 62120 558084 62172 558136
rect 35808 557540 35860 557592
rect 41512 557540 41564 557592
rect 673644 558288 673696 558340
rect 673644 557812 673696 557864
rect 673644 557676 673696 557728
rect 673552 557404 673604 557456
rect 35808 554752 35860 554804
rect 41696 554752 41748 554804
rect 35808 553392 35860 553444
rect 41328 553392 41380 553444
rect 41328 552032 41380 552084
rect 41696 552032 41748 552084
rect 651472 550604 651524 550656
rect 660304 550604 660356 550656
rect 41236 548088 41288 548140
rect 41696 548088 41748 548140
rect 31760 547816 31812 547868
rect 38476 547816 38528 547868
rect 675852 546456 675904 546508
rect 681004 546456 681056 546508
rect 47584 545096 47636 545148
rect 62120 545096 62172 545148
rect 33784 542988 33836 543040
rect 41512 542988 41564 543040
rect 38476 542308 38528 542360
rect 41696 542308 41748 542360
rect 651472 536800 651524 536852
rect 669412 536800 669464 536852
rect 50344 532720 50396 532772
rect 62120 532720 62172 532772
rect 651840 522996 651892 523048
rect 661868 522996 661920 523048
rect 676864 520276 676916 520328
rect 683120 520276 683172 520328
rect 54484 518916 54536 518968
rect 62120 518916 62172 518968
rect 675852 518780 675904 518832
rect 677876 518780 677928 518832
rect 651472 510620 651524 510672
rect 659108 510620 659160 510672
rect 46204 506472 46256 506524
rect 62120 506472 62172 506524
rect 676036 502324 676088 502376
rect 678244 502324 678296 502376
rect 675852 500896 675904 500948
rect 681004 500896 681056 500948
rect 652576 494708 652628 494760
rect 663248 494708 663300 494760
rect 48964 491920 49016 491972
rect 62120 491920 62172 491972
rect 677508 491104 677560 491156
rect 683304 491104 683356 491156
rect 651472 484440 651524 484492
rect 667204 484372 667256 484424
rect 681004 481516 681056 481568
rect 683120 481516 683172 481568
rect 51724 480224 51776 480276
rect 62120 480224 62172 480276
rect 651472 470568 651524 470620
rect 665824 470568 665876 470620
rect 51908 466420 51960 466472
rect 62120 466420 62172 466472
rect 652392 456764 652444 456816
rect 661684 456764 661736 456816
rect 673948 456152 674000 456204
rect 673828 455948 673880 456000
rect 673460 455812 673512 455864
rect 673598 455608 673650 455660
rect 673276 455336 673328 455388
rect 673388 455200 673440 455252
rect 672080 455064 672132 455116
rect 673046 454792 673098 454844
rect 672908 454656 672960 454708
rect 673164 454588 673216 454640
rect 672816 454180 672868 454232
rect 53104 454044 53156 454096
rect 62120 454044 62172 454096
rect 672724 453908 672776 453960
rect 651472 444456 651524 444508
rect 668584 444388 668636 444440
rect 50528 440240 50580 440292
rect 62120 440240 62172 440292
rect 651472 430584 651524 430636
rect 669964 430584 670016 430636
rect 54484 427796 54536 427848
rect 62120 427796 62172 427848
rect 651840 416780 651892 416832
rect 663064 416780 663116 416832
rect 33784 416032 33836 416084
rect 41696 416032 41748 416084
rect 651472 404336 651524 404388
rect 664444 404336 664496 404388
rect 55864 401616 55916 401668
rect 62120 401616 62172 401668
rect 675852 395700 675904 395752
rect 676404 395700 676456 395752
rect 652576 390532 652628 390584
rect 658924 390532 658976 390584
rect 47768 389240 47820 389292
rect 62120 389240 62172 389292
rect 35808 382508 35860 382560
rect 40040 382508 40092 382560
rect 35624 382372 35676 382424
rect 41696 382372 41748 382424
rect 35440 382236 35492 382288
rect 41512 382236 41564 382288
rect 35532 381012 35584 381064
rect 37924 381012 37976 381064
rect 35808 380876 35860 380928
rect 41328 380876 41380 380928
rect 652392 378156 652444 378208
rect 660304 378156 660356 378208
rect 35808 375980 35860 376032
rect 39580 375980 39632 376032
rect 51908 375368 51960 375420
rect 62120 375368 62172 375420
rect 651840 364352 651892 364404
rect 661868 364352 661920 364404
rect 50344 362924 50396 362976
rect 62120 362924 62172 362976
rect 44640 354968 44692 355020
rect 44824 354560 44876 354612
rect 44575 354492 44627 354544
rect 44799 354424 44851 354476
rect 44799 354288 44851 354340
rect 45192 353812 45244 353864
rect 45146 353676 45198 353728
rect 45359 353268 45411 353320
rect 652392 350548 652444 350600
rect 667204 350548 667256 350600
rect 46204 347012 46256 347064
rect 62120 347012 62172 347064
rect 35808 343612 35860 343664
rect 40224 343612 40276 343664
rect 35808 339464 35860 339516
rect 37556 339464 37608 339516
rect 54484 336744 54536 336796
rect 62120 336744 62172 336796
rect 651472 324300 651524 324352
rect 666652 324300 666704 324352
rect 51724 310496 51776 310548
rect 62120 310496 62172 310548
rect 651472 310496 651524 310548
rect 667388 310496 667440 310548
rect 45468 298120 45520 298172
rect 62120 298120 62172 298172
rect 675944 298052 675996 298104
rect 678980 298052 679032 298104
rect 676220 297032 676272 297084
rect 681004 297032 681056 297084
rect 41328 284928 41380 284980
rect 41696 284928 41748 284980
rect 39304 284724 39356 284776
rect 41696 284724 41748 284776
rect 651472 284316 651524 284368
rect 667572 284316 667624 284368
rect 482836 276632 482888 276684
rect 558828 276632 558880 276684
rect 103704 275952 103756 276004
rect 160744 275952 160796 276004
rect 166356 275952 166408 276004
rect 182088 275952 182140 276004
rect 188804 275952 188856 276004
rect 221464 275952 221516 276004
rect 410064 275952 410116 276004
rect 88340 275816 88392 275868
rect 146944 275816 146996 275868
rect 149796 275816 149848 275868
rect 187884 275816 187936 275868
rect 368848 275816 368900 275868
rect 373264 275816 373316 275868
rect 393780 275816 393832 275868
rect 411076 275816 411128 275868
rect 419540 275952 419592 276004
rect 439412 275952 439464 276004
rect 456064 275952 456116 276004
rect 466644 275952 466696 276004
rect 466828 275952 466880 276004
rect 523408 275952 523460 276004
rect 525800 275952 525852 276004
rect 607312 275952 607364 276004
rect 424048 275816 424100 275868
rect 432788 275816 432840 275868
rect 487896 275816 487948 275868
rect 504732 275816 504784 275868
rect 590752 275816 590804 275868
rect 220728 275748 220780 275800
rect 224960 275748 225012 275800
rect 249064 275748 249116 275800
rect 253480 275748 253532 275800
rect 277492 275748 277544 275800
rect 285128 275748 285180 275800
rect 96620 275680 96672 275732
rect 156604 275680 156656 275732
rect 174636 275680 174688 275732
rect 208400 275680 208452 275732
rect 212448 275680 212500 275732
rect 219900 275680 219952 275732
rect 232504 275680 232556 275732
rect 245660 275680 245712 275732
rect 373264 275680 373316 275732
rect 385040 275680 385092 275732
rect 400220 275680 400272 275732
rect 418160 275680 418212 275732
rect 418344 275680 418396 275732
rect 435916 275680 435968 275732
rect 259736 275612 259788 275664
rect 267004 275612 267056 275664
rect 85948 275544 86000 275596
rect 150808 275544 150860 275596
rect 160468 275544 160520 275596
rect 172428 275544 172480 275596
rect 181720 275544 181772 275596
rect 218612 275544 218664 275596
rect 225420 275544 225472 275596
rect 243544 275544 243596 275596
rect 244372 275544 244424 275596
rect 247040 275544 247092 275596
rect 283380 275544 283432 275596
rect 289084 275544 289136 275596
rect 367836 275544 367888 275596
rect 377956 275544 378008 275596
rect 382464 275544 382516 275596
rect 400404 275544 400456 275596
rect 403440 275544 403492 275596
rect 428832 275544 428884 275596
rect 435732 275544 435784 275596
rect 491484 275680 491536 275732
rect 493876 275680 493928 275732
rect 502064 275680 502116 275732
rect 505836 275680 505888 275732
rect 512736 275680 512788 275732
rect 516416 275680 516468 275732
rect 604920 275680 604972 275732
rect 605104 275680 605156 275732
rect 616788 275680 616840 275732
rect 441344 275544 441396 275596
rect 498568 275544 498620 275596
rect 510068 275544 510120 275596
rect 519820 275544 519872 275596
rect 523040 275544 523092 275596
rect 525616 275544 525668 275596
rect 525984 275544 526036 275596
rect 619088 275544 619140 275596
rect 625804 275544 625856 275596
rect 640432 275544 640484 275596
rect 76472 275408 76524 275460
rect 143264 275408 143316 275460
rect 148600 275408 148652 275460
rect 164148 275408 164200 275460
rect 167552 275408 167604 275460
rect 209044 275408 209096 275460
rect 218336 275408 218388 275460
rect 239404 275408 239456 275460
rect 253664 275408 253716 275460
rect 261484 275408 261536 275460
rect 284576 275408 284628 275460
rect 290096 275408 290148 275460
rect 349804 275408 349856 275460
rect 361396 275408 361448 275460
rect 362960 275408 363012 275460
rect 367284 275408 367336 275460
rect 376668 275408 376720 275460
rect 393320 275408 393372 275460
rect 395436 275408 395488 275460
rect 403992 275408 404044 275460
rect 407764 275408 407816 275460
rect 432328 275408 432380 275460
rect 438860 275408 438912 275460
rect 446496 275408 446548 275460
rect 450544 275408 450596 275460
rect 509148 275408 509200 275460
rect 512184 275408 512236 275460
rect 533988 275408 534040 275460
rect 535736 275408 535788 275460
rect 633348 275408 633400 275460
rect 70584 275272 70636 275324
rect 140136 275272 140188 275324
rect 156880 275272 156932 275324
rect 199292 275272 199344 275324
rect 211252 275272 211304 275324
rect 232688 275272 232740 275324
rect 246764 275272 246816 275324
rect 256700 275272 256752 275324
rect 260932 275272 260984 275324
rect 273536 275272 273588 275324
rect 273904 275272 273956 275324
rect 283288 275272 283340 275324
rect 328276 275272 328328 275324
rect 335360 275272 335412 275324
rect 347044 275272 347096 275324
rect 356704 275272 356756 275324
rect 359464 275272 359516 275324
rect 370872 275272 370924 275324
rect 377404 275272 377456 275324
rect 396908 275272 396960 275324
rect 400404 275272 400456 275324
rect 425244 275272 425296 275324
rect 427820 275272 427872 275324
rect 443000 275272 443052 275324
rect 453764 275272 453816 275324
rect 516232 275272 516284 275324
rect 523684 275272 523736 275324
rect 545856 275272 545908 275324
rect 546040 275272 546092 275324
rect 552940 275272 552992 275324
rect 553124 275272 553176 275324
rect 574192 275272 574244 275324
rect 110788 275136 110840 275188
rect 164976 275136 165028 275188
rect 171048 275136 171100 275188
rect 191012 275136 191064 275188
rect 428924 275136 428976 275188
rect 135628 275000 135680 275052
rect 167644 275000 167696 275052
rect 290464 275000 290516 275052
rect 294328 275000 294380 275052
rect 366364 275000 366416 275052
rect 369676 275000 369728 275052
rect 426256 275000 426308 275052
rect 477224 275000 477276 275052
rect 481548 275136 481600 275188
rect 544660 275136 544712 275188
rect 552664 275136 552716 275188
rect 560024 275136 560076 275188
rect 480812 275000 480864 275052
rect 487804 275000 487856 275052
rect 530492 275000 530544 275052
rect 530676 275000 530728 275052
rect 541072 275000 541124 275052
rect 542268 275000 542320 275052
rect 549352 275000 549404 275052
rect 551560 275000 551612 275052
rect 553124 275000 553176 275052
rect 559564 275000 559616 275052
rect 567108 275000 567160 275052
rect 81256 274932 81308 274984
rect 86224 274932 86276 274984
rect 129648 274864 129700 274916
rect 136088 274864 136140 274916
rect 142712 274864 142764 274916
rect 166264 274864 166316 274916
rect 469404 274864 469456 274916
rect 483204 274864 483256 274916
rect 490564 274864 490616 274916
rect 526904 274864 526956 274916
rect 543280 274864 543332 274916
rect 645124 274864 645176 274916
rect 199476 274796 199528 274848
rect 202236 274796 202288 274848
rect 208860 274796 208912 274848
rect 211068 274796 211120 274848
rect 257344 274796 257396 274848
rect 259920 274796 259972 274848
rect 357256 274796 357308 274848
rect 360200 274796 360252 274848
rect 369860 274796 369912 274848
rect 375564 274796 375616 274848
rect 146208 274728 146260 274780
rect 149704 274728 149756 274780
rect 150992 274728 151044 274780
rect 152740 274728 152792 274780
rect 163964 274728 164016 274780
rect 170404 274728 170456 274780
rect 172244 274728 172296 274780
rect 174360 274728 174412 274780
rect 387708 274728 387760 274780
rect 394516 274728 394568 274780
rect 397092 274728 397144 274780
rect 401508 274728 401560 274780
rect 415216 274728 415268 274780
rect 419356 274728 419408 274780
rect 446404 274728 446456 274780
rect 453580 274728 453632 274780
rect 483664 274728 483716 274780
rect 493876 274728 493928 274780
rect 498476 274728 498528 274780
rect 499764 274728 499816 274780
rect 501604 274728 501656 274780
rect 505652 274728 505704 274780
rect 506480 274728 506532 274780
rect 510344 274728 510396 274780
rect 510528 274728 510580 274780
rect 537300 274728 537352 274780
rect 537668 274728 537720 274780
rect 538772 274728 538824 274780
rect 539508 274728 539560 274780
rect 542084 274728 542136 274780
rect 71780 274660 71832 274712
rect 73804 274660 73856 274712
rect 74080 274660 74132 274712
rect 77208 274660 77260 274712
rect 210056 274660 210108 274712
rect 212264 274660 212316 274712
rect 243176 274660 243228 274712
rect 249064 274660 249116 274712
rect 289268 274660 289320 274712
rect 292764 274660 292816 274712
rect 296352 274660 296404 274712
rect 298376 274660 298428 274712
rect 298744 274660 298796 274712
rect 300124 274660 300176 274712
rect 324964 274660 325016 274712
rect 327080 274660 327132 274712
rect 338028 274660 338080 274712
rect 343640 274660 343692 274712
rect 344284 274660 344336 274712
rect 347228 274660 347280 274712
rect 347412 274660 347464 274712
rect 349620 274660 349672 274712
rect 360200 274660 360252 274712
rect 363788 274660 363840 274712
rect 478972 274660 479024 274712
rect 482008 274660 482060 274712
rect 619180 274660 619232 274712
rect 623872 274660 623924 274712
rect 120264 274592 120316 274644
rect 175280 274592 175332 274644
rect 384948 274592 385000 274644
rect 400220 274592 400272 274644
rect 403992 274592 404044 274644
rect 438860 274592 438912 274644
rect 445024 274592 445076 274644
rect 478420 274592 478472 274644
rect 482192 274592 482244 274644
rect 556436 274592 556488 274644
rect 559748 274592 559800 274644
rect 587164 274592 587216 274644
rect 114284 274456 114336 274508
rect 171600 274456 171652 274508
rect 179328 274456 179380 274508
rect 213184 274456 213236 274508
rect 213644 274456 213696 274508
rect 240416 274456 240468 274508
rect 378784 274456 378836 274508
rect 93032 274320 93084 274372
rect 95884 274320 95936 274372
rect 97724 274320 97776 274372
rect 158812 274320 158864 274372
rect 180524 274320 180576 274372
rect 216956 274320 217008 274372
rect 368296 274320 368348 274372
rect 387708 274320 387760 274372
rect 95424 274184 95476 274236
rect 157616 274184 157668 274236
rect 165620 274184 165672 274236
rect 205732 274184 205784 274236
rect 206560 274184 206612 274236
rect 234620 274184 234672 274236
rect 245660 274184 245712 274236
rect 254032 274184 254084 274236
rect 351184 274184 351236 274236
rect 362592 274184 362644 274236
rect 77668 274048 77720 274100
rect 145104 274048 145156 274100
rect 145288 274048 145340 274100
rect 189816 274048 189868 274100
rect 191196 274048 191248 274100
rect 224776 274048 224828 274100
rect 224960 274048 225012 274100
rect 245752 274048 245804 274100
rect 253480 274048 253532 274100
rect 265256 274048 265308 274100
rect 339132 274048 339184 274100
rect 353116 274048 353168 274100
rect 362776 274048 362828 274100
rect 386236 274184 386288 274236
rect 400128 274456 400180 274508
rect 419540 274456 419592 274508
rect 420736 274456 420788 274508
rect 470140 274456 470192 274508
rect 474372 274456 474424 274508
rect 523684 274456 523736 274508
rect 537484 274456 537536 274508
rect 613200 274456 613252 274508
rect 397276 274320 397328 274372
rect 418344 274320 418396 274372
rect 419172 274320 419224 274372
rect 467840 274320 467892 274372
rect 408684 274184 408736 274236
rect 427452 274184 427504 274236
rect 479340 274320 479392 274372
rect 479524 274320 479576 274372
rect 481548 274320 481600 274372
rect 487068 274320 487120 274372
rect 563520 274320 563572 274372
rect 563704 274320 563756 274372
rect 612004 274320 612056 274372
rect 471980 274184 472032 274236
rect 385684 274048 385736 274100
rect 395160 274048 395212 274100
rect 395620 274048 395672 274100
rect 426440 274048 426492 274100
rect 446588 274048 446640 274100
rect 468944 274048 468996 274100
rect 469128 274048 469180 274100
rect 75276 273912 75328 273964
rect 142160 273912 142212 273964
rect 147404 273912 147456 273964
rect 193312 273912 193364 273964
rect 193496 273912 193548 273964
rect 222844 273912 222896 273964
rect 223120 273912 223172 273964
rect 130844 273776 130896 273828
rect 181444 273776 181496 273828
rect 247040 273912 247092 273964
rect 262220 273912 262272 273964
rect 265624 273912 265676 273964
rect 276848 273912 276900 273964
rect 322756 273912 322808 273964
rect 330668 273912 330720 273964
rect 333796 273912 333848 273964
rect 344836 273912 344888 273964
rect 247040 273776 247092 273828
rect 344652 273776 344704 273828
rect 349804 273776 349856 273828
rect 350356 273776 350408 273828
rect 366364 273912 366416 273964
rect 367008 273912 367060 273964
rect 376668 273912 376720 273964
rect 376576 273776 376628 273828
rect 407488 273912 407540 273964
rect 409236 273912 409288 273964
rect 446404 273912 446456 273964
rect 468484 273912 468536 273964
rect 471980 273912 472032 273964
rect 475568 274048 475620 274100
rect 479524 274048 479576 274100
rect 481364 274184 481416 274236
rect 482192 274184 482244 274236
rect 500868 274184 500920 274236
rect 583668 274184 583720 274236
rect 494980 274048 495032 274100
rect 533436 274048 533488 274100
rect 630956 274048 631008 274100
rect 532792 273912 532844 273964
rect 542084 273912 542136 273964
rect 642732 273912 642784 273964
rect 431684 273776 431736 273828
rect 485504 273776 485556 273828
rect 488356 273776 488408 273828
rect 559564 273776 559616 273828
rect 124956 273640 125008 273692
rect 148416 273640 148468 273692
rect 155684 273640 155736 273692
rect 198096 273640 198148 273692
rect 457444 273640 457496 273692
rect 484308 273640 484360 273692
rect 484492 273640 484544 273692
rect 552664 273640 552716 273692
rect 439320 273504 439372 273556
rect 471336 273504 471388 273556
rect 473084 273504 473136 273556
rect 475568 273504 475620 273556
rect 478788 273504 478840 273556
rect 546040 273504 546092 273556
rect 552664 273504 552716 273556
rect 580080 273504 580132 273556
rect 464804 273368 464856 273420
rect 469128 273368 469180 273420
rect 475936 273368 475988 273420
rect 542268 273368 542320 273420
rect 330484 273232 330536 273284
rect 333060 273232 333112 273284
rect 127348 273164 127400 273216
rect 179880 273164 179932 273216
rect 401508 273164 401560 273216
rect 427820 273164 427872 273216
rect 438124 273164 438176 273216
rect 464252 273164 464304 273216
rect 471612 273164 471664 273216
rect 543464 273164 543516 273216
rect 111984 273028 112036 273080
rect 168380 273028 168432 273080
rect 182088 273028 182140 273080
rect 207296 273028 207348 273080
rect 382004 273028 382056 273080
rect 414572 273028 414624 273080
rect 429844 273028 429896 273080
rect 447692 273028 447744 273080
rect 451096 273028 451148 273080
rect 513932 273028 513984 273080
rect 520096 273028 520148 273080
rect 610808 273028 610860 273080
rect 102508 272892 102560 272944
rect 162124 272892 162176 272944
rect 190000 272892 190052 272944
rect 94228 272756 94280 272808
rect 155960 272756 156012 272808
rect 187608 272756 187660 272808
rect 212540 272756 212592 272808
rect 217140 272892 217192 272944
rect 242992 272892 243044 272944
rect 286876 272892 286928 272944
rect 287704 272892 287756 272944
rect 388812 272892 388864 272944
rect 400404 272892 400456 272944
rect 406844 272892 406896 272944
rect 450084 272892 450136 272944
rect 457996 272892 458048 272944
rect 522212 272892 522264 272944
rect 524052 272892 524104 272944
rect 617984 272892 618036 272944
rect 217416 272756 217468 272808
rect 219900 272756 219952 272808
rect 239220 272756 239272 272808
rect 252652 272756 252704 272808
rect 267832 272756 267884 272808
rect 343548 272756 343600 272808
rect 359004 272756 359056 272808
rect 360844 272756 360896 272808
rect 381544 272756 381596 272808
rect 394332 272756 394384 272808
rect 407764 272756 407816 272808
rect 408408 272756 408460 272808
rect 452108 272756 452160 272808
rect 452292 272756 452344 272808
rect 515128 272756 515180 272808
rect 517336 272756 517388 272808
rect 525800 272756 525852 272808
rect 526812 272756 526864 272808
rect 621480 272756 621532 272808
rect 82360 272620 82412 272672
rect 148232 272620 148284 272672
rect 161572 272620 161624 272672
rect 203064 272620 203116 272672
rect 203248 272620 203300 272672
rect 233240 272620 233292 272672
rect 239588 272620 239640 272672
rect 254584 272620 254636 272672
rect 280988 272620 281040 272672
rect 286324 272620 286376 272672
rect 349804 272620 349856 272672
rect 366088 272620 366140 272672
rect 370964 272620 371016 272672
rect 399208 272620 399260 272672
rect 412272 272620 412324 272672
rect 457168 272620 457220 272672
rect 461952 272620 462004 272672
rect 529296 272620 529348 272672
rect 529756 272620 529808 272672
rect 625068 272620 625120 272672
rect 65892 272484 65944 272536
rect 136824 272484 136876 272536
rect 137928 272484 137980 272536
rect 187700 272484 187752 272536
rect 192300 272484 192352 272536
rect 225512 272484 225564 272536
rect 236092 272484 236144 272536
rect 253204 272484 253256 272536
rect 255044 272484 255096 272536
rect 269304 272484 269356 272536
rect 270224 272484 270276 272536
rect 280344 272484 280396 272536
rect 331036 272484 331088 272536
rect 342444 272484 342496 272536
rect 356888 272484 356940 272536
rect 376852 272484 376904 272536
rect 380808 272484 380860 272536
rect 411996 272484 412048 272536
rect 413928 272484 413980 272536
rect 460664 272484 460716 272536
rect 467748 272484 467800 272536
rect 536380 272484 536432 272536
rect 539324 272484 539376 272536
rect 639236 272484 639288 272536
rect 128544 272348 128596 272400
rect 181260 272348 181312 272400
rect 212540 272348 212592 272400
rect 218796 272348 218848 272400
rect 457812 272348 457864 272400
rect 466828 272348 466880 272400
rect 470508 272348 470560 272400
rect 539876 272348 539928 272400
rect 541624 272348 541676 272400
rect 603724 272348 603776 272400
rect 116676 272212 116728 272264
rect 166080 272212 166132 272264
rect 166264 272212 166316 272264
rect 191840 272212 191892 272264
rect 424968 272212 425020 272264
rect 474924 272212 474976 272264
rect 479708 272212 479760 272264
rect 548156 272212 548208 272264
rect 152188 272076 152240 272128
rect 192484 272076 192536 272128
rect 447784 272076 447836 272128
rect 506848 272076 506900 272128
rect 514024 272076 514076 272128
rect 565912 272076 565964 272128
rect 121368 271804 121420 271856
rect 176752 271804 176804 271856
rect 185216 271804 185268 271856
rect 186964 271804 187016 271856
rect 187884 271804 187936 271856
rect 196440 271804 196492 271856
rect 276296 271804 276348 271856
rect 278044 271804 278096 271856
rect 288072 271804 288124 271856
rect 292948 271804 293000 271856
rect 293224 271804 293276 271856
rect 295800 271804 295852 271856
rect 375288 271804 375340 271856
rect 395436 271804 395488 271856
rect 434444 271804 434496 271856
rect 490288 271804 490340 271856
rect 496544 271804 496596 271856
rect 578884 271804 578936 271856
rect 318616 271736 318668 271788
rect 324780 271736 324832 271788
rect 104900 271668 104952 271720
rect 163320 271668 163372 271720
rect 164148 271668 164200 271720
rect 194784 271668 194836 271720
rect 197084 271668 197136 271720
rect 224224 271668 224276 271720
rect 224592 271668 224644 271720
rect 247776 271668 247828 271720
rect 363604 271668 363656 271720
rect 374368 271668 374420 271720
rect 384764 271668 384816 271720
rect 415216 271668 415268 271720
rect 418804 271668 418856 271720
rect 429660 271668 429712 271720
rect 437204 271668 437256 271720
rect 493692 271668 493744 271720
rect 499488 271668 499540 271720
rect 582472 271668 582524 271720
rect 106004 271532 106056 271584
rect 164792 271532 164844 271584
rect 178132 271532 178184 271584
rect 184204 271532 184256 271584
rect 184480 271532 184532 271584
rect 215944 271532 215996 271584
rect 216312 271532 216364 271584
rect 242072 271532 242124 271584
rect 248420 271532 248472 271584
rect 264336 271532 264388 271584
rect 340604 271532 340656 271584
rect 355140 271532 355192 271584
rect 355324 271532 355376 271584
rect 368480 271532 368532 271584
rect 369492 271532 369544 271584
rect 377404 271532 377456 271584
rect 379336 271532 379388 271584
rect 393780 271532 393832 271584
rect 395528 271532 395580 271584
rect 427636 271532 427688 271584
rect 89536 271396 89588 271448
rect 152372 271396 152424 271448
rect 162768 271396 162820 271448
rect 204720 271396 204772 271448
rect 205364 271396 205416 271448
rect 234988 271396 235040 271448
rect 241888 271396 241940 271448
rect 260288 271396 260340 271448
rect 334624 271396 334676 271448
rect 341340 271396 341392 271448
rect 348884 271396 348936 271448
rect 362960 271396 363012 271448
rect 366364 271396 366416 271448
rect 379152 271396 379204 271448
rect 387616 271396 387668 271448
rect 421656 271396 421708 271448
rect 425704 271396 425756 271448
rect 432972 271396 433024 271448
rect 437940 271396 437992 271448
rect 68192 271260 68244 271312
rect 138480 271260 138532 271312
rect 139124 271260 139176 271312
rect 141608 271260 141660 271312
rect 141792 271260 141844 271312
rect 189632 271260 189684 271312
rect 195704 271260 195756 271312
rect 227904 271260 227956 271312
rect 228824 271260 228876 271312
rect 236828 271260 236880 271312
rect 237288 271260 237340 271312
rect 256976 271260 257028 271312
rect 259920 271260 259972 271312
rect 270960 271260 271012 271312
rect 271512 271260 271564 271312
rect 280896 271260 280948 271312
rect 315764 271260 315816 271312
rect 319996 271260 320048 271312
rect 329748 271260 329800 271312
rect 338948 271260 339000 271312
rect 341524 271260 341576 271312
rect 348424 271260 348476 271312
rect 354588 271260 354640 271312
rect 369860 271260 369912 271312
rect 372528 271260 372580 271312
rect 382464 271260 382516 271312
rect 383384 271260 383436 271312
rect 416964 271260 417016 271312
rect 421564 271260 421616 271312
rect 437020 271260 437072 271312
rect 442908 271532 442960 271584
rect 500500 271532 500552 271584
rect 501972 271532 502024 271584
rect 585600 271532 585652 271584
rect 585784 271532 585836 271584
rect 608508 271532 608560 271584
rect 439964 271396 440016 271448
rect 497004 271396 497056 271448
rect 504916 271396 504968 271448
rect 589556 271396 589608 271448
rect 592684 271396 592736 271448
rect 622676 271396 622728 271448
rect 72976 271124 73028 271176
rect 142344 271124 142396 271176
rect 143264 271124 143316 271176
rect 144368 271124 144420 271176
rect 154304 271124 154356 271176
rect 197912 271124 197964 271176
rect 198280 271124 198332 271176
rect 229560 271124 229612 271176
rect 231400 271124 231452 271176
rect 252744 271124 252796 271176
rect 263232 271124 263284 271176
rect 275284 271124 275336 271176
rect 279792 271124 279844 271176
rect 287152 271124 287204 271176
rect 325516 271124 325568 271176
rect 334164 271124 334216 271176
rect 339316 271124 339368 271176
rect 354312 271124 354364 271176
rect 362684 271124 362736 271176
rect 387156 271124 387208 271176
rect 391756 271124 391808 271176
rect 403440 271124 403492 271176
rect 405004 271124 405056 271176
rect 445668 271260 445720 271312
rect 504456 271260 504508 271312
rect 509148 271260 509200 271312
rect 596640 271260 596692 271312
rect 596824 271260 596876 271312
rect 629760 271260 629812 271312
rect 83556 270988 83608 271040
rect 123484 270988 123536 271040
rect 123760 270988 123812 271040
rect 177488 270988 177540 271040
rect 448888 271124 448940 271176
rect 449808 271124 449860 271176
rect 511540 271124 511592 271176
rect 511908 271124 511960 271176
rect 600228 271124 600280 271176
rect 602344 271124 602396 271176
rect 643928 271124 643980 271176
rect 434720 270988 434772 271040
rect 434904 270988 434956 271040
rect 486700 270988 486752 271040
rect 495256 270988 495308 271040
rect 575388 270988 575440 271040
rect 576124 270988 576176 271040
rect 594340 270988 594392 271040
rect 134432 270852 134484 270904
rect 184940 270852 184992 270904
rect 418068 270852 418120 270904
rect 456064 270852 456116 270904
rect 492588 270852 492640 270904
rect 571800 270852 571852 270904
rect 113180 270716 113232 270768
rect 154028 270716 154080 270768
rect 175832 270716 175884 270768
rect 206284 270716 206336 270768
rect 404176 270716 404228 270768
rect 445300 270716 445352 270768
rect 459192 270716 459244 270768
rect 523040 270716 523092 270768
rect 526444 270716 526496 270768
rect 576584 270716 576636 270768
rect 414480 270580 414532 270632
rect 432972 270580 433024 270632
rect 433156 270580 433208 270632
rect 434904 270580 434956 270632
rect 456064 270580 456116 270632
rect 507952 270580 508004 270632
rect 509700 270580 509752 270632
rect 510528 270580 510580 270632
rect 100668 270444 100720 270496
rect 119804 270444 119856 270496
rect 122748 270444 122800 270496
rect 176200 270444 176252 270496
rect 176936 270444 176988 270496
rect 214748 270444 214800 270496
rect 219532 270444 219584 270496
rect 78864 270308 78916 270360
rect 132592 270308 132644 270360
rect 133788 270308 133840 270360
rect 183652 270308 183704 270360
rect 186412 270308 186464 270360
rect 201592 270308 201644 270360
rect 204168 270308 204220 270360
rect 220268 270308 220320 270360
rect 230388 270444 230440 270496
rect 252100 270444 252152 270496
rect 275100 270444 275152 270496
rect 276020 270444 276072 270496
rect 278688 270444 278740 270496
rect 285956 270444 286008 270496
rect 291660 270444 291712 270496
rect 295524 270444 295576 270496
rect 297916 270444 297968 270496
rect 299572 270444 299624 270496
rect 299940 270444 299992 270496
rect 300860 270444 300912 270496
rect 327080 270444 327132 270496
rect 328460 270444 328512 270496
rect 244924 270308 244976 270360
rect 336004 270308 336056 270360
rect 347412 270308 347464 270360
rect 85488 270172 85540 270224
rect 149428 270172 149480 270224
rect 153292 270172 153344 270224
rect 169852 270172 169904 270224
rect 170036 270172 170088 270224
rect 210148 270172 210200 270224
rect 211068 270172 211120 270224
rect 237472 270172 237524 270224
rect 258540 270172 258592 270224
rect 268016 270172 268068 270224
rect 321100 270172 321152 270224
rect 327448 270172 327500 270224
rect 345940 270172 345992 270224
rect 360200 270444 360252 270496
rect 377036 270444 377088 270496
rect 387892 270444 387944 270496
rect 400588 270444 400640 270496
rect 441620 270444 441672 270496
rect 453856 270444 453908 270496
rect 516600 270444 516652 270496
rect 517704 270444 517756 270496
rect 597560 270444 597612 270496
rect 359188 270308 359240 270360
rect 382280 270308 382332 270360
rect 390376 270308 390428 270360
rect 405740 270308 405792 270360
rect 407212 270308 407264 270360
rect 451464 270308 451516 270360
rect 456432 270308 456484 270360
rect 520280 270308 520332 270360
rect 523132 270308 523184 270360
rect 605104 270308 605156 270360
rect 360200 270172 360252 270224
rect 383660 270172 383712 270224
rect 388168 270172 388220 270224
rect 410064 270172 410116 270224
rect 410800 270172 410852 270224
rect 455420 270172 455472 270224
rect 461400 270172 461452 270224
rect 527180 270172 527232 270224
rect 528100 270172 528152 270224
rect 619180 270172 619232 270224
rect 309784 270104 309836 270156
rect 311348 270104 311400 270156
rect 67548 270036 67600 270088
rect 75920 270036 75972 270088
rect 80060 270036 80112 270088
rect 146392 270036 146444 270088
rect 158628 270036 158680 270088
rect 201040 270036 201092 270088
rect 202236 270036 202288 270088
rect 230848 270036 230900 270088
rect 233700 270036 233752 270088
rect 242716 270036 242768 270088
rect 245476 270036 245528 270088
rect 263140 270036 263192 270088
rect 266820 270036 266872 270088
rect 274640 270036 274692 270088
rect 316960 270036 317012 270088
rect 321560 270036 321612 270088
rect 323584 270036 323636 270088
rect 331220 270036 331272 270088
rect 346768 270036 346820 270088
rect 364340 270036 364392 270088
rect 364984 270036 365036 270088
rect 390560 270036 390612 270088
rect 409696 270036 409748 270088
rect 454040 270036 454092 270088
rect 455052 270036 455104 270088
rect 473360 270036 473412 270088
rect 525616 270036 525668 270088
rect 619640 270036 619692 270088
rect 77208 269900 77260 269952
rect 143908 269900 143960 269952
rect 144092 269900 144144 269952
rect 190828 269900 190880 269952
rect 201776 269900 201828 269952
rect 232504 269900 232556 269952
rect 234804 269900 234856 269952
rect 255688 269900 255740 269952
rect 262036 269900 262088 269952
rect 272524 269900 272576 269952
rect 273076 269900 273128 269952
rect 282184 269900 282236 269952
rect 285772 269900 285824 269952
rect 291292 269900 291344 269952
rect 329380 269900 329432 269952
rect 339500 269900 339552 269952
rect 341800 269900 341852 269952
rect 357440 269900 357492 269952
rect 364156 269900 364208 269952
rect 389180 269900 389232 269952
rect 390192 269900 390244 269952
rect 412640 269900 412692 269952
rect 414664 269900 414716 269952
rect 460940 269900 460992 269952
rect 463516 269900 463568 269952
rect 531320 269900 531372 269952
rect 531688 269900 531740 269952
rect 627920 269900 627972 269952
rect 69388 269764 69440 269816
rect 139768 269764 139820 269816
rect 140688 269764 140740 269816
rect 188620 269764 188672 269816
rect 194600 269764 194652 269816
rect 227260 269764 227312 269816
rect 119068 269628 119120 269680
rect 173348 269628 173400 269680
rect 174360 269628 174412 269680
rect 210976 269628 211028 269680
rect 226616 269628 226668 269680
rect 249892 269764 249944 269816
rect 250260 269764 250312 269816
rect 266452 269764 266504 269816
rect 268200 269764 268252 269816
rect 278872 269764 278924 269816
rect 314476 269764 314528 269816
rect 318984 269764 319036 269816
rect 326896 269764 326948 269816
rect 335544 269764 335596 269816
rect 336924 269764 336976 269816
rect 350540 269764 350592 269816
rect 351736 269764 351788 269816
rect 371240 269764 371292 269816
rect 374920 269764 374972 269816
rect 404360 269764 404412 269816
rect 412456 269764 412508 269816
rect 458180 269764 458232 269816
rect 458548 269764 458600 269816
rect 524420 269764 524472 269816
rect 535552 269764 535604 269816
rect 633532 269764 633584 269816
rect 387432 269628 387484 269680
rect 401692 269628 401744 269680
rect 401876 269628 401928 269680
rect 419724 269628 419776 269680
rect 422116 269628 422168 269680
rect 472164 269628 472216 269680
rect 474648 269628 474700 269680
rect 546500 269628 546552 269680
rect 126888 269492 126940 269544
rect 178684 269492 178736 269544
rect 183468 269492 183520 269544
rect 204168 269492 204220 269544
rect 383660 269492 383712 269544
rect 391940 269492 391992 269544
rect 392124 269492 392176 269544
rect 409880 269492 409932 269544
rect 424600 269492 424652 269544
rect 476120 269492 476172 269544
rect 476764 269492 476816 269544
rect 549904 269492 549956 269544
rect 136088 269356 136140 269408
rect 180892 269356 180944 269408
rect 419816 269356 419868 269408
rect 465080 269356 465132 269408
rect 507860 269356 507912 269408
rect 560300 269356 560352 269408
rect 251456 269220 251508 269272
rect 258080 269220 258132 269272
rect 294052 269220 294104 269272
rect 297088 269220 297140 269272
rect 441620 269220 441672 269272
rect 462320 269220 462372 269272
rect 466000 269220 466052 269272
rect 534172 269220 534224 269272
rect 146944 269152 146996 269204
rect 153844 269152 153896 269204
rect 282828 269084 282880 269136
rect 288808 269084 288860 269136
rect 295340 269084 295392 269136
rect 297916 269084 297968 269136
rect 319444 269084 319496 269136
rect 325700 269084 325752 269136
rect 331864 269084 331916 269136
rect 338028 269084 338080 269136
rect 342260 269084 342312 269136
rect 345112 269084 345164 269136
rect 115848 269016 115900 269068
rect 171232 269016 171284 269068
rect 413008 269016 413060 269068
rect 459744 269016 459796 269068
rect 469220 269016 469272 269068
rect 495440 269016 495492 269068
rect 495808 269016 495860 269068
rect 576860 269016 576912 269068
rect 108948 268880 109000 268932
rect 166264 268880 166316 268932
rect 172428 268880 172480 268932
rect 204352 268880 204404 268932
rect 208400 268880 208452 268932
rect 214288 268880 214340 268932
rect 428740 268880 428792 268932
rect 478972 268880 479024 268932
rect 498292 268880 498344 268932
rect 581000 268880 581052 268932
rect 582196 268880 582248 268932
rect 600412 268880 600464 268932
rect 99288 268744 99340 268796
rect 91008 268608 91060 268660
rect 99288 268608 99340 268660
rect 110236 268744 110288 268796
rect 167920 268744 167972 268796
rect 173808 268744 173860 268796
rect 212632 268744 212684 268796
rect 215208 268744 215260 268796
rect 223488 268744 223540 268796
rect 227720 268744 227772 268796
rect 250720 268744 250772 268796
rect 372344 268744 372396 268796
rect 397092 268744 397144 268796
rect 398748 268744 398800 268796
rect 422300 268744 422352 268796
rect 433708 268744 433760 268796
rect 488540 268744 488592 268796
rect 500684 268744 500736 268796
rect 584128 268744 584180 268796
rect 160468 268608 160520 268660
rect 168656 268608 168708 268660
rect 208492 268608 208544 268660
rect 212264 268608 212316 268660
rect 238300 268608 238352 268660
rect 256700 268608 256752 268660
rect 263968 268608 264020 268660
rect 326068 268608 326120 268660
rect 328276 268608 328328 268660
rect 355876 268608 355928 268660
rect 367836 268608 367888 268660
rect 382372 268608 382424 268660
rect 415400 268608 415452 268660
rect 416688 268608 416740 268660
rect 433340 268608 433392 268660
rect 436192 268608 436244 268660
rect 491852 268608 491904 268660
rect 92388 268472 92440 268524
rect 155500 268472 155552 268524
rect 160008 268472 160060 268524
rect 200396 268472 200448 268524
rect 208216 268472 208268 268524
rect 236644 268472 236696 268524
rect 241428 268472 241480 268524
rect 256700 268472 256752 268524
rect 269120 268472 269172 268524
rect 279700 268472 279752 268524
rect 343364 268472 343416 268524
rect 357256 268472 357308 268524
rect 357532 268472 357584 268524
rect 379520 268472 379572 268524
rect 393136 268472 393188 268524
rect 430580 268472 430632 268524
rect 441160 268472 441212 268524
rect 498476 268608 498528 268660
rect 503260 268608 503312 268660
rect 587900 268608 587952 268660
rect 492220 268472 492272 268524
rect 87144 268336 87196 268388
rect 152188 268336 152240 268388
rect 152740 268336 152792 268388
rect 196072 268336 196124 268388
rect 200580 268336 200632 268388
rect 231676 268336 231728 268388
rect 238668 268336 238720 268388
rect 256148 268336 256200 268388
rect 256516 268336 256568 268388
rect 270592 268336 270644 268388
rect 327724 268336 327776 268388
rect 336740 268336 336792 268388
rect 337660 268336 337712 268388
rect 352104 268336 352156 268388
rect 352564 268336 352616 268388
rect 368848 268336 368900 268388
rect 369952 268336 370004 268388
rect 397460 268336 397512 268388
rect 399760 268336 399812 268388
rect 440240 268336 440292 268388
rect 443644 268336 443696 268388
rect 502340 268336 502392 268388
rect 510712 268472 510764 268524
rect 598940 268472 598992 268524
rect 517888 268336 517940 268388
rect 534724 268336 534776 268388
rect 535736 268336 535788 268388
rect 536380 268336 536432 268388
rect 634820 268336 634872 268388
rect 118608 268200 118660 268252
rect 174544 268200 174596 268252
rect 429568 268200 429620 268252
rect 469404 268200 469456 268252
rect 137008 268064 137060 268116
rect 183008 268064 183060 268116
rect 422300 268064 422352 268116
rect 443276 268064 443328 268116
rect 459560 268064 459612 268116
rect 492128 268200 492180 268252
rect 492312 268200 492364 268252
rect 569960 268200 570012 268252
rect 489184 267928 489236 267980
rect 567384 268064 567436 268116
rect 490840 267928 490892 267980
rect 492312 267928 492364 267980
rect 493324 267928 493376 267980
rect 551560 267928 551612 267980
rect 132408 267656 132460 267708
rect 99288 267520 99340 267572
rect 154672 267520 154724 267572
rect 160744 267520 160796 267572
rect 164608 267520 164660 267572
rect 166448 267520 166500 267572
rect 172888 267520 172940 267572
rect 184204 267656 184256 267708
rect 193128 267792 193180 267844
rect 448612 267792 448664 267844
rect 506480 267792 506532 267844
rect 193128 267656 193180 267708
rect 204168 267656 204220 267708
rect 218428 267656 218480 267708
rect 218796 267656 218848 267708
rect 222568 267656 222620 267708
rect 377772 267656 377824 267708
rect 385684 267656 385736 267708
rect 387248 267656 387300 267708
rect 398748 267656 398800 267708
rect 404728 267656 404780 267708
rect 429844 267656 429896 267708
rect 436744 267656 436796 267708
rect 441620 267656 441672 267708
rect 442724 267656 442776 267708
rect 483664 267656 483716 267708
rect 483848 267656 483900 267708
rect 184480 267520 184532 267572
rect 186964 267520 187016 267572
rect 107660 267384 107712 267436
rect 167092 267384 167144 267436
rect 167644 267384 167696 267436
rect 186964 267384 187016 267436
rect 189908 267384 189960 267436
rect 192760 267384 192812 267436
rect 216772 267520 216824 267572
rect 217416 267520 217468 267572
rect 223028 267520 223080 267572
rect 224224 267520 224276 267572
rect 229192 267520 229244 267572
rect 373264 267520 373316 267572
rect 387432 267520 387484 267572
rect 402244 267520 402296 267572
rect 422300 267520 422352 267572
rect 430396 267520 430448 267572
rect 457444 267520 457496 267572
rect 462688 267520 462740 267572
rect 468944 267520 468996 267572
rect 475108 267520 475160 267572
rect 479708 267520 479760 267572
rect 484032 267520 484084 267572
rect 487804 267520 487856 267572
rect 490012 267656 490064 267708
rect 497280 267656 497332 267708
rect 499672 267656 499724 267708
rect 526444 267656 526496 267708
rect 527272 267656 527324 267708
rect 592684 267656 592736 267708
rect 507860 267520 507912 267572
rect 508228 267520 508280 267572
rect 522396 267520 522448 267572
rect 523684 267520 523736 267572
rect 530676 267520 530728 267572
rect 532240 267520 532292 267572
rect 596824 267520 596876 267572
rect 221740 267384 221792 267436
rect 232688 267384 232740 267436
rect 239128 267384 239180 267436
rect 261484 267384 261536 267436
rect 268936 267384 268988 267436
rect 340972 267384 341024 267436
rect 347044 267384 347096 267436
rect 350908 267384 350960 267436
rect 359464 267384 359516 267436
rect 361120 267384 361172 267436
rect 373080 267384 373132 267436
rect 375748 267384 375800 267436
rect 390376 267384 390428 267436
rect 390652 267384 390704 267436
rect 395528 267384 395580 267436
rect 397092 267384 397144 267436
rect 421564 267384 421616 267436
rect 436560 267384 436612 267436
rect 445024 267384 445076 267436
rect 450268 267384 450320 267436
rect 505836 267384 505888 267436
rect 507400 267384 507452 267436
rect 576124 267384 576176 267436
rect 95884 267248 95936 267300
rect 157156 267248 157208 267300
rect 170404 267248 170456 267300
rect 86224 267112 86276 267164
rect 148048 267112 148100 267164
rect 149704 267112 149756 267164
rect 194416 267112 194468 267164
rect 198188 267112 198240 267164
rect 200212 267112 200264 267164
rect 206284 267248 206336 267300
rect 213460 267248 213512 267300
rect 215944 267248 215996 267300
rect 220084 267248 220136 267300
rect 220268 267248 220320 267300
rect 234160 267248 234212 267300
rect 236828 267248 236880 267300
rect 251548 267248 251600 267300
rect 286324 267248 286376 267300
rect 287980 267248 288032 267300
rect 313648 267248 313700 267300
rect 317420 267248 317472 267300
rect 335176 267248 335228 267300
rect 341524 267248 341576 267300
rect 363328 267248 363380 267300
rect 377036 267248 377088 267300
rect 394792 267248 394844 267300
rect 416688 267248 416740 267300
rect 419632 267248 419684 267300
rect 446588 267248 446640 267300
rect 455236 267248 455288 267300
rect 507860 267248 507912 267300
rect 509884 267248 509936 267300
rect 517704 267248 517756 267300
rect 206836 267112 206888 267164
rect 207020 267112 207072 267164
rect 220912 267112 220964 267164
rect 223488 267112 223540 267164
rect 241612 267112 241664 267164
rect 242716 267112 242768 267164
rect 254860 267112 254912 267164
rect 267004 267112 267056 267164
rect 273076 267112 273128 267164
rect 276020 267112 276072 267164
rect 283840 267112 283892 267164
rect 324412 267112 324464 267164
rect 330484 267112 330536 267164
rect 334348 267112 334400 267164
rect 344284 267112 344336 267164
rect 353392 267112 353444 267164
rect 363604 267112 363656 267164
rect 365812 267112 365864 267164
rect 73804 266976 73856 267028
rect 141424 266976 141476 267028
rect 146944 266976 146996 267028
rect 189448 266976 189500 267028
rect 191012 266976 191064 267028
rect 211804 266976 211856 267028
rect 222016 266976 222068 267028
rect 246580 266976 246632 267028
rect 249064 266976 249116 267028
rect 261484 266976 261536 267028
rect 264980 266976 265032 267028
rect 276388 266976 276440 267028
rect 278044 266976 278096 267028
rect 284668 266976 284720 267028
rect 333520 266976 333572 267028
rect 342260 266976 342312 267028
rect 368112 266976 368164 267028
rect 377772 266976 377824 267028
rect 119804 266840 119856 266892
rect 161756 266840 161808 266892
rect 169852 266840 169904 266892
rect 199108 266840 199160 266892
rect 199292 266840 199344 266892
rect 201868 266840 201920 266892
rect 243544 266840 243596 266892
rect 249064 266840 249116 266892
rect 254584 266840 254636 266892
rect 259000 266840 259052 266892
rect 274640 266840 274692 266892
rect 278044 266840 278096 266892
rect 317788 266840 317840 266892
rect 322940 266840 322992 266892
rect 349252 266840 349304 266892
rect 355324 266840 355376 266892
rect 356704 266840 356756 266892
rect 366364 266840 366416 266892
rect 132592 266704 132644 266756
rect 147220 266704 147272 266756
rect 148508 266704 148560 266756
rect 179512 266704 179564 266756
rect 201592 266704 201644 266756
rect 207020 266704 207072 266756
rect 321928 266704 321980 266756
rect 327080 266704 327132 266756
rect 385684 267112 385736 267164
rect 401876 267112 401928 267164
rect 415492 267112 415544 267164
rect 436744 267112 436796 267164
rect 445300 267112 445352 267164
rect 450728 267112 450780 267164
rect 452568 267112 452620 267164
rect 456064 267112 456116 267164
rect 378968 266976 379020 267028
rect 392124 266976 392176 267028
rect 392308 266976 392360 267028
rect 418804 266976 418856 267028
rect 422944 266976 422996 267028
rect 455052 266976 455104 267028
rect 455420 266976 455472 267028
rect 459560 266976 459612 267028
rect 380624 266840 380676 266892
rect 390192 266840 390244 266892
rect 405556 266840 405608 266892
rect 425704 266840 425756 266892
rect 426072 266840 426124 266892
rect 436560 266840 436612 266892
rect 438676 266840 438728 266892
rect 469128 267112 469180 267164
rect 469312 267112 469364 267164
rect 470508 267112 470560 267164
rect 473268 267112 473320 267164
rect 512184 267112 512236 267164
rect 512368 267112 512420 267164
rect 582196 267248 582248 267300
rect 520648 267112 520700 267164
rect 524236 267112 524288 267164
rect 383660 266704 383712 266756
rect 398104 266704 398156 266756
rect 414480 266704 414532 266756
rect 423772 266704 423824 266756
rect 424968 266704 425020 266756
rect 425428 266704 425480 266756
rect 426256 266704 426308 266756
rect 427912 266704 427964 266756
rect 428924 266704 428976 266756
rect 437848 266704 437900 266756
rect 468484 266976 468536 267028
rect 468944 266976 468996 267028
rect 484032 266976 484084 267028
rect 465172 266840 465224 266892
rect 466828 266704 466880 266756
rect 467748 266704 467800 266756
rect 470140 266840 470192 266892
rect 523684 266976 523736 267028
rect 615500 267112 615552 267164
rect 487528 266840 487580 266892
rect 514024 266840 514076 266892
rect 514392 266840 514444 266892
rect 517520 266840 517572 266892
rect 518992 266840 519044 266892
rect 520096 266840 520148 266892
rect 522304 266840 522356 266892
rect 524236 266840 524288 266892
rect 528928 266840 528980 266892
rect 529756 266840 529808 266892
rect 537208 266976 537260 267028
rect 636200 266976 636252 267028
rect 537484 266840 537536 266892
rect 540980 266840 541032 266892
rect 541624 266840 541676 266892
rect 541900 266840 541952 266892
rect 602344 266840 602396 266892
rect 473268 266704 473320 266756
rect 473452 266704 473504 266756
rect 474372 266704 474424 266756
rect 477592 266704 477644 266756
rect 478604 266704 478656 266756
rect 483388 266704 483440 266756
rect 484308 266704 484360 266756
rect 485872 266704 485924 266756
rect 487068 266704 487120 266756
rect 494980 266704 495032 266756
rect 499672 266704 499724 266756
rect 499856 266704 499908 266756
rect 501604 266704 501656 266756
rect 502432 266704 502484 266756
rect 559748 266704 559800 266756
rect 258080 266636 258132 266688
rect 267280 266636 267332 266688
rect 312820 266636 312872 266688
rect 316408 266636 316460 266688
rect 389824 266636 389876 266688
rect 395344 266636 395396 266688
rect 123484 266568 123536 266620
rect 150532 266568 150584 266620
rect 154028 266568 154080 266620
rect 170404 266568 170456 266620
rect 416320 266568 416372 266620
rect 438124 266568 438176 266620
rect 446956 266568 447008 266620
rect 452568 266568 452620 266620
rect 452752 266568 452804 266620
rect 453672 266568 453724 266620
rect 454408 266568 454460 266620
rect 455420 266568 455472 266620
rect 456892 266568 456944 266620
rect 457996 266568 458048 266620
rect 460204 266568 460256 266620
rect 490564 266568 490616 266620
rect 491668 266568 491720 266620
rect 492588 266568 492640 266620
rect 494152 266568 494204 266620
rect 495256 266568 495308 266620
rect 497464 266568 497516 266620
rect 552664 266568 552716 266620
rect 222844 266500 222896 266552
rect 226708 266500 226760 266552
rect 253204 266500 253256 266552
rect 256516 266500 256568 266552
rect 256700 266500 256752 266552
rect 259828 266500 259880 266552
rect 308680 266500 308732 266552
rect 310888 266500 310940 266552
rect 311164 266500 311216 266552
rect 313280 266500 313332 266552
rect 320272 266500 320324 266552
rect 324964 266500 325016 266552
rect 330208 266500 330260 266552
rect 334624 266500 334676 266552
rect 345112 266500 345164 266552
rect 351184 266500 351236 266552
rect 395620 266500 395672 266552
rect 405004 266500 405056 266552
rect 141608 266432 141660 266484
rect 146944 266432 146996 266484
rect 421288 266432 421340 266484
rect 156604 266364 156656 266416
rect 159640 266364 159692 266416
rect 162124 266364 162176 266416
rect 162952 266364 163004 266416
rect 165068 266364 165120 266416
rect 169576 266364 169628 266416
rect 181536 266364 181588 266416
rect 182824 266364 182876 266416
rect 183008 266364 183060 266416
rect 186136 266364 186188 266416
rect 192484 266364 192536 266416
rect 197728 266364 197780 266416
rect 200396 266364 200448 266416
rect 202696 266364 202748 266416
rect 213184 266364 213236 266416
rect 215944 266364 215996 266416
rect 221464 266364 221516 266416
rect 224224 266364 224276 266416
rect 239496 266364 239548 266416
rect 244096 266364 244148 266416
rect 256148 266364 256200 266416
rect 258172 266364 258224 266416
rect 268016 266364 268068 266416
rect 272248 266364 272300 266416
rect 272524 266364 272576 266416
rect 274732 266364 274784 266416
rect 287704 266364 287756 266416
rect 292120 266364 292172 266416
rect 301044 266364 301096 266416
rect 302056 266364 302108 266416
rect 307852 266364 307904 266416
rect 309508 266364 309560 266416
rect 310336 266364 310388 266416
rect 311900 266364 311952 266416
rect 312360 266364 312412 266416
rect 314660 266364 314712 266416
rect 316132 266364 316184 266416
rect 320548 266364 320600 266416
rect 328552 266364 328604 266416
rect 329748 266364 329800 266416
rect 332692 266364 332744 266416
rect 333796 266364 333848 266416
rect 342628 266364 342680 266416
rect 343548 266364 343600 266416
rect 347596 266364 347648 266416
rect 349804 266364 349856 266416
rect 355048 266364 355100 266416
rect 356888 266364 356940 266416
rect 358360 266364 358412 266416
rect 360844 266364 360896 266416
rect 361672 266364 361724 266416
rect 362868 266364 362920 266416
rect 367468 266364 367520 266416
rect 368296 266364 368348 266416
rect 371608 266364 371660 266416
rect 372528 266364 372580 266416
rect 374092 266364 374144 266416
rect 375288 266364 375340 266416
rect 377404 266364 377456 266416
rect 378784 266364 378836 266416
rect 379888 266364 379940 266416
rect 380808 266364 380860 266416
rect 384028 266364 384080 266416
rect 384948 266364 385000 266416
rect 386512 266364 386564 266416
rect 387616 266364 387668 266416
rect 396448 266364 396500 266416
rect 397276 266364 397328 266416
rect 398932 266364 398984 266416
rect 400128 266364 400180 266416
rect 403072 266364 403124 266416
rect 404176 266364 404228 266416
rect 411352 266364 411404 266416
rect 412272 266364 412324 266416
rect 417148 266364 417200 266416
rect 419816 266364 419868 266416
rect 450728 266432 450780 266484
rect 499764 266432 499816 266484
rect 499948 266432 500000 266484
rect 500868 266432 500920 266484
rect 504088 266432 504140 266484
rect 504916 266432 504968 266484
rect 506572 266432 506624 266484
rect 507676 266432 507728 266484
rect 507860 266432 507912 266484
rect 510068 266432 510120 266484
rect 514852 266432 514904 266484
rect 516048 266432 516100 266484
rect 516508 266432 516560 266484
rect 517336 266432 517388 266484
rect 517520 266432 517572 266484
rect 540980 266432 541032 266484
rect 541348 266432 541400 266484
rect 542084 266432 542136 266484
rect 432052 266364 432104 266416
rect 433156 266364 433208 266416
rect 439320 266364 439372 266416
rect 440332 266364 440384 266416
rect 441344 266364 441396 266416
rect 441988 266364 442040 266416
rect 442908 266364 442960 266416
rect 444472 266364 444524 266416
rect 445668 266364 445720 266416
rect 446128 266364 446180 266416
rect 447784 266364 447836 266416
rect 448152 266364 448204 266416
rect 450544 266364 450596 266416
rect 480076 266296 480128 266348
rect 554780 266296 554832 266348
rect 485044 266160 485096 266212
rect 561680 266160 561732 266212
rect 486700 266024 486752 266076
rect 564440 266024 564492 266076
rect 142160 265888 142212 265940
rect 142804 265888 142856 265940
rect 234620 265888 234672 265940
rect 235540 265888 235592 265940
rect 292764 265888 292816 265940
rect 293500 265888 293552 265940
rect 492496 265888 492548 265940
rect 572720 265888 572772 265940
rect 515680 265752 515732 265804
rect 605840 265752 605892 265804
rect 518164 265616 518216 265668
rect 608692 265616 608744 265668
rect 481732 265480 481784 265532
rect 557540 265480 557592 265532
rect 479248 265344 479300 265396
rect 553400 265344 553452 265396
rect 577504 261604 577556 261656
rect 648620 261604 648672 261656
rect 570604 261468 570656 261520
rect 645860 261468 645912 261520
rect 554412 260856 554464 260908
rect 568580 260856 568632 260908
rect 675852 260176 675904 260228
rect 676404 260176 676456 260228
rect 554320 259428 554372 259480
rect 560944 259428 560996 259480
rect 553952 256708 554004 256760
rect 559564 256708 559616 256760
rect 35808 252696 35860 252748
rect 41696 252696 41748 252748
rect 35624 252560 35676 252612
rect 40684 252560 40736 252612
rect 554412 252560 554464 252612
rect 562324 252560 562376 252612
rect 675852 252220 675904 252272
rect 678244 252220 678296 252272
rect 35808 251200 35860 251252
rect 37924 251200 37976 251252
rect 554136 251200 554188 251252
rect 556804 251200 556856 251252
rect 675484 251200 675536 251252
rect 675484 250928 675536 250980
rect 553492 249024 553544 249076
rect 571340 249024 571392 249076
rect 553860 246304 553912 246356
rect 632704 246304 632756 246356
rect 554412 245624 554464 245676
rect 592684 245624 592736 245676
rect 553400 244264 553452 244316
rect 555424 244264 555476 244316
rect 37924 242836 37976 242888
rect 41696 242836 41748 242888
rect 34428 242156 34480 242208
rect 41696 242156 41748 242208
rect 558184 242156 558236 242208
rect 647240 242156 647292 242208
rect 553952 241476 554004 241528
rect 621664 241476 621716 241528
rect 554320 238688 554372 238740
rect 577504 238688 577556 238740
rect 671068 237804 671120 237856
rect 671712 237532 671764 237584
rect 668768 237396 668820 237448
rect 671344 237124 671396 237176
rect 671528 236988 671580 237040
rect 673092 236716 673144 236768
rect 673414 236852 673466 236904
rect 673528 236852 673580 236904
rect 672540 236444 672592 236496
rect 673752 236240 673804 236292
rect 673460 236104 673512 236156
rect 554504 236036 554556 236088
rect 558184 236036 558236 236088
rect 673460 235900 673512 235952
rect 674088 235628 674140 235680
rect 673368 235492 673420 235544
rect 674104 235084 674156 235136
rect 672540 234948 672592 235000
rect 554412 234540 554464 234592
rect 570604 234540 570656 234592
rect 668124 234540 668176 234592
rect 674196 234812 674248 234864
rect 674536 234948 674588 235000
rect 669596 234336 669648 234388
rect 675852 234336 675904 234388
rect 681004 234336 681056 234388
rect 673828 234200 673880 234252
rect 671712 233996 671764 234048
rect 670976 233860 671028 233912
rect 674748 233860 674800 233912
rect 675096 233860 675148 233912
rect 675236 233860 675288 233912
rect 672954 233656 673006 233708
rect 674840 233656 674892 233708
rect 675852 233724 675904 233776
rect 675116 233588 675168 233640
rect 675852 233588 675904 233640
rect 677692 233588 677744 233640
rect 670792 233316 670844 233368
rect 675852 233452 675904 233504
rect 676036 233316 676088 233368
rect 677876 233316 677928 233368
rect 683120 233384 683172 233436
rect 684500 233248 684552 233300
rect 673000 233180 673052 233232
rect 673948 233180 674000 233232
rect 669044 232976 669096 233028
rect 670240 232976 670292 233028
rect 669780 232840 669832 232892
rect 673368 232840 673420 232892
rect 661868 232500 661920 232552
rect 675852 232500 675904 232552
rect 683488 232500 683540 232552
rect 675484 232432 675536 232484
rect 665088 232160 665140 232212
rect 673460 231956 673512 232008
rect 675180 231684 675232 231736
rect 674172 231616 674224 231668
rect 674472 231616 674524 231668
rect 675070 231480 675122 231532
rect 662236 231072 662288 231124
rect 673460 231276 673512 231328
rect 674956 231276 675008 231328
rect 667940 231140 667992 231192
rect 675852 231072 675904 231124
rect 678612 231072 678664 231124
rect 129648 230868 129700 230920
rect 199108 230868 199160 230920
rect 674732 230868 674784 230920
rect 104808 230732 104860 230784
rect 179144 230732 179196 230784
rect 97908 230596 97960 230648
rect 173992 230596 174044 230648
rect 91008 230460 91060 230512
rect 168840 230460 168892 230512
rect 511816 230460 511868 230512
rect 196072 230392 196124 230444
rect 198464 230392 198516 230444
rect 207664 230392 207716 230444
rect 251272 230392 251324 230444
rect 256608 230392 256660 230444
rect 297640 230392 297692 230444
rect 311900 230392 311952 230444
rect 340144 230392 340196 230444
rect 441896 230392 441948 230444
rect 443552 230392 443604 230444
rect 444472 230392 444524 230444
rect 447600 230392 447652 230444
rect 476120 230392 476172 230444
rect 478604 230392 478656 230444
rect 387432 230324 387484 230376
rect 388444 230324 388496 230376
rect 439320 230324 439372 230376
rect 440332 230324 440384 230376
rect 449624 230324 449676 230376
rect 450544 230324 450596 230376
rect 451556 230324 451608 230376
rect 453304 230324 453356 230376
rect 455420 230324 455472 230376
rect 457168 230324 457220 230376
rect 463792 230324 463844 230376
rect 465724 230324 465776 230376
rect 481824 230324 481876 230376
rect 486516 230324 486568 230376
rect 503720 230324 503772 230376
rect 507124 230324 507176 230376
rect 510804 230324 510856 230376
rect 511816 230324 511868 230376
rect 133696 230256 133748 230308
rect 202328 230256 202380 230308
rect 126888 230120 126940 230172
rect 197176 230120 197228 230172
rect 197452 230120 197504 230172
rect 201040 230120 201092 230172
rect 202144 230120 202196 230172
rect 240968 230256 241020 230308
rect 242532 230256 242584 230308
rect 287336 230256 287388 230308
rect 305644 230256 305696 230308
rect 334992 230256 335044 230308
rect 376024 230256 376076 230308
rect 380716 230256 380768 230308
rect 531136 230460 531188 230512
rect 526904 230392 526956 230444
rect 520464 230324 520516 230376
rect 521568 230324 521620 230376
rect 518900 230256 518952 230308
rect 413836 230188 413888 230240
rect 420000 230188 420052 230240
rect 443828 230188 443880 230240
rect 444656 230188 444708 230240
rect 452844 230188 452896 230240
rect 454316 230188 454368 230240
rect 465448 230188 465500 230240
rect 469404 230188 469456 230240
rect 477960 230188 478012 230240
rect 478788 230188 478840 230240
rect 499856 230188 499908 230240
rect 504364 230188 504416 230240
rect 530124 230324 530176 230376
rect 531228 230324 531280 230376
rect 674472 230800 674524 230852
rect 674610 230664 674662 230716
rect 674396 230596 674448 230648
rect 534816 230188 534868 230240
rect 230480 230120 230532 230172
rect 277032 230120 277084 230172
rect 294604 230120 294656 230172
rect 323400 230120 323452 230172
rect 323584 230120 323636 230172
rect 324688 230120 324740 230172
rect 354864 230120 354916 230172
rect 371056 230120 371108 230172
rect 505652 230120 505704 230172
rect 513840 230120 513892 230172
rect 515312 230120 515364 230172
rect 525156 230120 525208 230172
rect 535460 230256 535512 230308
rect 539600 230256 539652 230308
rect 668124 230256 668176 230308
rect 673828 230256 673880 230308
rect 674396 230256 674448 230308
rect 543648 230120 543700 230172
rect 454132 230052 454184 230104
rect 455328 230052 455380 230104
rect 86224 229984 86276 230036
rect 155960 229984 156012 230036
rect 160192 229984 160244 230036
rect 220360 229984 220412 230036
rect 224960 229984 225012 230036
rect 271880 229984 271932 230036
rect 300124 229984 300176 230036
rect 329840 229984 329892 230036
rect 337844 229984 337896 230036
rect 360752 229984 360804 230036
rect 457352 229984 457404 230036
rect 464068 229984 464120 230036
rect 476672 229984 476724 230036
rect 480720 229984 480772 230036
rect 501788 229984 501840 230036
rect 509884 229984 509936 230036
rect 519176 229984 519228 230036
rect 528560 229984 528612 230036
rect 534632 229984 534684 230036
rect 552756 229984 552808 230036
rect 559564 229984 559616 230036
rect 567200 229984 567252 230036
rect 672156 229984 672208 230036
rect 672540 229984 672592 230036
rect 673276 229984 673328 230036
rect 675852 229984 675904 230036
rect 676496 229984 676548 230036
rect 453488 229916 453540 229968
rect 455788 229916 455840 229968
rect 117228 229848 117280 229900
rect 189448 229848 189500 229900
rect 189724 229848 189776 229900
rect 235816 229848 235868 229900
rect 283564 229848 283616 229900
rect 318248 229848 318300 229900
rect 324964 229848 325016 229900
rect 350448 229848 350500 229900
rect 361212 229848 361264 229900
rect 378784 229848 378836 229900
rect 389916 229848 389968 229900
rect 399392 229848 399444 229900
rect 410800 229848 410852 229900
rect 417424 229848 417476 229900
rect 479248 229848 479300 229900
rect 490564 229848 490616 229900
rect 494060 229848 494112 229900
rect 506112 229848 506164 229900
rect 517244 229848 517296 229900
rect 525984 229848 526036 229900
rect 528836 229848 528888 229900
rect 535460 229848 535512 229900
rect 536564 229848 536616 229900
rect 559748 229848 559800 229900
rect 433524 229780 433576 229832
rect 434168 229780 434220 229832
rect 438676 229780 438728 229832
rect 439320 229780 439372 229832
rect 673828 229780 673880 229832
rect 110328 229712 110380 229764
rect 184296 229712 184348 229764
rect 184480 229712 184532 229764
rect 225512 229712 225564 229764
rect 270132 229712 270184 229764
rect 307944 229712 307996 229764
rect 318064 229712 318116 229764
rect 345296 229712 345348 229764
rect 345664 229712 345716 229764
rect 355600 229712 355652 229764
rect 357072 229712 357124 229764
rect 376208 229712 376260 229764
rect 380716 229712 380768 229764
rect 394240 229712 394292 229764
rect 399852 229712 399904 229764
rect 409696 229712 409748 229764
rect 469588 229712 469640 229764
rect 476764 229712 476816 229764
rect 484768 229712 484820 229764
rect 496820 229712 496872 229764
rect 507584 229712 507636 229764
rect 516784 229712 516836 229764
rect 523040 229712 523092 229764
rect 534632 229712 534684 229764
rect 538496 229712 538548 229764
rect 565084 229712 565136 229764
rect 95240 229576 95292 229628
rect 161112 229576 161164 229628
rect 161296 229576 161348 229628
rect 217784 229576 217836 229628
rect 251732 229576 251784 229628
rect 292488 229576 292540 229628
rect 490196 229576 490248 229628
rect 493968 229576 494020 229628
rect 513656 229576 513708 229628
rect 522488 229576 522540 229628
rect 676036 229576 676088 229628
rect 677416 229576 677468 229628
rect 673948 229508 674000 229560
rect 144184 229440 144236 229492
rect 148876 229440 148928 229492
rect 150440 229440 150492 229492
rect 215208 229440 215260 229492
rect 217324 229440 217376 229492
rect 266728 229440 266780 229492
rect 276664 229440 276716 229492
rect 302792 229440 302844 229492
rect 673460 229440 673512 229492
rect 675852 229440 675904 229492
rect 676680 229440 676732 229492
rect 448980 229372 449032 229424
rect 451372 229372 451424 229424
rect 509516 229372 509568 229424
rect 518164 229372 518216 229424
rect 133880 229304 133932 229356
rect 146300 229304 146352 229356
rect 148692 229304 148744 229356
rect 210056 229304 210108 229356
rect 210424 229304 210476 229356
rect 261300 229304 261352 229356
rect 261484 229304 261536 229356
rect 282184 229304 282236 229356
rect 288716 229304 288768 229356
rect 313096 229304 313148 229356
rect 450268 229236 450320 229288
rect 451832 229236 451884 229288
rect 493416 229236 493468 229288
rect 500224 229236 500276 229288
rect 532700 229236 532752 229288
rect 536748 229236 536800 229288
rect 673460 229236 673512 229288
rect 94504 229168 94556 229220
rect 145656 229168 145708 229220
rect 146208 229168 146260 229220
rect 207480 229168 207532 229220
rect 213092 229168 213144 229220
rect 256424 229168 256476 229220
rect 419632 229100 419684 229152
rect 421932 229100 421984 229152
rect 423496 229100 423548 229152
rect 427728 229100 427780 229152
rect 441252 229100 441304 229152
rect 442080 229100 442132 229152
rect 446404 229100 446456 229152
rect 126428 229032 126480 229084
rect 195244 229032 195296 229084
rect 205272 229032 205324 229084
rect 257068 229032 257120 229084
rect 265624 229032 265676 229084
rect 274456 229032 274508 229084
rect 274640 229032 274692 229084
rect 309232 229032 309284 229084
rect 309692 229032 309744 229084
rect 320824 229032 320876 229084
rect 327724 229032 327776 229084
rect 337568 229032 337620 229084
rect 450912 229100 450964 229152
rect 452752 229100 452804 229152
rect 497924 229100 497976 229152
rect 524972 229100 525024 229152
rect 514852 229032 514904 229084
rect 448520 228964 448572 229016
rect 119804 228896 119856 228948
rect 190092 228896 190144 228948
rect 193128 228896 193180 228948
rect 246764 228896 246816 228948
rect 257804 228896 257856 228948
rect 299572 228896 299624 228948
rect 312912 228896 312964 228948
rect 340788 228896 340840 228948
rect 349988 228896 350040 228948
rect 369124 228896 369176 228948
rect 377956 228896 378008 228948
rect 390376 228896 390428 228948
rect 549536 228896 549588 228948
rect 673598 228896 673650 228948
rect 466000 228828 466052 228880
rect 469864 228828 469916 228880
rect 673368 228828 673420 228880
rect 100668 228760 100720 228812
rect 174636 228760 174688 228812
rect 176476 228760 176528 228812
rect 233884 228760 233936 228812
rect 234528 228760 234580 228812
rect 278320 228760 278372 228812
rect 285588 228760 285640 228812
rect 318892 228760 318944 228812
rect 320824 228760 320876 228812
rect 327264 228760 327316 228812
rect 335084 228760 335136 228812
rect 356888 228760 356940 228812
rect 373816 228760 373868 228812
rect 387156 228760 387208 228812
rect 447048 228760 447100 228812
rect 450176 228760 450228 228812
rect 518532 228760 518584 228812
rect 541256 228760 541308 228812
rect 106188 228624 106240 228676
rect 179788 228624 179840 228676
rect 183468 228624 183520 228676
rect 239036 228624 239088 228676
rect 246304 228624 246356 228676
rect 289268 228624 289320 228676
rect 304908 228624 304960 228676
rect 333704 228624 333756 228676
rect 340144 228624 340196 228676
rect 362684 228624 362736 228676
rect 371056 228624 371108 228676
rect 385224 228624 385276 228676
rect 403992 228624 404044 228676
rect 411076 228624 411128 228676
rect 485044 228624 485096 228676
rect 498844 228624 498896 228676
rect 514024 228624 514076 228676
rect 535736 228624 535788 228676
rect 535920 228624 535972 228676
rect 563060 228624 563112 228676
rect 93768 228488 93820 228540
rect 169484 228488 169536 228540
rect 169944 228488 169996 228540
rect 228732 228488 228784 228540
rect 235724 228488 235776 228540
rect 280252 228488 280304 228540
rect 288348 228488 288400 228540
rect 322756 228488 322808 228540
rect 326804 228488 326856 228540
rect 351092 228488 351144 228540
rect 362592 228488 362644 228540
rect 379428 228488 379480 228540
rect 390192 228488 390244 228540
rect 400036 228488 400088 228540
rect 57244 228352 57296 228404
rect 141148 228352 141200 228404
rect 146024 228352 146076 228404
rect 210700 228352 210752 228404
rect 215024 228352 215076 228404
rect 266084 228352 266136 228404
rect 271788 228352 271840 228404
rect 308588 228352 308640 228404
rect 309048 228352 309100 228404
rect 336280 228352 336332 228404
rect 336648 228352 336700 228404
rect 358820 228352 358872 228404
rect 359924 228352 359976 228404
rect 376852 228352 376904 228404
rect 378968 228352 379020 228404
rect 393596 228352 393648 228404
rect 400036 228352 400088 228404
rect 407764 228488 407816 228540
rect 411076 228488 411128 228540
rect 416136 228488 416188 228540
rect 478972 228488 479024 228540
rect 490748 228488 490800 228540
rect 491484 228488 491536 228540
rect 506480 228488 506532 228540
rect 510160 228488 510212 228540
rect 530952 228488 531004 228540
rect 531412 228488 531464 228540
rect 558368 228488 558420 228540
rect 673388 228488 673440 228540
rect 409604 228352 409656 228404
rect 415492 228352 415544 228404
rect 470232 228352 470284 228404
rect 479524 228352 479576 228404
rect 486976 228352 487028 228404
rect 501328 228352 501380 228404
rect 502432 228352 502484 228404
rect 521292 228352 521344 228404
rect 521752 228352 521804 228404
rect 545764 228352 545816 228404
rect 554044 228352 554096 228404
rect 581644 228352 581696 228404
rect 673276 228284 673328 228336
rect 133604 228216 133656 228268
rect 200396 228216 200448 228268
rect 210884 228216 210936 228268
rect 260288 228216 260340 228268
rect 398748 228216 398800 228268
rect 409052 228216 409104 228268
rect 139308 228080 139360 228132
rect 205548 228080 205600 228132
rect 222016 228080 222068 228132
rect 269948 228080 270000 228132
rect 140504 227944 140556 227996
rect 146208 227944 146260 227996
rect 152924 227944 152976 227996
rect 215852 227944 215904 227996
rect 252284 227944 252336 227996
rect 293132 227944 293184 227996
rect 671160 227944 671212 227996
rect 673046 228080 673098 228132
rect 393964 227876 394016 227928
rect 401324 227876 401376 227928
rect 402244 227876 402296 227928
rect 143172 227808 143224 227860
rect 148692 227808 148744 227860
rect 169484 227808 169536 227860
rect 169944 227808 169996 227860
rect 200672 227808 200724 227860
rect 230664 227808 230716 227860
rect 280804 227808 280856 227860
rect 284760 227808 284812 227860
rect 297364 227808 297416 227860
rect 305368 227808 305420 227860
rect 396724 227740 396776 227792
rect 397460 227740 397512 227792
rect 400864 227740 400916 227792
rect 402612 227740 402664 227792
rect 403256 227740 403308 227792
rect 409144 227740 409196 227792
rect 410340 227740 410392 227792
rect 411904 227740 411956 227792
rect 413560 227740 413612 227792
rect 416688 227740 416740 227792
rect 420644 227740 420696 227792
rect 474740 227740 474792 227792
rect 482744 227740 482796 227792
rect 659568 227740 659620 227792
rect 665272 227740 665324 227792
rect 117044 227672 117096 227724
rect 187516 227672 187568 227724
rect 200028 227672 200080 227724
rect 252008 227672 252060 227724
rect 263416 227672 263468 227724
rect 301504 227672 301556 227724
rect 516600 227672 516652 227724
rect 538864 227672 538916 227724
rect 672954 227672 673006 227724
rect 671620 227604 671672 227656
rect 109868 227536 109920 227588
rect 182364 227536 182416 227588
rect 182824 227536 182876 227588
rect 236460 227536 236512 227588
rect 242716 227536 242768 227588
rect 285404 227536 285456 227588
rect 293684 227536 293736 227588
rect 325332 227536 325384 227588
rect 512092 227536 512144 227588
rect 533160 227536 533212 227588
rect 103244 227400 103296 227452
rect 177212 227400 177264 227452
rect 185400 227400 185452 227452
rect 192668 227400 192720 227452
rect 198464 227400 198516 227452
rect 253204 227400 253256 227452
rect 259368 227400 259420 227452
rect 298284 227400 298336 227452
rect 301964 227400 302016 227452
rect 331128 227400 331180 227452
rect 333888 227400 333940 227452
rect 356244 227400 356296 227452
rect 493968 227400 494020 227452
rect 505652 227400 505704 227452
rect 521108 227400 521160 227452
rect 544568 227400 544620 227452
rect 672172 227400 672224 227452
rect 81348 227264 81400 227316
rect 95240 227264 95292 227316
rect 96528 227264 96580 227316
rect 172060 227264 172112 227316
rect 173164 227264 173216 227316
rect 185584 227264 185636 227316
rect 188988 227264 189040 227316
rect 244188 227264 244240 227316
rect 251088 227264 251140 227316
rect 294420 227264 294472 227316
rect 308864 227264 308916 227316
rect 339500 227264 339552 227316
rect 351184 227264 351236 227316
rect 363328 227264 363380 227316
rect 363604 227264 363656 227316
rect 368480 227264 368532 227316
rect 467656 227264 467708 227316
rect 476580 227264 476632 227316
rect 481180 227264 481232 227316
rect 492680 227264 492732 227316
rect 495348 227264 495400 227316
rect 511448 227264 511500 227316
rect 528192 227264 528244 227316
rect 553676 227264 553728 227316
rect 671804 227196 671856 227248
rect 68192 227128 68244 227180
rect 143724 227128 143776 227180
rect 156604 227128 156656 227180
rect 213276 227128 213328 227180
rect 224776 227128 224828 227180
rect 273812 227128 273864 227180
rect 274456 227128 274508 227180
rect 312452 227128 312504 227180
rect 319812 227128 319864 227180
rect 345848 227128 345900 227180
rect 346032 227128 346084 227180
rect 366548 227128 366600 227180
rect 369768 227128 369820 227180
rect 384580 227128 384632 227180
rect 391388 227128 391440 227180
rect 400680 227128 400732 227180
rect 401324 227128 401376 227180
rect 408408 227128 408460 227180
rect 474096 227128 474148 227180
rect 484860 227128 484912 227180
rect 488908 227128 488960 227180
rect 503260 227128 503312 227180
rect 506296 227128 506348 227180
rect 526444 227128 526496 227180
rect 533344 227128 533396 227180
rect 561312 227128 561364 227180
rect 56508 226992 56560 227044
rect 142436 226992 142488 227044
rect 143356 226992 143408 227044
rect 208124 226992 208176 227044
rect 122748 226856 122800 226908
rect 185400 226856 185452 226908
rect 185584 226856 185636 226908
rect 226156 226992 226208 227044
rect 228732 226992 228784 227044
rect 275100 226992 275152 227044
rect 284944 226992 284996 227044
rect 320180 226992 320232 227044
rect 325516 226992 325568 227044
rect 349160 226992 349212 227044
rect 357256 226992 357308 227044
rect 374276 226992 374328 227044
rect 376484 226992 376536 227044
rect 389732 226992 389784 227044
rect 395712 226992 395764 227044
rect 406476 226992 406528 227044
rect 412548 226992 412600 227044
rect 419356 226992 419408 227044
rect 477316 226992 477368 227044
rect 489000 226992 489052 227044
rect 499212 226992 499264 227044
rect 516416 226992 516468 227044
rect 523684 226992 523736 227044
rect 548524 226992 548576 227044
rect 555424 226992 555476 227044
rect 633716 226992 633768 227044
rect 672264 226992 672316 227044
rect 212356 226856 212408 226908
rect 262220 226856 262272 226908
rect 275468 226856 275520 226908
rect 311164 226856 311216 226908
rect 384764 226856 384816 226908
rect 395528 226856 395580 226908
rect 419448 226856 419500 226908
rect 424508 226856 424560 226908
rect 672264 226856 672316 226908
rect 129464 226720 129516 226772
rect 197820 226720 197872 226772
rect 224592 226720 224644 226772
rect 270592 226720 270644 226772
rect 150072 226584 150124 226636
rect 156604 226584 156656 226636
rect 160008 226584 160060 226636
rect 221004 226584 221056 226636
rect 671804 226584 671856 226636
rect 177304 226448 177356 226500
rect 231308 226448 231360 226500
rect 670700 226448 670752 226500
rect 385684 226312 385736 226364
rect 391664 226312 391716 226364
rect 407764 226312 407816 226364
rect 411628 226312 411680 226364
rect 63408 226244 63460 226296
rect 133972 226244 134024 226296
rect 135168 226244 135220 226296
rect 204260 226244 204312 226296
rect 219164 226244 219216 226296
rect 267372 226244 267424 226296
rect 286968 226244 287020 226296
rect 319536 226244 319588 226296
rect 518900 226244 518952 226296
rect 531964 226244 532016 226296
rect 99104 226108 99156 226160
rect 175924 226108 175976 226160
rect 205456 226108 205508 226160
rect 258356 226108 258408 226160
rect 296628 226108 296680 226160
rect 329196 226108 329248 226160
rect 330484 226108 330536 226160
rect 351920 226108 351972 226160
rect 352564 226108 352616 226160
rect 358176 226108 358228 226160
rect 501144 226108 501196 226160
rect 519268 226108 519320 226160
rect 525984 226108 526036 226160
rect 539784 226244 539836 226296
rect 671712 226244 671764 226296
rect 84108 225972 84160 226024
rect 161756 225972 161808 226024
rect 186044 225972 186096 226024
rect 241612 225972 241664 226024
rect 255136 225972 255188 226024
rect 296996 225972 297048 226024
rect 303252 225972 303304 226024
rect 333060 225972 333112 226024
rect 480720 225972 480772 226024
rect 487804 225972 487856 226024
rect 517888 225972 517940 226024
rect 540612 226108 540664 226160
rect 671804 226040 671856 226092
rect 539600 225972 539652 226024
rect 555332 225972 555384 226024
rect 350356 225904 350408 225956
rect 354864 225904 354916 225956
rect 70124 225836 70176 225888
rect 151452 225836 151504 225888
rect 155776 225836 155828 225888
rect 219716 225836 219768 225888
rect 220636 225836 220688 225888
rect 268016 225836 268068 225888
rect 268844 225836 268896 225888
rect 306012 225836 306064 225888
rect 319996 225836 320048 225888
rect 347228 225836 347280 225888
rect 355324 225836 355376 225888
rect 372344 225836 372396 225888
rect 388444 225836 388496 225888
rect 396540 225836 396592 225888
rect 486516 225836 486568 225888
rect 494796 225836 494848 225888
rect 495992 225836 496044 225888
rect 512276 225836 512328 225888
rect 525616 225836 525668 225888
rect 551008 225836 551060 225888
rect 458640 225768 458692 225820
rect 462596 225768 462648 225820
rect 60004 225700 60056 225752
rect 141792 225700 141844 225752
rect 142068 225700 142120 225752
rect 209412 225700 209464 225752
rect 209596 225700 209648 225752
rect 259644 225700 259696 225752
rect 264704 225700 264756 225752
rect 304724 225700 304776 225752
rect 306104 225700 306156 225752
rect 336924 225700 336976 225752
rect 340696 225700 340748 225752
rect 361488 225700 361540 225752
rect 365536 225700 365588 225752
rect 380072 225700 380124 225752
rect 380256 225700 380308 225752
rect 391020 225700 391072 225752
rect 472164 225700 472216 225752
rect 480812 225700 480864 225752
rect 487988 225700 488040 225752
rect 501512 225700 501564 225752
rect 505008 225700 505060 225752
rect 524144 225700 524196 225752
rect 537852 225700 537904 225752
rect 566096 225700 566148 225752
rect 671820 225700 671872 225752
rect 667940 225632 667992 225684
rect 61844 225564 61896 225616
rect 144368 225564 144420 225616
rect 158444 225564 158496 225616
rect 222292 225564 222344 225616
rect 239404 225564 239456 225616
rect 284116 225564 284168 225616
rect 288164 225564 288216 225616
rect 321468 225564 321520 225616
rect 324044 225564 324096 225616
rect 348516 225564 348568 225616
rect 349068 225564 349120 225616
rect 367192 225564 367244 225616
rect 375288 225564 375340 225616
rect 387800 225564 387852 225616
rect 391756 225564 391808 225616
rect 403532 225564 403584 225616
rect 469404 225564 469456 225616
rect 473544 225564 473596 225616
rect 478604 225564 478656 225616
rect 485872 225564 485924 225616
rect 491300 225564 491352 225616
rect 505928 225564 505980 225616
rect 508228 225564 508280 225616
rect 527364 225564 527416 225616
rect 535276 225564 535328 225616
rect 563520 225564 563572 225616
rect 132224 225428 132276 225480
rect 201684 225428 201736 225480
rect 202604 225428 202656 225480
rect 254492 225428 254544 225480
rect 254952 225428 255004 225480
rect 295708 225428 295760 225480
rect 670700 225428 670752 225480
rect 506112 225360 506164 225412
rect 510344 225360 510396 225412
rect 138848 225292 138900 225344
rect 206376 225292 206428 225344
rect 206560 225292 206612 225344
rect 228088 225292 228140 225344
rect 245568 225292 245620 225344
rect 287980 225292 288032 225344
rect 463148 225224 463200 225276
rect 467104 225224 467156 225276
rect 671160 225224 671212 225276
rect 155592 225156 155644 225208
rect 218428 225156 218480 225208
rect 225512 225156 225564 225208
rect 246120 225156 246172 225208
rect 166080 225020 166132 225072
rect 186872 225020 186924 225072
rect 195888 225020 195940 225072
rect 249340 225020 249392 225072
rect 670700 225020 670752 225072
rect 260104 224952 260156 225004
rect 264152 224952 264204 225004
rect 367744 224952 367796 225004
rect 373632 224952 373684 225004
rect 404176 224952 404228 225004
rect 412272 224952 412324 225004
rect 529848 224952 529900 225004
rect 619640 224952 619692 225004
rect 118608 224884 118660 224936
rect 185584 224884 185636 224936
rect 191472 224884 191524 224936
rect 248052 224884 248104 224936
rect 266268 224884 266320 224936
rect 303436 224884 303488 224936
rect 321468 224884 321520 224936
rect 346584 224884 346636 224936
rect 426440 224884 426492 224936
rect 426992 224884 427044 224936
rect 466368 224816 466420 224868
rect 471244 224816 471296 224868
rect 669044 224816 669096 224868
rect 112904 224748 112956 224800
rect 185860 224748 185912 224800
rect 105728 224612 105780 224664
rect 181076 224612 181128 224664
rect 185768 224612 185820 224664
rect 242900 224748 242952 224800
rect 271328 224748 271380 224800
rect 309876 224748 309928 224800
rect 313096 224748 313148 224800
rect 342076 224748 342128 224800
rect 186320 224612 186372 224664
rect 240324 224612 240376 224664
rect 249616 224612 249668 224664
rect 290556 224612 290608 224664
rect 295156 224612 295208 224664
rect 325976 224612 326028 224664
rect 347044 224612 347096 224664
rect 365904 224748 365956 224800
rect 534632 224748 534684 224800
rect 547420 224748 547472 224800
rect 551836 224748 551888 224800
rect 558184 224748 558236 224800
rect 558368 224748 558420 224800
rect 562048 224748 562100 224800
rect 85488 224476 85540 224528
rect 165620 224476 165672 224528
rect 172336 224476 172388 224528
rect 232596 224476 232648 224528
rect 233148 224476 233200 224528
rect 277676 224476 277728 224528
rect 282552 224476 282604 224528
rect 316316 224476 316368 224528
rect 316868 224476 316920 224528
rect 342996 224476 343048 224528
rect 343364 224476 343416 224528
rect 363972 224612 364024 224664
rect 493048 224612 493100 224664
rect 508596 224612 508648 224664
rect 598388 224612 598440 224664
rect 670884 224612 670936 224664
rect 363788 224476 363840 224528
rect 378140 224476 378192 224528
rect 394516 224476 394568 224528
rect 404544 224476 404596 224528
rect 506940 224476 506992 224528
rect 525800 224476 525852 224528
rect 526260 224476 526312 224528
rect 551284 224476 551336 224528
rect 552756 224476 552808 224528
rect 558000 224476 558052 224528
rect 558184 224476 558236 224528
rect 625252 224476 625304 224528
rect 76564 224340 76616 224392
rect 157800 224340 157852 224392
rect 165344 224340 165396 224392
rect 227444 224340 227496 224392
rect 241244 224340 241296 224392
rect 286692 224340 286744 224392
rect 291108 224340 291160 224392
rect 323860 224340 323912 224392
rect 341892 224340 341944 224392
rect 365260 224340 365312 224392
rect 368204 224340 368256 224392
rect 382556 224340 382608 224392
rect 382924 224340 382976 224392
rect 396172 224340 396224 224392
rect 436376 224340 436428 224392
rect 436836 224340 436888 224392
rect 480536 224340 480588 224392
rect 492864 224340 492916 224392
rect 497280 224340 497332 224392
rect 514024 224340 514076 224392
rect 519820 224340 519872 224392
rect 542544 224340 542596 224392
rect 549536 224340 549588 224392
rect 625436 224340 625488 224392
rect 63224 224204 63276 224256
rect 147588 224204 147640 224256
rect 151728 224204 151780 224256
rect 217140 224204 217192 224256
rect 223304 224204 223356 224256
rect 224960 224204 225012 224256
rect 231584 224204 231636 224256
rect 278964 224204 279016 224256
rect 281264 224204 281316 224256
rect 317604 224204 317656 224256
rect 322572 224204 322624 224256
rect 349804 224204 349856 224256
rect 351644 224204 351696 224256
rect 369584 224204 369636 224256
rect 372344 224204 372396 224256
rect 387432 224204 387484 224256
rect 387708 224204 387760 224256
rect 398104 224204 398156 224256
rect 405464 224204 405516 224256
rect 414204 224204 414256 224256
rect 420828 224204 420880 224256
rect 425152 224204 425204 224256
rect 427820 224204 427872 224256
rect 428740 224204 428792 224256
rect 436284 224204 436336 224256
rect 437020 224204 437072 224256
rect 438952 224204 439004 224256
rect 439596 224204 439648 224256
rect 451372 224204 451424 224256
rect 452016 224204 452068 224256
rect 456156 224204 456208 224256
rect 459744 224204 459796 224256
rect 462412 224204 462464 224256
rect 469680 224204 469732 224256
rect 470876 224204 470928 224256
rect 477500 224204 477552 224256
rect 489552 224204 489604 224256
rect 504088 224204 504140 224256
rect 504640 224204 504692 224256
rect 523040 224204 523092 224256
rect 527548 224204 527600 224256
rect 552020 224204 552072 224256
rect 556804 224204 556856 224256
rect 570328 224204 570380 224256
rect 115664 224068 115716 224120
rect 188804 224068 188856 224120
rect 189908 224068 189960 224120
rect 212632 224068 212684 224120
rect 216588 224068 216640 224120
rect 264428 224068 264480 224120
rect 275836 224068 275888 224120
rect 288716 224068 288768 224120
rect 510344 224000 510396 224052
rect 615500 224000 615552 224052
rect 122288 223932 122340 223984
rect 193956 223932 194008 223984
rect 196808 223932 196860 223984
rect 222936 223932 222988 223984
rect 226156 223932 226208 223984
rect 272524 223932 272576 223984
rect 289084 223864 289136 223916
rect 294788 223864 294840 223916
rect 514852 223864 514904 223916
rect 515220 223864 515272 223916
rect 616880 223864 616932 223916
rect 140044 223796 140096 223848
rect 171416 223796 171468 223848
rect 175188 223796 175240 223848
rect 235172 223796 235224 223848
rect 514668 223728 514720 223780
rect 536380 223728 536432 223780
rect 539784 223728 539836 223780
rect 622400 223728 622452 223780
rect 181904 223660 181956 223712
rect 102048 223524 102100 223576
rect 178500 223524 178552 223576
rect 185584 223660 185636 223712
rect 191012 223660 191064 223712
rect 227444 223660 227496 223712
rect 273168 223660 273220 223712
rect 415308 223660 415360 223712
rect 419632 223660 419684 223712
rect 460572 223660 460624 223712
rect 462964 223660 463016 223712
rect 670516 223660 670568 223712
rect 670930 224068 670982 224120
rect 543648 223592 543700 223644
rect 557448 223592 557500 223644
rect 626540 223592 626592 223644
rect 654968 223592 655020 223644
rect 656716 223592 656768 223644
rect 186320 223524 186372 223576
rect 194324 223524 194376 223576
rect 247408 223524 247460 223576
rect 253756 223524 253808 223576
rect 293500 223524 293552 223576
rect 307024 223524 307076 223576
rect 315396 223524 315448 223576
rect 454776 223524 454828 223576
rect 460112 223524 460164 223576
rect 473728 223524 473780 223576
rect 480996 223524 481048 223576
rect 670332 223524 670384 223576
rect 88248 223388 88300 223440
rect 164976 223388 165028 223440
rect 166448 223388 166500 223440
rect 192024 223388 192076 223440
rect 197268 223388 197320 223440
rect 249984 223388 250036 223440
rect 267372 223388 267424 223440
rect 307300 223388 307352 223440
rect 322848 223388 322900 223440
rect 332416 223388 332468 223440
rect 498568 223388 498620 223440
rect 515772 223388 515824 223440
rect 516784 223388 516836 223440
rect 527180 223388 527232 223440
rect 528560 223388 528612 223440
rect 542360 223388 542412 223440
rect 78404 223252 78456 223304
rect 81164 223116 81216 223168
rect 154304 223116 154356 223168
rect 157064 223252 157116 223304
rect 160192 223252 160244 223304
rect 157248 223116 157300 223168
rect 159272 223116 159324 223168
rect 181720 223252 181772 223304
rect 191656 223252 191708 223304
rect 244832 223252 244884 223304
rect 262128 223252 262180 223304
rect 300860 223252 300912 223304
rect 315672 223252 315724 223304
rect 341432 223252 341484 223304
rect 342076 223252 342128 223304
rect 362040 223252 362092 223304
rect 366916 223252 366968 223304
rect 382004 223252 382056 223304
rect 407028 223252 407080 223304
rect 414848 223252 414900 223304
rect 503444 223252 503496 223304
rect 521752 223252 521804 223304
rect 522488 223252 522540 223304
rect 534908 223252 534960 223304
rect 536748 223252 536800 223304
rect 559932 223252 559984 223304
rect 567752 223252 567804 223304
rect 670608 223252 670660 223304
rect 168288 223116 168340 223168
rect 226800 223116 226852 223168
rect 248144 223116 248196 223168
rect 291844 223116 291896 223168
rect 300768 223116 300820 223168
rect 330116 223116 330168 223168
rect 336464 223116 336516 223168
rect 359740 223116 359792 223168
rect 366732 223116 366784 223168
rect 383936 223116 383988 223168
rect 483112 223116 483164 223168
rect 495808 223116 495860 223168
rect 515956 223116 516008 223168
rect 538312 223116 538364 223168
rect 539048 223116 539100 223168
rect 75828 222980 75880 223032
rect 154672 222980 154724 223032
rect 164056 222980 164108 223032
rect 224224 222980 224276 223032
rect 238668 222980 238720 223032
rect 282828 222980 282880 223032
rect 292488 222980 292540 223032
rect 326620 222980 326672 223032
rect 329748 222980 329800 223032
rect 353668 222980 353720 223032
rect 355784 222980 355836 223032
rect 375564 222980 375616 223032
rect 382096 222980 382148 223032
rect 392952 222980 393004 223032
rect 479892 222980 479944 223032
rect 491944 222980 491996 223032
rect 500500 222980 500552 223032
rect 518440 222980 518492 223032
rect 518808 222980 518860 223032
rect 618260 222980 618312 223032
rect 68928 222844 68980 222896
rect 149520 222844 149572 222896
rect 154488 222844 154540 222896
rect 216220 222844 216272 222896
rect 217784 222844 217836 222896
rect 268660 222844 268712 222896
rect 278412 222844 278464 222896
rect 313740 222844 313792 222896
rect 315856 222844 315908 222896
rect 344652 222844 344704 222896
rect 346216 222844 346268 222896
rect 367468 222844 367520 222896
rect 386328 222844 386380 222896
rect 398380 222844 398432 222896
rect 398564 222844 398616 222896
rect 405832 222844 405884 222896
rect 459928 222844 459980 222896
rect 466736 222844 466788 222896
rect 467288 222844 467340 222896
rect 475016 222844 475068 222896
rect 486332 222844 486384 222896
rect 499856 222844 499908 222896
rect 508872 222844 508924 222896
rect 528928 222844 528980 222896
rect 537208 222844 537260 222896
rect 565636 222844 565688 222896
rect 571616 222844 571668 222896
rect 131028 222708 131080 222760
rect 196072 222708 196124 222760
rect 208124 222708 208176 222760
rect 260932 222708 260984 222760
rect 290924 222708 290976 222760
rect 321836 222708 321888 222760
rect 525156 222708 525208 222760
rect 537576 222708 537628 222760
rect 146024 222572 146076 222624
rect 211988 222572 212040 222624
rect 213828 222572 213880 222624
rect 262864 222572 262916 222624
rect 542360 222708 542412 222760
rect 622584 222708 622636 222760
rect 622768 222572 622820 222624
rect 134708 222436 134760 222488
rect 197452 222436 197504 222488
rect 204168 222436 204220 222488
rect 254768 222436 254820 222488
rect 527180 222436 527232 222488
rect 620008 222436 620060 222488
rect 416504 222368 416556 222420
rect 422208 222368 422260 222420
rect 154304 222300 154356 222352
rect 159824 222300 159876 222352
rect 178684 222300 178736 222352
rect 204904 222300 204956 222352
rect 244004 222300 244056 222352
rect 286048 222300 286100 222352
rect 524788 222300 524840 222352
rect 619824 222300 619876 222352
rect 529480 222164 529532 222216
rect 555700 222164 555752 222216
rect 567752 222164 567804 222216
rect 627092 222164 627144 222216
rect 670332 222164 670384 222216
rect 670792 222164 670844 222216
rect 111432 222096 111484 222148
rect 182548 222096 182600 222148
rect 184020 222096 184072 222148
rect 239220 222096 239272 222148
rect 267096 222096 267148 222148
rect 303804 222096 303856 222148
rect 330852 222096 330904 222148
rect 345664 222096 345716 222148
rect 424968 222096 425020 222148
rect 429292 222096 429344 222148
rect 462136 222096 462188 222148
rect 468484 222096 468536 222148
rect 471888 222096 471940 222148
rect 479248 222096 479300 222148
rect 509884 222096 509936 222148
rect 518808 222096 518860 222148
rect 519820 222096 519872 222148
rect 533344 222028 533396 222080
rect 538680 222028 538732 222080
rect 104624 221960 104676 222012
rect 177488 221960 177540 222012
rect 195152 221960 195204 222012
rect 250168 221960 250220 222012
rect 269948 221960 270000 222012
rect 306564 221960 306616 222012
rect 306840 221960 306892 222012
rect 335452 221960 335504 222012
rect 513748 221960 513800 222012
rect 524788 221960 524840 222012
rect 539048 221960 539100 222012
rect 604460 221960 604512 222012
rect 101496 221824 101548 221876
rect 175464 221824 175516 221876
rect 189448 221824 189500 221876
rect 245108 221824 245160 221876
rect 258080 221824 258132 221876
rect 269212 221824 269264 221876
rect 277860 221824 277912 221876
rect 314844 221824 314896 221876
rect 344928 221824 344980 221876
rect 364524 221824 364576 221876
rect 484308 221824 484360 221876
rect 496912 221824 496964 221876
rect 523960 221824 524012 221876
rect 548984 221824 549036 221876
rect 560760 221824 560812 221876
rect 561312 221824 561364 221876
rect 565084 221824 565136 221876
rect 567292 221824 567344 221876
rect 60648 221688 60700 221740
rect 94504 221688 94556 221740
rect 94872 221688 94924 221740
rect 161480 221688 161532 221740
rect 74172 221552 74224 221604
rect 86224 221552 86276 221604
rect 91560 221552 91612 221604
rect 167276 221688 167328 221740
rect 177672 221688 177724 221740
rect 234160 221688 234212 221740
rect 247132 221688 247184 221740
rect 253388 221688 253440 221740
rect 253572 221688 253624 221740
rect 258632 221688 258684 221740
rect 260472 221688 260524 221740
rect 298376 221688 298428 221740
rect 298560 221688 298612 221740
rect 328552 221688 328604 221740
rect 331680 221688 331732 221740
rect 353944 221688 353996 221740
rect 362316 221688 362368 221740
rect 376024 221688 376076 221740
rect 84936 221416 84988 221468
rect 162032 221552 162084 221604
rect 178500 221552 178552 221604
rect 237380 221552 237432 221604
rect 238852 221552 238904 221604
rect 248604 221552 248656 221604
rect 250536 221552 250588 221604
rect 291384 221552 291436 221604
rect 296444 221552 296496 221604
rect 327540 221552 327592 221604
rect 328368 221552 328420 221604
rect 351368 221552 351420 221604
rect 353392 221552 353444 221604
rect 369952 221552 370004 221604
rect 370504 221552 370556 221604
rect 382740 221688 382792 221740
rect 494336 221688 494388 221740
rect 510712 221688 510764 221740
rect 522856 221688 522908 221740
rect 546500 221688 546552 221740
rect 548524 221688 548576 221740
rect 607220 221688 607272 221740
rect 382740 221552 382792 221604
rect 394884 221552 394936 221604
rect 397092 221552 397144 221604
rect 407304 221552 407356 221604
rect 456708 221552 456760 221604
rect 461768 221552 461820 221604
rect 468760 221552 468812 221604
rect 474280 221552 474332 221604
rect 478788 221552 478840 221604
rect 489184 221552 489236 221604
rect 496176 221552 496228 221604
rect 513472 221552 513524 221604
rect 533712 221552 533764 221604
rect 535460 221552 535512 221604
rect 538496 221552 538548 221604
rect 538680 221552 538732 221604
rect 603080 221552 603132 221604
rect 161940 221416 161992 221468
rect 224408 221416 224460 221468
rect 234344 221416 234396 221468
rect 281724 221416 281776 221468
rect 284024 221416 284076 221468
rect 289912 221416 289964 221468
rect 292304 221416 292356 221468
rect 299756 221416 299808 221468
rect 302700 221416 302752 221468
rect 334072 221416 334124 221468
rect 335268 221416 335320 221468
rect 357532 221416 357584 221468
rect 358176 221416 358228 221468
rect 374552 221416 374604 221468
rect 375472 221416 375524 221468
rect 386512 221416 386564 221468
rect 390468 221416 390520 221468
rect 401692 221416 401744 221468
rect 408408 221416 408460 221468
rect 416872 221416 416924 221468
rect 452568 221416 452620 221468
rect 456708 221416 456760 221468
rect 484032 221416 484084 221468
rect 534632 221416 534684 221468
rect 560760 221416 560812 221468
rect 560944 221348 560996 221400
rect 568672 221348 568724 221400
rect 121368 221280 121420 221332
rect 190644 221280 190696 221332
rect 201408 221280 201460 221332
rect 255412 221280 255464 221332
rect 282828 221280 282880 221332
rect 283564 221280 283616 221332
rect 530952 221212 531004 221264
rect 603356 221212 603408 221264
rect 667940 221212 667992 221264
rect 670792 221212 670844 221264
rect 148692 221144 148744 221196
rect 214104 221144 214156 221196
rect 215208 221144 215260 221196
rect 263140 221144 263192 221196
rect 374000 221144 374052 221196
rect 381084 221144 381136 221196
rect 527364 221076 527416 221128
rect 528008 221076 528060 221128
rect 603540 221076 603592 221128
rect 141240 221008 141292 221060
rect 205824 221008 205876 221060
rect 222568 221008 222620 221060
rect 270868 221008 270920 221060
rect 387156 220940 387208 220992
rect 389916 220940 389968 220992
rect 526444 220940 526496 220992
rect 601792 220940 601844 220992
rect 161480 220872 161532 220924
rect 169760 220872 169812 220924
rect 172520 220872 172572 220924
rect 194968 220872 195020 220924
rect 228180 220872 228232 220924
rect 276112 220872 276164 220924
rect 420644 220804 420696 220856
rect 423864 220804 423916 220856
rect 521292 220804 521344 220856
rect 600412 220804 600464 220856
rect 108120 220736 108172 220788
rect 179972 220736 180024 220788
rect 187608 220736 187660 220788
rect 241796 220736 241848 220788
rect 261300 220736 261352 220788
rect 301780 220736 301832 220788
rect 313924 220736 313976 220788
rect 320364 220736 320416 220788
rect 338948 220736 339000 220788
rect 342444 220736 342496 220788
rect 455328 220736 455380 220788
rect 458548 220736 458600 220788
rect 465724 220736 465776 220788
rect 469312 220736 469364 220788
rect 476764 220736 476816 220788
rect 478420 220736 478472 220788
rect 518164 220668 518216 220720
rect 529848 220668 529900 220720
rect 534632 220668 534684 220720
rect 66720 220600 66772 220652
rect 144184 220600 144236 220652
rect 144552 220600 144604 220652
rect 208584 220600 208636 220652
rect 216404 220600 216456 220652
rect 217324 220600 217376 220652
rect 217508 220600 217560 220652
rect 265072 220600 265124 220652
rect 277032 220600 277084 220652
rect 311440 220600 311492 220652
rect 311624 220600 311676 220652
rect 338580 220600 338632 220652
rect 535092 220668 535144 220720
rect 543740 220668 543792 220720
rect 544476 220668 544528 220720
rect 551836 220668 551888 220720
rect 558000 220668 558052 220720
rect 558552 220668 558604 220720
rect 559748 220668 559800 220720
rect 563520 220668 563572 220720
rect 563704 220600 563756 220652
rect 535460 220532 535512 220584
rect 535736 220532 535788 220584
rect 553308 220532 553360 220584
rect 553492 220532 553544 220584
rect 558920 220532 558972 220584
rect 86592 220464 86644 220516
rect 164332 220464 164384 220516
rect 180708 220464 180760 220516
rect 79784 220328 79836 220380
rect 158904 220328 158956 220380
rect 171048 220328 171100 220380
rect 229100 220328 229152 220380
rect 231860 220464 231912 220516
rect 238024 220464 238076 220516
rect 246948 220464 247000 220516
rect 288532 220464 288584 220516
rect 310152 220464 310204 220516
rect 338212 220464 338264 220516
rect 342720 220464 342772 220516
rect 352380 220464 352432 220516
rect 353208 220464 353260 220516
rect 371424 220464 371476 220516
rect 432236 220464 432288 220516
rect 434812 220464 434864 220516
rect 482928 220464 482980 220516
rect 495348 220464 495400 220516
rect 500224 220464 500276 220516
rect 509240 220464 509292 220516
rect 513288 220464 513340 220516
rect 534632 220464 534684 220516
rect 562508 220464 562560 220516
rect 571340 220464 571392 220516
rect 571616 220600 571668 220652
rect 611360 220600 611412 220652
rect 610532 220464 610584 220516
rect 543740 220396 543792 220448
rect 552020 220396 552072 220448
rect 552756 220396 552808 220448
rect 236644 220328 236696 220380
rect 240600 220328 240652 220380
rect 283104 220328 283156 220380
rect 299204 220328 299256 220380
rect 331404 220328 331456 220380
rect 338028 220328 338080 220380
rect 359004 220328 359056 220380
rect 372528 220328 372580 220380
rect 385408 220328 385460 220380
rect 469128 220328 469180 220380
rect 476120 220328 476172 220380
rect 485688 220328 485740 220380
rect 499120 220328 499172 220380
rect 504364 220328 504416 220380
rect 517704 220328 517756 220380
rect 518808 220328 518860 220380
rect 521568 220328 521620 220380
rect 608692 220328 608744 220380
rect 76380 220192 76432 220244
rect 156144 220192 156196 220244
rect 161480 220192 161532 220244
rect 73068 220056 73120 220108
rect 153752 220056 153804 220108
rect 157800 220056 157852 220108
rect 218612 220056 218664 220108
rect 220820 220192 220872 220244
rect 233424 220192 233476 220244
rect 237288 220192 237340 220244
rect 280528 220192 280580 220244
rect 283656 220192 283708 220244
rect 316592 220192 316644 220244
rect 329196 220192 329248 220244
rect 354680 220192 354732 220244
rect 361488 220192 361540 220244
rect 376852 220192 376904 220244
rect 377036 220192 377088 220244
rect 388628 220192 388680 220244
rect 459468 220192 459520 220244
rect 465172 220192 465224 220244
rect 473268 220192 473320 220244
rect 481732 220192 481784 220244
rect 488172 220192 488224 220244
rect 502432 220192 502484 220244
rect 507124 220192 507176 220244
rect 521936 220192 521988 220244
rect 531228 220192 531280 220244
rect 556252 220260 556304 220312
rect 558552 220192 558604 220244
rect 609428 220192 609480 220244
rect 548708 220124 548760 220176
rect 221280 220056 221332 220108
rect 230204 220056 230256 220108
rect 275284 220056 275336 220108
rect 280068 220056 280120 220108
rect 313740 220056 313792 220108
rect 318432 220056 318484 220108
rect 114468 219920 114520 219972
rect 185124 219920 185176 219972
rect 200856 219920 200908 219972
rect 252744 219920 252796 219972
rect 257160 219920 257212 219972
rect 295984 219920 296036 219972
rect 343640 220056 343692 220108
rect 347872 220056 347924 220108
rect 354312 220056 354364 220108
rect 372804 220056 372856 220108
rect 379428 220056 379480 220108
rect 392124 220056 392176 220108
rect 395988 220056 396040 220108
rect 404728 220056 404780 220108
rect 421932 220056 421984 220108
rect 426808 220056 426860 220108
rect 475936 220056 475988 220108
rect 485872 220056 485924 220108
rect 491668 220056 491720 220108
rect 507768 220056 507820 220108
rect 511816 220056 511868 220108
rect 531504 220056 531556 220108
rect 532516 220056 532568 220108
rect 414480 219988 414532 220040
rect 418344 219988 418396 220040
rect 553492 219988 553544 220040
rect 592684 220056 592736 220108
rect 633440 220056 633492 220108
rect 636476 220056 636528 220108
rect 653404 220056 653456 220108
rect 675852 220056 675904 220108
rect 676496 220056 676548 220108
rect 582564 219988 582616 220040
rect 343824 219920 343876 219972
rect 528560 219920 528612 219972
rect 534264 219920 534316 219972
rect 542544 219852 542596 219904
rect 543096 219852 543148 219904
rect 605840 219852 605892 219904
rect 127992 219784 128044 219836
rect 195612 219784 195664 219836
rect 207480 219784 207532 219836
rect 257344 219784 257396 219836
rect 288532 219784 288584 219836
rect 310520 219784 310572 219836
rect 543740 219716 543792 219768
rect 548708 219716 548760 219768
rect 551008 219716 551060 219768
rect 607772 219716 607824 219768
rect 137928 219648 137980 219700
rect 203156 219648 203208 219700
rect 236460 219648 236512 219700
rect 261484 219648 261536 219700
rect 464988 219580 465040 219632
rect 471980 219580 472032 219632
rect 545764 219580 545816 219632
rect 606668 219580 606720 219632
rect 179512 219512 179564 219564
rect 232044 219512 232096 219564
rect 235908 219512 235960 219564
rect 243084 219512 243136 219564
rect 273076 219512 273128 219564
rect 279240 219512 279292 219564
rect 406200 219512 406252 219564
rect 412732 219512 412784 219564
rect 108304 219376 108356 219428
rect 146852 219376 146904 219428
rect 153660 219376 153712 219428
rect 160744 219376 160796 219428
rect 163596 219376 163648 219428
rect 184204 219376 184256 219428
rect 192944 219376 192996 219428
rect 233884 219376 233936 219428
rect 253020 219376 253072 219428
rect 93584 219104 93636 219156
rect 140044 219240 140096 219292
rect 147036 219240 147088 219292
rect 189908 219240 189960 219292
rect 209688 219240 209740 219292
rect 210424 219240 210476 219292
rect 214380 219240 214432 219292
rect 253572 219240 253624 219292
rect 123852 219104 123904 219156
rect 87420 218968 87472 219020
rect 106924 218968 106976 219020
rect 107292 218968 107344 219020
rect 100484 218832 100536 218884
rect 108304 218832 108356 218884
rect 113916 218968 113968 219020
rect 166080 218968 166132 219020
rect 159272 218832 159324 218884
rect 183100 219104 183152 219156
rect 189724 219104 189776 219156
rect 199844 219104 199896 219156
rect 247132 219104 247184 219156
rect 272524 219376 272576 219428
rect 297364 219376 297416 219428
rect 323400 219376 323452 219428
rect 324044 219376 324096 219428
rect 324228 219376 324280 219428
rect 324872 219376 324924 219428
rect 325056 219376 325108 219428
rect 325516 219376 325568 219428
rect 259184 219240 259236 219292
rect 292304 219240 292356 219292
rect 307668 219240 307720 219292
rect 327724 219376 327776 219428
rect 373632 219376 373684 219428
rect 377036 219376 377088 219428
rect 417792 219376 417844 219428
rect 421012 219444 421064 219496
rect 428280 219376 428332 219428
rect 432052 219512 432104 219564
rect 521936 219444 521988 219496
rect 522580 219444 522632 219496
rect 528744 219512 528796 219564
rect 540612 219444 540664 219496
rect 606024 219444 606076 219496
rect 430212 219376 430264 219428
rect 432696 219376 432748 219428
rect 676220 219376 676272 219428
rect 678612 219376 678664 219428
rect 504548 219308 504600 219360
rect 327540 219240 327592 219292
rect 342720 219240 342772 219292
rect 354588 219240 354640 219292
rect 355324 219240 355376 219292
rect 457996 219240 458048 219292
rect 461124 219240 461176 219292
rect 166632 218968 166684 219020
rect 173164 218968 173216 219020
rect 173532 218968 173584 219020
rect 172520 218832 172572 218884
rect 174912 218832 174964 218884
rect 178684 218832 178736 218884
rect 179328 218968 179380 219020
rect 182824 218968 182876 219020
rect 186780 218968 186832 219020
rect 235908 218968 235960 219020
rect 238116 218968 238168 219020
rect 239404 218968 239456 219020
rect 239772 218968 239824 219020
rect 246488 218968 246540 219020
rect 249248 218968 249300 219020
rect 284024 218968 284076 219020
rect 300584 219104 300636 219156
rect 322848 219104 322900 219156
rect 325608 219104 325660 219156
rect 330484 219104 330536 219156
rect 363972 219104 364024 219156
rect 374000 219104 374052 219156
rect 388812 219104 388864 219156
rect 393964 219104 394016 219156
rect 419264 219104 419316 219156
rect 422668 219104 422720 219156
rect 496912 219104 496964 219156
rect 504732 219104 504784 219156
rect 289084 218968 289136 219020
rect 294420 218968 294472 219020
rect 309784 218968 309836 219020
rect 314292 218968 314344 219020
rect 338948 218968 339000 219020
rect 340512 218968 340564 219020
rect 351184 218968 351236 219020
rect 383568 218968 383620 219020
rect 388444 218968 388496 219020
rect 407580 218968 407632 219020
rect 411904 218968 411956 219020
rect 499856 218900 499908 218952
rect 214564 218832 214616 218884
rect 232964 218832 233016 218884
rect 273076 218832 273128 218884
rect 286140 218832 286192 218884
rect 313924 218832 313976 218884
rect 59820 218696 59872 218748
rect 68192 218696 68244 218748
rect 83924 218696 83976 218748
rect 160192 218696 160244 218748
rect 162768 218696 162820 218748
rect 169024 218696 169076 218748
rect 174360 218696 174412 218748
rect 179512 218696 179564 218748
rect 180156 218696 180208 218748
rect 231860 218696 231912 218748
rect 233884 218696 233936 218748
rect 238852 218696 238904 218748
rect 244740 218696 244792 218748
rect 246304 218696 246356 218748
rect 246488 218696 246540 218748
rect 280804 218696 280856 218748
rect 291936 218696 291988 218748
rect 323584 218696 323636 218748
rect 120540 218560 120592 218612
rect 166448 218560 166500 218612
rect 170220 218560 170272 218612
rect 200672 218560 200724 218612
rect 206652 218560 206704 218612
rect 214380 218560 214432 218612
rect 214748 218560 214800 218612
rect 260104 218560 260156 218612
rect 262956 218560 263008 218612
rect 276664 218560 276716 218612
rect 279516 218560 279568 218612
rect 137100 218424 137152 218476
rect 174912 218424 174964 218476
rect 176292 218424 176344 218476
rect 183100 218424 183152 218476
rect 183284 218424 183336 218476
rect 202144 218424 202196 218476
rect 203340 218424 203392 218476
rect 213092 218424 213144 218476
rect 214564 218424 214616 218476
rect 220820 218424 220872 218476
rect 225972 218424 226024 218476
rect 265624 218424 265676 218476
rect 266084 218424 266136 218476
rect 272524 218424 272576 218476
rect 272892 218424 272944 218476
rect 288532 218424 288584 218476
rect 320916 218560 320968 218612
rect 343640 218832 343692 218884
rect 347412 218832 347464 218884
rect 363604 218832 363656 218884
rect 402060 218832 402112 218884
rect 407764 218832 407816 218884
rect 411996 218832 412048 218884
rect 412548 218832 412600 218884
rect 333704 218696 333756 218748
rect 352564 218696 352616 218748
rect 354036 218696 354088 218748
rect 367744 218696 367796 218748
rect 386144 218696 386196 218748
rect 396724 218696 396776 218748
rect 402704 218696 402756 218748
rect 409144 218696 409196 218748
rect 412548 218696 412600 218748
rect 417148 218696 417200 218748
rect 484860 218696 484912 218748
rect 506296 218696 506348 218748
rect 392952 218560 393004 218612
rect 400864 218560 400916 218612
rect 504732 218560 504784 218612
rect 505284 218560 505336 218612
rect 534080 219308 534132 219360
rect 543924 219308 543976 219360
rect 553124 219308 553176 219360
rect 582472 219308 582524 219360
rect 596824 219308 596876 219360
rect 579436 219240 579488 219292
rect 579712 219240 579764 219292
rect 524052 219172 524104 219224
rect 528468 219172 528520 219224
rect 544660 219172 544712 219224
rect 558368 219172 558420 219224
rect 563244 219172 563296 219224
rect 563704 219172 563756 219224
rect 564440 219172 564492 219224
rect 565176 219172 565228 219224
rect 583116 219172 583168 219224
rect 534264 219104 534316 219156
rect 544292 219104 544344 219156
rect 562784 219104 562836 219156
rect 563060 219104 563112 219156
rect 567016 219104 567068 219156
rect 577504 219104 577556 219156
rect 547420 219036 547472 219088
rect 558184 219036 558236 219088
rect 514760 218900 514812 218952
rect 524052 218900 524104 218952
rect 534080 218900 534132 218952
rect 543648 218900 543700 218952
rect 543924 218900 543976 218952
rect 528284 218832 528336 218884
rect 529020 218832 529072 218884
rect 543464 218764 543516 218816
rect 543924 218764 543976 218816
rect 552572 218900 552624 218952
rect 553860 218900 553912 218952
rect 555332 218900 555384 218952
rect 567476 218968 567528 219020
rect 567660 218968 567712 219020
rect 572168 218968 572220 219020
rect 558736 218832 558788 218884
rect 568120 218832 568172 218884
rect 568304 218832 568356 218884
rect 572444 218832 572496 218884
rect 576216 218832 576268 218884
rect 553308 218764 553360 218816
rect 523960 218696 524012 218748
rect 531964 218696 532016 218748
rect 532608 218696 532660 218748
rect 528284 218628 528336 218680
rect 514944 218560 514996 218612
rect 534264 218560 534316 218612
rect 469864 218492 469916 218544
rect 470968 218492 471020 218544
rect 307024 218424 307076 218476
rect 365352 218424 365404 218476
rect 370504 218424 370556 218476
rect 523776 218424 523828 218476
rect 528468 218424 528520 218476
rect 528652 218424 528704 218476
rect 534448 218424 534500 218476
rect 553492 218696 553544 218748
rect 563060 218696 563112 218748
rect 543464 218560 543516 218612
rect 544108 218560 544160 218612
rect 544292 218560 544344 218612
rect 552940 218560 552992 218612
rect 553124 218560 553176 218612
rect 553860 218560 553912 218612
rect 558184 218560 558236 218612
rect 576216 218696 576268 218748
rect 576584 218968 576636 219020
rect 577688 218968 577740 219020
rect 576584 218832 576636 218884
rect 582380 218832 582432 218884
rect 595904 218832 595956 218884
rect 597560 218832 597612 218884
rect 611820 218696 611872 218748
rect 567752 218560 567804 218612
rect 577872 218560 577924 218612
rect 578056 218424 578108 218476
rect 582380 218424 582432 218476
rect 596088 218424 596140 218476
rect 450544 218356 450596 218408
rect 453580 218356 453632 218408
rect 57612 218288 57664 218340
rect 64144 218288 64196 218340
rect 68744 218288 68796 218340
rect 72424 218288 72476 218340
rect 159824 218288 159876 218340
rect 196808 218288 196860 218340
rect 199200 218288 199252 218340
rect 200028 218288 200080 218340
rect 203892 218288 203944 218340
rect 207664 218288 207716 218340
rect 213276 218288 213328 218340
rect 214748 218288 214800 218340
rect 219900 218288 219952 218340
rect 258080 218288 258132 218340
rect 344100 218288 344152 218340
rect 347044 218288 347096 218340
rect 370596 218288 370648 218340
rect 375472 218288 375524 218340
rect 377220 218288 377272 218340
rect 385684 218288 385736 218340
rect 426808 218288 426860 218340
rect 429568 218288 429620 218340
rect 479524 218288 479576 218340
rect 480352 218288 480404 218340
rect 534908 218288 534960 218340
rect 567752 218288 567804 218340
rect 568120 218288 568172 218340
rect 55956 218152 56008 218204
rect 56508 218152 56560 218204
rect 64236 218152 64288 218204
rect 65524 218152 65576 218204
rect 67548 218152 67600 218204
rect 71044 218152 71096 218204
rect 75644 218152 75696 218204
rect 76564 218152 76616 218204
rect 130476 218152 130528 218204
rect 167552 218152 167604 218204
rect 168104 218152 168156 218204
rect 170588 218152 170640 218204
rect 172152 218152 172204 218204
rect 177304 218152 177356 218204
rect 190092 218152 190144 218204
rect 225512 218152 225564 218204
rect 246396 218152 246448 218204
rect 249248 218152 249300 218204
rect 249432 218152 249484 218204
rect 251824 218152 251876 218204
rect 289452 218152 289504 218204
rect 294604 218152 294656 218204
rect 332508 218152 332560 218204
rect 335268 218152 335320 218204
rect 339132 218152 339184 218204
rect 340144 218152 340196 218204
rect 348884 218152 348936 218204
rect 353392 218152 353444 218204
rect 358728 218152 358780 218204
rect 363788 218152 363840 218204
rect 375104 218152 375156 218204
rect 380164 218152 380216 218204
rect 381912 218152 381964 218204
rect 382924 218152 382976 218204
rect 394332 218152 394384 218204
rect 402244 218152 402296 218204
rect 424416 218152 424468 218204
rect 426992 218152 427044 218204
rect 433248 218152 433300 218204
rect 435272 218152 435324 218204
rect 436008 218152 436060 218204
rect 436836 218152 436888 218204
rect 461952 218152 462004 218204
rect 466000 218152 466052 218204
rect 505652 218152 505704 218204
rect 558184 218152 558236 218204
rect 558368 218152 558420 218204
rect 567016 218152 567068 218204
rect 567476 218152 567528 218204
rect 594984 218152 595036 218204
rect 613016 218152 613068 218204
rect 56508 218016 56560 218068
rect 57244 218016 57296 218068
rect 58440 218016 58492 218068
rect 60004 218016 60056 218068
rect 62580 218016 62632 218068
rect 63224 218016 63276 218068
rect 65892 218016 65944 218068
rect 66904 218016 66956 218068
rect 68376 218016 68428 218068
rect 68928 218016 68980 218068
rect 72516 218016 72568 218068
rect 73804 218016 73856 218068
rect 75000 218016 75052 218068
rect 75828 218016 75880 218068
rect 79048 218016 79100 218068
rect 79968 218016 80020 218068
rect 80796 218016 80848 218068
rect 81348 218016 81400 218068
rect 83280 218016 83332 218068
rect 84108 218016 84160 218068
rect 93216 218016 93268 218068
rect 93768 218016 93820 218068
rect 97356 218016 97408 218068
rect 97908 218016 97960 218068
rect 99840 218016 99892 218068
rect 100668 218016 100720 218068
rect 103980 218016 104032 218068
rect 104808 218016 104860 218068
rect 112260 218016 112312 218068
rect 112904 218016 112956 218068
rect 116400 218016 116452 218068
rect 117044 218016 117096 218068
rect 128636 218016 128688 218068
rect 129648 218016 129700 218068
rect 132960 218016 133012 218068
rect 133604 218016 133656 218068
rect 142896 218016 142948 218068
rect 143356 218016 143408 218068
rect 145380 218016 145432 218068
rect 146024 218016 146076 218068
rect 149520 218016 149572 218068
rect 150072 218016 150124 218068
rect 155316 218016 155368 218068
rect 155776 218016 155828 218068
rect 159456 218016 159508 218068
rect 160008 218016 160060 218068
rect 160192 218016 160244 218068
rect 163228 218016 163280 218068
rect 166080 218016 166132 218068
rect 166632 218016 166684 218068
rect 167736 218016 167788 218068
rect 168288 218016 168340 218068
rect 171876 218016 171928 218068
rect 172336 218016 172388 218068
rect 176016 218016 176068 218068
rect 176476 218016 176528 218068
rect 182640 218016 182692 218068
rect 183468 218016 183520 218068
rect 184848 218016 184900 218068
rect 185584 218016 185636 218068
rect 188436 218016 188488 218068
rect 189448 218016 189500 218068
rect 190920 218016 190972 218068
rect 191656 218016 191708 218068
rect 192576 218016 192628 218068
rect 193128 218016 193180 218068
rect 196716 218016 196768 218068
rect 203892 218016 203944 218068
rect 204996 218016 205048 218068
rect 205456 218016 205508 218068
rect 211620 218016 211672 218068
rect 215208 218016 215260 218068
rect 215760 218016 215812 218068
rect 216588 218016 216640 218068
rect 221556 218016 221608 218068
rect 222568 218016 222620 218068
rect 224040 218016 224092 218068
rect 224592 218016 224644 218068
rect 225696 218016 225748 218068
rect 226156 218016 226208 218068
rect 229836 218016 229888 218068
rect 230388 218016 230440 218068
rect 232320 218016 232372 218068
rect 233148 218016 233200 218068
rect 233976 218016 234028 218068
rect 234528 218016 234580 218068
rect 242256 218016 242308 218068
rect 242716 218016 242768 218068
rect 248880 218016 248932 218068
rect 249616 218016 249668 218068
rect 254676 218016 254728 218068
rect 255136 218016 255188 218068
rect 258816 218016 258868 218068
rect 259368 218016 259420 218068
rect 265440 218016 265492 218068
rect 266268 218016 266320 218068
rect 269580 218016 269632 218068
rect 270132 218016 270184 218068
rect 273720 218016 273772 218068
rect 274272 218016 274324 218068
rect 282000 218016 282052 218068
rect 282552 218016 282604 218068
rect 284208 218016 284260 218068
rect 284944 218016 284996 218068
rect 287796 218016 287848 218068
rect 288348 218016 288400 218068
rect 290280 218016 290332 218068
rect 290924 218016 290976 218068
rect 296076 218016 296128 218068
rect 296628 218016 296680 218068
rect 297732 218016 297784 218068
rect 300032 218016 300084 218068
rect 300216 218016 300268 218068
rect 300768 218016 300820 218068
rect 304356 218016 304408 218068
rect 305644 218016 305696 218068
rect 308496 218016 308548 218068
rect 309048 218016 309100 218068
rect 310980 218016 311032 218068
rect 311808 218016 311860 218068
rect 312636 218016 312688 218068
rect 313096 218016 313148 218068
rect 315120 218016 315172 218068
rect 315672 218016 315724 218068
rect 317328 218016 317380 218068
rect 318064 218016 318116 218068
rect 319260 218016 319312 218068
rect 319996 218016 320048 218068
rect 333336 218016 333388 218068
rect 333888 218016 333940 218068
rect 335820 218016 335872 218068
rect 336464 218016 336516 218068
rect 339960 218016 340012 218068
rect 340696 218016 340748 218068
rect 341616 218016 341668 218068
rect 342076 218016 342128 218068
rect 345756 218016 345808 218068
rect 346216 218016 346268 218068
rect 348240 218016 348292 218068
rect 349068 218016 349120 218068
rect 352380 218016 352432 218068
rect 354312 218016 354364 218068
rect 356520 218016 356572 218068
rect 357256 218016 357308 218068
rect 360660 218016 360712 218068
rect 361304 218016 361356 218068
rect 364800 218016 364852 218068
rect 365536 218016 365588 218068
rect 366456 218016 366508 218068
rect 366916 218016 366968 218068
rect 368940 218016 368992 218068
rect 372528 218016 372580 218068
rect 372988 218016 373040 218068
rect 373816 218016 373868 218068
rect 374736 218016 374788 218068
rect 375288 218016 375340 218068
rect 381360 218016 381412 218068
rect 382096 218016 382148 218068
rect 385500 218016 385552 218068
rect 386328 218016 386380 218068
rect 389640 218016 389692 218068
rect 390192 218016 390244 218068
rect 393780 218016 393832 218068
rect 394516 218016 394568 218068
rect 397920 218016 397972 218068
rect 398564 218016 398616 218068
rect 399576 218016 399628 218068
rect 400036 218016 400088 218068
rect 403716 218016 403768 218068
rect 404176 218016 404228 218068
rect 410340 218016 410392 218068
rect 410892 218016 410944 218068
rect 416136 218016 416188 218068
rect 416688 218016 416740 218068
rect 418620 218016 418672 218068
rect 419448 218016 419500 218068
rect 420276 218016 420328 218068
rect 420828 218016 420880 218068
rect 422760 218016 422812 218068
rect 425428 218016 425480 218068
rect 426072 218016 426124 218068
rect 428464 218016 428516 218068
rect 429108 218016 429160 218068
rect 430672 218016 430724 218068
rect 432696 218016 432748 218068
rect 433800 218016 433852 218068
rect 434996 218016 435048 218068
rect 436284 218016 436336 218068
rect 436468 218016 436520 218068
rect 437480 218016 437532 218068
rect 438492 218016 438544 218068
rect 438952 218016 439004 218068
rect 440148 218016 440200 218068
rect 440700 218016 440752 218068
rect 453304 218016 453356 218068
rect 455420 218016 455472 218068
rect 462964 218016 463016 218068
rect 464344 218016 464396 218068
rect 467104 218016 467156 218068
rect 467840 218016 467892 218068
rect 471244 218016 471296 218068
rect 472624 218016 472676 218068
rect 480996 218016 481048 218068
rect 482560 218016 482612 218068
rect 482744 218016 482796 218068
rect 485044 218016 485096 218068
rect 495348 218016 495400 218068
rect 500224 218016 500276 218068
rect 502432 218016 502484 218068
rect 648252 218016 648304 218068
rect 654784 218016 654836 218068
rect 614488 217948 614540 218000
rect 565176 217880 565228 217932
rect 568304 217880 568356 217932
rect 572168 217880 572220 217932
rect 576032 217880 576084 217932
rect 576216 217880 576268 217932
rect 447140 217812 447192 217864
rect 447784 217812 447836 217864
rect 525800 217812 525852 217864
rect 526444 217812 526496 217864
rect 555700 217812 555752 217864
rect 562876 217812 562928 217864
rect 572352 217744 572404 217796
rect 576584 217744 576636 217796
rect 578240 217744 578292 217796
rect 561128 217676 561180 217728
rect 563244 217676 563296 217728
rect 605104 217676 605156 217728
rect 614120 217676 614172 217728
rect 553216 217540 553268 217592
rect 554228 217540 554280 217592
rect 563060 217540 563112 217592
rect 577320 217608 577372 217660
rect 597560 217540 597612 217592
rect 613384 217540 613436 217592
rect 576584 217472 576636 217524
rect 576952 217472 577004 217524
rect 591580 217472 591632 217524
rect 595720 217472 595772 217524
rect 611820 217404 611872 217456
rect 628288 217404 628340 217456
rect 571708 217336 571760 217388
rect 577136 217336 577188 217388
rect 594984 217268 595036 217320
rect 626080 217268 626132 217320
rect 563060 217200 563112 217252
rect 562692 217064 562744 217116
rect 572536 217064 572588 217116
rect 582380 217200 582432 217252
rect 591948 217200 592000 217252
rect 591764 217064 591816 217116
rect 595168 217064 595220 217116
rect 582564 216724 582616 216776
rect 663248 216112 663300 216164
rect 664444 216112 664496 216164
rect 622952 216044 623004 216096
rect 629944 216044 629996 216096
rect 577688 215908 577740 215960
rect 628840 215908 628892 215960
rect 655428 215296 655480 215348
rect 656164 215296 656216 215348
rect 577320 215092 577372 215144
rect 612280 215092 612332 215144
rect 675852 215092 675904 215144
rect 676864 215092 676916 215144
rect 577872 214956 577924 215008
rect 621848 214956 621900 215008
rect 578056 214820 578108 214872
rect 621112 214820 621164 214872
rect 621664 214820 621716 214872
rect 632888 214820 632940 214872
rect 578240 214684 578292 214736
rect 624424 214684 624476 214736
rect 648436 214684 648488 214736
rect 658924 214684 658976 214736
rect 577504 214548 577556 214600
rect 599032 214412 599084 214464
rect 599584 214412 599636 214464
rect 600412 214412 600464 214464
rect 601240 214412 601292 214464
rect 615500 214412 615552 214464
rect 616144 214412 616196 214464
rect 616880 214548 616932 214600
rect 617340 214548 617392 214600
rect 619640 214548 619692 214600
rect 620560 214548 620612 214600
rect 622584 214548 622636 214600
rect 623320 214548 623372 214600
rect 623780 214548 623832 214600
rect 623872 214412 623924 214464
rect 625252 214548 625304 214600
rect 625620 214548 625672 214600
rect 636292 214548 636344 214600
rect 639604 214548 639656 214600
rect 652760 214548 652812 214600
rect 665824 214548 665876 214600
rect 631600 214412 631652 214464
rect 675852 214412 675904 214464
rect 677416 214412 677468 214464
rect 600504 214276 600556 214328
rect 600872 214276 600924 214328
rect 41328 213936 41380 213988
rect 41696 213936 41748 213988
rect 638316 213868 638368 213920
rect 640616 213868 640668 213920
rect 648620 213868 648672 213920
rect 649264 213868 649316 213920
rect 650460 213868 650512 213920
rect 653128 213868 653180 213920
rect 660396 213868 660448 213920
rect 660948 213868 661000 213920
rect 641628 213732 641680 213784
rect 650644 213732 650696 213784
rect 660948 213732 661000 213784
rect 662972 213732 663024 213784
rect 640248 213596 640300 213648
rect 649724 213596 649776 213648
rect 651840 213596 651892 213648
rect 657544 213596 657596 213648
rect 676036 213528 676088 213580
rect 677048 213528 677100 213580
rect 635556 213460 635608 213512
rect 652392 213460 652444 213512
rect 638868 213324 638920 213376
rect 660212 213324 660264 213376
rect 642180 213188 642232 213240
rect 661500 213120 661552 213172
rect 666284 213120 666336 213172
rect 613016 212848 613068 212900
rect 615040 212848 615092 212900
rect 664260 212984 664312 213036
rect 665088 212984 665140 213036
rect 665456 212848 665508 212900
rect 632704 212712 632756 212764
rect 634360 212712 634412 212764
rect 658740 212712 658792 212764
rect 659568 212712 659620 212764
rect 601792 212372 601844 212424
rect 602344 212372 602396 212424
rect 603080 212372 603132 212424
rect 604000 212372 604052 212424
rect 604460 212372 604512 212424
rect 605104 212372 605156 212424
rect 41328 211284 41380 211336
rect 41696 211284 41748 211336
rect 41144 211148 41196 211200
rect 41512 211148 41564 211200
rect 578516 211148 578568 211200
rect 580908 211148 580960 211200
rect 603264 211012 603316 211064
rect 603632 211012 603684 211064
rect 605840 210060 605892 210112
rect 606208 210060 606260 210112
rect 622400 210060 622452 210112
rect 622768 210060 622820 210112
rect 578424 209788 578476 209840
rect 580080 209788 580132 209840
rect 580264 208564 580316 208616
rect 632152 209516 632204 209568
rect 652208 209652 652260 209704
rect 652024 209516 652076 209568
rect 666836 209176 666888 209228
rect 667020 209040 667072 209092
rect 578884 208292 578936 208344
rect 589464 208292 589516 208344
rect 580080 207612 580132 207664
rect 589648 207612 589700 207664
rect 580908 206864 580960 206916
rect 589464 206864 589516 206916
rect 579528 205776 579580 205828
rect 582380 205776 582432 205828
rect 579712 204212 579764 204264
rect 589464 204212 589516 204264
rect 578516 202920 578568 202972
rect 580448 202920 580500 202972
rect 582380 202784 582432 202836
rect 589464 202784 589516 202836
rect 578792 200132 578844 200184
rect 590384 200132 590436 200184
rect 580448 199996 580500 200048
rect 589464 199996 589516 200048
rect 579528 198704 579580 198756
rect 589464 198704 589516 198756
rect 578516 195984 578568 196036
rect 589280 195984 589332 196036
rect 579528 194556 579580 194608
rect 589464 194556 589516 194608
rect 668032 192448 668084 192500
rect 669320 192448 669372 192500
rect 579528 191836 579580 191888
rect 589464 191836 589516 191888
rect 579528 190476 579580 190528
rect 590568 190476 590620 190528
rect 669136 188436 669188 188488
rect 669320 188164 669372 188216
rect 579528 187688 579580 187740
rect 589464 187688 589516 187740
rect 579528 186260 579580 186312
rect 589648 186260 589700 186312
rect 579528 184832 579580 184884
rect 589464 184832 589516 184884
rect 667940 184492 667992 184544
rect 669596 184492 669648 184544
rect 579528 182112 579580 182164
rect 589464 182112 589516 182164
rect 578792 180752 578844 180804
rect 590568 180752 590620 180804
rect 578792 178032 578844 178084
rect 589464 178032 589516 178084
rect 579528 177896 579580 177948
rect 589648 177896 589700 177948
rect 582380 175244 582432 175296
rect 589464 175312 589516 175364
rect 667940 174836 667992 174888
rect 669780 174836 669832 174888
rect 578424 174496 578476 174548
rect 589648 174496 589700 174548
rect 578240 173204 578292 173256
rect 582380 173204 582432 173256
rect 578424 172456 578476 172508
rect 589464 172524 589516 172576
rect 579804 171096 579856 171148
rect 589464 171096 589516 171148
rect 668032 169668 668084 169720
rect 670332 169668 670384 169720
rect 582380 167016 582432 167068
rect 589464 167016 589516 167068
rect 579528 166268 579580 166320
rect 589188 166268 589240 166320
rect 667940 165180 667992 165232
rect 670148 165180 670200 165232
rect 579344 164840 579396 164892
rect 589832 164840 589884 164892
rect 580908 162868 580960 162920
rect 589464 162868 589516 162920
rect 578240 162528 578292 162580
rect 582380 162528 582432 162580
rect 675852 162528 675904 162580
rect 681004 162528 681056 162580
rect 578424 162120 578476 162172
rect 589648 162120 589700 162172
rect 582380 160080 582432 160132
rect 589464 160080 589516 160132
rect 667940 160012 667992 160064
rect 669964 160012 670016 160064
rect 583760 159332 583812 159384
rect 590568 159332 590620 159384
rect 578516 157564 578568 157616
rect 580908 157564 580960 157616
rect 587164 157360 587216 157412
rect 589280 157360 589332 157412
rect 585784 154572 585836 154624
rect 589464 154572 589516 154624
rect 578700 154164 578752 154216
rect 583760 154164 583812 154216
rect 584404 153212 584456 153264
rect 589464 153212 589516 153264
rect 578240 152600 578292 152652
rect 582380 152600 582432 152652
rect 583024 151784 583076 151836
rect 589464 151784 589516 151836
rect 578332 151036 578384 151088
rect 588544 151036 588596 151088
rect 668308 150220 668360 150272
rect 670792 150220 670844 150272
rect 579528 148316 579580 148368
rect 587164 148316 587216 148368
rect 585968 146276 586020 146328
rect 589464 146276 589516 146328
rect 578884 145528 578936 145580
rect 589188 145528 589240 145580
rect 579436 144644 579488 144696
rect 585784 144644 585836 144696
rect 587164 143556 587216 143608
rect 589464 143556 589516 143608
rect 579528 143420 579580 143472
rect 584404 143420 584456 143472
rect 583208 140768 583260 140820
rect 589464 140768 589516 140820
rect 579528 140564 579580 140616
rect 583024 140564 583076 140616
rect 584404 139408 584456 139460
rect 589464 139408 589516 139460
rect 578608 139272 578660 139324
rect 589924 139272 589976 139324
rect 579528 138116 579580 138168
rect 585968 138116 586020 138168
rect 580448 137368 580500 137420
rect 589648 137368 589700 137420
rect 579068 137232 579120 137284
rect 588728 137232 588780 137284
rect 585968 135260 586020 135312
rect 589464 135260 589516 135312
rect 581828 131860 581880 131912
rect 590292 131860 590344 131912
rect 578700 131724 578752 131776
rect 587164 131724 587216 131776
rect 587532 131112 587584 131164
rect 590108 131112 590160 131164
rect 578516 127984 578568 128036
rect 580448 127984 580500 128036
rect 579068 126964 579120 127016
rect 589464 126964 589516 127016
rect 580632 125604 580684 125656
rect 589464 125604 589516 125656
rect 579528 125332 579580 125384
rect 583208 125332 583260 125384
rect 583024 124856 583076 124908
rect 589280 124856 589332 124908
rect 579252 124108 579304 124160
rect 584404 124108 584456 124160
rect 584588 122816 584640 122868
rect 589464 122816 589516 122868
rect 578884 122204 578936 122256
rect 587532 122204 587584 122256
rect 580448 122068 580500 122120
rect 589740 122068 589792 122120
rect 587348 121456 587400 121508
rect 589280 121456 589332 121508
rect 578516 121320 578568 121372
rect 588544 121320 588596 121372
rect 667940 120708 667992 120760
rect 669780 120708 669832 120760
rect 579528 118396 579580 118448
rect 585968 118396 586020 118448
rect 667940 118056 667992 118108
rect 670148 118056 670200 118108
rect 585784 117308 585836 117360
rect 589464 117308 589516 117360
rect 675852 117240 675904 117292
rect 679624 117240 679676 117292
rect 579344 117172 579396 117224
rect 581828 117172 581880 117224
rect 585968 115948 586020 116000
rect 589464 115948 589516 116000
rect 578516 114452 578568 114504
rect 580264 114452 580316 114504
rect 588544 113704 588596 113756
rect 589556 113704 589608 113756
rect 579528 113092 579580 113144
rect 589924 113092 589976 113144
rect 667940 111392 667992 111444
rect 669964 111392 670016 111444
rect 583208 111052 583260 111104
rect 590292 111052 590344 111104
rect 581828 109692 581880 109744
rect 589372 109692 589424 109744
rect 578332 108672 578384 108724
rect 580632 108672 580684 108724
rect 583760 107652 583812 107704
rect 589464 107652 589516 107704
rect 580264 106292 580316 106344
rect 589464 106292 589516 106344
rect 668400 106156 668452 106208
rect 670792 106156 670844 106208
rect 579436 105136 579488 105188
rect 583760 105136 583812 105188
rect 587164 104864 587216 104916
rect 589832 104864 589884 104916
rect 579252 103300 579304 103352
rect 583024 103300 583076 103352
rect 578332 101668 578384 101720
rect 584588 101668 584640 101720
rect 584404 101396 584456 101448
rect 590292 101396 590344 101448
rect 624792 100104 624844 100156
rect 667940 100104 667992 100156
rect 614856 99900 614908 99952
rect 668124 99968 668176 100020
rect 578608 99288 578660 99340
rect 580448 99288 580500 99340
rect 622308 99288 622360 99340
rect 630772 99288 630824 99340
rect 623688 99152 623740 99204
rect 633532 99152 633584 99204
rect 625068 99016 625120 99068
rect 636292 99016 636344 99068
rect 627552 98880 627604 98932
rect 640708 98880 640760 98932
rect 579252 98744 579304 98796
rect 587348 98744 587400 98796
rect 629024 98744 629076 98796
rect 643652 98744 643704 98796
rect 580632 98608 580684 98660
rect 590108 98608 590160 98660
rect 647148 98608 647200 98660
rect 661960 98608 662012 98660
rect 630496 98472 630548 98524
rect 646596 98472 646648 98524
rect 631416 98200 631468 98252
rect 642180 98200 642232 98252
rect 581644 97928 581696 97980
rect 595260 98064 595312 98116
rect 592684 97928 592736 97980
rect 597560 97928 597612 97980
rect 618720 97928 618772 97980
rect 625804 97928 625856 97980
rect 629760 97928 629812 97980
rect 645308 97996 645360 98048
rect 592868 97792 592920 97844
rect 598204 97792 598256 97844
rect 628288 97792 628340 97844
rect 631416 97792 631468 97844
rect 633348 97792 633400 97844
rect 650552 97792 650604 97844
rect 653956 97792 654008 97844
rect 655060 97792 655112 97844
rect 659200 97792 659252 97844
rect 663892 97792 663944 97844
rect 590108 97656 590160 97708
rect 600412 97656 600464 97708
rect 626080 97656 626132 97708
rect 637764 97656 637816 97708
rect 643008 97656 643060 97708
rect 659752 97656 659804 97708
rect 659936 97656 659988 97708
rect 665364 97656 665416 97708
rect 583024 97520 583076 97572
rect 596180 97520 596232 97572
rect 623136 97520 623188 97572
rect 632060 97520 632112 97572
rect 634728 97520 634780 97572
rect 649080 97520 649132 97572
rect 651840 97520 651892 97572
rect 659568 97520 659620 97572
rect 577688 97384 577740 97436
rect 596732 97384 596784 97436
rect 605472 97384 605524 97436
rect 613384 97384 613436 97436
rect 620192 97384 620244 97436
rect 625988 97384 626040 97436
rect 632704 97384 632756 97436
rect 650184 97384 650236 97436
rect 658188 97384 658240 97436
rect 663064 97384 663116 97436
rect 577504 97248 577556 97300
rect 601884 97248 601936 97300
rect 612648 97248 612700 97300
rect 620284 97248 620336 97300
rect 621664 97248 621716 97300
rect 629300 97248 629352 97300
rect 631876 97248 631928 97300
rect 648620 97248 648672 97300
rect 650368 97248 650420 97300
rect 658280 97248 658332 97300
rect 634176 97112 634228 97164
rect 647608 97112 647660 97164
rect 656808 97112 656860 97164
rect 661408 97112 661460 97164
rect 615040 96976 615092 97028
rect 616144 96976 616196 97028
rect 626816 96976 626868 97028
rect 639236 96976 639288 97028
rect 644296 96976 644348 97028
rect 658832 96976 658884 97028
rect 612096 96908 612148 96960
rect 612648 96908 612700 96960
rect 617248 96908 617300 96960
rect 618168 96908 618220 96960
rect 613568 96840 613620 96892
rect 615040 96840 615092 96892
rect 624608 96840 624660 96892
rect 635004 96840 635056 96892
rect 654784 96840 654836 96892
rect 655428 96840 655480 96892
rect 660672 96840 660724 96892
rect 663248 96840 663300 96892
rect 615776 96772 615828 96824
rect 618904 96772 618956 96824
rect 606208 96704 606260 96756
rect 607128 96704 607180 96756
rect 610624 96704 610676 96756
rect 611176 96704 611228 96756
rect 638592 96704 638644 96756
rect 647240 96704 647292 96756
rect 655244 96704 655296 96756
rect 662512 96704 662564 96756
rect 639052 96568 639104 96620
rect 649264 96568 649316 96620
rect 653312 96568 653364 96620
rect 665180 96568 665232 96620
rect 640064 96432 640116 96484
rect 645124 96432 645176 96484
rect 645768 96432 645820 96484
rect 652024 96432 652076 96484
rect 652576 96432 652628 96484
rect 664168 96432 664220 96484
rect 640524 96296 640576 96348
rect 648436 96296 648488 96348
rect 648896 96296 648948 96348
rect 664352 96296 664404 96348
rect 637580 96160 637632 96212
rect 660672 96160 660724 96212
rect 641536 96024 641588 96076
rect 663708 96024 663760 96076
rect 609152 95888 609204 95940
rect 621664 95888 621716 95940
rect 644940 95888 644992 95940
rect 648068 95888 648120 95940
rect 648436 95888 648488 95940
rect 664536 95888 664588 95940
rect 645124 95752 645176 95804
rect 652208 95752 652260 95804
rect 646412 95616 646464 95668
rect 653404 95616 653456 95668
rect 648068 95480 648120 95532
rect 656164 95752 656216 95804
rect 631232 95412 631284 95464
rect 643468 95412 643520 95464
rect 647884 95412 647936 95464
rect 647148 95208 647200 95260
rect 579252 95140 579304 95192
rect 588728 95140 588780 95192
rect 620928 95140 620980 95192
rect 626448 95140 626500 95192
rect 647608 95140 647660 95192
rect 650000 95140 650052 95192
rect 616512 95004 616564 95056
rect 623228 95004 623280 95056
rect 648252 94732 648304 94784
rect 654784 94732 654836 94784
rect 596824 94528 596876 94580
rect 598940 94528 598992 94580
rect 607680 94460 607732 94512
rect 620928 94460 620980 94512
rect 619548 93780 619600 93832
rect 626448 93780 626500 93832
rect 651288 93508 651340 93560
rect 655428 93508 655480 93560
rect 579344 93100 579396 93152
rect 585784 93100 585836 93152
rect 611176 93100 611228 93152
rect 622400 93100 622452 93152
rect 617984 92420 618036 92472
rect 626448 92420 626500 92472
rect 578240 91808 578292 91860
rect 585968 91808 586020 91860
rect 606944 91740 606996 91792
rect 626264 91740 626316 91792
rect 647240 91672 647292 91724
rect 654692 91672 654744 91724
rect 610992 90992 611044 91044
rect 617524 90992 617576 91044
rect 618168 90992 618220 91044
rect 626448 90992 626500 91044
rect 649264 90652 649316 90704
rect 655428 90652 655480 90704
rect 584588 90312 584640 90364
rect 590108 90312 590160 90364
rect 620928 89632 620980 89684
rect 625436 89632 625488 89684
rect 623228 89496 623280 89548
rect 626448 89496 626500 89548
rect 649724 88748 649776 88800
rect 658556 88748 658608 88800
rect 662328 88748 662380 88800
rect 663892 88748 663944 88800
rect 579344 88272 579396 88324
rect 588544 88272 588596 88324
rect 617524 88272 617576 88324
rect 626448 88272 626500 88324
rect 655244 88272 655296 88324
rect 658464 88272 658516 88324
rect 659568 86912 659620 86964
rect 663248 86912 663300 86964
rect 653404 86844 653456 86896
rect 657176 86844 657228 86896
rect 647884 86708 647936 86760
rect 661408 86708 661460 86760
rect 656164 86572 656216 86624
rect 660672 86572 660724 86624
rect 578792 86436 578844 86488
rect 580632 86436 580684 86488
rect 652208 86436 652260 86488
rect 660120 86436 660172 86488
rect 622400 86300 622452 86352
rect 626448 86300 626500 86352
rect 654876 86300 654928 86352
rect 662512 86300 662564 86352
rect 652024 86164 652076 86216
rect 657728 86164 657780 86216
rect 609888 85484 609940 85536
rect 626448 85484 626500 85536
rect 621664 85348 621716 85400
rect 625252 85348 625304 85400
rect 608508 84124 608560 84176
rect 625804 84124 625856 84176
rect 579344 83988 579396 84040
rect 581828 83988 581880 84040
rect 581644 83444 581696 83496
rect 589924 83444 589976 83496
rect 578700 82764 578752 82816
rect 583208 82764 583260 82816
rect 578884 82084 578936 82136
rect 587164 82084 587216 82136
rect 628748 80928 628800 80980
rect 642456 80928 642508 80980
rect 618904 80792 618956 80844
rect 648988 80792 649040 80844
rect 595444 80656 595496 80708
rect 636752 80656 636804 80708
rect 629208 79976 629260 80028
rect 633440 79976 633492 80028
rect 614028 79432 614080 79484
rect 646044 79432 646096 79484
rect 588544 79296 588596 79348
rect 592868 79296 592920 79348
rect 612648 79296 612700 79348
rect 646320 79296 646372 79348
rect 578608 78208 578660 78260
rect 580264 78208 580316 78260
rect 633440 78208 633492 78260
rect 645308 78208 645360 78260
rect 631048 78072 631100 78124
rect 643100 78072 643152 78124
rect 615040 77936 615092 77988
rect 649172 77936 649224 77988
rect 622032 77256 622084 77308
rect 631048 77392 631100 77444
rect 628472 77256 628524 77308
rect 632796 77256 632848 77308
rect 578700 77188 578752 77240
rect 584588 77188 584640 77240
rect 616144 76644 616196 76696
rect 646872 76644 646924 76696
rect 579068 76508 579120 76560
rect 666560 76508 666612 76560
rect 621664 75896 621716 75948
rect 628472 75896 628524 75948
rect 618904 75624 618956 75676
rect 622032 75624 622084 75676
rect 620284 75420 620336 75472
rect 648804 75420 648856 75472
rect 607128 75284 607180 75336
rect 646504 75284 646556 75336
rect 613384 75148 613436 75200
rect 662604 75148 662656 75200
rect 579528 73108 579580 73160
rect 584404 73108 584456 73160
rect 579252 71476 579304 71528
rect 581644 71476 581696 71528
rect 579528 66240 579580 66292
rect 623044 66240 623096 66292
rect 578516 62024 578568 62076
rect 612004 62024 612056 62076
rect 579528 60664 579580 60716
rect 624424 60664 624476 60716
rect 579528 57876 579580 57928
rect 614856 57876 614908 57928
rect 579528 56516 579580 56568
rect 621664 56516 621716 56568
rect 576124 53048 576176 53100
rect 617524 53048 617576 53100
rect 464988 52776 465040 52828
rect 467012 52776 467064 52828
rect 463608 52640 463660 52692
rect 466828 52640 466880 52692
rect 464068 52504 464120 52556
rect 466460 52504 466512 52556
rect 459468 52368 459520 52420
rect 464988 52368 465040 52420
rect 465448 52368 465500 52420
rect 475384 52368 475436 52420
rect 475568 52368 475620 52420
rect 577688 52368 577740 52420
rect 457720 52232 457772 52284
rect 459744 52232 459796 52284
rect 462228 52232 462280 52284
rect 457904 52096 457956 52148
rect 460848 52096 460900 52148
rect 463148 52096 463200 52148
rect 465908 52232 465960 52284
rect 572076 52232 572128 52284
rect 625804 52232 625856 52284
rect 50344 51960 50396 52012
rect 130384 51960 130436 52012
rect 458088 51960 458140 52012
rect 460204 51960 460256 52012
rect 464528 51960 464580 52012
rect 49148 51824 49200 51876
rect 129372 51824 129424 51876
rect 47584 51688 47636 51740
rect 129004 51688 129056 51740
rect 145380 51688 145432 51740
rect 306012 51688 306064 51740
rect 576124 52096 576176 52148
rect 576308 52096 576360 52148
rect 583024 52096 583076 52148
rect 571708 52028 571760 52080
rect 464988 51960 465040 52012
rect 475200 51892 475252 51944
rect 475384 51892 475436 51944
rect 572076 51892 572128 51944
rect 600320 51756 600372 51808
rect 592684 51552 592736 51604
rect 466460 51416 466512 51468
rect 475200 51416 475252 51468
rect 475568 51280 475620 51332
rect 571708 51416 571760 51468
rect 578884 51416 578936 51468
rect 576308 51280 576360 51332
rect 467012 51008 467064 51060
rect 596824 51008 596876 51060
rect 466828 50872 466880 50924
rect 588544 50872 588596 50924
rect 50528 50600 50580 50652
rect 128452 50600 128504 50652
rect 47768 50464 47820 50516
rect 131028 50464 131080 50516
rect 318340 50464 318392 50516
rect 458272 50464 458324 50516
rect 46204 50328 46256 50380
rect 128636 50328 128688 50380
rect 314016 50328 314068 50380
rect 458456 50328 458508 50380
rect 521108 50328 521160 50380
rect 544016 50328 544068 50380
rect 467012 49376 467064 49428
rect 577504 49376 577556 49428
rect 48964 49240 49016 49292
rect 129556 49240 129608 49292
rect 466644 49240 466696 49292
rect 599124 49240 599176 49292
rect 45468 49104 45520 49156
rect 128820 49104 128872 49156
rect 466460 49104 466512 49156
rect 601700 49104 601752 49156
rect 46388 48968 46440 49020
rect 130476 48968 130528 49020
rect 466828 48968 466880 49020
rect 618904 48968 618956 49020
rect 128452 48084 128504 48136
rect 131948 48084 132000 48136
rect 128636 47812 128688 47864
rect 131764 47812 131816 47864
rect 623044 46452 623096 46504
rect 661592 46452 661644 46504
rect 129556 45024 129608 45076
rect 129004 44888 129056 44940
rect 129188 44752 129240 44804
rect 129372 44616 129424 44668
rect 131764 44684 131816 44736
rect 131948 44532 132000 44584
rect 132592 44276 132644 44328
rect 128820 44208 128872 44260
rect 130660 44072 130712 44124
rect 131028 43936 131080 43988
rect 43628 42780 43680 42832
rect 187332 43528 187384 43580
rect 431224 43596 431276 43648
rect 439596 43596 439648 43648
rect 441620 43596 441672 43648
rect 310428 42712 310480 42764
rect 431224 42712 431276 42764
rect 456064 42712 456116 42764
rect 463056 42712 463108 42764
rect 404452 42304 404504 42356
rect 405556 42304 405608 42356
rect 420736 42304 420788 42356
rect 427084 42304 427136 42356
rect 662420 42173 662472 42225
rect 431224 42032 431276 42084
rect 456064 42032 456116 42084
rect 404452 41420 404504 41472
rect 420736 41420 420788 41472
rect 427084 41420 427136 41472
rect 459192 41420 459244 41472
<< metal2 >>
rect 110170 1029098 110262 1029126
rect 212934 1029098 213026 1029126
rect 264362 1029098 264454 1029126
rect 315974 1029098 316066 1029126
rect 366390 1029098 366482 1029126
rect 433734 1029098 433826 1029126
rect 510738 1029098 510830 1029126
rect 562166 1029098 562258 1029126
rect 110170 1028622 110262 1028650
rect 212934 1028622 213026 1028650
rect 264362 1028622 264454 1028650
rect 315974 1028622 316066 1028650
rect 366390 1028622 366482 1028650
rect 433734 1028622 433826 1028650
rect 510738 1028622 510830 1028650
rect 562166 1028622 562258 1028650
rect 110170 1028177 110262 1028205
rect 212934 1028177 213026 1028205
rect 264362 1028177 264454 1028205
rect 315974 1028177 316066 1028205
rect 366390 1028177 366482 1028205
rect 433734 1028177 433826 1028205
rect 510738 1028177 510830 1028205
rect 562166 1028177 562258 1028205
rect 366180 1027880 366232 1027886
rect 366180 1027822 366232 1027828
rect 366548 1027880 366600 1027886
rect 366548 1027822 366600 1027828
rect 110170 1027738 110262 1027766
rect 212934 1027738 213026 1027766
rect 264362 1027738 264454 1027766
rect 315974 1027738 316066 1027766
rect 366192 1027752 366220 1027822
rect 366560 1027752 366588 1027822
rect 433734 1027738 433826 1027766
rect 510738 1027738 510830 1027766
rect 562166 1027738 562258 1027766
rect 110170 1027262 110262 1027290
rect 212934 1027262 213026 1027290
rect 264362 1027262 264454 1027290
rect 315974 1027262 316066 1027290
rect 366390 1027262 366482 1027290
rect 433734 1027262 433826 1027290
rect 510738 1027262 510830 1027290
rect 562166 1027262 562258 1027290
rect 110170 1026786 110262 1026814
rect 212934 1026786 213026 1026814
rect 264362 1026786 264454 1026814
rect 315974 1026786 316066 1026814
rect 366390 1026786 366482 1026814
rect 433734 1026786 433826 1026814
rect 510738 1026786 510830 1026814
rect 562166 1026786 562258 1026814
rect 110170 1026310 110262 1026338
rect 212934 1026310 213026 1026338
rect 264362 1026310 264454 1026338
rect 315974 1026310 316066 1026338
rect 366284 1026202 366312 1026324
rect 366468 1026202 366496 1026324
rect 433734 1026310 433826 1026338
rect 510738 1026310 510830 1026338
rect 562166 1026310 562258 1026338
rect 366284 1026174 366496 1026202
rect 366284 1026038 366496 1026066
rect 110170 1025902 110262 1025930
rect 212934 1025902 213026 1025930
rect 264362 1025902 264454 1025930
rect 315974 1025902 316066 1025930
rect 366284 1025916 366312 1026038
rect 366468 1025916 366496 1026038
rect 433734 1025902 433826 1025930
rect 510738 1025902 510830 1025930
rect 562166 1025902 562258 1025930
rect 110170 1025426 110262 1025454
rect 212934 1025426 213026 1025454
rect 264362 1025426 264454 1025454
rect 315974 1025426 316066 1025454
rect 366390 1025426 366482 1025454
rect 433734 1025426 433826 1025454
rect 510738 1025426 510830 1025454
rect 562166 1025426 562258 1025454
rect 110170 1024950 110262 1024978
rect 212934 1024950 213026 1024978
rect 264362 1024950 264454 1024978
rect 315974 1024950 316066 1024978
rect 366390 1024950 366482 1024978
rect 433734 1024950 433826 1024978
rect 510738 1024950 510830 1024978
rect 562166 1024950 562258 1024978
rect 110170 1024474 110262 1024502
rect 212934 1024474 213026 1024502
rect 264362 1024474 264454 1024502
rect 315974 1024474 316066 1024502
rect 366192 1024418 366220 1024488
rect 366560 1024418 366588 1024488
rect 433734 1024474 433826 1024502
rect 510738 1024474 510830 1024502
rect 562166 1024474 562258 1024502
rect 366180 1024412 366232 1024418
rect 366180 1024354 366232 1024360
rect 366548 1024412 366600 1024418
rect 366548 1024354 366600 1024360
rect 110170 1024037 110262 1024065
rect 212934 1024037 213026 1024065
rect 264362 1024037 264454 1024065
rect 315974 1024037 316066 1024065
rect 366390 1024037 366482 1024065
rect 433734 1024037 433826 1024065
rect 510738 1024037 510830 1024065
rect 562166 1024037 562258 1024065
rect 110170 1023590 110262 1023618
rect 212934 1023590 213026 1023618
rect 264362 1023590 264454 1023618
rect 315974 1023590 316066 1023618
rect 366390 1023590 366482 1023618
rect 433734 1023590 433826 1023618
rect 510738 1023590 510830 1023618
rect 562166 1023590 562258 1023618
rect 202694 1007448 202750 1007457
rect 200028 1007412 200080 1007418
rect 202694 1007383 202696 1007392
rect 200028 1007354 200080 1007360
rect 202748 1007383 202750 1007392
rect 202696 1007354 202748 1007360
rect 153750 1006632 153806 1006641
rect 145748 1006596 145800 1006602
rect 153750 1006567 153752 1006576
rect 145748 1006538 145800 1006544
rect 153804 1006567 153806 1006576
rect 153752 1006538 153804 1006544
rect 102322 1006496 102378 1006505
rect 93308 1006460 93360 1006466
rect 102322 1006431 102324 1006440
rect 93308 1006402 93360 1006408
rect 102376 1006431 102378 1006440
rect 145564 1006460 145616 1006466
rect 102324 1006402 102376 1006408
rect 145564 1006402 145616 1006408
rect 93124 1006052 93176 1006058
rect 93124 1005994 93176 1006000
rect 92664 1002516 92716 1002522
rect 92664 1002458 92716 1002464
rect 92296 998436 92348 998442
rect 92296 998378 92348 998384
rect 81254 995752 81310 995761
rect 81310 995710 81374 995738
rect 81254 995687 81310 995696
rect 86498 995616 86554 995625
rect 86342 995574 86498 995602
rect 87786 995616 87842 995625
rect 87538 995574 87786 995602
rect 86498 995551 86554 995560
rect 90178 995616 90234 995625
rect 90022 995574 90178 995602
rect 87786 995551 87842 995560
rect 90178 995551 90234 995560
rect 77050 995438 77248 995466
rect 77220 995353 77248 995438
rect 77206 995344 77262 995353
rect 77206 995279 77262 995288
rect 77680 994702 77708 995452
rect 77668 994696 77720 994702
rect 77668 994638 77720 994644
rect 78324 994566 78352 995452
rect 80164 994838 80192 995452
rect 80152 994832 80204 994838
rect 80152 994774 80204 994780
rect 78312 994560 78364 994566
rect 78312 994502 78364 994508
rect 80716 994430 80744 995452
rect 82004 994809 82032 995452
rect 84488 995081 84516 995452
rect 84474 995072 84530 995081
rect 84474 995007 84530 995016
rect 81990 994800 82046 994809
rect 81990 994735 82046 994744
rect 85040 994537 85068 995452
rect 85026 994528 85082 994537
rect 85026 994463 85082 994472
rect 80704 994424 80756 994430
rect 80704 994366 80756 994372
rect 85684 994265 85712 995452
rect 88734 995438 89024 995466
rect 88996 994294 89024 995438
rect 89364 995081 89392 995452
rect 91218 995438 91692 995466
rect 91664 995330 91692 995438
rect 92308 995330 92336 998378
rect 92480 997620 92532 997626
rect 92480 997562 92532 997568
rect 92492 997257 92520 997562
rect 92478 997248 92534 997257
rect 92478 997183 92534 997192
rect 92480 997008 92532 997014
rect 92676 996985 92704 1002458
rect 92480 996950 92532 996956
rect 92662 996976 92718 996985
rect 92492 996441 92520 996950
rect 92662 996911 92718 996920
rect 92478 996432 92534 996441
rect 92478 996367 92534 996376
rect 91664 995302 92336 995330
rect 89350 995072 89406 995081
rect 89350 995007 89406 995016
rect 93136 994430 93164 1005994
rect 93320 994702 93348 1006402
rect 101954 1006360 102010 1006369
rect 101954 1006295 101956 1006304
rect 102008 1006295 102010 1006304
rect 144184 1006324 144236 1006330
rect 101956 1006266 102008 1006272
rect 144184 1006266 144236 1006272
rect 103978 1006224 104034 1006233
rect 101404 1006188 101456 1006194
rect 103978 1006159 103980 1006168
rect 101404 1006130 101456 1006136
rect 104032 1006159 104034 1006168
rect 107658 1006224 107714 1006233
rect 107658 1006159 107660 1006168
rect 103980 1006130 104032 1006136
rect 107712 1006159 107714 1006168
rect 124864 1006188 124916 1006194
rect 107660 1006130 107712 1006136
rect 124864 1006130 124916 1006136
rect 98274 1006088 98330 1006097
rect 94504 1006052 94556 1006058
rect 98274 1006023 98276 1006032
rect 94504 1005994 94556 1006000
rect 98328 1006023 98330 1006032
rect 98276 1005994 98328 1006000
rect 94516 996713 94544 1005994
rect 100298 1002688 100354 1002697
rect 97448 1002652 97500 1002658
rect 100298 1002623 100300 1002632
rect 97448 1002594 97500 1002600
rect 100352 1002623 100354 1002632
rect 100300 1002594 100352 1002600
rect 97264 1002380 97316 1002386
rect 97264 1002322 97316 1002328
rect 95884 1002108 95936 1002114
rect 95884 1002050 95936 1002056
rect 95148 999184 95200 999190
rect 95148 999126 95200 999132
rect 94502 996704 94558 996713
rect 94502 996639 94558 996648
rect 93308 994696 93360 994702
rect 93308 994638 93360 994644
rect 93124 994424 93176 994430
rect 93124 994366 93176 994372
rect 88984 994288 89036 994294
rect 85670 994256 85726 994265
rect 95160 994265 95188 999126
rect 88984 994230 89036 994236
rect 95146 994256 95202 994265
rect 85670 994191 85726 994200
rect 95146 994191 95202 994200
rect 51724 993200 51776 993206
rect 51724 993142 51776 993148
rect 50344 993064 50396 993070
rect 50344 993006 50396 993012
rect 47584 991772 47636 991778
rect 47584 991714 47636 991720
rect 44824 990140 44876 990146
rect 44824 990082 44876 990088
rect 43444 975724 43496 975730
rect 43444 975666 43496 975672
rect 42168 968833 42196 969272
rect 42154 968824 42210 968833
rect 42154 968759 42210 968768
rect 42168 967609 42196 968048
rect 42154 967600 42210 967609
rect 42154 967535 42210 967544
rect 42798 967600 42854 967609
rect 42798 967535 42854 967544
rect 41984 967201 42012 967405
rect 41970 967192 42026 967201
rect 41970 967127 42026 967136
rect 42430 966784 42486 966793
rect 42182 966742 42430 966770
rect 42430 966719 42486 966728
rect 42812 966014 42840 967535
rect 43456 966793 43484 975666
rect 44546 968824 44602 968833
rect 44546 968759 44602 968768
rect 43442 966784 43498 966793
rect 43442 966719 43498 966728
rect 42720 965986 42840 966014
rect 42182 965551 42472 965579
rect 42444 964753 42472 965551
rect 42430 964744 42486 964753
rect 42430 964679 42486 964688
rect 42182 964362 42472 964390
rect 42444 963937 42472 964362
rect 42430 963928 42486 963937
rect 42430 963863 42486 963872
rect 42182 963711 42472 963739
rect 42444 963393 42472 963711
rect 42720 963506 42748 965986
rect 44362 964744 44418 964753
rect 44362 964679 44418 964688
rect 44178 963928 44234 963937
rect 44178 963863 44234 963872
rect 42720 963478 42840 963506
rect 42430 963384 42486 963393
rect 42430 963319 42486 963328
rect 42812 963234 42840 963478
rect 43166 963384 43222 963393
rect 43166 963319 43222 963328
rect 42720 963206 42840 963234
rect 42430 963112 42486 963121
rect 42182 963070 42430 963098
rect 42430 963047 42486 963056
rect 41800 962169 41828 962540
rect 41786 962160 41842 962169
rect 41786 962095 41842 962104
rect 41800 959857 41828 960024
rect 41786 959848 41842 959857
rect 41786 959783 41842 959792
rect 41800 959177 41828 959412
rect 41786 959168 41842 959177
rect 42720 959114 42748 963206
rect 42982 963112 43038 963121
rect 42982 963047 43038 963056
rect 41786 959103 41842 959112
rect 42628 959086 42748 959114
rect 42168 958854 42288 958882
rect 42168 958732 42196 958854
rect 42260 958746 42288 958854
rect 42430 958760 42486 958769
rect 42260 958718 42430 958746
rect 42430 958695 42486 958704
rect 42076 957953 42104 958188
rect 42062 957944 42118 957953
rect 42062 957879 42118 957888
rect 42182 956338 42380 956366
rect 41800 955505 41828 955740
rect 41786 955496 41842 955505
rect 41786 955431 41842 955440
rect 42168 955182 42288 955210
rect 42168 955060 42196 955182
rect 42260 953594 42288 955182
rect 41708 953566 42288 953594
rect 28538 952912 28594 952921
rect 28538 952847 28594 952856
rect 8588 944180 8616 944316
rect 9048 944180 9076 944316
rect 9508 944180 9536 944316
rect 9968 944180 9996 944316
rect 10428 944180 10456 944316
rect 10888 944180 10916 944316
rect 11348 944180 11376 944316
rect 11808 944180 11836 944316
rect 12268 944180 12296 944316
rect 12728 944180 12756 944316
rect 13188 944180 13216 944316
rect 13648 944180 13676 944316
rect 14108 944180 14136 944316
rect 28552 942721 28580 952847
rect 41708 952474 41736 953566
rect 36544 952468 36596 952474
rect 36544 952410 36596 952416
rect 41696 952468 41748 952474
rect 41696 952410 41748 952416
rect 28538 942712 28594 942721
rect 28538 942647 28594 942656
rect 36556 938471 36584 952410
rect 42352 952354 42380 956338
rect 42628 953594 42656 959086
rect 42628 953566 42748 953594
rect 41708 952326 42380 952354
rect 41708 952270 41736 952326
rect 37924 952264 37976 952270
rect 41696 952264 41748 952270
rect 37924 952206 37976 952212
rect 39302 952232 39358 952241
rect 37936 939049 37964 952206
rect 41696 952206 41748 952212
rect 39302 952167 39358 952176
rect 37922 939040 37978 939049
rect 37922 938975 37978 938984
rect 36542 938462 36598 938471
rect 36542 938397 36598 938406
rect 39316 937417 39344 952167
rect 42062 951960 42118 951969
rect 42062 951895 42118 951904
rect 40038 951824 40094 951833
rect 40038 951759 40094 951768
rect 39302 937408 39358 937417
rect 39302 937343 39358 937352
rect 40052 934561 40080 951759
rect 41418 951688 41474 951697
rect 41418 951623 41474 951632
rect 41234 943120 41290 943129
rect 41234 943055 41290 943064
rect 41248 942614 41276 943055
rect 41236 942608 41288 942614
rect 41236 942550 41288 942556
rect 41234 941896 41290 941905
rect 41234 941831 41290 941840
rect 41248 941254 41276 941831
rect 41236 941248 41288 941254
rect 41236 941190 41288 941196
rect 41142 939448 41198 939457
rect 41142 939383 41198 939392
rect 40960 938664 41012 938670
rect 40960 938606 41012 938612
rect 40972 938471 41000 938606
rect 40958 938462 41014 938471
rect 41156 938466 41184 939383
rect 41432 938670 41460 951623
rect 41696 942608 41748 942614
rect 41748 942556 41920 942562
rect 41696 942550 41920 942556
rect 41708 942534 41920 942550
rect 41696 941248 41748 941254
rect 41696 941190 41748 941196
rect 41420 938664 41472 938670
rect 41420 938606 41472 938612
rect 40958 938397 41014 938406
rect 41144 938460 41196 938466
rect 41144 938402 41196 938408
rect 41512 938460 41564 938466
rect 41512 938402 41564 938408
rect 40038 934552 40094 934561
rect 40038 934487 40094 934496
rect 41524 911713 41552 938402
rect 41708 911985 41736 941190
rect 41892 937034 41920 942534
rect 42076 937825 42104 951895
rect 42720 943934 42748 953566
rect 42260 943906 42748 943934
rect 42062 937816 42118 937825
rect 42062 937751 42118 937760
rect 41892 937006 42104 937034
rect 42076 935785 42104 937006
rect 42062 935776 42118 935785
rect 42062 935711 42118 935720
rect 42260 932929 42288 943906
rect 42996 934153 43024 963047
rect 43180 934969 43208 963319
rect 43444 961920 43496 961926
rect 43444 961862 43496 961868
rect 43456 952921 43484 961862
rect 43718 958760 43774 958769
rect 43718 958695 43774 958704
rect 43442 952912 43498 952921
rect 43442 952847 43498 952856
rect 43534 940264 43590 940273
rect 43534 940199 43590 940208
rect 43166 934960 43222 934969
rect 43166 934895 43222 934904
rect 42982 934144 43038 934153
rect 42982 934079 43038 934088
rect 42246 932920 42302 932929
rect 42246 932855 42302 932864
rect 43350 932104 43406 932113
rect 43350 932039 43406 932048
rect 41694 911976 41750 911985
rect 41694 911911 41750 911920
rect 41510 911704 41566 911713
rect 41510 911639 41566 911648
rect 42936 892528 42992 892537
rect 42936 892463 42992 892472
rect 42950 892328 42978 892463
rect 42938 892322 42990 892328
rect 42938 892264 42990 892270
rect 43074 891984 43130 891993
rect 43074 891919 43076 891928
rect 43128 891919 43130 891928
rect 43076 891890 43128 891896
rect 41602 885456 41658 885465
rect 41602 885391 41658 885400
rect 41418 885184 41474 885193
rect 41418 885119 41474 885128
rect 8588 818380 8616 818516
rect 9048 818380 9076 818516
rect 9508 818380 9536 818516
rect 9968 818380 9996 818516
rect 10428 818380 10456 818516
rect 10888 818380 10916 818516
rect 11348 818380 11376 818516
rect 11808 818380 11836 818516
rect 12268 818380 12296 818516
rect 12728 818380 12756 818516
rect 13188 818380 13216 818516
rect 13648 818380 13676 818516
rect 14108 818380 14136 818516
rect 41234 817320 41290 817329
rect 41234 817255 41290 817264
rect 41248 817086 41276 817255
rect 41236 817080 41288 817086
rect 41236 817022 41288 817028
rect 41234 816504 41290 816513
rect 41234 816439 41290 816448
rect 41248 815658 41276 816439
rect 41236 815652 41288 815658
rect 41236 815594 41288 815600
rect 41432 814042 41460 885119
rect 41616 823874 41644 885391
rect 42062 884640 42118 884649
rect 42062 884575 42118 884584
rect 42076 823874 42104 884575
rect 41524 823846 41644 823874
rect 41708 823846 42104 823874
rect 41524 815674 41552 823846
rect 41708 817086 41736 823846
rect 41696 817080 41748 817086
rect 41696 817022 41748 817028
rect 41524 815658 41644 815674
rect 41524 815652 41656 815658
rect 41524 815646 41604 815652
rect 41604 815594 41656 815600
rect 41786 814056 41842 814065
rect 41432 814014 41786 814042
rect 41786 813991 41842 814000
rect 40958 813240 41014 813249
rect 40958 813175 41014 813184
rect 40774 812832 40830 812841
rect 40774 812767 40830 812776
rect 39302 811608 39358 811617
rect 39302 811543 39358 811552
rect 33046 811200 33102 811209
rect 33046 811135 33102 811144
rect 33060 802466 33088 811135
rect 33048 802460 33100 802466
rect 33048 802402 33100 802408
rect 39316 801786 39344 811543
rect 40788 810762 40816 812767
rect 40776 810756 40828 810762
rect 40776 810698 40828 810704
rect 40972 805633 41000 813175
rect 41142 812424 41198 812433
rect 41142 812359 41198 812368
rect 41156 807430 41184 812359
rect 41696 810756 41748 810762
rect 41696 810698 41748 810704
rect 41708 809146 41736 810698
rect 42982 810384 43038 810393
rect 42982 810319 43038 810328
rect 41708 809118 42472 809146
rect 41970 808344 42026 808353
rect 41970 808279 42026 808288
rect 41144 807424 41196 807430
rect 41144 807366 41196 807372
rect 41604 807424 41656 807430
rect 41604 807366 41656 807372
rect 41616 807242 41644 807366
rect 41786 807256 41842 807265
rect 41616 807214 41786 807242
rect 41786 807191 41842 807200
rect 40958 805624 41014 805633
rect 40958 805559 41014 805568
rect 41984 805089 42012 808279
rect 42246 806712 42302 806721
rect 42246 806647 42302 806656
rect 41970 805080 42026 805089
rect 41970 805015 42026 805024
rect 41696 802460 41748 802466
rect 41696 802402 41748 802408
rect 41708 802346 41736 802402
rect 41708 802318 41828 802346
rect 39304 801780 39356 801786
rect 39304 801722 39356 801728
rect 41604 801712 41656 801718
rect 41602 801680 41604 801689
rect 41656 801680 41658 801689
rect 41602 801615 41658 801624
rect 41800 800329 41828 802318
rect 41786 800320 41842 800329
rect 41786 800255 41842 800264
rect 41786 799912 41842 799921
rect 41786 799847 41842 799856
rect 41800 799445 41828 799847
rect 42260 799354 42288 806647
rect 42444 801794 42472 809118
rect 42798 807936 42854 807945
rect 42798 807871 42854 807880
rect 42168 799326 42288 799354
rect 42352 801766 42472 801794
rect 42168 798946 42196 799326
rect 42168 798918 42288 798946
rect 42260 798266 42288 798918
rect 42182 798238 42288 798266
rect 42352 797619 42380 801766
rect 42614 801680 42670 801689
rect 42614 801615 42670 801624
rect 42182 797591 42380 797619
rect 42154 797328 42210 797337
rect 42154 797263 42210 797272
rect 42168 796960 42196 797263
rect 42154 796240 42210 796249
rect 42154 796175 42210 796184
rect 42168 795765 42196 796175
rect 42628 795682 42656 801615
rect 42812 796362 42840 807871
rect 42536 795654 42656 795682
rect 42720 796334 42840 796362
rect 42062 795016 42118 795025
rect 42062 794951 42118 794960
rect 42076 794580 42104 794951
rect 41786 794472 41842 794481
rect 41786 794407 41842 794416
rect 41800 793900 41828 794407
rect 41786 793792 41842 793801
rect 41786 793727 41842 793736
rect 41800 793288 41828 793727
rect 42536 792758 42564 795654
rect 42720 795025 42748 796334
rect 42706 795016 42762 795025
rect 42706 794951 42762 794960
rect 42996 794894 43024 810319
rect 43166 809568 43222 809577
rect 43166 809503 43222 809512
rect 43180 796249 43208 809503
rect 43166 796240 43222 796249
rect 43166 796175 43222 796184
rect 42182 792730 42564 792758
rect 42812 794866 43024 794894
rect 42246 792568 42302 792577
rect 42246 792503 42302 792512
rect 42260 790650 42288 792503
rect 42430 792296 42486 792305
rect 42430 792231 42486 792240
rect 42168 790622 42288 790650
rect 42168 790228 42196 790622
rect 42444 789630 42472 792231
rect 42182 789602 42472 789630
rect 42812 789449 42840 794866
rect 42154 789440 42210 789449
rect 42154 789375 42210 789384
rect 42798 789440 42854 789449
rect 42798 789375 42854 789384
rect 42168 788936 42196 789375
rect 42338 789168 42394 789177
rect 42338 789103 42394 789112
rect 42352 788406 42380 789103
rect 42614 788760 42670 788769
rect 42614 788695 42670 788704
rect 42182 788378 42380 788406
rect 42246 788216 42302 788225
rect 42246 788151 42302 788160
rect 42430 788216 42486 788225
rect 42430 788151 42486 788160
rect 42260 786570 42288 788151
rect 42182 786542 42288 786570
rect 42444 785958 42472 788151
rect 42168 785890 42196 785944
rect 42260 785930 42472 785958
rect 42260 785890 42288 785930
rect 42168 785862 42288 785890
rect 42628 785278 42656 788695
rect 42798 788624 42854 788633
rect 42798 788559 42854 788568
rect 42812 788406 42840 788559
rect 42182 785250 42656 785278
rect 42720 788378 42840 788406
rect 42720 779714 42748 788378
rect 41708 779686 42748 779714
rect 8588 775132 8616 775268
rect 9048 775132 9076 775268
rect 9508 775132 9536 775268
rect 9968 775132 9996 775268
rect 10428 775132 10456 775268
rect 10888 775132 10916 775268
rect 11348 775132 11376 775268
rect 11808 775132 11836 775268
rect 12268 775132 12296 775268
rect 12728 775132 12756 775268
rect 13188 775132 13216 775268
rect 13648 775132 13676 775268
rect 14108 775132 14136 775268
rect 35806 773936 35862 773945
rect 35806 773871 35862 773880
rect 35820 772886 35848 773871
rect 41708 772886 41736 779686
rect 35808 772880 35860 772886
rect 35808 772822 35860 772828
rect 41696 772880 41748 772886
rect 41696 772822 41748 772828
rect 35346 769448 35402 769457
rect 35346 769383 35402 769392
rect 35360 768738 35388 769383
rect 35530 769040 35586 769049
rect 35530 768975 35586 768984
rect 35806 769040 35862 769049
rect 35806 768975 35808 768984
rect 35544 768874 35572 768975
rect 35860 768975 35862 768984
rect 40040 769004 40092 769010
rect 35808 768946 35860 768952
rect 40040 768946 40092 768952
rect 35532 768868 35584 768874
rect 35532 768810 35584 768816
rect 39304 768868 39356 768874
rect 39304 768810 39356 768816
rect 35348 768732 35400 768738
rect 35348 768674 35400 768680
rect 35622 768224 35678 768233
rect 35622 768159 35678 768168
rect 31022 767816 31078 767825
rect 31022 767751 31078 767760
rect 31036 759694 31064 767751
rect 35636 767378 35664 768159
rect 35806 767816 35862 767825
rect 35806 767751 35862 767760
rect 35820 767514 35848 767751
rect 35808 767508 35860 767514
rect 35808 767450 35860 767456
rect 36544 767508 36596 767514
rect 36544 767450 36596 767456
rect 35624 767372 35676 767378
rect 35624 767314 35676 767320
rect 35162 767000 35218 767009
rect 35162 766935 35218 766944
rect 31024 759688 31076 759694
rect 31024 759630 31076 759636
rect 35176 758334 35204 766935
rect 35806 763328 35862 763337
rect 35806 763263 35808 763272
rect 35860 763263 35862 763272
rect 35808 763234 35860 763240
rect 36556 759121 36584 767450
rect 37924 763292 37976 763298
rect 37924 763234 37976 763240
rect 36542 759112 36598 759121
rect 36542 759047 36598 759056
rect 35164 758328 35216 758334
rect 35164 758270 35216 758276
rect 37936 757790 37964 763234
rect 37924 757784 37976 757790
rect 39316 757761 39344 768810
rect 40052 764794 40080 768946
rect 41696 768732 41748 768738
rect 41696 768674 41748 768680
rect 41328 767372 41380 767378
rect 41328 767314 41380 767320
rect 41340 765377 41368 767314
rect 41708 765914 41736 768674
rect 43074 766728 43130 766737
rect 43074 766663 43130 766672
rect 41708 765886 42288 765914
rect 41326 765368 41382 765377
rect 41326 765303 41382 765312
rect 40040 764788 40092 764794
rect 40040 764730 40092 764736
rect 41696 764788 41748 764794
rect 41696 764730 41748 764736
rect 41708 764266 41736 764730
rect 42260 764402 42288 765886
rect 42522 765368 42578 765377
rect 42522 765303 42578 765312
rect 42536 764402 42564 765303
rect 42798 764688 42854 764697
rect 42798 764623 42854 764632
rect 42260 764374 42380 764402
rect 42536 764374 42748 764402
rect 41708 764238 42288 764266
rect 42260 761774 42288 764238
rect 42168 761746 42288 761774
rect 41696 759688 41748 759694
rect 41696 759630 41748 759636
rect 40316 758328 40368 758334
rect 40316 758270 40368 758276
rect 40328 758033 40356 758270
rect 41708 758146 41736 759630
rect 41708 758118 42012 758146
rect 40314 758024 40370 758033
rect 40314 757959 40370 757968
rect 40316 757784 40368 757790
rect 37924 757726 37976 757732
rect 39302 757752 39358 757761
rect 40316 757726 40368 757732
rect 41984 757738 42012 758118
rect 42168 757897 42196 761746
rect 42352 761682 42380 764374
rect 42720 763154 42748 764374
rect 42628 763126 42748 763154
rect 42628 761774 42656 763126
rect 42628 761746 42748 761774
rect 42260 761654 42380 761682
rect 42260 759506 42288 761654
rect 42260 759478 42472 759506
rect 42154 757888 42210 757897
rect 42154 757823 42210 757832
rect 39302 757687 39358 757696
rect 40328 757489 40356 757726
rect 41984 757710 42288 757738
rect 40314 757480 40370 757489
rect 40314 757415 40370 757424
rect 42260 756254 42288 757710
rect 42168 756226 42288 756254
rect 41786 755440 41842 755449
rect 41786 755375 41842 755384
rect 41800 755072 41828 755375
rect 42444 754474 42472 759478
rect 42720 756922 42748 761746
rect 42352 754446 42472 754474
rect 42536 756894 42748 756922
rect 42352 754406 42380 754446
rect 42182 754378 42380 754406
rect 42062 754080 42118 754089
rect 42062 754015 42118 754024
rect 42076 753780 42104 754015
rect 42246 753672 42302 753681
rect 42246 753607 42302 753616
rect 41970 752992 42026 753001
rect 41970 752927 42026 752936
rect 41984 752556 42012 752927
rect 42260 752049 42288 753607
rect 42536 753522 42564 756894
rect 42352 753494 42564 753522
rect 42352 752162 42380 753494
rect 42614 753400 42670 753409
rect 42614 753335 42670 753344
rect 42352 752134 42564 752162
rect 42246 752040 42302 752049
rect 42246 751975 42302 751984
rect 42536 751890 42564 752134
rect 42260 751862 42564 751890
rect 42062 751768 42118 751777
rect 42062 751703 42118 751712
rect 42076 751369 42104 751703
rect 41786 751088 41842 751097
rect 41786 751023 41842 751032
rect 41800 750720 41828 751023
rect 41786 750408 41842 750417
rect 41786 750343 41842 750352
rect 41800 750108 41828 750343
rect 42260 749986 42288 751862
rect 42168 749958 42288 749986
rect 42168 749529 42196 749958
rect 42246 749456 42302 749465
rect 42246 749391 42302 749400
rect 42260 749170 42288 749391
rect 42430 749320 42486 749329
rect 42430 749255 42486 749264
rect 42260 749142 42380 749170
rect 42352 747062 42380 749142
rect 42182 747034 42380 747062
rect 42444 746722 42472 749255
rect 42076 746694 42472 746722
rect 42076 746401 42104 746694
rect 42246 746600 42302 746609
rect 42246 746535 42302 746544
rect 41970 746056 42026 746065
rect 41970 745991 42026 746000
rect 41984 745756 42012 745991
rect 42062 745512 42118 745521
rect 42062 745447 42118 745456
rect 42076 745212 42104 745447
rect 42260 743390 42288 746535
rect 42430 746328 42486 746337
rect 42430 746263 42486 746272
rect 42182 743362 42288 743390
rect 42168 742750 42288 742778
rect 42168 742696 42196 742750
rect 42260 742710 42288 742750
rect 42444 742710 42472 746263
rect 42628 745521 42656 753335
rect 42812 751777 42840 764623
rect 42798 751768 42854 751777
rect 42798 751703 42854 751712
rect 43088 749329 43116 766663
rect 43074 749320 43130 749329
rect 43074 749255 43130 749264
rect 42614 745512 42670 745521
rect 42614 745447 42670 745456
rect 42706 745104 42762 745113
rect 42260 742682 42472 742710
rect 42536 745062 42706 745090
rect 42536 742098 42564 745062
rect 42706 745039 42762 745048
rect 42706 743064 42762 743073
rect 42706 742999 42762 743008
rect 42182 742070 42564 742098
rect 42720 736934 42748 742999
rect 41708 736906 42748 736934
rect 8588 731884 8616 732020
rect 9048 731884 9076 732020
rect 9508 731884 9536 732020
rect 9968 731884 9996 732020
rect 10428 731884 10456 732020
rect 10888 731884 10916 732020
rect 11348 731884 11376 732020
rect 11808 731884 11836 732020
rect 12268 731884 12296 732020
rect 12728 731884 12756 732020
rect 13188 731884 13216 732020
rect 13648 731884 13676 732020
rect 14108 731884 14136 732020
rect 35806 730960 35862 730969
rect 35806 730895 35862 730904
rect 35820 730114 35848 730895
rect 41708 730114 41736 736906
rect 35808 730108 35860 730114
rect 35808 730050 35860 730056
rect 41696 730108 41748 730114
rect 41696 730050 41748 730056
rect 41326 726472 41382 726481
rect 41326 726407 41382 726416
rect 41142 726064 41198 726073
rect 41142 725999 41198 726008
rect 39302 725248 39358 725257
rect 39302 725183 39358 725192
rect 36542 724840 36598 724849
rect 36542 724775 36598 724784
rect 31666 724432 31722 724441
rect 31666 724367 31722 724376
rect 31680 715465 31708 724367
rect 34518 724024 34574 724033
rect 34518 723959 34574 723968
rect 34150 720352 34206 720361
rect 34150 720287 34152 720296
rect 34204 720287 34206 720296
rect 34152 720258 34204 720264
rect 34532 715562 34560 723959
rect 36556 717398 36584 724775
rect 38660 720316 38712 720322
rect 38660 720258 38712 720264
rect 36544 717392 36596 717398
rect 36544 717334 36596 717340
rect 34520 715556 34572 715562
rect 34520 715498 34572 715504
rect 31666 715456 31722 715465
rect 31666 715391 31722 715400
rect 38672 714513 38700 720258
rect 39316 716242 39344 725183
rect 40682 723208 40738 723217
rect 40682 723143 40738 723152
rect 39304 716236 39356 716242
rect 39304 716178 39356 716184
rect 40316 715556 40368 715562
rect 40316 715498 40368 715504
rect 40328 715193 40356 715498
rect 40314 715184 40370 715193
rect 40314 715119 40370 715128
rect 38658 714504 38714 714513
rect 38658 714439 38714 714448
rect 40696 714241 40724 723143
rect 41156 721777 41184 725999
rect 41340 725966 41368 726407
rect 41328 725960 41380 725966
rect 41328 725902 41380 725908
rect 41696 725960 41748 725966
rect 41748 725908 41920 725914
rect 41696 725902 41920 725908
rect 41708 725886 41920 725902
rect 41326 725656 41382 725665
rect 41326 725591 41382 725600
rect 41340 724810 41368 725591
rect 41328 724804 41380 724810
rect 41328 724746 41380 724752
rect 41696 724804 41748 724810
rect 41696 724746 41748 724752
rect 41142 721768 41198 721777
rect 41142 721703 41198 721712
rect 41708 719137 41736 724746
rect 41892 719545 41920 725886
rect 43074 719808 43130 719817
rect 43074 719743 43130 719752
rect 41878 719536 41934 719545
rect 41878 719471 41934 719480
rect 42522 719536 42578 719545
rect 42522 719471 42578 719480
rect 41694 719128 41750 719137
rect 41694 719063 41750 719072
rect 41696 717392 41748 717398
rect 41696 717334 41748 717340
rect 41512 716236 41564 716242
rect 41512 716178 41564 716184
rect 41524 714241 41552 716178
rect 41708 716122 41736 717334
rect 41616 716094 41736 716122
rect 41616 714854 41644 716094
rect 42338 715184 42394 715193
rect 42338 715119 42394 715128
rect 41616 714826 41736 714854
rect 41708 714626 41736 714826
rect 41708 714598 41828 714626
rect 40682 714232 40738 714241
rect 40682 714167 40738 714176
rect 41510 714232 41566 714241
rect 41510 714167 41566 714176
rect 41800 713969 41828 714598
rect 42062 714504 42118 714513
rect 42118 714462 42288 714490
rect 42062 714439 42118 714448
rect 41786 713960 41842 713969
rect 41786 713895 41842 713904
rect 41786 713552 41842 713561
rect 41786 713487 41842 713496
rect 41800 713048 41828 713487
rect 42260 712314 42288 714462
rect 42168 712286 42288 712314
rect 42168 711824 42196 712286
rect 42154 711376 42210 711385
rect 42154 711311 42210 711320
rect 42168 711212 42196 711311
rect 42154 711104 42210 711113
rect 42154 711039 42210 711048
rect 42168 710561 42196 711039
rect 42352 710002 42380 715119
rect 42536 714854 42564 719471
rect 42706 719128 42762 719137
rect 42706 719063 42762 719072
rect 42444 714826 42564 714854
rect 42444 714354 42472 714826
rect 42720 714490 42748 719063
rect 42720 714462 42840 714490
rect 42444 714326 42564 714354
rect 42536 711498 42564 714326
rect 42536 711470 42656 711498
rect 42628 711385 42656 711470
rect 42614 711376 42670 711385
rect 42614 711311 42670 711320
rect 42812 711090 42840 714462
rect 42628 711062 42840 711090
rect 42352 709974 42564 710002
rect 41786 709880 41842 709889
rect 41786 709815 41842 709824
rect 41800 709376 41828 709815
rect 42246 709200 42302 709209
rect 42246 709135 42302 709144
rect 42062 708520 42118 708529
rect 42062 708455 42118 708464
rect 42076 708152 42104 708455
rect 42062 707840 42118 707849
rect 42062 707775 42118 707784
rect 42076 707540 42104 707775
rect 42260 707418 42288 709135
rect 42168 707390 42288 707418
rect 42168 706860 42196 707390
rect 42062 706752 42118 706761
rect 42062 706687 42118 706696
rect 42076 706316 42104 706687
rect 42246 705528 42302 705537
rect 42246 705463 42302 705472
rect 41786 704304 41842 704313
rect 41786 704239 41842 704248
rect 41800 703868 41828 704239
rect 42260 703746 42288 705463
rect 42536 705194 42564 709974
rect 42076 703718 42288 703746
rect 42444 705166 42564 705194
rect 42628 705194 42656 711062
rect 42890 710832 42946 710841
rect 42890 710767 42946 710776
rect 42904 708529 42932 710767
rect 42890 708520 42946 708529
rect 42890 708455 42946 708464
rect 42628 705166 42748 705194
rect 42076 703188 42104 703718
rect 42444 702590 42472 705166
rect 42168 702522 42196 702576
rect 42260 702562 42472 702590
rect 42260 702522 42288 702562
rect 42168 702494 42288 702522
rect 42430 702400 42486 702409
rect 42430 702335 42486 702344
rect 42246 702128 42302 702137
rect 42246 702063 42302 702072
rect 42076 701865 42104 702032
rect 42062 701856 42118 701865
rect 42062 701791 42118 701800
rect 42260 700179 42288 702063
rect 42182 700151 42288 700179
rect 42444 699530 42472 702335
rect 42720 701865 42748 705166
rect 42706 701856 42762 701865
rect 42706 701791 42762 701800
rect 42614 701584 42670 701593
rect 42614 701519 42670 701528
rect 42182 699502 42472 699530
rect 42628 698918 42656 701519
rect 42168 698850 42196 698904
rect 42260 698890 42656 698918
rect 42260 698850 42288 698890
rect 42168 698822 42288 698850
rect 35622 691384 35678 691393
rect 35622 691319 35678 691328
rect 8588 688772 8616 688908
rect 9048 688772 9076 688908
rect 9508 688772 9536 688908
rect 9968 688772 9996 688908
rect 10428 688772 10456 688908
rect 10888 688772 10916 688908
rect 11348 688772 11376 688908
rect 11808 688772 11836 688908
rect 12268 688772 12296 688908
rect 12728 688772 12756 688908
rect 13188 688772 13216 688908
rect 13648 688772 13676 688908
rect 14108 688772 14136 688908
rect 35636 687313 35664 691319
rect 41418 689344 41474 689353
rect 41418 689279 41474 689288
rect 35806 687712 35862 687721
rect 35806 687647 35862 687656
rect 35622 687304 35678 687313
rect 35820 687274 35848 687647
rect 41432 687274 41460 689279
rect 35622 687239 35678 687248
rect 35808 687268 35860 687274
rect 35808 687210 35860 687216
rect 41420 687268 41472 687274
rect 41420 687210 41472 687216
rect 35806 683224 35862 683233
rect 35806 683159 35808 683168
rect 35860 683159 35862 683168
rect 41696 683188 41748 683194
rect 35808 683130 35860 683136
rect 41696 683130 41748 683136
rect 35438 682816 35494 682825
rect 35438 682751 35494 682760
rect 35452 681766 35480 682751
rect 35622 682408 35678 682417
rect 35622 682343 35678 682352
rect 35636 681902 35664 682343
rect 35808 682032 35860 682038
rect 35806 682000 35808 682009
rect 36544 682032 36596 682038
rect 35860 682000 35862 682009
rect 36544 681974 36596 681980
rect 41708 681986 41736 683130
rect 35806 681935 35862 681944
rect 35624 681896 35676 681902
rect 35624 681838 35676 681844
rect 35440 681760 35492 681766
rect 35440 681702 35492 681708
rect 32402 681592 32458 681601
rect 32402 681527 32458 681536
rect 31022 681184 31078 681193
rect 31022 681119 31078 681128
rect 31036 672761 31064 681119
rect 32416 672790 32444 681527
rect 35162 680776 35218 680785
rect 35162 680711 35218 680720
rect 32404 672784 32456 672790
rect 31022 672752 31078 672761
rect 32404 672726 32456 672732
rect 31022 672687 31078 672696
rect 35176 671362 35204 680711
rect 36556 671702 36584 681974
rect 41708 681958 42104 681986
rect 41696 681896 41748 681902
rect 41694 681864 41696 681873
rect 41748 681864 41750 681873
rect 41694 681799 41750 681808
rect 41604 681692 41656 681698
rect 41604 681634 41656 681640
rect 41616 678586 41644 681634
rect 41786 678600 41842 678609
rect 41616 678558 41786 678586
rect 41786 678535 41842 678544
rect 41326 677104 41382 677113
rect 41326 677039 41382 677048
rect 41340 672489 41368 677039
rect 42076 676214 42104 681958
rect 42522 681864 42578 681873
rect 42522 681799 42578 681808
rect 42536 678974 42564 681799
rect 42798 679960 42854 679969
rect 42798 679895 42854 679904
rect 42444 678946 42564 678974
rect 42444 676214 42472 678946
rect 42076 676186 42196 676214
rect 42444 676186 42564 676214
rect 41604 672784 41656 672790
rect 41656 672732 41828 672738
rect 41604 672726 41828 672732
rect 41616 672710 41828 672726
rect 41326 672480 41382 672489
rect 41326 672415 41382 672424
rect 36544 671696 36596 671702
rect 36544 671638 36596 671644
rect 39672 671696 39724 671702
rect 39672 671638 39724 671644
rect 35164 671356 35216 671362
rect 35164 671298 35216 671304
rect 39684 670993 39712 671638
rect 41328 671356 41380 671362
rect 41328 671298 41380 671304
rect 41340 671129 41368 671298
rect 41326 671120 41382 671129
rect 41326 671055 41382 671064
rect 39670 670984 39726 670993
rect 39670 670919 39726 670928
rect 41800 670721 41828 672710
rect 42168 672217 42196 676186
rect 42536 674834 42564 676186
rect 42352 674806 42564 674834
rect 42154 672208 42210 672217
rect 42154 672143 42210 672152
rect 42352 671242 42380 674806
rect 42260 671214 42380 671242
rect 41786 670712 41842 670721
rect 41786 670647 41842 670656
rect 41786 670304 41842 670313
rect 41786 670239 41842 670248
rect 41800 669868 41828 670239
rect 42260 670018 42288 671214
rect 42614 671120 42670 671129
rect 42614 671055 42670 671064
rect 42260 669990 42564 670018
rect 41786 669080 41842 669089
rect 41786 669015 41842 669024
rect 41800 668644 41828 669015
rect 42246 668944 42302 668953
rect 42246 668879 42302 668888
rect 42168 667978 42196 668032
rect 42260 667978 42288 668879
rect 42168 667950 42288 667978
rect 42246 667856 42302 667865
rect 42302 667814 42472 667842
rect 42246 667791 42302 667800
rect 41970 667720 42026 667729
rect 41970 667655 42026 667664
rect 41984 667352 42012 667655
rect 42246 667584 42302 667593
rect 42246 667519 42302 667528
rect 42260 667298 42288 667519
rect 42260 667270 42380 667298
rect 42062 667040 42118 667049
rect 42118 666998 42288 667026
rect 42062 666975 42118 666984
rect 42062 666632 42118 666641
rect 42062 666567 42118 666576
rect 42076 666165 42104 666567
rect 42062 665680 42118 665689
rect 42260 665666 42288 666998
rect 42118 665638 42288 665666
rect 42062 665615 42118 665624
rect 41786 665408 41842 665417
rect 41786 665343 41842 665352
rect 41800 664972 41828 665343
rect 42352 665258 42380 667270
rect 42168 665230 42380 665258
rect 42168 665145 42196 665230
rect 42154 665136 42210 665145
rect 42154 665071 42210 665080
rect 42154 664864 42210 664873
rect 42154 664799 42210 664808
rect 42168 664325 42196 664799
rect 41970 664048 42026 664057
rect 41970 663983 42026 663992
rect 41984 663680 42012 663983
rect 42444 663150 42472 667814
rect 42182 663122 42472 663150
rect 42536 662969 42564 669990
rect 42628 665174 42656 671055
rect 42812 667298 42840 679895
rect 43088 678974 43116 719743
rect 43088 678946 43300 678974
rect 43074 676696 43130 676705
rect 43074 676631 43130 676640
rect 43088 676546 43116 676631
rect 43088 676518 43208 676546
rect 43180 669314 43208 676518
rect 43088 669286 43208 669314
rect 42812 667270 42932 667298
rect 42904 666641 42932 667270
rect 42890 666632 42946 666641
rect 42890 666567 42946 666576
rect 42628 665146 42748 665174
rect 42522 662960 42578 662969
rect 42522 662895 42578 662904
rect 42720 662833 42748 665146
rect 43088 664442 43116 669286
rect 42904 664414 43116 664442
rect 42706 662824 42762 662833
rect 42706 662759 42762 662768
rect 42338 662552 42394 662561
rect 42338 662487 42394 662496
rect 42154 661056 42210 661065
rect 42154 660991 42210 661000
rect 42168 660620 42196 660991
rect 42154 660512 42210 660521
rect 42154 660447 42210 660456
rect 42168 660008 42196 660447
rect 42352 659654 42380 662487
rect 42706 659832 42762 659841
rect 42706 659767 42762 659776
rect 42260 659626 42380 659654
rect 42260 659371 42288 659626
rect 42182 659343 42288 659371
rect 42154 659016 42210 659025
rect 42154 658951 42210 658960
rect 42168 658784 42196 658951
rect 42338 658608 42394 658617
rect 42338 658543 42394 658552
rect 42154 657384 42210 657393
rect 42154 657319 42210 657328
rect 42168 656948 42196 657319
rect 42352 656350 42380 658543
rect 42522 658336 42578 658345
rect 42522 658271 42578 658280
rect 42182 656322 42380 656350
rect 42168 655710 42288 655738
rect 42168 655656 42196 655710
rect 42260 655670 42288 655710
rect 42536 655670 42564 658271
rect 42720 657393 42748 659767
rect 42706 657384 42762 657393
rect 42706 657319 42762 657328
rect 42260 655642 42564 655670
rect 35806 646776 35862 646785
rect 35806 646711 35862 646720
rect 8588 645524 8616 645660
rect 9048 645524 9076 645660
rect 9508 645524 9536 645660
rect 9968 645524 9996 645660
rect 10428 645524 10456 645660
rect 10888 645524 10916 645660
rect 11348 645524 11376 645660
rect 11808 645524 11836 645660
rect 12268 645524 12296 645660
rect 12728 645524 12756 645660
rect 13188 645524 13216 645660
rect 13648 645524 13676 645660
rect 14108 645524 14136 645660
rect 35820 644745 35848 646711
rect 35806 644736 35862 644745
rect 35806 644671 35862 644680
rect 41786 641676 41842 641685
rect 41786 641611 41842 641620
rect 41800 641209 41828 641611
rect 41786 641200 41842 641209
rect 41786 641135 41842 641144
rect 35622 639840 35678 639849
rect 35622 639775 35678 639784
rect 35636 638994 35664 639775
rect 35806 639432 35862 639441
rect 35806 639367 35862 639376
rect 35820 639130 35848 639367
rect 35808 639124 35860 639130
rect 35808 639066 35860 639072
rect 36544 639124 36596 639130
rect 36544 639066 36596 639072
rect 35624 638988 35676 638994
rect 35624 638930 35676 638936
rect 35806 638616 35862 638625
rect 35806 638551 35862 638560
rect 32402 638208 32458 638217
rect 32402 638143 32458 638152
rect 32416 629950 32444 638143
rect 35820 636886 35848 638551
rect 35808 636880 35860 636886
rect 35808 636822 35860 636828
rect 36556 630737 36584 639066
rect 41512 638988 41564 638994
rect 41512 638930 41564 638936
rect 41524 634814 41552 638930
rect 41696 636880 41748 636886
rect 41696 636822 41748 636828
rect 41708 636018 41736 636822
rect 41708 635990 42656 636018
rect 42628 634814 42656 635990
rect 41524 634786 42564 634814
rect 42628 634786 42748 634814
rect 42338 633856 42394 633865
rect 42338 633791 42394 633800
rect 36542 630728 36598 630737
rect 36542 630663 36598 630672
rect 32404 629944 32456 629950
rect 32404 629886 32456 629892
rect 41696 629944 41748 629950
rect 41748 629892 42288 629898
rect 41696 629886 42288 629892
rect 41708 629870 42288 629886
rect 42260 627178 42288 629870
rect 42168 627150 42288 627178
rect 42168 626620 42196 627150
rect 42352 625478 42380 633791
rect 42536 633706 42564 634786
rect 42444 633678 42564 633706
rect 42444 630674 42472 633678
rect 42444 630646 42564 630674
rect 42182 625450 42380 625478
rect 42536 624866 42564 630646
rect 42168 624838 42288 624866
rect 42168 624784 42196 624838
rect 42260 624798 42288 624838
rect 42444 624838 42564 624866
rect 42444 624798 42472 624838
rect 42260 624770 42472 624798
rect 42154 624472 42210 624481
rect 42154 624407 42210 624416
rect 42430 624472 42486 624481
rect 42430 624407 42486 624416
rect 42168 624172 42196 624407
rect 42246 623792 42302 623801
rect 42246 623727 42302 623736
rect 42062 623384 42118 623393
rect 42062 623319 42118 623328
rect 42076 622948 42104 623319
rect 42168 621738 42196 621792
rect 42260 621738 42288 623727
rect 42444 623642 42472 624407
rect 42168 621710 42288 621738
rect 42352 623614 42472 623642
rect 42352 621126 42380 623614
rect 42182 621098 42380 621126
rect 42720 621014 42748 634786
rect 42536 620986 42748 621014
rect 42062 620936 42118 620945
rect 42062 620871 42118 620880
rect 42076 620500 42104 620871
rect 42536 619970 42564 620986
rect 42706 620392 42762 620401
rect 42706 620327 42762 620336
rect 42168 619834 42196 619956
rect 42260 619942 42564 619970
rect 42260 619834 42288 619942
rect 42168 619806 42288 619834
rect 42246 619712 42302 619721
rect 42246 619647 42302 619656
rect 42260 618474 42288 619647
rect 42522 618624 42578 618633
rect 42522 618559 42578 618568
rect 42260 618446 42472 618474
rect 42062 618352 42118 618361
rect 42118 618310 42288 618338
rect 42062 618287 42118 618296
rect 42260 617681 42288 618310
rect 42246 617672 42302 617681
rect 42246 617607 42302 617616
rect 42444 617454 42472 618446
rect 42168 617386 42196 617440
rect 42352 617426 42472 617454
rect 42352 617386 42380 617426
rect 42168 617358 42380 617386
rect 42062 617128 42118 617137
rect 42062 617063 42118 617072
rect 42076 616828 42104 617063
rect 42536 616593 42564 618559
rect 42062 616584 42118 616593
rect 42062 616519 42118 616528
rect 42522 616584 42578 616593
rect 42522 616519 42578 616528
rect 42076 616148 42104 616519
rect 42154 615904 42210 615913
rect 42154 615839 42210 615848
rect 42168 615604 42196 615839
rect 42720 615618 42748 620327
rect 42904 616185 42932 664414
rect 43272 659654 43300 678946
rect 43088 659626 43300 659654
rect 42890 616176 42946 616185
rect 42890 616111 42946 616120
rect 42720 615590 42840 615618
rect 42614 615496 42670 615505
rect 42614 615431 42670 615440
rect 42246 615224 42302 615233
rect 42246 615159 42302 615168
rect 41786 614136 41842 614145
rect 41786 614071 41842 614080
rect 41800 613768 41828 614071
rect 42260 613135 42288 615159
rect 42182 613107 42288 613135
rect 42628 612490 42656 615431
rect 42812 615346 42840 615590
rect 42182 612462 42656 612490
rect 42720 615318 42840 615346
rect 42720 611354 42748 615318
rect 43088 611969 43116 659626
rect 43364 621014 43392 932039
rect 43548 814881 43576 940199
rect 43732 936193 43760 958695
rect 43718 936184 43774 936193
rect 43718 936119 43774 936128
rect 44192 933745 44220 963863
rect 44376 935377 44404 964679
rect 44560 937009 44588 968759
rect 44836 941497 44864 990082
rect 45560 946008 45612 946014
rect 45560 945950 45612 945956
rect 45572 943537 45600 945950
rect 45558 943528 45614 943537
rect 45558 943463 45614 943472
rect 44822 941488 44878 941497
rect 44822 941423 44878 941432
rect 44546 937000 44602 937009
rect 44546 936935 44602 936944
rect 44362 935368 44418 935377
rect 44362 935303 44418 935312
rect 44178 933736 44234 933745
rect 44178 933671 44234 933680
rect 46938 933328 46994 933337
rect 46938 933263 46994 933272
rect 44086 892800 44142 892809
rect 44086 892735 44088 892744
rect 44140 892735 44142 892744
rect 44088 892706 44140 892712
rect 44086 892256 44142 892265
rect 44086 892191 44142 892200
rect 44100 891886 44128 892191
rect 44088 891880 44140 891886
rect 44088 891822 44140 891828
rect 46204 870868 46256 870874
rect 46204 870810 46256 870816
rect 44178 816096 44234 816105
rect 44178 816031 44234 816040
rect 43534 814872 43590 814881
rect 43534 814807 43590 814816
rect 43534 807664 43590 807673
rect 43534 807599 43590 807608
rect 43272 620986 43392 621014
rect 43272 612950 43300 620986
rect 43260 612944 43312 612950
rect 43260 612886 43312 612892
rect 43548 612354 43576 807599
rect 43718 806304 43774 806313
rect 43718 806239 43774 806248
rect 43732 612542 43760 806239
rect 44192 773265 44220 816031
rect 45006 815280 45062 815289
rect 45006 815215 45062 815224
rect 44362 814464 44418 814473
rect 44362 814399 44418 814408
rect 44178 773256 44234 773265
rect 44178 773191 44234 773200
rect 44376 772154 44404 814399
rect 44638 813648 44694 813657
rect 44638 813583 44694 813592
rect 44284 772126 44404 772154
rect 44284 771633 44312 772126
rect 44454 772032 44510 772041
rect 44454 771967 44510 771976
rect 44270 771624 44326 771633
rect 44270 771559 44326 771568
rect 44270 770400 44326 770409
rect 44270 770335 44326 770344
rect 43902 763056 43958 763065
rect 43902 762991 43958 763000
rect 43720 612536 43772 612542
rect 43720 612478 43772 612484
rect 43548 612338 43622 612354
rect 43548 612332 43634 612338
rect 43548 612326 43582 612332
rect 43582 612274 43634 612280
rect 43916 612134 43944 762991
rect 44284 727705 44312 770335
rect 44468 729337 44496 771967
rect 44652 770817 44680 813583
rect 44822 809976 44878 809985
rect 44822 809911 44878 809920
rect 44836 792305 44864 809911
rect 44822 792296 44878 792305
rect 44822 792231 44878 792240
rect 44822 772848 44878 772857
rect 44822 772783 44878 772792
rect 44638 770808 44694 770817
rect 44638 770743 44694 770752
rect 44638 766320 44694 766329
rect 44638 766255 44694 766264
rect 44652 754905 44680 766255
rect 44638 754896 44694 754905
rect 44638 754831 44694 754840
rect 44836 730153 44864 772783
rect 45020 772449 45048 815215
rect 45190 810792 45246 810801
rect 45190 810727 45246 810736
rect 45204 788225 45232 810727
rect 45374 799096 45430 799105
rect 45374 799031 45430 799040
rect 45388 797337 45416 799031
rect 45374 797328 45430 797337
rect 45374 797263 45430 797272
rect 45190 788216 45246 788225
rect 45190 788151 45246 788160
rect 45006 772440 45062 772449
rect 45006 772375 45062 772384
rect 45006 771216 45062 771225
rect 45006 771151 45062 771160
rect 44822 730144 44878 730153
rect 44822 730079 44878 730088
rect 44638 729736 44694 729745
rect 44638 729671 44694 729680
rect 44454 729328 44510 729337
rect 44454 729263 44510 729272
rect 44270 727696 44326 727705
rect 44270 727631 44326 727640
rect 44454 723616 44510 723625
rect 44454 723551 44510 723560
rect 44178 722800 44234 722809
rect 44178 722735 44234 722744
rect 44192 707849 44220 722735
rect 44178 707840 44234 707849
rect 44178 707775 44234 707784
rect 44468 705537 44496 723551
rect 44454 705528 44510 705537
rect 44454 705463 44510 705472
rect 44652 686905 44680 729671
rect 45020 728521 45048 771151
rect 45558 764280 45614 764289
rect 45558 764215 45614 764224
rect 45190 728920 45246 728929
rect 45190 728855 45246 728864
rect 45006 728512 45062 728521
rect 45006 728447 45062 728456
rect 44914 721168 44970 721177
rect 44914 721103 44970 721112
rect 44638 686896 44694 686905
rect 44638 686831 44694 686840
rect 44362 686488 44418 686497
rect 44362 686423 44418 686432
rect 44178 679552 44234 679561
rect 44178 679487 44234 679496
rect 44192 667593 44220 679487
rect 44178 667584 44234 667593
rect 44178 667519 44234 667528
rect 44376 643657 44404 686423
rect 44546 679144 44602 679153
rect 44546 679079 44602 679088
rect 44560 661065 44588 679079
rect 44730 677920 44786 677929
rect 44730 677855 44786 677864
rect 44546 661056 44602 661065
rect 44546 660991 44602 661000
rect 44744 654134 44772 677855
rect 44744 654106 44864 654134
rect 44362 643648 44418 643657
rect 44362 643583 44418 643592
rect 44178 636576 44234 636585
rect 44008 636534 44178 636562
rect 44008 634814 44036 636534
rect 44178 636511 44234 636520
rect 44362 636304 44418 636313
rect 44362 636239 44418 636248
rect 44178 635352 44234 635361
rect 44178 635287 44234 635296
rect 44192 634814 44220 635287
rect 44008 634786 44128 634814
rect 44192 634786 44312 634814
rect 44100 625297 44128 634786
rect 44086 625288 44142 625297
rect 44086 625223 44142 625232
rect 44284 624594 44312 634786
rect 44192 624566 44312 624594
rect 44192 620945 44220 624566
rect 44376 624481 44404 636239
rect 44836 636154 44864 654106
rect 44652 636126 44864 636154
rect 44652 635882 44680 636126
rect 44652 635854 44772 635882
rect 44546 635760 44602 635769
rect 44546 635695 44602 635704
rect 44362 624472 44418 624481
rect 44362 624407 44418 624416
rect 44178 620936 44234 620945
rect 44178 620871 44234 620880
rect 44560 619721 44588 635695
rect 44546 619712 44602 619721
rect 44546 619647 44602 619656
rect 44086 616176 44142 616185
rect 44086 616111 44142 616120
rect 44100 615482 44128 616111
rect 44100 615454 44220 615482
rect 43904 612128 43956 612134
rect 43904 612070 43956 612076
rect 43074 611960 43130 611969
rect 43074 611895 43130 611904
rect 43929 611960 43985 611969
rect 43929 611895 43985 611904
rect 43943 611726 43971 611895
rect 43931 611720 43983 611726
rect 44192 611674 44220 615454
rect 43931 611662 43983 611668
rect 44167 611646 44220 611674
rect 44167 611386 44195 611646
rect 42536 611326 42748 611354
rect 44155 611380 44207 611386
rect 42536 611017 42564 611326
rect 44155 611322 44207 611328
rect 44744 611114 44772 635854
rect 44928 611522 44956 721103
rect 45204 686089 45232 728855
rect 45374 721576 45430 721585
rect 45374 721511 45430 721520
rect 45388 710841 45416 721511
rect 45374 710832 45430 710841
rect 45374 710767 45430 710776
rect 45190 686080 45246 686089
rect 45190 686015 45246 686024
rect 45282 685672 45338 685681
rect 45282 685607 45338 685616
rect 45098 643376 45154 643385
rect 45098 643311 45154 643320
rect 44916 611516 44968 611522
rect 44916 611458 44968 611464
rect 44732 611108 44784 611114
rect 44732 611050 44784 611056
rect 42522 611008 42578 611017
rect 42522 610943 42578 610952
rect 44500 611008 44556 611017
rect 44500 610943 44556 610952
rect 44514 610774 44542 610943
rect 44502 610768 44554 610774
rect 44502 610710 44554 610716
rect 8588 602276 8616 602412
rect 9048 602276 9076 602412
rect 9508 602276 9536 602412
rect 9968 602276 9996 602412
rect 10428 602276 10456 602412
rect 10888 602276 10916 602412
rect 11348 602276 11376 602412
rect 11808 602276 11836 602412
rect 12268 602276 12296 602412
rect 12728 602276 12756 602412
rect 13188 602276 13216 602412
rect 13648 602276 13676 602412
rect 14108 602276 14136 602412
rect 45112 600545 45140 643311
rect 45296 643113 45324 685607
rect 45282 643104 45338 643113
rect 45282 643039 45338 643048
rect 45374 642560 45430 642569
rect 45374 642495 45430 642504
rect 45388 634814 45416 642495
rect 45388 634786 45508 634814
rect 45480 621014 45508 634786
rect 45296 620986 45508 621014
rect 45296 611354 45324 620986
rect 45572 611930 45600 764215
rect 46216 754089 46244 870810
rect 46202 754080 46258 754089
rect 46202 754015 46258 754024
rect 45742 728104 45798 728113
rect 45742 728039 45798 728048
rect 45756 685273 45784 728039
rect 46110 727424 46166 727433
rect 46110 727359 46166 727368
rect 45742 685264 45798 685273
rect 45742 685199 45798 685208
rect 45926 684856 45982 684865
rect 45926 684791 45982 684800
rect 45742 684040 45798 684049
rect 45742 683975 45798 683984
rect 45756 641481 45784 683975
rect 45940 642297 45968 684791
rect 46124 684457 46152 727359
rect 46110 684448 46166 684457
rect 46110 684383 46166 684392
rect 46110 680368 46166 680377
rect 46110 680303 46166 680312
rect 46124 660521 46152 680303
rect 46110 660512 46166 660521
rect 46110 660447 46166 660456
rect 45926 642288 45982 642297
rect 45926 642223 45982 642232
rect 45742 641472 45798 641481
rect 45742 641407 45798 641416
rect 45926 641200 45982 641209
rect 45926 641135 45982 641144
rect 45742 633448 45798 633457
rect 45742 633383 45798 633392
rect 45560 611924 45612 611930
rect 45560 611866 45612 611872
rect 45296 611326 45416 611354
rect 45098 600536 45154 600545
rect 45098 600471 45154 600480
rect 44638 600128 44694 600137
rect 44638 600063 44694 600072
rect 42982 597000 43038 597009
rect 42982 596935 43038 596944
rect 42154 596864 42210 596873
rect 42154 596799 42210 596808
rect 41234 596048 41290 596057
rect 41234 595983 41290 595992
rect 33046 595640 33102 595649
rect 33046 595575 33102 595584
rect 31022 594416 31078 594425
rect 31022 594351 31078 594360
rect 31036 585818 31064 594351
rect 33060 587178 33088 595575
rect 35162 595232 35218 595241
rect 35162 595167 35218 595176
rect 33048 587172 33100 587178
rect 33048 587114 33100 587120
rect 35176 585954 35204 595167
rect 40682 594824 40738 594833
rect 40682 594759 40738 594768
rect 40498 593192 40554 593201
rect 40498 593127 40554 593136
rect 40316 592340 40368 592346
rect 40316 592282 40368 592288
rect 39946 590744 40002 590753
rect 39946 590679 40002 590688
rect 39960 586158 39988 590679
rect 40328 589393 40356 592282
rect 40512 589665 40540 593127
rect 40498 589656 40554 589665
rect 40498 589591 40554 589600
rect 40314 589384 40370 589393
rect 40314 589319 40370 589328
rect 40408 587172 40460 587178
rect 40408 587114 40460 587120
rect 40420 586537 40448 587114
rect 40406 586528 40462 586537
rect 40406 586463 40462 586472
rect 39948 586152 40000 586158
rect 39948 586094 40000 586100
rect 35164 585948 35216 585954
rect 35164 585890 35216 585896
rect 31024 585812 31076 585818
rect 31024 585754 31076 585760
rect 40696 584633 40724 594759
rect 41248 594538 41276 595983
rect 41694 594552 41750 594561
rect 41248 594510 41694 594538
rect 41694 594487 41750 594496
rect 41786 593600 41842 593609
rect 41616 593558 41786 593586
rect 41616 592890 41644 593558
rect 41786 593535 41842 593544
rect 40868 592884 40920 592890
rect 40868 592826 40920 592832
rect 41604 592884 41656 592890
rect 41604 592826 41656 592832
rect 40682 584624 40738 584633
rect 40880 584594 40908 592826
rect 41786 592784 41842 592793
rect 41432 592742 41786 592770
rect 41432 592346 41460 592742
rect 41786 592719 41842 592728
rect 41786 592376 41842 592385
rect 41420 592340 41472 592346
rect 41786 592311 41842 592320
rect 41420 592282 41472 592288
rect 41800 589529 41828 592311
rect 41786 589520 41842 589529
rect 41786 589455 41842 589464
rect 42168 589274 42196 596799
rect 42614 594552 42670 594561
rect 42614 594487 42670 594496
rect 42628 592034 42656 594487
rect 42798 594008 42854 594017
rect 42798 593943 42854 593952
rect 42536 592006 42656 592034
rect 42536 589274 42564 592006
rect 42076 589246 42196 589274
rect 42260 589246 42564 589274
rect 42076 586809 42104 589246
rect 42062 586800 42118 586809
rect 42062 586735 42118 586744
rect 42260 586650 42288 589246
rect 42260 586622 42380 586650
rect 41696 586152 41748 586158
rect 42352 586140 42380 586622
rect 42522 586528 42578 586537
rect 42578 586486 42748 586514
rect 42522 586463 42578 586472
rect 42352 586112 42656 586140
rect 41748 586100 41920 586106
rect 41696 586094 41920 586100
rect 41708 586078 41920 586094
rect 41892 585970 41920 586078
rect 41696 585948 41748 585954
rect 41892 585942 42380 585970
rect 41696 585890 41748 585896
rect 41708 585834 41736 585890
rect 41708 585806 42288 585834
rect 41696 585744 41748 585750
rect 41696 585686 41748 585692
rect 41708 584905 41736 585686
rect 41694 584896 41750 584905
rect 41694 584831 41750 584840
rect 40682 584559 40738 584568
rect 40868 584588 40920 584594
rect 40868 584530 40920 584536
rect 41604 584588 41656 584594
rect 41604 584530 41656 584536
rect 41616 584474 41644 584530
rect 41616 584446 41828 584474
rect 41800 584361 41828 584446
rect 41786 584352 41842 584361
rect 41786 584287 41842 584296
rect 42260 583930 42288 585806
rect 42168 583902 42288 583930
rect 42168 583440 42196 583902
rect 42352 583386 42380 585942
rect 42260 583358 42380 583386
rect 42260 582374 42288 583358
rect 42168 582346 42288 582374
rect 42168 582249 42196 582346
rect 42338 581768 42394 581777
rect 42338 581703 42394 581712
rect 41984 581505 42012 581604
rect 41970 581496 42026 581505
rect 41970 581431 42026 581440
rect 42352 580975 42380 581703
rect 42182 580947 42380 580975
rect 42246 580816 42302 580825
rect 42246 580751 42302 580760
rect 42430 580816 42486 580825
rect 42430 580751 42486 580760
rect 41970 580272 42026 580281
rect 41970 580207 42026 580216
rect 41984 579768 42012 580207
rect 42260 578626 42288 580751
rect 42444 579578 42472 580751
rect 42628 579578 42656 586112
rect 42168 578598 42288 578626
rect 42352 579550 42472 579578
rect 42536 579550 42656 579578
rect 42168 578544 42196 578598
rect 41786 578232 41842 578241
rect 42352 578234 42380 579550
rect 42536 578234 42564 579550
rect 41786 578167 41842 578176
rect 42260 578206 42380 578234
rect 42444 578206 42564 578234
rect 41800 577932 41828 578167
rect 41786 577552 41842 577561
rect 41786 577487 41842 577496
rect 41800 577281 41828 577487
rect 42260 577266 42288 578206
rect 42260 577238 42380 577266
rect 42154 577144 42210 577153
rect 42154 577079 42210 577088
rect 42168 576708 42196 577079
rect 41970 576600 42026 576609
rect 42026 576558 42196 576586
rect 41970 576535 42026 576544
rect 42168 576450 42196 576558
rect 42168 576422 42288 576450
rect 42260 574274 42288 576422
rect 42182 574246 42288 574274
rect 42154 574152 42210 574161
rect 42154 574087 42210 574096
rect 42168 573580 42196 574087
rect 42352 572982 42380 577238
rect 42182 572954 42380 572982
rect 42444 572438 42472 578206
rect 42720 577561 42748 586486
rect 42812 578234 42840 593943
rect 42996 579614 43024 596935
rect 44454 591968 44510 591977
rect 44454 591903 44510 591912
rect 43442 591560 43498 591569
rect 43442 591495 43498 591504
rect 43166 584896 43222 584905
rect 43166 584831 43222 584840
rect 43180 580825 43208 584831
rect 43166 580816 43222 580825
rect 43166 580751 43222 580760
rect 42996 579586 43116 579614
rect 42812 578206 42932 578234
rect 42904 577969 42932 578206
rect 42890 577960 42946 577969
rect 42890 577895 42946 577904
rect 42706 577552 42762 577561
rect 42706 577487 42762 577496
rect 43088 577266 43116 579586
rect 42904 577238 43116 577266
rect 42904 574818 42932 577238
rect 42904 574790 43024 574818
rect 42614 573336 42670 573345
rect 42614 573271 42670 573280
rect 42168 572370 42196 572424
rect 42260 572410 42472 572438
rect 42260 572370 42288 572410
rect 42168 572342 42288 572370
rect 42628 572234 42656 573271
rect 42352 572206 42656 572234
rect 42352 571010 42380 572206
rect 42522 572112 42578 572121
rect 42522 572047 42578 572056
rect 42076 570982 42380 571010
rect 42076 570588 42104 570982
rect 41786 570208 41842 570217
rect 41786 570143 41842 570152
rect 41800 569908 41828 570143
rect 42536 569514 42564 572047
rect 42076 569486 42564 569514
rect 42076 569296 42104 569486
rect 42338 569256 42394 569265
rect 42338 569191 42394 569200
rect 42352 567194 42380 569191
rect 41524 567166 42380 567194
rect 8588 559164 8616 559300
rect 9048 559164 9076 559300
rect 9508 559164 9536 559300
rect 9968 559164 9996 559300
rect 10428 559164 10456 559300
rect 10888 559164 10916 559300
rect 11348 559164 11376 559300
rect 11808 559164 11836 559300
rect 12268 559164 12296 559300
rect 12728 559164 12756 559300
rect 13188 559164 13216 559300
rect 13648 559164 13676 559300
rect 14108 559164 14136 559300
rect 35806 558104 35862 558113
rect 35806 558039 35862 558048
rect 35820 557598 35848 558039
rect 41524 557598 41552 567166
rect 42062 558512 42118 558521
rect 42062 558447 42118 558456
rect 35808 557592 35860 557598
rect 35808 557534 35860 557540
rect 41512 557592 41564 557598
rect 42076 557569 42104 558447
rect 41512 557534 41564 557540
rect 42062 557560 42118 557569
rect 42996 557534 43024 574790
rect 42062 557495 42118 557504
rect 42812 557506 43024 557534
rect 35806 554840 35862 554849
rect 42812 554826 42840 557506
rect 41708 554810 42840 554826
rect 35806 554775 35808 554784
rect 35860 554775 35862 554784
rect 41696 554804 42840 554810
rect 35808 554746 35860 554752
rect 41748 554798 42840 554804
rect 41696 554746 41748 554752
rect 35806 553616 35862 553625
rect 35806 553551 35862 553560
rect 35820 553450 35848 553551
rect 35808 553444 35860 553450
rect 41328 553444 41380 553450
rect 35808 553386 35860 553392
rect 41156 553392 41328 553394
rect 41156 553386 41380 553392
rect 41156 553366 41368 553386
rect 33782 551984 33838 551993
rect 33782 551919 33838 551928
rect 31758 548142 31814 548151
rect 31758 548077 31814 548086
rect 31772 547874 31800 548077
rect 31760 547868 31812 547874
rect 31760 547810 31812 547816
rect 33796 543046 33824 551919
rect 41156 550610 41184 553366
rect 41326 552800 41382 552809
rect 41326 552735 41382 552744
rect 41340 552090 41368 552735
rect 41328 552084 41380 552090
rect 41328 552026 41380 552032
rect 41696 552084 41748 552090
rect 41696 552026 41748 552032
rect 41708 551857 41736 552026
rect 41694 551848 41750 551857
rect 41694 551783 41750 551792
rect 43074 551576 43130 551585
rect 43074 551511 43130 551520
rect 41786 550760 41842 550769
rect 41786 550695 41842 550704
rect 41800 550634 41828 550695
rect 41156 550582 41460 550610
rect 40498 549944 40554 549953
rect 40498 549879 40554 549888
rect 38476 547868 38528 547874
rect 38476 547810 38528 547816
rect 33784 543040 33836 543046
rect 33784 542982 33836 542988
rect 38488 542366 38516 547810
rect 40512 545465 40540 549879
rect 41234 548142 41290 548151
rect 41234 548077 41290 548086
rect 41432 547874 41460 550582
rect 41708 550606 41828 550634
rect 41708 550474 41736 550606
rect 41708 550446 41828 550474
rect 41800 548457 41828 550446
rect 41970 550352 42026 550361
rect 41970 550287 42026 550296
rect 41786 548448 41842 548457
rect 41786 548383 41842 548392
rect 41694 548176 41750 548185
rect 41694 548111 41696 548120
rect 41748 548111 41750 548120
rect 41696 548082 41748 548088
rect 41432 547846 41736 547874
rect 40498 545456 40554 545465
rect 40498 545391 40554 545400
rect 41708 543734 41736 547846
rect 41984 545737 42012 550287
rect 42890 548448 42946 548457
rect 42890 548383 42946 548392
rect 41970 545728 42026 545737
rect 41970 545663 42026 545672
rect 41708 543706 42472 543734
rect 41512 543040 41564 543046
rect 41512 542982 41564 542988
rect 38476 542360 38528 542366
rect 38476 542302 38528 542308
rect 41524 542178 41552 542982
rect 41696 542360 41748 542366
rect 41748 542308 42288 542314
rect 41696 542302 42288 542308
rect 41708 542286 42288 542302
rect 41524 542150 41828 542178
rect 41800 541113 41828 542150
rect 41786 541104 41842 541113
rect 41786 541039 41842 541048
rect 42260 540818 42288 542286
rect 42260 540790 42380 540818
rect 41786 540696 41842 540705
rect 41786 540631 41842 540640
rect 41800 540260 41828 540631
rect 42352 539050 42380 540790
rect 42182 539022 42380 539050
rect 42444 538506 42472 543706
rect 42614 540288 42670 540297
rect 42614 540223 42670 540232
rect 42352 538478 42472 538506
rect 42352 538438 42380 538478
rect 42168 538370 42196 538424
rect 42260 538410 42380 538438
rect 42260 538370 42288 538410
rect 42168 538342 42288 538370
rect 42246 538248 42302 538257
rect 42246 538183 42302 538192
rect 42260 538098 42288 538183
rect 42260 538070 42380 538098
rect 42062 537976 42118 537985
rect 42062 537911 42118 537920
rect 42076 537744 42104 537911
rect 42352 537758 42380 538070
rect 42628 537985 42656 540223
rect 42614 537976 42670 537985
rect 42614 537911 42670 537920
rect 42260 537730 42380 537758
rect 42168 536466 42196 536588
rect 42260 536466 42288 537730
rect 42614 537432 42670 537441
rect 42614 537367 42670 537376
rect 42168 536438 42288 536466
rect 42246 536344 42302 536353
rect 42246 536279 42302 536288
rect 42260 535378 42288 536279
rect 42182 535350 42288 535378
rect 41786 535256 41842 535265
rect 41786 535191 41842 535200
rect 41800 534752 41828 535191
rect 42628 534426 42656 537367
rect 42352 534398 42656 534426
rect 42352 534086 42380 534398
rect 42522 534304 42578 534313
rect 42522 534239 42578 534248
rect 42182 534058 42380 534086
rect 42536 534074 42564 534239
rect 42904 534074 42932 548383
rect 43088 534074 43116 551511
rect 42444 534046 42564 534074
rect 42812 534046 42932 534074
rect 42996 534046 43116 534074
rect 42444 533542 42472 534046
rect 42182 533514 42472 533542
rect 42430 533352 42486 533361
rect 42430 533287 42486 533296
rect 42444 531059 42472 533287
rect 42812 532794 42840 534046
rect 42182 531031 42472 531059
rect 42536 532766 42840 532794
rect 42536 530414 42564 532766
rect 42706 532672 42762 532681
rect 42706 532607 42762 532616
rect 42182 530386 42564 530414
rect 42430 530224 42486 530233
rect 42430 530159 42486 530168
rect 42062 529952 42118 529961
rect 42062 529887 42118 529896
rect 42076 529757 42104 529887
rect 41878 529408 41934 529417
rect 41878 529343 41934 529352
rect 41892 529205 41920 529343
rect 42168 527462 42288 527490
rect 42168 527340 42196 527462
rect 42260 527354 42288 527462
rect 42444 527354 42472 530159
rect 42720 529961 42748 532607
rect 42706 529952 42762 529961
rect 42706 529887 42762 529896
rect 42996 529802 43024 534046
rect 42260 527326 42472 527354
rect 42536 529774 43024 529802
rect 42536 526742 42564 529774
rect 42706 529680 42762 529689
rect 42706 529615 42762 529624
rect 42182 526714 42564 526742
rect 42720 526091 42748 529615
rect 42182 526063 42748 526091
rect 8588 431596 8616 431664
rect 9048 431596 9076 431664
rect 9508 431596 9536 431664
rect 9968 431596 9996 431664
rect 10428 431596 10456 431664
rect 10888 431596 10916 431664
rect 11348 431596 11376 431664
rect 11808 431596 11836 431664
rect 12268 431596 12296 431664
rect 12728 431596 12756 431664
rect 13188 431596 13216 431664
rect 13648 431596 13676 431664
rect 14108 431596 14136 431664
rect 41326 426048 41382 426057
rect 41326 425983 41382 425992
rect 40958 425640 41014 425649
rect 40958 425575 41014 425584
rect 33782 424416 33838 424425
rect 33782 424351 33838 424360
rect 33796 416090 33824 424351
rect 40972 422226 41000 425575
rect 41340 424266 41368 425983
rect 41340 424238 41552 424266
rect 41524 424130 41552 424238
rect 41524 424102 42012 424130
rect 41786 422784 41842 422793
rect 41786 422719 41842 422728
rect 40972 422198 41184 422226
rect 41156 418849 41184 422198
rect 41142 418840 41198 418849
rect 41142 418775 41198 418784
rect 41800 418577 41828 422719
rect 41786 418568 41842 418577
rect 41786 418503 41842 418512
rect 41984 418154 42012 424102
rect 42798 424008 42854 424017
rect 42798 423943 42854 423952
rect 42522 419928 42578 419937
rect 42522 419863 42578 419872
rect 41984 418126 42472 418154
rect 33784 416084 33836 416090
rect 33784 416026 33836 416032
rect 41696 416084 41748 416090
rect 41696 416026 41748 416032
rect 41708 415970 41736 416026
rect 41708 415942 42288 415970
rect 42260 413114 42288 415942
rect 42444 415394 42472 418126
rect 42168 413086 42288 413114
rect 42352 415366 42472 415394
rect 42536 415394 42564 419863
rect 42536 415366 42656 415394
rect 42168 412624 42196 413086
rect 42062 411904 42118 411913
rect 42062 411839 42118 411848
rect 42076 411468 42104 411839
rect 42352 411074 42380 415366
rect 42628 411913 42656 415366
rect 42614 411904 42670 411913
rect 42614 411839 42670 411848
rect 42168 411046 42380 411074
rect 42168 410788 42196 411046
rect 42182 410162 42472 410190
rect 41786 409456 41842 409465
rect 41786 409391 41842 409400
rect 41800 408952 41828 409391
rect 42444 408513 42472 410162
rect 42430 408504 42486 408513
rect 42430 408439 42486 408448
rect 42430 407824 42486 407833
rect 42168 407674 42196 407796
rect 42260 407782 42430 407810
rect 42260 407674 42288 407782
rect 42430 407759 42486 407768
rect 42168 407646 42288 407674
rect 42182 407102 42472 407130
rect 42062 406736 42118 406745
rect 42062 406671 42118 406680
rect 42076 406504 42104 406671
rect 41786 406328 41842 406337
rect 41786 406263 41842 406272
rect 41800 405929 41828 406263
rect 42444 405657 42472 407102
rect 42430 405648 42486 405657
rect 42430 405583 42486 405592
rect 41786 403880 41842 403889
rect 41786 403815 41842 403824
rect 41800 403444 41828 403815
rect 42338 402928 42394 402937
rect 42168 402886 42338 402914
rect 42168 402801 42196 402886
rect 42338 402863 42394 402872
rect 42430 402520 42486 402529
rect 42430 402455 42486 402464
rect 42444 402166 42472 402455
rect 42182 402138 42472 402166
rect 41786 401976 41842 401985
rect 41786 401911 41842 401920
rect 41800 401608 41828 401911
rect 42430 399800 42486 399809
rect 42182 399758 42430 399786
rect 42430 399735 42486 399744
rect 42812 399135 42840 423943
rect 43258 420744 43314 420753
rect 43258 420679 43314 420688
rect 43074 419248 43130 419257
rect 43074 419183 43130 419192
rect 42182 399107 42840 399135
rect 41786 398848 41842 398857
rect 41786 398783 41842 398792
rect 41800 398480 41828 398783
rect 8588 388348 8616 388484
rect 9048 388348 9076 388484
rect 9508 388348 9536 388484
rect 9968 388348 9996 388484
rect 10428 388348 10456 388484
rect 10888 388348 10916 388484
rect 11348 388348 11376 388484
rect 11808 388348 11836 388484
rect 12268 388348 12296 388484
rect 12728 388348 12756 388484
rect 13188 388348 13216 388484
rect 13648 388348 13676 388484
rect 14108 388348 14136 388484
rect 42062 387696 42118 387705
rect 42062 387631 42118 387640
rect 41878 387288 41934 387297
rect 41878 387223 41934 387232
rect 41142 387152 41198 387161
rect 41142 387087 41198 387096
rect 41156 386322 41184 387087
rect 41892 386481 41920 387223
rect 42076 386753 42104 387631
rect 42062 386744 42118 386753
rect 42062 386679 42118 386688
rect 41878 386472 41934 386481
rect 41878 386407 41934 386416
rect 42062 386472 42118 386481
rect 42062 386407 42118 386416
rect 42076 386322 42104 386407
rect 41156 386294 42104 386322
rect 35438 383072 35494 383081
rect 35438 383007 35494 383016
rect 35452 382294 35480 383007
rect 35622 382664 35678 382673
rect 35622 382599 35678 382608
rect 35636 382430 35664 382599
rect 35808 382560 35860 382566
rect 35808 382502 35860 382508
rect 40040 382560 40092 382566
rect 40040 382502 40092 382508
rect 35624 382424 35676 382430
rect 35624 382366 35676 382372
rect 35440 382288 35492 382294
rect 35820 382265 35848 382502
rect 35440 382230 35492 382236
rect 35806 382256 35862 382265
rect 35806 382191 35862 382200
rect 35530 381440 35586 381449
rect 35530 381375 35586 381384
rect 35806 381440 35862 381449
rect 35806 381375 35862 381384
rect 35544 381070 35572 381375
rect 35532 381064 35584 381070
rect 35532 381006 35584 381012
rect 35820 380934 35848 381375
rect 37924 381064 37976 381070
rect 37924 381006 37976 381012
rect 35808 380928 35860 380934
rect 35808 380870 35860 380876
rect 35806 376544 35862 376553
rect 35806 376479 35862 376488
rect 35820 376038 35848 376479
rect 35808 376032 35860 376038
rect 35808 375974 35860 375980
rect 37936 371385 37964 381006
rect 40052 376961 40080 382502
rect 41696 382424 41748 382430
rect 41696 382366 41748 382372
rect 41512 382288 41564 382294
rect 41510 382256 41512 382265
rect 41564 382256 41566 382265
rect 41510 382191 41566 382200
rect 41328 380928 41380 380934
rect 41328 380870 41380 380876
rect 41340 378593 41368 380870
rect 41708 379514 41736 382366
rect 42798 382256 42854 382265
rect 42798 382191 42854 382200
rect 41708 379486 42564 379514
rect 41326 378584 41382 378593
rect 41326 378519 41382 378528
rect 42338 378584 42394 378593
rect 42338 378519 42394 378528
rect 40038 376952 40094 376961
rect 40038 376887 40094 376896
rect 42352 376754 42380 378519
rect 42352 376726 42472 376754
rect 39580 376032 39632 376038
rect 39580 375974 39632 375980
rect 39592 375737 39620 375974
rect 39578 375728 39634 375737
rect 39578 375663 39634 375672
rect 37922 371376 37978 371385
rect 37922 371311 37978 371320
rect 42444 369458 42472 376726
rect 42182 369430 42472 369458
rect 41786 368656 41842 368665
rect 41786 368591 41842 368600
rect 41800 368249 41828 368591
rect 42536 367622 42564 379486
rect 42182 367594 42564 367622
rect 42430 367024 42486 367033
rect 42182 366968 42430 366975
rect 42182 366959 42486 366968
rect 42182 366947 42472 366959
rect 42430 365800 42486 365809
rect 42182 365758 42430 365786
rect 42430 365735 42486 365744
rect 41800 364313 41828 364548
rect 41786 364304 41842 364313
rect 41786 364239 41842 364248
rect 42430 364304 42486 364313
rect 42430 364239 42486 364248
rect 42444 363950 42472 364239
rect 42182 363922 42472 363950
rect 41786 363760 41842 363769
rect 41786 363695 41842 363704
rect 41800 363256 41828 363695
rect 41786 362944 41842 362953
rect 41786 362879 41842 362888
rect 41800 362712 41828 362879
rect 41800 360097 41828 360264
rect 41786 360088 41842 360097
rect 41786 360023 41842 360032
rect 42154 359952 42210 359961
rect 42154 359887 42210 359896
rect 42168 359584 42196 359887
rect 42182 358958 42472 358986
rect 41786 358728 41842 358737
rect 41786 358663 41842 358672
rect 41800 358428 41828 358663
rect 42444 357377 42472 358958
rect 42430 357368 42486 357377
rect 42430 357303 42486 357312
rect 42812 356674 42840 382191
rect 42536 356646 42840 356674
rect 42536 356606 42564 356646
rect 42168 356538 42196 356592
rect 42260 356578 42564 356606
rect 42260 356538 42288 356578
rect 42168 356510 42288 356538
rect 42338 356008 42394 356017
rect 42168 355966 42338 355994
rect 42168 355912 42196 355966
rect 42338 355943 42394 355952
rect 41878 355736 41934 355745
rect 41878 355671 41934 355680
rect 41892 355300 41920 355671
rect 43088 355609 43116 419183
rect 43074 355600 43130 355609
rect 43074 355535 43130 355544
rect 43272 353705 43300 420679
rect 43456 379514 43484 591495
rect 43626 590336 43682 590345
rect 43626 590271 43682 590280
rect 43456 379486 43576 379514
rect 43548 354226 43576 379486
rect 43640 354362 43668 590271
rect 44468 581097 44496 591903
rect 44454 581088 44510 581097
rect 44454 581023 44510 581032
rect 44652 557297 44680 600063
rect 45388 599729 45416 611326
rect 45756 610910 45784 633383
rect 45744 610904 45796 610910
rect 45744 610846 45796 610852
rect 45374 599720 45430 599729
rect 45374 599655 45430 599664
rect 44822 599312 44878 599321
rect 44822 599247 44878 599256
rect 44638 557288 44694 557297
rect 44638 557223 44694 557232
rect 44836 556481 44864 599247
rect 45940 598913 45968 641135
rect 46110 640928 46166 640937
rect 46110 640863 46166 640872
rect 45926 598904 45982 598913
rect 45926 598839 45982 598848
rect 45006 598496 45062 598505
rect 45006 598431 45062 598440
rect 44822 556472 44878 556481
rect 44822 556407 44878 556416
rect 45020 555665 45048 598431
rect 46124 598097 46152 640863
rect 46952 612746 46980 933263
rect 47596 891993 47624 991714
rect 48964 991636 49016 991642
rect 48964 991578 49016 991584
rect 48976 942313 49004 991578
rect 48962 942304 49018 942313
rect 48962 942239 49018 942248
rect 50356 940681 50384 993006
rect 50342 940672 50398 940681
rect 50342 940607 50398 940616
rect 51736 939865 51764 993142
rect 55864 992928 55916 992934
rect 55864 992870 55916 992876
rect 54484 991500 54536 991506
rect 54484 991442 54536 991448
rect 53288 988780 53340 988786
rect 53288 988722 53340 988728
rect 51722 939856 51778 939865
rect 51722 939791 51778 939800
rect 53104 923296 53156 923302
rect 53104 923238 53156 923244
rect 50344 909492 50396 909498
rect 50344 909434 50396 909440
rect 47768 897048 47820 897054
rect 47768 896990 47820 896996
rect 47582 891984 47638 891993
rect 47582 891919 47638 891928
rect 47584 818372 47636 818378
rect 47584 818314 47636 818320
rect 47596 711113 47624 818314
rect 47780 817737 47808 896990
rect 47766 817728 47822 817737
rect 47766 817663 47822 817672
rect 50356 816921 50384 909434
rect 51724 858424 51776 858430
rect 51724 858366 51776 858372
rect 50342 816912 50398 816921
rect 50342 816847 50398 816856
rect 50344 805996 50396 806002
rect 50344 805938 50396 805944
rect 48964 767372 49016 767378
rect 48964 767314 49016 767320
rect 47582 711104 47638 711113
rect 47582 711039 47638 711048
rect 48976 669361 49004 767314
rect 50356 730561 50384 805938
rect 51736 773537 51764 858366
rect 53116 799105 53144 923238
rect 53300 892265 53328 988722
rect 54496 892537 54524 991442
rect 55876 892809 55904 992870
rect 73436 990276 73488 990282
rect 73436 990218 73488 990224
rect 73448 983620 73476 990218
rect 95896 988786 95924 1002050
rect 96068 1001972 96120 1001978
rect 96068 1001914 96120 1001920
rect 96080 991778 96108 1001914
rect 97276 994537 97304 1002322
rect 97460 994809 97488 1002594
rect 99470 1002552 99526 1002561
rect 99470 1002487 99472 1002496
rect 99524 1002487 99526 1002496
rect 100024 1002516 100076 1002522
rect 99472 1002458 99524 1002464
rect 100024 1002458 100076 1002464
rect 98828 1002244 98880 1002250
rect 98828 1002186 98880 1002192
rect 98274 1002008 98330 1002017
rect 98274 1001943 98276 1001952
rect 98328 1001943 98330 1001952
rect 98644 1001972 98696 1001978
rect 98276 1001914 98328 1001920
rect 98644 1001914 98696 1001920
rect 98000 1000544 98052 1000550
rect 98000 1000486 98052 1000492
rect 98012 998442 98040 1000486
rect 98000 998436 98052 998442
rect 98000 998378 98052 998384
rect 98656 995897 98684 1001914
rect 98840 999190 98868 1002186
rect 99102 1002144 99158 1002153
rect 99102 1002079 99104 1002088
rect 99156 1002079 99158 1002088
rect 99104 1002050 99156 1002056
rect 98828 999184 98880 999190
rect 98828 999126 98880 999132
rect 100036 997626 100064 1002458
rect 100298 1002416 100354 1002425
rect 100298 1002351 100300 1002360
rect 100352 1002351 100354 1002360
rect 100300 1002322 100352 1002328
rect 101126 1002280 101182 1002289
rect 101126 1002215 101128 1002224
rect 101180 1002215 101182 1002224
rect 101128 1002186 101180 1002192
rect 101126 1002008 101182 1002017
rect 100208 1001972 100260 1001978
rect 100208 1001914 100260 1001920
rect 100772 1001966 101126 1001994
rect 100220 1000550 100248 1001914
rect 100208 1000544 100260 1000550
rect 100208 1000486 100260 1000492
rect 100024 997620 100076 997626
rect 100024 997562 100076 997568
rect 100772 997014 100800 1001966
rect 101126 1001943 101182 1001952
rect 100760 997008 100812 997014
rect 100760 996950 100812 996956
rect 98642 995888 98698 995897
rect 98642 995823 98698 995832
rect 101416 995353 101444 1006130
rect 104806 1006088 104862 1006097
rect 102784 1006052 102836 1006058
rect 104806 1006023 104808 1006032
rect 102784 1005994 102836 1006000
rect 104860 1006023 104862 1006032
rect 108486 1006088 108542 1006097
rect 108486 1006023 108488 1006032
rect 104808 1005994 104860 1006000
rect 108540 1006023 108542 1006032
rect 108488 1005994 108540 1006000
rect 101954 1002144 102010 1002153
rect 101954 1002079 101956 1002088
rect 102008 1002079 102010 1002088
rect 101956 1002050 102008 1002056
rect 101402 995344 101458 995353
rect 101402 995279 101458 995288
rect 97446 994800 97502 994809
rect 97446 994735 97502 994744
rect 102796 994566 102824 1005994
rect 106830 1002688 106886 1002697
rect 106830 1002623 106832 1002632
rect 106884 1002623 106886 1002632
rect 109500 1002652 109552 1002658
rect 106832 1002594 106884 1002600
rect 109500 1002594 109552 1002600
rect 103150 1002552 103206 1002561
rect 103150 1002487 103152 1002496
rect 103204 1002487 103206 1002496
rect 108026 1002552 108082 1002561
rect 108026 1002487 108028 1002496
rect 103152 1002458 103204 1002464
rect 108080 1002487 108082 1002496
rect 108028 1002458 108080 1002464
rect 106002 1002416 106058 1002425
rect 106002 1002351 106004 1002360
rect 106056 1002351 106058 1002360
rect 108304 1002380 108356 1002386
rect 106004 1002322 106056 1002328
rect 108304 1002322 108356 1002328
rect 105634 1002280 105690 1002289
rect 105634 1002215 105636 1002224
rect 105688 1002215 105690 1002224
rect 107936 1002244 107988 1002250
rect 105636 1002186 105688 1002192
rect 107936 1002186 107988 1002192
rect 106830 1002144 106886 1002153
rect 106830 1002079 106832 1002088
rect 106884 1002079 106886 1002088
rect 106832 1002050 106884 1002056
rect 103150 1002008 103206 1002017
rect 103978 1002008 104034 1002017
rect 103150 1001943 103152 1001952
rect 103204 1001943 103206 1001952
rect 103532 1001966 103978 1001994
rect 103152 1001914 103204 1001920
rect 103532 994838 103560 1001966
rect 103978 1001943 104034 1001952
rect 106002 1002008 106058 1002017
rect 106002 1001943 106004 1001952
rect 106056 1001943 106058 1001952
rect 107752 1001972 107804 1001978
rect 106004 1001914 106056 1001920
rect 107752 1001914 107804 1001920
rect 106924 997076 106976 997082
rect 106924 997018 106976 997024
rect 103520 994832 103572 994838
rect 103520 994774 103572 994780
rect 104900 994696 104952 994702
rect 104900 994638 104952 994644
rect 102784 994560 102836 994566
rect 97262 994528 97318 994537
rect 102784 994502 102836 994508
rect 97262 994463 97318 994472
rect 96068 991772 96120 991778
rect 96068 991714 96120 991720
rect 95884 988780 95936 988786
rect 95884 988722 95936 988728
rect 104912 986678 104940 994638
rect 104900 986672 104952 986678
rect 104900 986614 104952 986620
rect 105820 986672 105872 986678
rect 105820 986614 105872 986620
rect 89628 985992 89680 985998
rect 89628 985934 89680 985940
rect 89640 983620 89668 985934
rect 105832 983620 105860 986614
rect 106936 985998 106964 997018
rect 107764 993070 107792 1001914
rect 107948 993206 107976 1002186
rect 108316 997762 108344 1002322
rect 108854 1002280 108910 1002289
rect 108854 1002215 108856 1002224
rect 108908 1002215 108910 1002224
rect 108856 1002186 108908 1002192
rect 109040 1002108 109092 1002114
rect 109040 1002050 109092 1002056
rect 108854 1002008 108910 1002017
rect 108854 1001943 108856 1001952
rect 108908 1001943 108910 1001952
rect 108856 1001914 108908 1001920
rect 108304 997756 108356 997762
rect 108304 997698 108356 997704
rect 107936 993200 107988 993206
rect 107936 993142 107988 993148
rect 107752 993064 107804 993070
rect 107752 993006 107804 993012
rect 109052 990146 109080 1002050
rect 109512 997626 109540 1002594
rect 110696 1002516 110748 1002522
rect 110696 1002458 110748 1002464
rect 109682 1002144 109738 1002153
rect 109682 1002079 109684 1002088
rect 109736 1002079 109738 1002088
rect 109684 1002050 109736 1002056
rect 110512 1001972 110564 1001978
rect 110512 1001914 110564 1001920
rect 109500 997620 109552 997626
rect 109500 997562 109552 997568
rect 110524 994702 110552 1001914
rect 110512 994696 110564 994702
rect 110512 994638 110564 994644
rect 110708 991642 110736 1002458
rect 112076 1002244 112128 1002250
rect 112076 1002186 112128 1002192
rect 111892 1002108 111944 1002114
rect 111892 1002050 111944 1002056
rect 111904 997082 111932 1002050
rect 111892 997076 111944 997082
rect 111892 997018 111944 997024
rect 110696 991636 110748 991642
rect 110696 991578 110748 991584
rect 112088 990282 112116 1002186
rect 116308 997756 116360 997762
rect 116308 997698 116360 997704
rect 116320 996985 116348 997698
rect 117228 997620 117280 997626
rect 117228 997562 117280 997568
rect 117240 997257 117268 997562
rect 117226 997248 117282 997257
rect 117226 997183 117282 997192
rect 116306 996976 116362 996985
rect 116306 996911 116362 996920
rect 124876 995081 124904 1006130
rect 126244 1006052 126296 1006058
rect 126244 1005994 126296 1006000
rect 126256 995353 126284 1005994
rect 144000 1002108 144052 1002114
rect 144000 1002050 144052 1002056
rect 143724 998436 143776 998442
rect 143724 998378 143776 998384
rect 143736 997914 143764 998378
rect 143644 997886 143764 997914
rect 136468 995858 136496 995860
rect 137756 995858 137784 995860
rect 136456 995852 136508 995858
rect 136456 995794 136508 995800
rect 137744 995852 137796 995858
rect 137744 995794 137796 995800
rect 143644 995761 143672 997886
rect 143816 997756 143868 997762
rect 143816 997698 143868 997704
rect 143828 997257 143856 997698
rect 143814 997248 143870 997257
rect 143814 997183 143870 997192
rect 143816 996736 143868 996742
rect 144012 996713 144040 1002050
rect 144196 1001894 144224 1006266
rect 144736 1006188 144788 1006194
rect 144736 1006130 144788 1006136
rect 144748 1001894 144776 1006130
rect 144196 1001866 144408 1001894
rect 144184 997892 144236 997898
rect 144184 997834 144236 997840
rect 143816 996678 143868 996684
rect 143998 996704 144054 996713
rect 143828 995994 143856 996678
rect 143998 996639 144054 996648
rect 143998 996160 144054 996169
rect 143998 996095 144000 996104
rect 144052 996095 144054 996104
rect 144000 996066 144052 996072
rect 143816 995988 143868 995994
rect 143816 995930 143868 995936
rect 140410 995752 140466 995761
rect 140162 995710 140410 995738
rect 141054 995752 141110 995761
rect 140806 995710 141054 995738
rect 140410 995687 140466 995696
rect 141054 995687 141110 995696
rect 143630 995752 143686 995761
rect 143630 995687 143686 995696
rect 136270 995616 136326 995625
rect 135930 995574 136270 995602
rect 144196 995586 144224 997834
rect 136270 995551 136326 995560
rect 143448 995580 143500 995586
rect 143448 995522 143500 995528
rect 144184 995580 144236 995586
rect 144184 995522 144236 995528
rect 141698 995480 141754 995489
rect 126242 995344 126298 995353
rect 126242 995279 126298 995288
rect 124862 995072 124918 995081
rect 124862 995007 124918 995016
rect 128464 994838 128492 995452
rect 128452 994832 128504 994838
rect 129108 994809 129136 995452
rect 128452 994774 128504 994780
rect 129094 994800 129150 994809
rect 129094 994735 129150 994744
rect 129752 994566 129780 995452
rect 131592 994702 131620 995452
rect 131580 994696 131632 994702
rect 131580 994638 131632 994644
rect 129740 994560 129792 994566
rect 129740 994502 129792 994508
rect 132144 994430 132172 995452
rect 132132 994424 132184 994430
rect 132132 994366 132184 994372
rect 121736 994288 121788 994294
rect 132788 994265 132816 995452
rect 133446 995438 133828 995466
rect 133800 995058 133828 995438
rect 133800 995030 133920 995058
rect 121736 994230 121788 994236
rect 132774 994256 132830 994265
rect 112076 990276 112128 990282
rect 112076 990218 112128 990224
rect 109040 990140 109092 990146
rect 109040 990082 109092 990088
rect 106924 985992 106976 985998
rect 106924 985934 106976 985940
rect 121748 983634 121776 994230
rect 132774 994191 132830 994200
rect 133892 993721 133920 995030
rect 137112 994537 137140 995452
rect 138966 995438 139348 995466
rect 141450 995438 141698 995466
rect 139320 995058 139348 995438
rect 142646 995438 143028 995466
rect 141698 995415 141754 995424
rect 141514 995344 141570 995353
rect 142066 995344 142122 995353
rect 141570 995302 142066 995330
rect 141514 995279 141570 995288
rect 143000 995330 143028 995438
rect 143460 995330 143488 995522
rect 143000 995302 143488 995330
rect 142066 995279 142122 995288
rect 139320 995030 139440 995058
rect 137098 994528 137154 994537
rect 137098 994463 137154 994472
rect 139412 993993 139440 995030
rect 142066 994528 142122 994537
rect 142066 994463 142122 994472
rect 139398 993984 139454 993993
rect 142080 993954 142108 994463
rect 142342 993984 142398 993993
rect 139398 993919 139454 993928
rect 142068 993948 142120 993954
rect 142342 993919 142344 993928
rect 142068 993890 142120 993896
rect 142396 993919 142398 993928
rect 142344 993890 142396 993896
rect 142068 993744 142120 993750
rect 133878 993712 133934 993721
rect 133878 993647 133934 993656
rect 142066 993712 142068 993721
rect 144380 993721 144408 1001866
rect 144656 1001866 144776 1001894
rect 144656 995858 144684 1001866
rect 144828 997620 144880 997626
rect 144828 997562 144880 997568
rect 144840 996985 144868 997562
rect 144826 996976 144882 996985
rect 144826 996911 144882 996920
rect 144644 995852 144696 995858
rect 144644 995794 144696 995800
rect 145576 993993 145604 1006402
rect 145760 994430 145788 1006538
rect 152094 1006496 152150 1006505
rect 152094 1006431 152096 1006440
rect 152148 1006431 152150 1006440
rect 157430 1006496 157486 1006505
rect 157430 1006431 157432 1006440
rect 152096 1006402 152148 1006408
rect 157484 1006431 157486 1006440
rect 166264 1006460 166316 1006466
rect 157432 1006402 157484 1006408
rect 166264 1006402 166316 1006408
rect 171784 1006460 171836 1006466
rect 171784 1006402 171836 1006408
rect 151726 1006360 151782 1006369
rect 151726 1006295 151728 1006304
rect 151780 1006295 151782 1006304
rect 158258 1006360 158314 1006369
rect 158258 1006295 158260 1006304
rect 151728 1006266 151780 1006272
rect 158312 1006295 158314 1006304
rect 158260 1006266 158312 1006272
rect 150898 1006224 150954 1006233
rect 150898 1006159 150900 1006168
rect 150952 1006159 150954 1006168
rect 160282 1006224 160338 1006233
rect 166276 1006194 166304 1006402
rect 160282 1006159 160284 1006168
rect 150900 1006130 150952 1006136
rect 160336 1006159 160338 1006168
rect 164884 1006188 164936 1006194
rect 160284 1006130 160336 1006136
rect 164884 1006130 164936 1006136
rect 166264 1006188 166316 1006194
rect 166264 1006130 166316 1006136
rect 150070 1006088 150126 1006097
rect 147588 1006052 147640 1006058
rect 150070 1006023 150072 1006032
rect 147588 1005994 147640 1006000
rect 150124 1006023 150126 1006032
rect 159454 1006088 159510 1006097
rect 159454 1006023 159456 1006032
rect 150072 1005994 150124 1006000
rect 159508 1006023 159510 1006032
rect 159456 1005994 159508 1006000
rect 147600 1002114 147628 1005994
rect 152922 1005408 152978 1005417
rect 149704 1005372 149756 1005378
rect 152922 1005343 152924 1005352
rect 149704 1005314 149756 1005320
rect 152976 1005343 152978 1005352
rect 152924 1005314 152976 1005320
rect 148508 1002244 148560 1002250
rect 148508 1002186 148560 1002192
rect 147588 1002108 147640 1002114
rect 147588 1002050 147640 1002056
rect 148324 1002108 148376 1002114
rect 148324 1002050 148376 1002056
rect 146944 1001972 146996 1001978
rect 146944 1001914 146996 1001920
rect 145748 994424 145800 994430
rect 145748 994366 145800 994372
rect 145562 993984 145618 993993
rect 145562 993919 145618 993928
rect 142120 993712 142122 993721
rect 142066 993647 142122 993656
rect 142250 993712 142306 993721
rect 142250 993647 142252 993656
rect 142304 993647 142306 993656
rect 144366 993712 144422 993721
rect 144366 993647 144422 993656
rect 142252 993618 142304 993624
rect 146956 992934 146984 1001914
rect 147678 996432 147734 996441
rect 147678 996367 147734 996376
rect 147692 992934 147720 996367
rect 146944 992928 146996 992934
rect 146944 992870 146996 992876
rect 147680 992928 147732 992934
rect 147680 992870 147732 992876
rect 138296 991636 138348 991642
rect 138296 991578 138348 991584
rect 121748 983606 122130 983634
rect 138308 983620 138336 991578
rect 148336 991506 148364 1002050
rect 148520 996742 148548 1002186
rect 149242 1002008 149298 1002017
rect 149242 1001943 149244 1001952
rect 149296 1001943 149298 1001952
rect 149244 1001914 149296 1001920
rect 148508 996736 148560 996742
rect 148508 996678 148560 996684
rect 149716 994537 149744 1005314
rect 152922 1005136 152978 1005145
rect 149888 1005100 149940 1005106
rect 152922 1005071 152924 1005080
rect 149888 1005042 149940 1005048
rect 152976 1005071 152978 1005080
rect 152924 1005042 152976 1005048
rect 149702 994528 149758 994537
rect 149702 994463 149758 994472
rect 149900 994265 149928 1005042
rect 153750 1005000 153806 1005009
rect 151084 1004964 151136 1004970
rect 153750 1004935 153752 1004944
rect 151084 1004906 151136 1004912
rect 153804 1004935 153806 1004944
rect 158626 1005000 158682 1005009
rect 158626 1004935 158628 1004944
rect 153752 1004906 153804 1004912
rect 158680 1004935 158682 1004944
rect 162124 1004964 162176 1004970
rect 158628 1004906 158680 1004912
rect 162124 1004906 162176 1004912
rect 150898 1002144 150954 1002153
rect 150898 1002079 150900 1002088
rect 150952 1002079 150954 1002088
rect 150900 1002050 150952 1002056
rect 151096 994809 151124 1004906
rect 160650 1004864 160706 1004873
rect 160650 1004799 160652 1004808
rect 160704 1004799 160706 1004808
rect 160652 1004770 160704 1004776
rect 154118 1004728 154174 1004737
rect 151268 1004692 151320 1004698
rect 154118 1004663 154120 1004672
rect 151268 1004634 151320 1004640
rect 154172 1004663 154174 1004672
rect 161110 1004728 161166 1004737
rect 161110 1004663 161112 1004672
rect 154120 1004634 154172 1004640
rect 161164 1004663 161166 1004672
rect 161112 1004634 161164 1004640
rect 151280 997898 151308 1004634
rect 155774 1002552 155830 1002561
rect 153844 1002516 153896 1002522
rect 155774 1002487 155776 1002496
rect 153844 1002458 153896 1002464
rect 155828 1002487 155830 1002496
rect 155776 1002458 155828 1002464
rect 151726 1002280 151782 1002289
rect 151726 1002215 151728 1002224
rect 151780 1002215 151782 1002224
rect 151728 1002186 151780 1002192
rect 152464 1001972 152516 1001978
rect 152464 1001914 152516 1001920
rect 151268 997892 151320 997898
rect 151268 997834 151320 997840
rect 152476 995858 152504 1001914
rect 153856 998442 153884 1002458
rect 156602 1002416 156658 1002425
rect 156602 1002351 156604 1002360
rect 156656 1002351 156658 1002360
rect 158720 1002380 158772 1002386
rect 156604 1002322 156656 1002328
rect 158720 1002322 158772 1002328
rect 155774 1002280 155830 1002289
rect 155774 1002215 155776 1002224
rect 155828 1002215 155830 1002224
rect 157340 1002244 157392 1002250
rect 155776 1002186 155828 1002192
rect 157340 1002186 157392 1002192
rect 156602 1002144 156658 1002153
rect 155224 1002108 155276 1002114
rect 156602 1002079 156604 1002088
rect 155224 1002050 155276 1002056
rect 156656 1002079 156658 1002088
rect 156604 1002050 156656 1002056
rect 154578 1002008 154634 1002017
rect 154578 1001943 154580 1001952
rect 154632 1001943 154634 1001952
rect 154946 1002008 155002 1002017
rect 154946 1001943 154948 1001952
rect 154580 1001914 154632 1001920
rect 155000 1001943 155002 1001952
rect 154948 1001914 155000 1001920
rect 155236 1001894 155264 1002050
rect 155960 1001972 156012 1001978
rect 155960 1001914 156012 1001920
rect 155236 1001866 155356 1001894
rect 153844 998436 153896 998442
rect 153844 998378 153896 998384
rect 152464 995852 152516 995858
rect 152464 995794 152516 995800
rect 155130 995616 155186 995625
rect 155130 995551 155186 995560
rect 155144 995081 155172 995551
rect 155130 995072 155186 995081
rect 155130 995007 155186 995016
rect 151082 994800 151138 994809
rect 151082 994735 151138 994744
rect 155328 994566 155356 1001866
rect 155972 994702 156000 1001914
rect 157352 994838 157380 1002186
rect 157798 1002008 157854 1002017
rect 157798 1001943 157800 1001952
rect 157852 1001943 157854 1001952
rect 157800 1001914 157852 1001920
rect 158732 997626 158760 1002322
rect 160100 1001972 160152 1001978
rect 160100 1001914 160152 1001920
rect 160112 997762 160140 1001914
rect 162136 997762 162164 1004906
rect 163136 1004828 163188 1004834
rect 163136 1004770 163188 1004776
rect 162952 1004692 163004 1004698
rect 162952 1004634 163004 1004640
rect 160100 997756 160152 997762
rect 160100 997698 160152 997704
rect 162124 997756 162176 997762
rect 162124 997698 162176 997704
rect 158720 997620 158772 997626
rect 158720 997562 158772 997568
rect 162964 997218 162992 1004634
rect 160744 997212 160796 997218
rect 160744 997154 160796 997160
rect 162952 997212 163004 997218
rect 162952 997154 163004 997160
rect 157340 994832 157392 994838
rect 157340 994774 157392 994780
rect 155960 994696 156012 994702
rect 155960 994638 156012 994644
rect 155316 994560 155368 994566
rect 155316 994502 155368 994508
rect 149886 994256 149942 994265
rect 149886 994191 149942 994200
rect 148324 991500 148376 991506
rect 148324 991442 148376 991448
rect 160756 985726 160784 997154
rect 163148 991642 163176 1004770
rect 163136 991636 163188 991642
rect 163136 991578 163188 991584
rect 164896 990894 164924 1006130
rect 170312 997756 170364 997762
rect 170312 997698 170364 997704
rect 170324 997257 170352 997698
rect 170310 997248 170366 997257
rect 170310 997183 170366 997192
rect 171796 996130 171824 1006402
rect 175924 1006188 175976 1006194
rect 175924 1006130 175976 1006136
rect 171784 996124 171836 996130
rect 171784 996066 171836 996072
rect 175936 995994 175964 1006130
rect 177304 1006052 177356 1006058
rect 177304 1005994 177356 1006000
rect 196808 1006052 196860 1006058
rect 196808 1005994 196860 1006000
rect 169392 995988 169444 995994
rect 169392 995930 169444 995936
rect 171508 995988 171560 995994
rect 171508 995930 171560 995936
rect 175924 995988 175976 995994
rect 175924 995930 175976 995936
rect 169404 994770 169432 995930
rect 170680 995852 170732 995858
rect 170680 995794 170732 995800
rect 169392 994764 169444 994770
rect 169392 994706 169444 994712
rect 170692 994158 170720 995794
rect 171048 995580 171100 995586
rect 171048 995522 171100 995528
rect 170864 994881 170916 994887
rect 170864 994823 170916 994829
rect 170680 994152 170732 994158
rect 170680 994094 170732 994100
rect 170876 993682 170904 994823
rect 171060 994634 171088 995522
rect 171520 995223 171548 995930
rect 177316 995858 177344 1005994
rect 196624 998844 196676 998850
rect 196624 998786 196676 998792
rect 195244 998436 195296 998442
rect 195244 998378 195296 998384
rect 195058 996432 195114 996441
rect 195058 996367 195114 996376
rect 171692 995852 171744 995858
rect 171692 995794 171744 995800
rect 177304 995852 177356 995858
rect 177304 995794 177356 995800
rect 171704 995335 171732 995794
rect 189446 995752 189502 995761
rect 189152 995710 189446 995738
rect 190458 995752 190514 995761
rect 190348 995710 190458 995738
rect 189446 995687 189502 995696
rect 190458 995687 190514 995696
rect 179860 995438 180196 995466
rect 172426 995344 172482 995353
rect 171692 995329 171744 995335
rect 172426 995279 172482 995288
rect 171692 995271 171744 995277
rect 171508 995217 171560 995223
rect 171508 995159 171560 995165
rect 172440 995110 172468 995279
rect 172428 995104 172480 995110
rect 172428 995046 172480 995052
rect 171232 994881 171284 994887
rect 171232 994823 171284 994829
rect 171048 994628 171100 994634
rect 171048 994570 171100 994576
rect 171244 993818 171272 994823
rect 180168 994498 180196 995438
rect 180490 995246 180518 995452
rect 181148 995438 181484 995466
rect 180708 995376 180760 995382
rect 180708 995318 180760 995324
rect 180478 995240 180530 995246
rect 180478 995182 180530 995188
rect 180720 994974 180748 995318
rect 181456 995110 181484 995438
rect 182652 995438 182988 995466
rect 183540 995438 183876 995466
rect 184184 995438 184520 995466
rect 184828 995438 184888 995466
rect 187312 995438 187648 995466
rect 187864 995438 188200 995466
rect 188508 995438 189028 995466
rect 191544 995438 191788 995466
rect 192188 995438 192524 995466
rect 192832 995438 193168 995466
rect 194028 995438 194364 995466
rect 182652 995382 182680 995438
rect 182640 995376 182692 995382
rect 182640 995318 182692 995324
rect 181444 995104 181496 995110
rect 181444 995046 181496 995052
rect 180708 994968 180760 994974
rect 180708 994910 180760 994916
rect 180156 994492 180208 994498
rect 180156 994434 180208 994440
rect 171232 993812 171284 993818
rect 171232 993754 171284 993760
rect 170864 993676 170916 993682
rect 170864 993618 170916 993624
rect 183848 993585 183876 995438
rect 184492 995081 184520 995438
rect 184664 995240 184716 995246
rect 184664 995182 184716 995188
rect 184478 995072 184534 995081
rect 184478 995007 184534 995016
rect 184676 994362 184704 995182
rect 184860 994809 184888 995438
rect 187620 995353 187648 995438
rect 187606 995344 187662 995353
rect 187606 995279 187662 995288
rect 184846 994800 184902 994809
rect 184846 994735 184902 994744
rect 188172 994537 188200 995438
rect 189000 995058 189028 995438
rect 190368 995240 190420 995246
rect 190368 995182 190420 995188
rect 190552 995240 190604 995246
rect 190552 995182 190604 995188
rect 190380 995081 190408 995182
rect 190564 995081 190592 995182
rect 190366 995072 190422 995081
rect 189000 995030 189120 995058
rect 188158 994528 188214 994537
rect 188158 994463 188214 994472
rect 184664 994356 184716 994362
rect 184664 994298 184716 994304
rect 189092 994265 189120 995030
rect 190366 995007 190422 995016
rect 190550 995072 190606 995081
rect 191760 995058 191788 995438
rect 192496 995246 192524 995438
rect 193140 995382 193168 995438
rect 193128 995376 193180 995382
rect 193128 995318 193180 995324
rect 194336 995246 194364 995438
rect 195072 995382 195100 996367
rect 195060 995376 195112 995382
rect 195060 995318 195112 995324
rect 195256 995246 195284 998378
rect 195796 998028 195848 998034
rect 195796 997970 195848 997976
rect 195428 997892 195480 997898
rect 195428 997834 195480 997840
rect 195440 996713 195468 997834
rect 195612 997756 195664 997762
rect 195612 997698 195664 997704
rect 195426 996704 195482 996713
rect 195426 996639 195482 996648
rect 195624 996418 195652 997698
rect 195440 996390 195652 996418
rect 192484 995240 192536 995246
rect 192484 995182 192536 995188
rect 194140 995240 194192 995246
rect 194140 995182 194192 995188
rect 194324 995240 194376 995246
rect 194324 995182 194376 995188
rect 195244 995240 195296 995246
rect 195244 995182 195296 995188
rect 194152 995058 194180 995182
rect 195440 995058 195468 996390
rect 195612 996260 195664 996266
rect 195612 996202 195664 996208
rect 191760 995030 191880 995058
rect 194152 995030 195468 995058
rect 190550 995007 190606 995016
rect 189078 994256 189134 994265
rect 189078 994191 189134 994200
rect 183834 993576 183890 993585
rect 183834 993511 183890 993520
rect 186504 992928 186556 992934
rect 191852 992905 191880 995030
rect 195624 993682 195652 996202
rect 195808 993818 195836 997970
rect 196636 994265 196664 998786
rect 196820 996441 196848 1005994
rect 198004 998708 198056 998714
rect 198004 998650 198056 998656
rect 196806 996432 196862 996441
rect 196806 996367 196862 996376
rect 198016 994537 198044 998650
rect 199384 998164 199436 998170
rect 199384 998106 199436 998112
rect 199396 996402 199424 998106
rect 200040 997898 200068 1007354
rect 505374 1007176 505430 1007185
rect 505374 1007111 505376 1007120
rect 505428 1007111 505430 1007120
rect 513840 1007140 513892 1007146
rect 505376 1007082 505428 1007088
rect 513840 1007082 513892 1007088
rect 428004 1006936 428056 1006942
rect 357714 1006904 357770 1006913
rect 428002 1006904 428004 1006913
rect 505376 1006936 505428 1006942
rect 428056 1006904 428058 1006913
rect 357714 1006839 357716 1006848
rect 357768 1006839 357770 1006848
rect 369860 1006868 369912 1006874
rect 357716 1006810 357768 1006816
rect 428002 1006839 428058 1006848
rect 505374 1006904 505376 1006913
rect 505428 1006904 505430 1006913
rect 505374 1006839 505430 1006848
rect 369860 1006810 369912 1006816
rect 360198 1006768 360254 1006777
rect 360198 1006703 360200 1006712
rect 360252 1006703 360254 1006712
rect 360200 1006674 360252 1006680
rect 210054 1006496 210110 1006505
rect 206192 1006460 206244 1006466
rect 306930 1006496 306986 1006505
rect 210054 1006431 210056 1006440
rect 206192 1006402 206244 1006408
rect 210108 1006431 210110 1006440
rect 300308 1006460 300360 1006466
rect 210056 1006402 210108 1006408
rect 306930 1006431 306932 1006440
rect 300308 1006402 300360 1006408
rect 306984 1006431 306986 1006440
rect 306932 1006402 306984 1006408
rect 201038 1006088 201094 1006097
rect 201038 1006023 201040 1006032
rect 201092 1006023 201094 1006032
rect 201040 1005994 201092 1006000
rect 203524 1002108 203576 1002114
rect 203524 1002050 203576 1002056
rect 202694 998744 202750 998753
rect 202694 998679 202696 998688
rect 202748 998679 202750 998688
rect 202696 998650 202748 998656
rect 201040 998572 201092 998578
rect 201040 998514 201092 998520
rect 200670 998064 200726 998073
rect 200670 997999 200672 998008
rect 200724 997999 200726 998008
rect 200672 997970 200724 997976
rect 200028 997892 200080 997898
rect 200028 997834 200080 997840
rect 201052 997754 201080 998514
rect 201866 998200 201922 998209
rect 201866 998135 201868 998144
rect 201920 998135 201922 998144
rect 201868 998106 201920 998112
rect 202328 998028 202380 998034
rect 202328 997970 202380 997976
rect 202144 997892 202196 997898
rect 202144 997834 202196 997840
rect 200960 997726 201080 997754
rect 200212 997280 200264 997286
rect 200210 997248 200212 997257
rect 200264 997248 200266 997257
rect 200210 997183 200266 997192
rect 200764 996736 200816 996742
rect 200764 996678 200816 996684
rect 199384 996396 199436 996402
rect 199384 996338 199436 996344
rect 200776 994809 200804 996678
rect 200960 995761 200988 997726
rect 200946 995752 201002 995761
rect 200946 995687 201002 995696
rect 200762 994800 200818 994809
rect 200762 994735 200818 994744
rect 198002 994528 198058 994537
rect 198002 994463 198058 994472
rect 196622 994256 196678 994265
rect 196622 994191 196678 994200
rect 195796 993812 195848 993818
rect 195796 993754 195848 993760
rect 195612 993676 195664 993682
rect 195612 993618 195664 993624
rect 202156 993585 202184 997834
rect 202340 994362 202368 997970
rect 202512 996736 202564 996742
rect 202512 996678 202564 996684
rect 202524 995897 202552 996678
rect 202510 995888 202566 995897
rect 202510 995823 202566 995832
rect 203536 995353 203564 1002050
rect 205546 1002008 205602 1002017
rect 204168 1001972 204220 1001978
rect 205546 1001943 205548 1001952
rect 204168 1001914 204220 1001920
rect 205600 1001943 205602 1001952
rect 205548 1001914 205600 1001920
rect 203890 998880 203946 998889
rect 203890 998815 203892 998824
rect 203944 998815 203946 998824
rect 203892 998786 203944 998792
rect 203890 998608 203946 998617
rect 203890 998543 203892 998552
rect 203944 998543 203946 998552
rect 203892 998514 203944 998520
rect 204180 998442 204208 1001914
rect 204168 998436 204220 998442
rect 204168 998378 204220 998384
rect 205546 998064 205602 998073
rect 205546 997999 205548 998008
rect 205600 997999 205602 998008
rect 205548 997970 205600 997976
rect 204718 997928 204774 997937
rect 204718 997863 204720 997872
rect 204772 997863 204774 997872
rect 204720 997834 204772 997840
rect 206204 997286 206232 1006402
rect 210422 1006360 210478 1006369
rect 256146 1006360 256202 1006369
rect 210422 1006295 210424 1006304
rect 210476 1006295 210478 1006304
rect 228364 1006324 228416 1006330
rect 210424 1006266 210476 1006272
rect 228364 1006266 228416 1006272
rect 249248 1006324 249300 1006330
rect 256146 1006295 256148 1006304
rect 249248 1006266 249300 1006272
rect 256200 1006295 256202 1006304
rect 298928 1006324 298980 1006330
rect 256148 1006266 256200 1006272
rect 298928 1006266 298980 1006272
rect 208398 1006224 208454 1006233
rect 208398 1006159 208400 1006168
rect 208452 1006159 208454 1006168
rect 208400 1006130 208452 1006136
rect 209226 1006088 209282 1006097
rect 209226 1006023 209228 1006032
rect 209280 1006023 209282 1006032
rect 211804 1006052 211856 1006058
rect 209228 1005994 209280 1006000
rect 211804 1005994 211856 1006000
rect 208400 1005168 208452 1005174
rect 208398 1005136 208400 1005145
rect 209872 1005168 209924 1005174
rect 208452 1005136 208454 1005145
rect 209872 1005110 209924 1005116
rect 208398 1005071 208454 1005080
rect 207572 1005032 207624 1005038
rect 207570 1005000 207572 1005009
rect 207624 1005000 207626 1005009
rect 207570 1004935 207626 1004944
rect 209226 1004864 209282 1004873
rect 209226 1004799 209228 1004808
rect 209280 1004799 209282 1004808
rect 209228 1004770 209280 1004776
rect 207202 1002552 207258 1002561
rect 207258 1002510 207428 1002538
rect 207202 1002487 207258 1002496
rect 207202 1002280 207258 1002289
rect 207032 1002238 207202 1002266
rect 206374 1002144 206430 1002153
rect 206374 1002079 206376 1002088
rect 206428 1002079 206430 1002088
rect 206376 1002050 206428 1002056
rect 206742 1002008 206798 1002017
rect 206742 1001943 206744 1001952
rect 206796 1001943 206798 1001952
rect 206744 1001914 206796 1001920
rect 207032 997762 207060 1002238
rect 207202 1002215 207258 1002224
rect 207020 997756 207072 997762
rect 207020 997698 207072 997704
rect 206192 997280 206244 997286
rect 206192 997222 206244 997228
rect 203522 995344 203578 995353
rect 203522 995279 203578 995288
rect 207400 994498 207428 1002510
rect 208400 1001972 208452 1001978
rect 208400 1001914 208452 1001920
rect 208412 994974 208440 1001914
rect 209884 995994 209912 1005110
rect 210056 1005032 210108 1005038
rect 210056 1004974 210108 1004980
rect 209872 995988 209924 995994
rect 209872 995930 209924 995936
rect 210068 995110 210096 1004974
rect 211160 1004828 211212 1004834
rect 211160 1004770 211212 1004776
rect 211172 1002674 211200 1004770
rect 211080 1002646 211200 1002674
rect 210882 1002144 210938 1002153
rect 211080 1002130 211108 1002646
rect 211250 1002552 211306 1002561
rect 211250 1002487 211252 1002496
rect 211304 1002487 211306 1002496
rect 211252 1002458 211304 1002464
rect 211250 1002280 211306 1002289
rect 211250 1002215 211252 1002224
rect 211304 1002215 211306 1002224
rect 211252 1002186 211304 1002192
rect 211080 1002102 211200 1002130
rect 210882 1002079 210884 1002088
rect 210936 1002079 210938 1002088
rect 210884 1002050 210936 1002056
rect 211172 996130 211200 1002102
rect 211816 996130 211844 1005994
rect 212538 1004728 212594 1004737
rect 212538 1004663 212540 1004672
rect 212592 1004663 212594 1004672
rect 217324 1004692 217376 1004698
rect 212540 1004634 212592 1004640
rect 217324 1004634 217376 1004640
rect 215944 1002516 215996 1002522
rect 215944 1002458 215996 1002464
rect 213184 1002244 213236 1002250
rect 213184 1002186 213236 1002192
rect 212540 1002108 212592 1002114
rect 212540 1002050 212592 1002056
rect 212078 1002008 212134 1002017
rect 212078 1001943 212080 1001952
rect 212132 1001943 212134 1001952
rect 212080 1001914 212132 1001920
rect 211160 996124 211212 996130
rect 211160 996066 211212 996072
rect 211804 996124 211856 996130
rect 211804 996066 211856 996072
rect 212552 995858 212580 1002050
rect 213196 995994 213224 1002186
rect 213920 1001972 213972 1001978
rect 213920 1001914 213972 1001920
rect 213184 995988 213236 995994
rect 213184 995930 213236 995936
rect 212540 995852 212592 995858
rect 212540 995794 212592 995800
rect 210056 995104 210108 995110
rect 210056 995046 210108 995052
rect 208400 994968 208452 994974
rect 208400 994910 208452 994916
rect 207388 994492 207440 994498
rect 207388 994434 207440 994440
rect 202328 994356 202380 994362
rect 202328 994298 202380 994304
rect 202142 993576 202198 993585
rect 202142 993511 202198 993520
rect 213932 992934 213960 1001914
rect 202880 992928 202932 992934
rect 186504 992870 186556 992876
rect 191838 992896 191894 992905
rect 164884 990888 164936 990894
rect 164884 990830 164936 990836
rect 170772 990888 170824 990894
rect 170772 990830 170824 990836
rect 154488 985720 154540 985726
rect 154488 985662 154540 985668
rect 160744 985720 160796 985726
rect 160744 985662 160796 985668
rect 154500 983620 154528 985662
rect 170784 983620 170812 990830
rect 186516 983634 186544 992870
rect 202880 992870 202932 992876
rect 213920 992928 213972 992934
rect 213920 992870 213972 992876
rect 191838 992831 191894 992840
rect 202892 983634 202920 992870
rect 215956 985998 215984 1002458
rect 217336 986678 217364 1004634
rect 228376 995081 228404 1006266
rect 249064 1006188 249116 1006194
rect 249064 1006130 249116 1006136
rect 229744 1006052 229796 1006058
rect 229744 1005994 229796 1006000
rect 247040 1006052 247092 1006058
rect 247040 1005994 247092 1006000
rect 229756 995858 229784 1005994
rect 247052 997898 247080 1005994
rect 247224 998300 247276 998306
rect 247224 998242 247276 998248
rect 246580 997892 246632 997898
rect 246580 997834 246632 997840
rect 247040 997892 247092 997898
rect 247040 997834 247092 997840
rect 229744 995852 229796 995858
rect 229744 995794 229796 995800
rect 246592 995761 246620 997834
rect 247236 997754 247264 998242
rect 247684 997824 247736 997830
rect 247684 997766 247736 997772
rect 247144 997726 247264 997754
rect 246948 997688 247000 997694
rect 246948 997630 247000 997636
rect 246764 997552 246816 997558
rect 246764 997494 246816 997500
rect 240874 995752 240930 995761
rect 240580 995710 240874 995738
rect 240874 995687 240930 995696
rect 244094 995752 244150 995761
rect 246578 995752 246634 995761
rect 244150 995710 244260 995738
rect 244094 995687 244150 995696
rect 246578 995687 246634 995696
rect 246212 995580 246264 995586
rect 246212 995522 246264 995528
rect 241978 995480 242034 995489
rect 231288 995438 231624 995466
rect 231932 995438 232268 995466
rect 232576 995438 232912 995466
rect 234416 995438 234568 995466
rect 228362 995072 228418 995081
rect 228362 995007 228418 995016
rect 231596 994362 231624 995438
rect 231584 994356 231636 994362
rect 231584 994298 231636 994304
rect 232240 994022 232268 995438
rect 232884 994974 232912 995438
rect 234540 995110 234568 995438
rect 234954 995246 234982 995452
rect 235612 995438 235948 995466
rect 236256 995438 236592 995466
rect 234942 995240 234994 995246
rect 234942 995182 234994 995188
rect 234528 995104 234580 995110
rect 234528 995046 234580 995052
rect 232872 994968 232924 994974
rect 232872 994910 232924 994916
rect 235920 994498 235948 995438
rect 236564 994809 236592 995438
rect 238680 995438 238740 995466
rect 239292 995438 239628 995466
rect 239936 995438 240088 995466
rect 241776 995438 241978 995466
rect 236550 994800 236606 994809
rect 236550 994735 236606 994744
rect 235908 994492 235960 994498
rect 235908 994434 235960 994440
rect 238680 994265 238708 995438
rect 239600 994537 239628 995438
rect 239586 994528 239642 994537
rect 239586 994463 239642 994472
rect 238666 994256 238722 994265
rect 238666 994191 238722 994200
rect 232228 994016 232280 994022
rect 240060 993993 240088 995438
rect 243818 995480 243874 995489
rect 242972 995438 243400 995466
rect 243616 995438 243818 995466
rect 241978 995415 242034 995424
rect 243372 995330 243400 995438
rect 245456 995438 245608 995466
rect 243818 995415 243874 995424
rect 245580 995382 245608 995438
rect 245568 995376 245620 995382
rect 244002 995344 244058 995353
rect 243372 995302 244002 995330
rect 245568 995318 245620 995324
rect 244002 995279 244058 995288
rect 243728 994492 243780 994498
rect 243728 994434 243780 994440
rect 243360 994356 243412 994362
rect 243360 994298 243412 994304
rect 243544 994356 243596 994362
rect 243544 994298 243596 994304
rect 232228 993958 232280 993964
rect 240046 993984 240102 993993
rect 240046 993919 240102 993928
rect 243372 993886 243400 994298
rect 243556 994022 243584 994298
rect 243740 994022 243768 994434
rect 243544 994016 243596 994022
rect 243544 993958 243596 993964
rect 243728 994016 243780 994022
rect 243728 993958 243780 993964
rect 246224 993886 246252 995522
rect 246776 995382 246804 997494
rect 246960 996441 246988 997630
rect 246946 996432 247002 996441
rect 246946 996367 247002 996376
rect 246948 996260 247000 996266
rect 246948 996202 247000 996208
rect 246764 995376 246816 995382
rect 246764 995318 246816 995324
rect 246960 994537 246988 996202
rect 247144 995353 247172 997726
rect 247130 995344 247186 995353
rect 247130 995279 247186 995288
rect 247696 994770 247724 997766
rect 247684 994764 247736 994770
rect 247684 994706 247736 994712
rect 246946 994528 247002 994537
rect 246946 994463 247002 994472
rect 249076 993993 249104 1006130
rect 249260 994022 249288 1006266
rect 255318 1006224 255374 1006233
rect 255318 1006159 255320 1006168
rect 255372 1006159 255374 1006168
rect 261850 1006224 261906 1006233
rect 261850 1006159 261852 1006168
rect 255320 1006130 255372 1006136
rect 261904 1006159 261906 1006168
rect 279424 1006188 279476 1006194
rect 261852 1006130 261904 1006136
rect 279424 1006130 279476 1006136
rect 252466 1006088 252522 1006097
rect 252466 1006023 252468 1006032
rect 252520 1006023 252522 1006032
rect 260194 1006088 260250 1006097
rect 260194 1006023 260196 1006032
rect 252468 1005994 252520 1006000
rect 260248 1006023 260250 1006032
rect 260196 1005994 260248 1006000
rect 263046 1005000 263102 1005009
rect 263046 1004935 263048 1004944
rect 263100 1004935 263102 1004944
rect 268384 1004964 268436 1004970
rect 263048 1004906 263100 1004912
rect 268384 1004906 268436 1004912
rect 256146 1002688 256202 1002697
rect 253204 1002652 253256 1002658
rect 256146 1002623 256148 1002632
rect 253204 1002594 253256 1002600
rect 256200 1002623 256202 1002632
rect 256148 1002594 256200 1002600
rect 251824 1002516 251876 1002522
rect 251824 1002458 251876 1002464
rect 250444 998164 250496 998170
rect 250444 998106 250496 998112
rect 250456 996033 250484 998106
rect 250628 997960 250680 997966
rect 250628 997902 250680 997908
rect 250640 997257 250668 997902
rect 250626 997248 250682 997257
rect 250626 997183 250682 997192
rect 251640 996736 251692 996742
rect 251638 996704 251640 996713
rect 251692 996704 251694 996713
rect 251638 996639 251694 996648
rect 250442 996024 250498 996033
rect 250442 995959 250498 995968
rect 251836 994809 251864 1002458
rect 252008 1002108 252060 1002114
rect 252008 1002050 252060 1002056
rect 252020 996266 252048 1002050
rect 252468 997824 252520 997830
rect 252466 997792 252468 997801
rect 252520 997792 252522 997801
rect 252466 997727 252522 997736
rect 252008 996260 252060 996266
rect 252008 996202 252060 996208
rect 253216 995246 253244 1002594
rect 254490 1002552 254546 1002561
rect 254490 1002487 254492 1002496
rect 254544 1002487 254546 1002496
rect 254492 1002458 254544 1002464
rect 261022 1002416 261078 1002425
rect 261022 1002351 261024 1002360
rect 261076 1002351 261078 1002360
rect 264244 1002380 264296 1002386
rect 261024 1002322 261076 1002328
rect 264244 1002322 264296 1002328
rect 262678 1002280 262734 1002289
rect 262678 1002215 262680 1002224
rect 262732 1002215 262734 1002224
rect 262680 1002186 262732 1002192
rect 254122 1002144 254178 1002153
rect 254122 1002079 254124 1002088
rect 254176 1002079 254178 1002088
rect 263874 1002144 263930 1002153
rect 263874 1002079 263876 1002088
rect 254124 1002050 254176 1002056
rect 263928 1002079 263930 1002088
rect 263876 1002050 263928 1002056
rect 255318 1002008 255374 1002017
rect 253388 1001972 253440 1001978
rect 255318 1001943 255320 1001952
rect 253388 1001914 253440 1001920
rect 255372 1001943 255374 1001952
rect 263506 1002008 263562 1002017
rect 263506 1001943 263508 1001952
rect 255320 1001914 255372 1001920
rect 263560 1001943 263562 1001952
rect 263508 1001914 263560 1001920
rect 253400 996742 253428 1001914
rect 259366 998336 259422 998345
rect 259366 998271 259368 998280
rect 259420 998271 259422 998280
rect 260932 998300 260984 998306
rect 259368 998242 259420 998248
rect 260932 998242 260984 998248
rect 253662 998200 253718 998209
rect 253662 998135 253664 998144
rect 253716 998135 253718 998144
rect 258170 998200 258226 998209
rect 258170 998135 258172 998144
rect 253664 998106 253716 998112
rect 258224 998135 258226 998144
rect 259460 998164 259512 998170
rect 258172 998106 258224 998112
rect 259460 998106 259512 998112
rect 254768 998096 254820 998102
rect 257344 998096 257396 998102
rect 254768 998038 254820 998044
rect 257342 998064 257344 998073
rect 257396 998064 257398 998073
rect 253664 997960 253716 997966
rect 253662 997928 253664 997937
rect 254584 997960 254636 997966
rect 253716 997928 253718 997937
rect 254584 997902 254636 997908
rect 253662 997863 253718 997872
rect 253388 996736 253440 996742
rect 253388 996678 253440 996684
rect 253204 995240 253256 995246
rect 253204 995182 253256 995188
rect 251822 994800 251878 994809
rect 251822 994735 251878 994744
rect 254596 994362 254624 997902
rect 254584 994356 254636 994362
rect 254584 994298 254636 994304
rect 254780 994265 254808 998038
rect 257342 997999 257398 998008
rect 256516 997960 256568 997966
rect 256514 997928 256516 997937
rect 256568 997928 256570 997937
rect 258170 997928 258226 997937
rect 256514 997863 256570 997872
rect 257356 997886 258170 997914
rect 256974 997792 257030 997801
rect 255976 997750 256974 997778
rect 255976 997558 256004 997750
rect 256974 997727 257030 997736
rect 255964 997552 256016 997558
rect 255964 997494 256016 997500
rect 257356 995586 257384 997886
rect 258170 997863 258226 997872
rect 258998 997792 259054 997801
rect 258092 997750 258998 997778
rect 258092 997694 258120 997750
rect 258998 997727 259054 997736
rect 258080 997688 258132 997694
rect 258080 997630 258132 997636
rect 257344 995580 257396 995586
rect 257344 995522 257396 995528
rect 259472 995110 259500 998106
rect 259828 998096 259880 998102
rect 259826 998064 259828 998073
rect 259880 998064 259882 998073
rect 259826 997999 259882 998008
rect 260196 997960 260248 997966
rect 260194 997928 260196 997937
rect 260248 997928 260250 997937
rect 260194 997863 260250 997872
rect 259460 995104 259512 995110
rect 259460 995046 259512 995052
rect 260944 994974 260972 998242
rect 262312 998096 262364 998102
rect 262312 998038 262364 998044
rect 261850 997792 261906 997801
rect 261128 997736 261850 997754
rect 261128 997727 261906 997736
rect 261128 997726 261892 997727
rect 261128 995994 261156 997726
rect 261116 995988 261168 995994
rect 261116 995930 261168 995936
rect 262324 995858 262352 998038
rect 262496 997960 262548 997966
rect 262496 997902 262548 997908
rect 262508 996130 262536 997902
rect 262496 996124 262548 996130
rect 262496 996066 262548 996072
rect 264256 995858 264284 1002322
rect 265808 1002244 265860 1002250
rect 265808 1002186 265860 1002192
rect 265624 1001972 265676 1001978
rect 265624 1001914 265676 1001920
rect 262312 995852 262364 995858
rect 262312 995794 262364 995800
rect 264244 995852 264296 995858
rect 264244 995794 264296 995800
rect 260932 994968 260984 994974
rect 260932 994910 260984 994916
rect 254766 994256 254822 994265
rect 254766 994191 254822 994200
rect 249248 994016 249300 994022
rect 249062 993984 249118 993993
rect 249248 993958 249300 993964
rect 249062 993919 249118 993928
rect 243360 993880 243412 993886
rect 243360 993822 243412 993828
rect 246212 993880 246264 993886
rect 246212 993822 246264 993828
rect 251454 992896 251510 992905
rect 251454 992831 251510 992840
rect 217324 986672 217376 986678
rect 217324 986614 217376 986620
rect 219440 986672 219492 986678
rect 219440 986614 219492 986620
rect 215944 985992 215996 985998
rect 215944 985934 215996 985940
rect 186516 983606 186990 983634
rect 202892 983606 203182 983634
rect 219452 983620 219480 986614
rect 235632 985992 235684 985998
rect 235632 985934 235684 985940
rect 235644 983620 235672 985934
rect 251468 983634 251496 992831
rect 265636 990894 265664 1001914
rect 265820 996130 265848 1002186
rect 267004 1002108 267056 1002114
rect 267004 1002050 267056 1002056
rect 265808 996124 265860 996130
rect 265808 996066 265860 996072
rect 267016 991506 267044 1002050
rect 267004 991500 267056 991506
rect 267004 991442 267056 991448
rect 265624 990888 265676 990894
rect 265624 990830 265676 990836
rect 267648 990888 267700 990894
rect 267648 990830 267700 990836
rect 267660 985334 267688 990830
rect 268396 985998 268424 1004906
rect 278136 997824 278188 997830
rect 278136 997766 278188 997772
rect 278148 994430 278176 997766
rect 279436 995081 279464 1006130
rect 280804 1006052 280856 1006058
rect 280804 1005994 280856 1006000
rect 298744 1006052 298796 1006058
rect 298744 1005994 298796 1006000
rect 280816 995994 280844 1005994
rect 298756 1001894 298784 1005994
rect 298572 1001866 298784 1001894
rect 298098 997928 298154 997937
rect 298098 997863 298154 997872
rect 280804 995988 280856 995994
rect 280804 995930 280856 995936
rect 282734 995752 282790 995761
rect 287978 995752 288034 995761
rect 282790 995710 282854 995738
rect 287822 995710 287978 995738
rect 282734 995687 282790 995696
rect 291750 995752 291806 995761
rect 291502 995710 291750 995738
rect 287978 995687 288034 995696
rect 293498 995752 293554 995761
rect 293342 995710 293498 995738
rect 291750 995687 291806 995696
rect 293498 995687 293554 995696
rect 295062 995752 295118 995761
rect 298112 995738 298140 997863
rect 298376 997076 298428 997082
rect 298376 997018 298428 997024
rect 295118 995710 295182 995738
rect 297836 995710 298140 995738
rect 295062 995687 295118 995696
rect 296166 995616 296222 995625
rect 295826 995574 296166 995602
rect 296166 995551 296222 995560
rect 283484 995110 283512 995452
rect 283472 995104 283524 995110
rect 279422 995072 279478 995081
rect 283472 995046 283524 995052
rect 279422 995007 279478 995016
rect 284128 994974 284156 995452
rect 285982 995438 286272 995466
rect 286244 995353 286272 995438
rect 286230 995344 286286 995353
rect 286230 995279 286286 995288
rect 284116 994968 284168 994974
rect 284116 994910 284168 994916
rect 278136 994424 278188 994430
rect 278136 994366 278188 994372
rect 286520 994022 286548 995452
rect 287164 994838 287192 995452
rect 287152 994832 287204 994838
rect 290292 994809 290320 995452
rect 287152 994774 287204 994780
rect 290278 994800 290334 994809
rect 290278 994735 290334 994744
rect 290844 994265 290872 995452
rect 292146 995438 292528 995466
rect 292500 995246 292528 995438
rect 294156 995438 294538 995466
rect 297022 995438 297404 995466
rect 292488 995240 292540 995246
rect 292488 995182 292540 995188
rect 294156 994294 294184 995438
rect 297376 995330 297404 995438
rect 297836 995330 297864 995710
rect 297376 995302 297864 995330
rect 294144 994288 294196 994294
rect 290830 994256 290886 994265
rect 294144 994230 294196 994236
rect 290830 994191 290886 994200
rect 298388 994022 298416 997018
rect 298572 994634 298600 1001866
rect 298744 997756 298796 997762
rect 298744 997698 298796 997704
rect 298756 996985 298784 997698
rect 298742 996976 298798 996985
rect 298742 996911 298798 996920
rect 298940 995858 298968 1006266
rect 300124 1006188 300176 1006194
rect 300124 1006130 300176 1006136
rect 299388 997620 299440 997626
rect 299388 997562 299440 997568
rect 299400 996577 299428 997562
rect 299386 996568 299442 996577
rect 299386 996503 299442 996512
rect 299386 996296 299442 996305
rect 299386 996231 299442 996240
rect 298928 995852 298980 995858
rect 298928 995794 298980 995800
rect 299400 995761 299428 996231
rect 299846 996024 299902 996033
rect 299584 995982 299846 996010
rect 299386 995752 299442 995761
rect 299386 995687 299442 995696
rect 299202 995616 299258 995625
rect 299584 995602 299612 995982
rect 299846 995959 299902 995968
rect 299258 995574 299612 995602
rect 299202 995551 299258 995560
rect 298560 994628 298612 994634
rect 298560 994570 298612 994576
rect 300136 994265 300164 1006130
rect 300320 996441 300348 1006402
rect 361394 1006360 361450 1006369
rect 311808 1006324 311860 1006330
rect 361394 1006295 361396 1006304
rect 311808 1006266 311860 1006272
rect 361448 1006295 361450 1006304
rect 361396 1006266 361448 1006272
rect 306102 1006224 306158 1006233
rect 306102 1006159 306104 1006168
rect 306156 1006159 306158 1006168
rect 306104 1006130 306156 1006136
rect 311820 1006097 311848 1006266
rect 357346 1006224 357402 1006233
rect 357346 1006159 357348 1006168
rect 357400 1006159 357402 1006168
rect 362224 1006188 362276 1006194
rect 357348 1006130 357400 1006136
rect 362224 1006130 362276 1006136
rect 301686 1006088 301742 1006097
rect 301686 1006023 301742 1006032
rect 303250 1006088 303306 1006097
rect 303250 1006023 303252 1006032
rect 301504 1002108 301556 1002114
rect 301504 1002050 301556 1002056
rect 300306 996432 300362 996441
rect 300306 996367 300362 996376
rect 300122 994256 300178 994265
rect 300122 994191 300178 994200
rect 301516 994158 301544 1002050
rect 301700 996033 301728 1006023
rect 303304 1006023 303306 1006032
rect 304078 1006088 304134 1006097
rect 304078 1006023 304080 1006032
rect 303252 1005994 303304 1006000
rect 304132 1006023 304134 1006032
rect 311806 1006088 311862 1006097
rect 311806 1006023 311862 1006032
rect 314658 1006088 314714 1006097
rect 354862 1006088 354918 1006097
rect 314658 1006023 314660 1006032
rect 304080 1005994 304132 1006000
rect 314712 1006023 314714 1006032
rect 319444 1006052 319496 1006058
rect 314660 1005994 314712 1006000
rect 354862 1006023 354918 1006032
rect 356886 1006088 356942 1006097
rect 356886 1006023 356888 1006032
rect 319444 1005994 319496 1006000
rect 304080 1005848 304132 1005854
rect 304078 1005816 304080 1005825
rect 304132 1005816 304134 1005825
rect 304078 1005751 304134 1005760
rect 313830 1005000 313886 1005009
rect 313830 1004935 313832 1004944
rect 313884 1004935 313886 1004944
rect 316040 1004964 316092 1004970
rect 313832 1004906 313884 1004912
rect 316040 1004906 316092 1004912
rect 314658 1004864 314714 1004873
rect 314658 1004799 314660 1004808
rect 314712 1004799 314714 1004808
rect 314660 1004770 314712 1004776
rect 315486 1004728 315542 1004737
rect 315486 1004663 315488 1004672
rect 315540 1004663 315542 1004672
rect 315488 1004634 315540 1004640
rect 304906 1002144 304962 1002153
rect 304906 1002079 304908 1002088
rect 304960 1002079 304962 1002088
rect 310150 1002144 310206 1002153
rect 310150 1002079 310152 1002088
rect 304908 1002050 304960 1002056
rect 310204 1002079 310206 1002088
rect 311900 1002108 311952 1002114
rect 310152 1002050 310204 1002056
rect 311900 1002050 311952 1002056
rect 310978 1002008 311034 1002017
rect 310978 1001943 310980 1001952
rect 311032 1001943 311034 1001952
rect 310980 1001914 311032 1001920
rect 308954 998608 309010 998617
rect 303252 998572 303304 998578
rect 308954 998543 308956 998552
rect 303252 998514 303304 998520
rect 309008 998543 309010 998552
rect 308956 998514 309008 998520
rect 302884 998300 302936 998306
rect 302884 998242 302936 998248
rect 301686 996024 301742 996033
rect 301686 995959 301742 995968
rect 302896 995761 302924 998242
rect 303264 997937 303292 998514
rect 307298 998472 307354 998481
rect 304264 998436 304316 998442
rect 307298 998407 307300 998416
rect 304264 998378 304316 998384
rect 307352 998407 307354 998416
rect 307300 998378 307352 998384
rect 303250 997928 303306 997937
rect 303068 997892 303120 997898
rect 303250 997863 303306 997872
rect 303068 997834 303120 997840
rect 302882 995752 302938 995761
rect 302882 995687 302938 995696
rect 303080 995246 303108 997834
rect 303252 997280 303304 997286
rect 303250 997248 303252 997257
rect 303304 997248 303306 997257
rect 303250 997183 303306 997192
rect 303068 995240 303120 995246
rect 303068 995182 303120 995188
rect 304276 994838 304304 998378
rect 306102 998336 306158 998345
rect 306102 998271 306104 998280
rect 306156 998271 306158 998280
rect 306104 998242 306156 998248
rect 308126 998200 308182 998209
rect 305644 998164 305696 998170
rect 308126 998135 308128 998144
rect 305644 998106 305696 998112
rect 308180 998135 308182 998144
rect 308128 998106 308180 998112
rect 304448 998028 304500 998034
rect 304448 997970 304500 997976
rect 304460 997286 304488 997970
rect 305274 997928 305330 997937
rect 305274 997863 305276 997872
rect 305328 997863 305330 997872
rect 305276 997834 305328 997840
rect 304448 997280 304500 997286
rect 304448 997222 304500 997228
rect 305656 995110 305684 998106
rect 306930 998064 306986 998073
rect 310610 998064 310666 998073
rect 306930 997999 306932 998008
rect 306984 997999 306986 998008
rect 308404 998028 308456 998034
rect 306932 997970 306984 997976
rect 310610 997999 310612 998008
rect 308404 997970 308456 997976
rect 310664 997999 310666 998008
rect 310612 997970 310664 997976
rect 307024 997892 307076 997898
rect 307024 997834 307076 997840
rect 305644 995104 305696 995110
rect 305644 995046 305696 995052
rect 304264 994832 304316 994838
rect 307036 994809 307064 997834
rect 307758 997792 307814 997801
rect 307220 997750 307758 997778
rect 307220 997082 307248 997750
rect 307758 997727 307814 997736
rect 307208 997076 307260 997082
rect 307208 997018 307260 997024
rect 308416 994974 308444 997970
rect 308954 997928 309010 997937
rect 308954 997863 308956 997872
rect 309008 997863 309010 997872
rect 308956 997834 309008 997840
rect 310610 997792 310666 997801
rect 310532 997736 310610 997754
rect 311912 997762 311940 1002050
rect 313280 1001972 313332 1001978
rect 313280 1001914 313332 1001920
rect 310532 997727 310666 997736
rect 311900 997756 311952 997762
rect 310532 997726 310652 997727
rect 310532 997626 310560 997726
rect 311900 997698 311952 997704
rect 310520 997620 310572 997626
rect 310520 997562 310572 997568
rect 313292 995994 313320 1001914
rect 316052 996130 316080 1004906
rect 316684 1004828 316736 1004834
rect 316684 1004770 316736 1004776
rect 316040 996124 316092 996130
rect 316040 996066 316092 996072
rect 313280 995988 313332 995994
rect 313280 995930 313332 995936
rect 308404 994968 308456 994974
rect 308404 994910 308456 994916
rect 304264 994774 304316 994780
rect 307022 994800 307078 994809
rect 307022 994735 307078 994744
rect 316408 994424 316460 994430
rect 316408 994366 316460 994372
rect 301504 994152 301556 994158
rect 301504 994094 301556 994100
rect 286508 994016 286560 994022
rect 286508 993958 286560 993964
rect 298376 994016 298428 994022
rect 298376 993958 298428 993964
rect 284300 991500 284352 991506
rect 284300 991442 284352 991448
rect 268384 985992 268436 985998
rect 268384 985934 268436 985940
rect 267660 985306 267780 985334
rect 267752 983634 267780 985306
rect 251468 983606 251850 983634
rect 267752 983606 268134 983634
rect 284312 983620 284340 991442
rect 300492 985992 300544 985998
rect 300492 985934 300544 985940
rect 300504 983620 300532 985934
rect 316420 983634 316448 994366
rect 316696 992934 316724 1004770
rect 318064 1004692 318116 1004698
rect 318064 1004634 318116 1004640
rect 316684 992928 316736 992934
rect 316684 992870 316736 992876
rect 318076 991506 318104 1004634
rect 318064 991500 318116 991506
rect 318064 991442 318116 991448
rect 319456 990146 319484 1005994
rect 353208 1004828 353260 1004834
rect 353208 1004770 353260 1004776
rect 351828 1001972 351880 1001978
rect 351828 1001914 351880 1001920
rect 351840 998442 351868 1001914
rect 353220 1001230 353248 1004770
rect 354404 1004692 354456 1004698
rect 354404 1004634 354456 1004640
rect 354034 1002008 354090 1002017
rect 354034 1001943 354036 1001952
rect 354088 1001943 354090 1001952
rect 354036 1001914 354088 1001920
rect 353208 1001224 353260 1001230
rect 353208 1001166 353260 1001172
rect 351828 998436 351880 998442
rect 351828 998378 351880 998384
rect 354416 994498 354444 1004634
rect 354876 1001366 354904 1006023
rect 356940 1006023 356942 1006032
rect 360844 1006052 360896 1006058
rect 356888 1005994 356940 1006000
rect 360844 1005994 360896 1006000
rect 360568 1005576 360620 1005582
rect 360566 1005544 360568 1005553
rect 360620 1005544 360622 1005553
rect 360566 1005479 360622 1005488
rect 358544 1005440 358596 1005446
rect 358542 1005408 358544 1005417
rect 358596 1005408 358598 1005417
rect 358542 1005343 358598 1005352
rect 357716 1005304 357768 1005310
rect 357714 1005272 357716 1005281
rect 357768 1005272 357770 1005281
rect 357714 1005207 357770 1005216
rect 355690 1004864 355746 1004873
rect 355690 1004799 355692 1004808
rect 355744 1004799 355746 1004808
rect 355692 1004770 355744 1004776
rect 356518 1004728 356574 1004737
rect 356518 1004663 356520 1004672
rect 356572 1004663 356574 1004672
rect 356520 1004634 356572 1004640
rect 360568 1003944 360620 1003950
rect 360566 1003912 360568 1003921
rect 360620 1003912 360622 1003921
rect 360566 1003847 360622 1003856
rect 355690 1003368 355746 1003377
rect 355690 1003303 355692 1003312
rect 355744 1003303 355746 1003312
rect 355692 1003274 355744 1003280
rect 358544 1002584 358596 1002590
rect 358542 1002552 358544 1002561
rect 358596 1002552 358598 1002561
rect 358542 1002487 358598 1002496
rect 359370 1002280 359426 1002289
rect 357348 1002244 357400 1002250
rect 359370 1002215 359372 1002224
rect 357348 1002186 357400 1002192
rect 359424 1002215 359426 1002224
rect 359372 1002186 359424 1002192
rect 354864 1001360 354916 1001366
rect 354864 1001302 354916 1001308
rect 357360 997082 357388 1002186
rect 359370 1002008 359426 1002017
rect 358728 1001972 358780 1001978
rect 359370 1001943 359372 1001952
rect 358728 1001914 358780 1001920
rect 359424 1001943 359426 1001952
rect 359372 1001914 359424 1001920
rect 357348 997076 357400 997082
rect 357348 997018 357400 997024
rect 358740 995042 358768 1001914
rect 360856 995178 360884 1005994
rect 361394 1005000 361450 1005009
rect 361394 1004935 361396 1004944
rect 361448 1004935 361450 1004944
rect 361396 1004906 361448 1004912
rect 362236 997218 362264 1006130
rect 363418 1006088 363474 1006097
rect 363418 1006023 363420 1006032
rect 363472 1006023 363474 1006032
rect 363420 1005994 363472 1006000
rect 364892 1004964 364944 1004970
rect 364892 1004906 364944 1004912
rect 362590 1004864 362646 1004873
rect 362590 1004799 362592 1004808
rect 362644 1004799 362646 1004808
rect 362592 1004770 362644 1004776
rect 364246 1004728 364302 1004737
rect 364246 1004663 364248 1004672
rect 364300 1004663 364302 1004672
rect 364248 1004634 364300 1004640
rect 363604 1003332 363656 1003338
rect 363604 1003274 363656 1003280
rect 362224 997212 362276 997218
rect 362224 997154 362276 997160
rect 360844 995172 360896 995178
rect 360844 995114 360896 995120
rect 358728 995036 358780 995042
rect 358728 994978 358780 994984
rect 363616 994634 363644 1003274
rect 364904 995858 364932 1004906
rect 365260 1004828 365312 1004834
rect 365260 1004770 365312 1004776
rect 365076 1002312 365128 1002318
rect 365074 1002280 365076 1002289
rect 365128 1002280 365130 1002289
rect 365074 1002215 365130 1002224
rect 365076 1002040 365128 1002046
rect 365074 1002008 365076 1002017
rect 365128 1002008 365130 1002017
rect 365074 1001943 365130 1001952
rect 365272 997626 365300 1004770
rect 366364 1004692 366416 1004698
rect 366364 1004634 366416 1004640
rect 365904 1002176 365956 1002182
rect 365902 1002144 365904 1002153
rect 365956 1002144 365958 1002153
rect 365902 1002079 365958 1002088
rect 365260 997620 365312 997626
rect 365260 997562 365312 997568
rect 366376 995994 366404 1004634
rect 367928 1002312 367980 1002318
rect 367928 1002254 367980 1002260
rect 367744 1002040 367796 1002046
rect 367744 1001982 367796 1001988
rect 366364 995988 366416 995994
rect 366364 995930 366416 995936
rect 364892 995852 364944 995858
rect 364892 995794 364944 995800
rect 363604 994628 363656 994634
rect 363604 994570 363656 994576
rect 354404 994492 354456 994498
rect 354404 994434 354456 994440
rect 364984 992928 365036 992934
rect 364984 992870 365036 992876
rect 349160 991500 349212 991506
rect 349160 991442 349212 991448
rect 319444 990140 319496 990146
rect 319444 990082 319496 990088
rect 332968 990140 333020 990146
rect 332968 990082 333020 990088
rect 316420 983606 316802 983634
rect 332980 983620 333008 990082
rect 349172 983620 349200 991442
rect 364996 983634 365024 992870
rect 367756 991506 367784 1001982
rect 367940 992934 367968 1002254
rect 369124 1002176 369176 1002182
rect 369124 1002118 369176 1002124
rect 367928 992928 367980 992934
rect 367928 992870 367980 992876
rect 367744 991500 367796 991506
rect 367744 991442 367796 991448
rect 369136 990146 369164 1002118
rect 369872 1002046 369900 1006810
rect 430856 1006800 430908 1006806
rect 430854 1006768 430856 1006777
rect 434628 1006800 434680 1006806
rect 430908 1006768 430910 1006777
rect 373264 1006732 373316 1006738
rect 506204 1006800 506256 1006806
rect 434628 1006742 434680 1006748
rect 506202 1006768 506204 1006777
rect 506256 1006768 506258 1006777
rect 430854 1006703 430910 1006712
rect 373264 1006674 373316 1006680
rect 371884 1005440 371936 1005446
rect 371884 1005382 371936 1005388
rect 371148 1002584 371200 1002590
rect 371148 1002526 371200 1002532
rect 369860 1002040 369912 1002046
rect 369860 1001982 369912 1001988
rect 371160 997762 371188 1002526
rect 371896 998578 371924 1005382
rect 371884 998572 371936 998578
rect 371884 998514 371936 998520
rect 373276 998345 373304 1006674
rect 430028 1006528 430080 1006534
rect 430026 1006496 430028 1006505
rect 433984 1006528 434036 1006534
rect 430080 1006496 430082 1006505
rect 431682 1006496 431738 1006505
rect 430026 1006431 430082 1006440
rect 431512 1006454 431682 1006482
rect 429198 1006360 429254 1006369
rect 375012 1006324 375064 1006330
rect 375012 1006266 375064 1006272
rect 402244 1006324 402296 1006330
rect 429198 1006295 429200 1006304
rect 402244 1006266 402296 1006272
rect 429252 1006295 429254 1006304
rect 429200 1006266 429252 1006272
rect 375024 1003270 375052 1006266
rect 382924 1006052 382976 1006058
rect 382924 1005994 382976 1006000
rect 400864 1006052 400916 1006058
rect 400864 1005994 400916 1006000
rect 378784 1005576 378836 1005582
rect 378784 1005518 378836 1005524
rect 376760 1005304 376812 1005310
rect 376760 1005246 376812 1005252
rect 375380 1003944 375432 1003950
rect 375380 1003886 375432 1003892
rect 375012 1003264 375064 1003270
rect 375012 1003206 375064 1003212
rect 374644 1002040 374696 1002046
rect 374644 1001982 374696 1001988
rect 373262 998336 373318 998345
rect 373262 998271 373318 998280
rect 371148 997756 371200 997762
rect 371148 997698 371200 997704
rect 372528 997756 372580 997762
rect 372528 997698 372580 997704
rect 372344 997620 372396 997626
rect 372344 997562 372396 997568
rect 372356 997257 372384 997562
rect 372342 997248 372398 997257
rect 372342 997183 372398 997192
rect 372344 997076 372396 997082
rect 372344 997018 372396 997024
rect 372356 996033 372384 997018
rect 372540 996441 372568 997698
rect 372712 997212 372764 997218
rect 372712 997154 372764 997160
rect 372526 996432 372582 996441
rect 372526 996367 372582 996376
rect 372342 996024 372398 996033
rect 372342 995959 372398 995968
rect 372724 994906 372752 997154
rect 374656 994945 374684 1001982
rect 375392 997762 375420 1003886
rect 376772 999190 376800 1005246
rect 377956 1001360 378008 1001366
rect 377956 1001302 378008 1001308
rect 376760 999184 376812 999190
rect 376760 999126 376812 999132
rect 377968 999002 377996 1001302
rect 377968 998974 378180 999002
rect 375380 997756 375432 997762
rect 375380 997698 375432 997704
rect 378152 995314 378180 998974
rect 378796 997830 378824 1005518
rect 379428 1003264 379480 1003270
rect 379428 1003206 379480 1003212
rect 379440 997966 379468 1003206
rect 380900 1001224 380952 1001230
rect 380900 1001166 380952 1001172
rect 379428 997960 379480 997966
rect 379428 997902 379480 997908
rect 378784 997824 378836 997830
rect 378784 997766 378836 997772
rect 378600 997756 378652 997762
rect 378600 997698 378652 997704
rect 378140 995308 378192 995314
rect 378140 995250 378192 995256
rect 374642 994936 374698 994945
rect 372712 994900 372764 994906
rect 374642 994871 374698 994880
rect 372712 994842 372764 994848
rect 378612 994770 378640 997698
rect 380912 995489 380940 1001166
rect 382740 998572 382792 998578
rect 382740 998514 382792 998520
rect 382280 998436 382332 998442
rect 382280 998378 382332 998384
rect 380898 995480 380954 995489
rect 380898 995415 380954 995424
rect 382292 995217 382320 998378
rect 382752 995586 382780 998514
rect 382936 996130 382964 1005994
rect 383384 999184 383436 999190
rect 383384 999126 383436 999132
rect 383200 997960 383252 997966
rect 383200 997902 383252 997908
rect 382924 996124 382976 996130
rect 382924 996066 382976 996072
rect 383212 995761 383240 997902
rect 383396 996713 383424 999126
rect 383568 997824 383620 997830
rect 383620 997772 383700 997778
rect 383568 997766 383700 997772
rect 383580 997750 383700 997766
rect 383382 996704 383438 996713
rect 383382 996639 383438 996648
rect 383198 995752 383254 995761
rect 383198 995687 383254 995696
rect 382740 995580 382792 995586
rect 382740 995522 382792 995528
rect 383672 995330 383700 997750
rect 399944 997756 399996 997762
rect 399944 997698 399996 997704
rect 399956 996985 399984 997698
rect 400128 997144 400180 997150
rect 400128 997086 400180 997092
rect 399942 996976 399998 996985
rect 399942 996911 399998 996920
rect 400140 996441 400168 997086
rect 400126 996432 400182 996441
rect 400126 996367 400182 996376
rect 400876 995994 400904 1005994
rect 400864 995988 400916 995994
rect 400864 995930 400916 995936
rect 402256 995858 402284 1006266
rect 431512 1006194 431540 1006454
rect 433984 1006470 434036 1006476
rect 431682 1006431 431738 1006440
rect 431684 1006256 431736 1006262
rect 431682 1006224 431684 1006233
rect 431736 1006224 431738 1006233
rect 431500 1006188 431552 1006194
rect 431682 1006159 431738 1006168
rect 431500 1006130 431552 1006136
rect 421838 1006088 421894 1006097
rect 421838 1006023 421894 1006032
rect 428370 1006088 428426 1006097
rect 428370 1006023 428372 1006032
rect 420644 1004828 420696 1004834
rect 420644 1004770 420696 1004776
rect 419448 1001972 419500 1001978
rect 419448 1001914 419500 1001920
rect 402244 995852 402296 995858
rect 402244 995794 402296 995800
rect 385682 995752 385738 995761
rect 386694 995752 386750 995761
rect 385738 995710 385986 995738
rect 385682 995687 385738 995696
rect 387890 995752 387946 995761
rect 387826 995710 387890 995738
rect 386694 995687 386750 995696
rect 387890 995687 387946 995696
rect 388166 995752 388222 995761
rect 391938 995752 391994 995761
rect 388222 995710 388378 995738
rect 388166 995687 388222 995696
rect 396538 995752 396594 995761
rect 391994 995710 392150 995738
rect 396382 995710 396538 995738
rect 391938 995687 391994 995696
rect 396538 995687 396594 995696
rect 416134 995752 416190 995761
rect 416134 995687 416190 995696
rect 384960 995586 385342 995602
rect 384948 995580 385342 995586
rect 385000 995574 385342 995580
rect 384948 995522 385000 995528
rect 386708 995518 386736 995687
rect 386696 995512 386748 995518
rect 384316 995438 384698 995466
rect 386696 995454 386748 995460
rect 388628 995512 388680 995518
rect 415398 995480 415454 995489
rect 388680 995460 389022 995466
rect 388628 995454 389022 995460
rect 388640 995438 389022 995454
rect 384316 995330 384344 995438
rect 383672 995302 384344 995330
rect 382278 995208 382334 995217
rect 389652 995178 389680 995452
rect 382278 995143 382334 995152
rect 389640 995172 389692 995178
rect 389640 995114 389692 995120
rect 378600 994764 378652 994770
rect 378600 994706 378652 994712
rect 392688 994498 392716 995452
rect 393332 994906 393360 995452
rect 393320 994900 393372 994906
rect 393320 994842 393372 994848
rect 393976 994634 394004 995452
rect 395172 994945 395200 995452
rect 395158 994936 395214 994945
rect 395158 994871 395214 994880
rect 397012 994770 397040 995452
rect 397656 995314 397684 995452
rect 397644 995308 397696 995314
rect 397644 995250 397696 995256
rect 398852 995042 398880 995452
rect 415398 995415 415400 995424
rect 415452 995415 415454 995424
rect 415400 995386 415452 995392
rect 416148 995293 416176 995687
rect 416136 995287 416188 995293
rect 416136 995229 416188 995235
rect 398840 995036 398892 995042
rect 398840 994978 398892 994984
rect 419460 994974 419488 1001914
rect 419448 994968 419500 994974
rect 419448 994910 419500 994916
rect 397000 994764 397052 994770
rect 397000 994706 397052 994712
rect 420656 994702 420684 1004770
rect 421852 1002726 421880 1006023
rect 428424 1006023 428426 1006032
rect 428372 1005994 428424 1006000
rect 425520 1005712 425572 1005718
rect 425518 1005680 425520 1005689
rect 425572 1005680 425574 1005689
rect 425518 1005615 425574 1005624
rect 427176 1005576 427228 1005582
rect 427174 1005544 427176 1005553
rect 427228 1005544 427230 1005553
rect 427174 1005479 427230 1005488
rect 428372 1005440 428424 1005446
rect 428370 1005408 428372 1005417
rect 428424 1005408 428426 1005417
rect 428370 1005343 428426 1005352
rect 423496 1005304 423548 1005310
rect 423494 1005272 423496 1005281
rect 423548 1005272 423550 1005281
rect 423494 1005207 423550 1005216
rect 431222 1005000 431278 1005009
rect 431222 1004935 431224 1004944
rect 431276 1004935 431278 1004944
rect 433524 1004964 433576 1004970
rect 431224 1004906 431276 1004912
rect 433524 1004906 433576 1004912
rect 422666 1004864 422722 1004873
rect 422666 1004799 422668 1004808
rect 422720 1004799 422722 1004808
rect 432050 1004864 432106 1004873
rect 432050 1004799 432052 1004808
rect 422668 1004770 422720 1004776
rect 432104 1004799 432106 1004808
rect 432052 1004770 432104 1004776
rect 430026 1004728 430082 1004737
rect 430026 1004663 430028 1004672
rect 430080 1004663 430082 1004672
rect 431960 1004692 432012 1004698
rect 430028 1004634 430080 1004640
rect 431960 1004634 432012 1004640
rect 424692 1004080 424744 1004086
rect 424690 1004048 424692 1004057
rect 424744 1004048 424746 1004057
rect 424690 1003983 424746 1003992
rect 426348 1003944 426400 1003950
rect 426346 1003912 426348 1003921
rect 426400 1003912 426402 1003921
rect 426346 1003847 426402 1003856
rect 421840 1002720 421892 1002726
rect 421840 1002662 421892 1002668
rect 423496 1002584 423548 1002590
rect 423494 1002552 423496 1002561
rect 423548 1002552 423550 1002561
rect 423494 1002487 423550 1002496
rect 425518 1002144 425574 1002153
rect 424508 1002108 424560 1002114
rect 425518 1002079 425520 1002088
rect 424508 1002050 424560 1002056
rect 425572 1002079 425574 1002088
rect 427542 1002144 427598 1002153
rect 427542 1002079 427544 1002088
rect 425520 1002050 425572 1002056
rect 427596 1002079 427598 1002088
rect 429844 1002108 429896 1002114
rect 427544 1002050 427596 1002056
rect 429844 1002050 429896 1002056
rect 423588 1002040 423640 1002046
rect 421470 1002008 421526 1002017
rect 424324 1002040 424376 1002046
rect 423588 1001982 423640 1001988
rect 424322 1002008 424324 1002017
rect 424376 1002008 424378 1002017
rect 421470 1001943 421472 1001952
rect 421524 1001943 421526 1001952
rect 421472 1001914 421524 1001920
rect 423600 998442 423628 1001982
rect 424322 1001943 424378 1001952
rect 424520 998578 424548 1002050
rect 425150 1002008 425206 1002017
rect 426346 1002008 426402 1002017
rect 425206 1001966 425744 1001994
rect 425150 1001943 425206 1001952
rect 424508 998572 424560 998578
rect 424508 998514 424560 998520
rect 423588 998436 423640 998442
rect 423588 998378 423640 998384
rect 425716 995110 425744 1001966
rect 429198 1002008 429254 1002017
rect 426402 1001966 427124 1001994
rect 426346 1001943 426402 1001952
rect 427096 998714 427124 1001966
rect 429198 1001943 429200 1001952
rect 429252 1001943 429254 1001952
rect 429200 1001914 429252 1001920
rect 429856 1001230 429884 1002050
rect 431224 1001972 431276 1001978
rect 431224 1001914 431276 1001920
rect 429844 1001224 429896 1001230
rect 429844 1001166 429896 1001172
rect 427084 998708 427136 998714
rect 427084 998650 427136 998656
rect 431236 997626 431264 1001914
rect 431972 997762 432000 1004634
rect 433338 1002144 433394 1002153
rect 433338 1002079 433340 1002088
rect 433392 1002079 433394 1002088
rect 433340 1002050 433392 1002056
rect 432878 1002008 432934 1002017
rect 432878 1001943 432880 1001952
rect 432932 1001943 432934 1001952
rect 432880 1001914 432932 1001920
rect 431960 997756 432012 997762
rect 431960 997698 432012 997704
rect 431224 997620 431276 997626
rect 431224 997562 431276 997568
rect 433536 996130 433564 1004906
rect 433524 996124 433576 996130
rect 433524 996066 433576 996072
rect 425704 995104 425756 995110
rect 425704 995046 425756 995052
rect 433996 994838 434024 1006470
rect 434640 1006330 434668 1006742
rect 506202 1006703 506258 1006712
rect 508226 1006496 508282 1006505
rect 447784 1006460 447836 1006466
rect 508226 1006431 508228 1006440
rect 447784 1006402 447836 1006408
rect 508280 1006431 508282 1006440
rect 508228 1006402 508280 1006408
rect 434628 1006324 434680 1006330
rect 434628 1006266 434680 1006272
rect 438124 1006052 438176 1006058
rect 438124 1005994 438176 1006000
rect 435548 1004828 435600 1004834
rect 435548 1004770 435600 1004776
rect 435364 1002108 435416 1002114
rect 435364 1002050 435416 1002056
rect 433984 994832 434036 994838
rect 433984 994774 434036 994780
rect 420644 994696 420696 994702
rect 420644 994638 420696 994644
rect 393964 994628 394016 994634
rect 393964 994570 394016 994576
rect 392676 994492 392728 994498
rect 392676 994434 392728 994440
rect 381176 994288 381228 994294
rect 381176 994230 381228 994236
rect 369124 990140 369176 990146
rect 369124 990082 369176 990088
rect 381188 983634 381216 994230
rect 429936 992928 429988 992934
rect 429936 992870 429988 992876
rect 397828 991500 397880 991506
rect 397828 991442 397880 991448
rect 364996 983606 365470 983634
rect 381188 983606 381662 983634
rect 397840 983620 397868 991442
rect 414112 990140 414164 990146
rect 414112 990082 414164 990088
rect 414124 983620 414152 990082
rect 429948 983634 429976 992870
rect 435376 991506 435404 1002050
rect 435560 992934 435588 1004770
rect 436744 1001972 436796 1001978
rect 436744 1001914 436796 1001920
rect 435548 992928 435600 992934
rect 435548 992870 435600 992876
rect 435364 991500 435416 991506
rect 435364 991442 435416 991448
rect 436756 985998 436784 1001914
rect 438136 997762 438164 1005994
rect 446036 1004080 446088 1004086
rect 446036 1004022 446088 1004028
rect 438124 997756 438176 997762
rect 438124 997698 438176 997704
rect 439872 997756 439924 997762
rect 439872 997698 439924 997704
rect 439688 997620 439740 997626
rect 439688 997562 439740 997568
rect 439700 996985 439728 997562
rect 439686 996976 439742 996985
rect 439686 996911 439742 996920
rect 439884 996441 439912 997698
rect 446048 997286 446076 1004022
rect 447140 1001224 447192 1001230
rect 447140 1001166 447192 1001172
rect 447152 1000074 447180 1001166
rect 447796 1000822 447824 1006402
rect 469864 1006324 469916 1006330
rect 469864 1006266 469916 1006272
rect 452568 1005712 452620 1005718
rect 452568 1005654 452620 1005660
rect 452580 1003950 452608 1005654
rect 458824 1005576 458876 1005582
rect 458824 1005518 458876 1005524
rect 449900 1003944 449952 1003950
rect 449900 1003886 449952 1003892
rect 452568 1003944 452620 1003950
rect 452568 1003886 452620 1003892
rect 449912 1001162 449940 1003886
rect 449900 1001156 449952 1001162
rect 449900 1001098 449952 1001104
rect 453764 1001156 453816 1001162
rect 453764 1001098 453816 1001104
rect 447784 1000816 447836 1000822
rect 447784 1000758 447836 1000764
rect 449900 1000816 449952 1000822
rect 449900 1000758 449952 1000764
rect 447140 1000068 447192 1000074
rect 447140 1000010 447192 1000016
rect 449912 998850 449940 1000758
rect 450084 1000068 450136 1000074
rect 450084 1000010 450136 1000016
rect 449900 998844 449952 998850
rect 449900 998786 449952 998792
rect 446036 997280 446088 997286
rect 446036 997222 446088 997228
rect 450096 997218 450124 1000010
rect 450084 997212 450136 997218
rect 450084 997154 450136 997160
rect 446128 997144 446180 997150
rect 446128 997086 446180 997092
rect 439870 996432 439926 996441
rect 439870 996367 439926 996376
rect 436744 985992 436796 985998
rect 436744 985934 436796 985940
rect 446140 983634 446168 997086
rect 453776 995858 453804 1001098
rect 453764 995852 453816 995858
rect 453764 995794 453816 995800
rect 458836 994537 458864 1005518
rect 465724 1005440 465776 1005446
rect 465724 1005382 465776 1005388
rect 460940 1003944 460992 1003950
rect 460940 1003886 460992 1003892
rect 460952 995625 460980 1003886
rect 462964 1002720 463016 1002726
rect 462964 1002662 463016 1002668
rect 460938 995616 460994 995625
rect 460938 995551 460994 995560
rect 462976 994566 463004 1002662
rect 462964 994560 463016 994566
rect 458822 994528 458878 994537
rect 462964 994502 463016 994508
rect 458822 994463 458878 994472
rect 465736 994430 465764 1005382
rect 467104 1005304 467156 1005310
rect 467104 1005246 467156 1005252
rect 467116 998209 467144 1005246
rect 468484 1002584 468536 1002590
rect 468484 1002526 468536 1002532
rect 467102 998200 467158 998209
rect 467102 998135 467158 998144
rect 465724 994424 465776 994430
rect 465724 994366 465776 994372
rect 468496 993993 468524 1002526
rect 469220 997076 469272 997082
rect 469220 997018 469272 997024
rect 469232 994809 469260 997018
rect 469876 995081 469904 1006266
rect 507030 1006224 507086 1006233
rect 507030 1006159 507032 1006168
rect 507084 1006159 507086 1006168
rect 507032 1006130 507084 1006136
rect 498842 1006088 498898 1006097
rect 471244 1006052 471296 1006058
rect 471244 1005994 471296 1006000
rect 496728 1006052 496780 1006058
rect 498842 1006023 498844 1006032
rect 496728 1005994 496780 1006000
rect 498896 1006023 498898 1006032
rect 502522 1006088 502578 1006097
rect 509054 1006088 509110 1006097
rect 502522 1006023 502524 1006032
rect 498844 1005994 498896 1006000
rect 502576 1006023 502578 1006032
rect 505744 1006052 505796 1006058
rect 502524 1005994 502576 1006000
rect 509054 1006023 509056 1006032
rect 505744 1005994 505796 1006000
rect 509108 1006023 509110 1006032
rect 509056 1005994 509108 1006000
rect 471256 996033 471284 1005994
rect 496544 1001972 496596 1001978
rect 496544 1001914 496596 1001920
rect 496556 1001230 496584 1001914
rect 496544 1001224 496596 1001230
rect 496544 1001166 496596 1001172
rect 496740 999138 496768 1005994
rect 505008 1005712 505060 1005718
rect 505006 1005680 505008 1005689
rect 505060 1005680 505062 1005689
rect 505006 1005615 505062 1005624
rect 502156 1005440 502208 1005446
rect 502154 1005408 502156 1005417
rect 502208 1005408 502210 1005417
rect 502154 1005343 502210 1005352
rect 499672 1005304 499724 1005310
rect 499670 1005272 499672 1005281
rect 499724 1005272 499726 1005281
rect 499670 1005207 499726 1005216
rect 500498 1005136 500554 1005145
rect 500498 1005071 500500 1005080
rect 500552 1005071 500554 1005080
rect 500500 1005042 500552 1005048
rect 500498 1004864 500554 1004873
rect 498108 1004828 498160 1004834
rect 500498 1004799 500500 1004808
rect 498108 1004770 498160 1004776
rect 500552 1004799 500554 1004808
rect 500500 1004770 500552 1004776
rect 496740 999110 496860 999138
rect 472624 998844 472676 998850
rect 472624 998786 472676 998792
rect 472440 998708 472492 998714
rect 472440 998650 472492 998656
rect 472256 998572 472308 998578
rect 472256 998514 472308 998520
rect 472072 998436 472124 998442
rect 472072 998378 472124 998384
rect 471888 997212 471940 997218
rect 471888 997154 471940 997160
rect 471242 996024 471298 996033
rect 471242 995959 471298 995968
rect 469862 995072 469918 995081
rect 469862 995007 469918 995016
rect 469218 994800 469274 994809
rect 469218 994735 469274 994744
rect 471900 994265 471928 997154
rect 472084 995330 472112 998378
rect 472268 996713 472296 998514
rect 472254 996704 472310 996713
rect 472254 996639 472310 996648
rect 472452 995761 472480 998650
rect 472438 995752 472494 995761
rect 472438 995687 472494 995696
rect 472636 995586 472664 998786
rect 489000 997756 489052 997762
rect 489000 997698 489052 997704
rect 489012 996985 489040 997698
rect 488998 996976 489054 996985
rect 488998 996911 489054 996920
rect 494058 996432 494114 996441
rect 494058 996367 494114 996376
rect 488908 995920 488960 995926
rect 488908 995862 488960 995868
rect 488920 995761 488948 995862
rect 474002 995752 474058 995761
rect 474738 995752 474794 995761
rect 474058 995710 474306 995738
rect 474002 995687 474058 995696
rect 477038 995752 477094 995761
rect 474794 995710 474950 995738
rect 474738 995687 474794 995696
rect 481454 995752 481510 995761
rect 477094 995710 477342 995738
rect 477038 995687 477094 995696
rect 482742 995752 482798 995761
rect 481510 995710 481666 995738
rect 481454 995687 481510 995696
rect 485594 995752 485650 995761
rect 482798 995710 482954 995738
rect 485346 995710 485594 995738
rect 482742 995687 482798 995696
rect 487986 995752 488042 995761
rect 487830 995710 487986 995738
rect 485594 995687 485650 995696
rect 487986 995687 488042 995696
rect 488906 995752 488962 995761
rect 488906 995687 488962 995696
rect 473372 995586 473662 995602
rect 472624 995580 472676 995586
rect 472624 995522 472676 995528
rect 473360 995580 473662 995586
rect 473412 995574 473662 995580
rect 473360 995522 473412 995528
rect 473820 995512 473872 995518
rect 478236 995512 478288 995518
rect 473820 995454 473872 995460
rect 477682 995480 477738 995489
rect 473832 995330 473860 995454
rect 472084 995302 473860 995330
rect 474648 994560 474700 994566
rect 474648 994502 474700 994508
rect 474660 994294 474688 994502
rect 474648 994288 474700 994294
rect 471886 994256 471942 994265
rect 476776 994265 476804 995452
rect 477738 995438 477986 995466
rect 478288 995460 478630 995466
rect 478236 995454 478630 995460
rect 478248 995438 478630 995454
rect 477682 995415 477738 995424
rect 474648 994230 474700 994236
rect 476762 994256 476818 994265
rect 471886 994191 471942 994200
rect 476762 994191 476818 994200
rect 481100 993993 481128 995452
rect 482296 994809 482324 995452
rect 484136 995110 484164 995452
rect 484124 995104 484176 995110
rect 484124 995046 484176 995052
rect 482282 994800 482338 994809
rect 482282 994735 482338 994744
rect 485976 994566 486004 995452
rect 485964 994560 486016 994566
rect 485964 994502 486016 994508
rect 486620 994430 486648 995452
rect 486608 994424 486660 994430
rect 486608 994366 486660 994372
rect 494072 994294 494100 996367
rect 496832 995586 496860 999110
rect 498120 997626 498148 1004770
rect 501326 1004728 501382 1004737
rect 499488 1004692 499540 1004698
rect 501326 1004663 501328 1004672
rect 499488 1004634 499540 1004640
rect 501380 1004663 501382 1004672
rect 501328 1004634 501380 1004640
rect 498474 1002008 498530 1002017
rect 498474 1001943 498476 1001952
rect 498528 1001943 498530 1001952
rect 498476 1001914 498528 1001920
rect 499500 1001366 499528 1004634
rect 504548 1003944 504600 1003950
rect 504546 1003912 504548 1003921
rect 504600 1003912 504602 1003921
rect 504546 1003847 504602 1003856
rect 503350 1002416 503406 1002425
rect 500868 1002380 500920 1002386
rect 503350 1002351 503352 1002360
rect 500868 1002322 500920 1002328
rect 503404 1002351 503406 1002360
rect 503352 1002322 503404 1002328
rect 499488 1001360 499540 1001366
rect 499488 1001302 499540 1001308
rect 498108 997620 498160 997626
rect 498108 997562 498160 997568
rect 500880 997082 500908 1002322
rect 504178 1002280 504234 1002289
rect 502248 1002244 502300 1002250
rect 504178 1002215 504180 1002224
rect 502248 1002186 502300 1002192
rect 504232 1002215 504234 1002224
rect 504180 1002186 504232 1002192
rect 501694 1002008 501750 1002017
rect 501694 1001943 501696 1001952
rect 501748 1001943 501750 1001952
rect 501696 1001914 501748 1001920
rect 502260 998578 502288 1002186
rect 502522 1002144 502578 1002153
rect 502522 1002079 502524 1002088
rect 502576 1002079 502578 1002088
rect 503720 1002108 503772 1002114
rect 502524 1002050 502576 1002056
rect 503720 1002050 503772 1002056
rect 503350 1002008 503406 1002017
rect 502984 1001972 503036 1001978
rect 503350 1001943 503352 1001952
rect 502984 1001914 503036 1001920
rect 503404 1001943 503406 1001952
rect 503352 1001914 503404 1001920
rect 502248 998572 502300 998578
rect 502248 998514 502300 998520
rect 500868 997076 500920 997082
rect 500868 997018 500920 997024
rect 502062 995616 502118 995625
rect 496820 995580 496872 995586
rect 502062 995551 502118 995560
rect 496820 995522 496872 995528
rect 502076 995081 502104 995551
rect 502062 995072 502118 995081
rect 502062 995007 502118 995016
rect 502996 994430 503024 1001914
rect 503732 998442 503760 1002050
rect 504364 1001972 504416 1001978
rect 504364 1001914 504416 1001920
rect 503720 998436 503772 998442
rect 503720 998378 503772 998384
rect 504376 997490 504404 1001914
rect 504364 997484 504416 997490
rect 504364 997426 504416 997432
rect 505756 995110 505784 1005994
rect 508504 1005100 508556 1005106
rect 508504 1005042 508556 1005048
rect 507858 1004864 507914 1004873
rect 507858 1004799 507860 1004808
rect 507912 1004799 507914 1004808
rect 507860 1004770 507912 1004776
rect 507398 1004728 507454 1004737
rect 507398 1004663 507400 1004672
rect 507452 1004663 507454 1004672
rect 507400 1004634 507452 1004640
rect 506202 1002008 506258 1002017
rect 506258 1001966 506520 1001994
rect 506202 1001943 506258 1001952
rect 506492 997762 506520 1001966
rect 506480 997756 506532 997762
rect 506480 997698 506532 997704
rect 505744 995104 505796 995110
rect 505744 995046 505796 995052
rect 508516 994566 508544 1005042
rect 509700 1004828 509752 1004834
rect 509700 1004770 509752 1004776
rect 509240 1004692 509292 1004698
rect 509240 1004634 509292 1004640
rect 509252 994838 509280 1004634
rect 509712 997762 509740 1004770
rect 513852 1003406 513880 1007082
rect 518164 1006936 518216 1006942
rect 554780 1006936 554832 1006942
rect 518164 1006878 518216 1006884
rect 554778 1006904 554780 1006913
rect 569224 1006936 569276 1006942
rect 554832 1006904 554834 1006913
rect 514024 1005984 514076 1005990
rect 514024 1005926 514076 1005932
rect 513840 1003400 513892 1003406
rect 513840 1003342 513892 1003348
rect 509882 1002144 509938 1002153
rect 509882 1002079 509884 1002088
rect 509936 1002079 509938 1002088
rect 512828 1002108 512880 1002114
rect 509884 1002050 509936 1002056
rect 512828 1002050 512880 1002056
rect 510342 1002008 510398 1002017
rect 510342 1001943 510344 1001952
rect 510396 1001943 510398 1001952
rect 512644 1001972 512696 1001978
rect 510344 1001914 510396 1001920
rect 512644 1001914 512696 1001920
rect 509700 997756 509752 997762
rect 509700 997698 509752 997704
rect 509240 994832 509292 994838
rect 509240 994774 509292 994780
rect 508504 994560 508556 994566
rect 508504 994502 508556 994508
rect 502984 994424 503036 994430
rect 502984 994366 503036 994372
rect 494060 994288 494112 994294
rect 494060 994230 494112 994236
rect 511080 994288 511132 994294
rect 511080 994230 511132 994236
rect 468482 993984 468538 993993
rect 468482 993919 468538 993928
rect 481086 993984 481142 993993
rect 481086 993919 481142 993928
rect 494704 992928 494756 992934
rect 494704 992870 494756 992876
rect 478972 991500 479024 991506
rect 478972 991442 479024 991448
rect 462780 985992 462832 985998
rect 462780 985934 462832 985940
rect 429948 983606 430330 983634
rect 446140 983606 446522 983634
rect 462792 983620 462820 985934
rect 478984 983620 479012 991442
rect 494716 983634 494744 992870
rect 511092 983634 511120 994230
rect 512656 991506 512684 1001914
rect 512840 992934 512868 1002050
rect 512828 992928 512880 992934
rect 512828 992870 512880 992876
rect 512644 991500 512696 991506
rect 512644 991442 512696 991448
rect 514036 985998 514064 1005926
rect 515404 1005712 515456 1005718
rect 515404 1005654 515456 1005660
rect 515416 998850 515444 1005654
rect 516784 1005304 516836 1005310
rect 516784 1005246 516836 1005252
rect 516796 1001894 516824 1005246
rect 516336 1001866 516824 1001894
rect 515404 998844 515456 998850
rect 515404 998786 515456 998792
rect 516336 993682 516364 1001866
rect 516968 1001360 517020 1001366
rect 516968 1001302 517020 1001308
rect 516980 998730 517008 1001302
rect 517152 998844 517204 998850
rect 517152 998786 517204 998792
rect 516980 998702 517100 998730
rect 516508 998572 516560 998578
rect 516508 998514 516560 998520
rect 516520 995330 516548 998514
rect 516876 997620 516928 997626
rect 516876 997562 516928 997568
rect 516692 997484 516744 997490
rect 516692 997426 516744 997432
rect 516704 996713 516732 997426
rect 516690 996704 516746 996713
rect 516690 996639 516746 996648
rect 516888 996441 516916 997562
rect 516874 996432 516930 996441
rect 516874 996367 516930 996376
rect 517072 996282 517100 998702
rect 516980 996254 517100 996282
rect 516980 995625 517008 996254
rect 517164 995897 517192 998786
rect 517336 997756 517388 997762
rect 517336 997698 517388 997704
rect 517348 996985 517376 997698
rect 517334 996976 517390 996985
rect 517334 996911 517390 996920
rect 517150 995888 517206 995897
rect 517150 995823 517206 995832
rect 516966 995616 517022 995625
rect 516966 995551 517022 995560
rect 516690 995344 516746 995353
rect 516520 995302 516690 995330
rect 516690 995279 516746 995288
rect 518176 994294 518204 1006878
rect 569224 1006878 569276 1006884
rect 554778 1006839 554834 1006848
rect 555976 1006800 556028 1006806
rect 555974 1006768 555976 1006777
rect 565820 1006800 565872 1006806
rect 556028 1006768 556030 1006777
rect 520924 1006732 520976 1006738
rect 565820 1006742 565872 1006748
rect 555974 1006703 556030 1006712
rect 520924 1006674 520976 1006680
rect 519544 1005440 519596 1005446
rect 519544 1005382 519596 1005388
rect 518900 1003400 518952 1003406
rect 518900 1003342 518952 1003348
rect 518912 996169 518940 1003342
rect 518898 996160 518954 996169
rect 518898 996095 518954 996104
rect 518164 994288 518216 994294
rect 518164 994230 518216 994236
rect 519556 994158 519584 1005382
rect 520280 1003944 520332 1003950
rect 520280 1003886 520332 1003892
rect 520292 997830 520320 1003886
rect 520280 997824 520332 997830
rect 520280 997766 520332 997772
rect 520188 995580 520240 995586
rect 520188 995522 520240 995528
rect 520200 994809 520228 995522
rect 520936 995081 520964 1006674
rect 559654 1006496 559710 1006505
rect 556988 1006460 557040 1006466
rect 559654 1006431 559656 1006440
rect 556988 1006402 557040 1006408
rect 559708 1006431 559710 1006440
rect 559656 1006402 559708 1006408
rect 522304 1006324 522356 1006330
rect 522304 1006266 522356 1006272
rect 522316 996130 522344 1006266
rect 556802 1006224 556858 1006233
rect 556802 1006159 556804 1006168
rect 556856 1006159 556858 1006168
rect 556804 1006130 556856 1006136
rect 551098 1006088 551154 1006097
rect 523684 1006052 523736 1006058
rect 551098 1006023 551154 1006032
rect 555146 1006088 555202 1006097
rect 555146 1006023 555148 1006032
rect 523684 1005994 523736 1006000
rect 522764 1001224 522816 1001230
rect 522764 1001166 522816 1001172
rect 522304 996124 522356 996130
rect 522304 996066 522356 996072
rect 520922 995072 520978 995081
rect 520922 995007 520978 995016
rect 520186 994800 520242 994809
rect 520186 994735 520242 994744
rect 519544 994152 519596 994158
rect 519544 994094 519596 994100
rect 522776 993818 522804 1001166
rect 522948 997076 523000 997082
rect 522948 997018 523000 997024
rect 522960 994022 522988 997018
rect 523696 995858 523724 1005994
rect 551112 1004086 551140 1006023
rect 555200 1006023 555202 1006032
rect 556436 1006052 556488 1006058
rect 555148 1005994 555200 1006000
rect 556436 1005994 556488 1006000
rect 556448 1005582 556476 1005994
rect 556436 1005576 556488 1005582
rect 556436 1005518 556488 1005524
rect 553124 1005440 553176 1005446
rect 553122 1005408 553124 1005417
rect 553176 1005408 553178 1005417
rect 553122 1005343 553178 1005352
rect 551468 1005304 551520 1005310
rect 551466 1005272 551468 1005281
rect 551520 1005272 551522 1005281
rect 551466 1005207 551522 1005216
rect 555974 1004864 556030 1004873
rect 555974 1004799 555976 1004808
rect 556028 1004799 556030 1004808
rect 555976 1004770 556028 1004776
rect 551100 1004080 551152 1004086
rect 551100 1004022 551152 1004028
rect 552296 1003944 552348 1003950
rect 552294 1003912 552296 1003921
rect 552348 1003912 552350 1003921
rect 552294 1003847 552350 1003856
rect 553950 1002280 554006 1002289
rect 553308 1002244 553360 1002250
rect 553950 1002215 553952 1002224
rect 553308 1002186 553360 1002192
rect 554004 1002215 554006 1002224
rect 553952 1002186 554004 1002192
rect 550272 1001224 550324 1001230
rect 550270 1001192 550272 1001201
rect 550324 1001192 550326 1001201
rect 550270 1001127 550326 1001136
rect 552294 998472 552350 998481
rect 524052 998436 524104 998442
rect 552294 998407 552296 998416
rect 524052 998378 524104 998384
rect 552348 998407 552350 998416
rect 552296 998378 552348 998384
rect 523868 997824 523920 997830
rect 523868 997766 523920 997772
rect 523684 995852 523736 995858
rect 523684 995794 523736 995800
rect 523880 994838 523908 997766
rect 524064 997257 524092 998378
rect 551466 998064 551522 998073
rect 549168 998028 549220 998034
rect 551466 997999 551468 998008
rect 549168 997970 549220 997976
rect 551520 997999 551522 998008
rect 551468 997970 551520 997976
rect 540888 997756 540940 997762
rect 540888 997698 540940 997704
rect 524050 997248 524106 997257
rect 524050 997183 524106 997192
rect 540900 996985 540928 997698
rect 540886 996976 540942 996985
rect 540886 996911 540942 996920
rect 524050 996704 524106 996713
rect 524050 996639 524106 996648
rect 524064 995586 524092 996639
rect 524786 995752 524842 995761
rect 532146 995752 532202 995761
rect 524842 995710 525090 995738
rect 524786 995687 524842 995696
rect 532790 995752 532846 995761
rect 532202 995710 532542 995738
rect 532146 995687 532202 995696
rect 535918 995752 535974 995761
rect 532846 995710 533094 995738
rect 535578 995710 535918 995738
rect 532790 995687 532846 995696
rect 535918 995687 535974 995696
rect 538218 995752 538274 995761
rect 538218 995687 538274 995696
rect 525352 995586 525734 995602
rect 524052 995580 524104 995586
rect 524052 995522 524104 995528
rect 525340 995580 525734 995586
rect 525392 995574 525734 995580
rect 525340 995522 525392 995528
rect 529572 995512 529624 995518
rect 523868 994832 523920 994838
rect 526364 994809 526392 995452
rect 527928 995438 528218 995466
rect 529414 995460 529572 995466
rect 530216 995512 530268 995518
rect 529414 995454 529624 995460
rect 529846 995480 529902 995489
rect 527928 994838 527956 995438
rect 528756 995110 528784 995452
rect 529414 995438 529612 995454
rect 530214 995480 530216 995489
rect 530268 995480 530270 995489
rect 529902 995438 530058 995466
rect 529846 995415 529902 995424
rect 530214 995415 530270 995424
rect 528744 995104 528796 995110
rect 528744 995046 528796 995052
rect 527916 994832 527968 994838
rect 523868 994774 523920 994780
rect 526350 994800 526406 994809
rect 527916 994774 527968 994780
rect 529020 994832 529072 994838
rect 529020 994774 529072 994780
rect 526350 994735 526406 994744
rect 529032 994158 529060 994774
rect 533724 994430 533752 995452
rect 534368 994566 534396 995452
rect 536760 994809 536788 995452
rect 537418 995438 537800 995466
rect 537772 995178 537800 995438
rect 537760 995172 537812 995178
rect 537760 995114 537812 995120
rect 536746 994800 536802 994809
rect 536746 994735 536802 994744
rect 534356 994560 534408 994566
rect 538048 994537 538076 995452
rect 538232 994838 538260 995687
rect 538404 995172 538456 995178
rect 538404 995114 538456 995120
rect 538220 994832 538272 994838
rect 538220 994774 538272 994780
rect 534356 994502 534408 994508
rect 538034 994528 538090 994537
rect 538034 994463 538090 994472
rect 533712 994424 533764 994430
rect 533712 994366 533764 994372
rect 529388 994288 529440 994294
rect 529388 994230 529440 994236
rect 529020 994152 529072 994158
rect 529020 994094 529072 994100
rect 529400 994022 529428 994230
rect 538416 994158 538444 995114
rect 539244 994294 539272 995452
rect 539232 994288 539284 994294
rect 539232 994230 539284 994236
rect 538404 994152 538456 994158
rect 538404 994094 538456 994100
rect 522948 994016 523000 994022
rect 522948 993958 523000 993964
rect 529388 994016 529440 994022
rect 529388 993958 529440 993964
rect 522764 993812 522816 993818
rect 522764 993754 522816 993760
rect 516324 993676 516376 993682
rect 516324 993618 516376 993624
rect 549180 993546 549208 997970
rect 553122 997928 553178 997937
rect 551560 997892 551612 997898
rect 553122 997863 553124 997872
rect 551560 997834 551612 997840
rect 553176 997863 553178 997872
rect 553124 997834 553176 997840
rect 551572 997354 551600 997834
rect 553320 997558 553348 1002186
rect 553950 1002008 554006 1002017
rect 553412 1001966 553950 1001994
rect 553412 1001894 553440 1001966
rect 553950 1001943 554006 1001952
rect 554778 1002008 554834 1002017
rect 554778 1001943 554834 1001952
rect 553412 1001866 553532 1001894
rect 553308 997552 553360 997558
rect 553308 997494 553360 997500
rect 551560 997348 551612 997354
rect 551560 997290 551612 997296
rect 553504 997218 553532 1001866
rect 553492 997212 553544 997218
rect 553492 997154 553544 997160
rect 549168 993540 549220 993546
rect 549168 993482 549220 993488
rect 554792 993410 554820 1001943
rect 557000 997762 557028 1006402
rect 557170 1006088 557226 1006097
rect 557170 1006023 557172 1006032
rect 557224 1006023 557226 1006032
rect 557172 1005994 557224 1006000
rect 558184 1004828 558236 1004834
rect 558184 1004770 558236 1004776
rect 557630 1004728 557686 1004737
rect 557630 1004663 557632 1004672
rect 557684 1004663 557686 1004672
rect 557632 1004634 557684 1004640
rect 557998 1002416 558054 1002425
rect 557998 1002351 558000 1002360
rect 558052 1002351 558054 1002360
rect 558000 1002322 558052 1002328
rect 556988 997756 557040 997762
rect 556988 997698 557040 997704
rect 558196 995994 558224 1004770
rect 560850 1004728 560906 1004737
rect 559564 1004692 559616 1004698
rect 560850 1004663 560852 1004672
rect 559564 1004634 559616 1004640
rect 560904 1004663 560906 1004672
rect 560852 1004634 560904 1004640
rect 558826 1002688 558882 1002697
rect 558826 1002623 558828 1002632
rect 558880 1002623 558882 1002632
rect 558828 1002594 558880 1002600
rect 558826 1002008 558882 1002017
rect 558826 1001943 558828 1001952
rect 558880 1001943 558882 1001952
rect 558828 1001914 558880 1001920
rect 558184 995988 558236 995994
rect 558184 995930 558236 995936
rect 554780 993404 554832 993410
rect 554780 993346 554832 993352
rect 527272 992928 527324 992934
rect 527272 992870 527324 992876
rect 514024 985992 514076 985998
rect 514024 985934 514076 985940
rect 527284 983634 527312 992870
rect 559576 991506 559604 1004634
rect 564440 1004080 564492 1004086
rect 564440 1004022 564492 1004028
rect 562508 1002652 562560 1002658
rect 562508 1002594 562560 1002600
rect 560850 1002552 560906 1002561
rect 560850 1002487 560852 1002496
rect 560904 1002487 560906 1002496
rect 560852 1002458 560904 1002464
rect 560944 1002380 560996 1002386
rect 560944 1002322 560996 1002328
rect 560482 1002280 560538 1002289
rect 560482 1002215 560484 1002224
rect 560536 1002215 560538 1002224
rect 560484 1002186 560536 1002192
rect 560022 1002144 560078 1002153
rect 560022 1002079 560024 1002088
rect 560076 1002079 560078 1002088
rect 560024 1002050 560076 1002056
rect 560300 1001972 560352 1001978
rect 560300 1001914 560352 1001920
rect 560312 995858 560340 1001914
rect 560300 995852 560352 995858
rect 560300 995794 560352 995800
rect 543832 991500 543884 991506
rect 543832 991442 543884 991448
rect 559564 991500 559616 991506
rect 559564 991442 559616 991448
rect 494716 983606 495190 983634
rect 511092 983606 511474 983634
rect 527284 983606 527666 983634
rect 543844 983620 543872 991442
rect 560956 990146 560984 1002322
rect 562324 1002108 562376 1002114
rect 562324 1002050 562376 1002056
rect 561678 1002008 561734 1002017
rect 561678 1001943 561680 1001952
rect 561732 1001943 561734 1001952
rect 561680 1001914 561732 1001920
rect 562336 990282 562364 1002050
rect 562520 992934 562548 1002594
rect 563060 1002244 563112 1002250
rect 563060 1002186 563112 1002192
rect 563072 996130 563100 1002186
rect 563704 1001972 563756 1001978
rect 563704 1001914 563756 1001920
rect 563060 996124 563112 996130
rect 563060 996066 563112 996072
rect 563716 993070 563744 1001914
rect 564452 999122 564480 1004022
rect 565832 1003678 565860 1006742
rect 567844 1006188 567896 1006194
rect 567844 1006130 567896 1006136
rect 566464 1004692 566516 1004698
rect 566464 1004634 566516 1004640
rect 565820 1003672 565872 1003678
rect 565820 1003614 565872 1003620
rect 565084 1002516 565136 1002522
rect 565084 1002458 565136 1002464
rect 564440 999116 564492 999122
rect 564440 999058 564492 999064
rect 563704 993064 563756 993070
rect 563704 993006 563756 993012
rect 562508 992928 562560 992934
rect 562508 992870 562560 992876
rect 562324 990276 562376 990282
rect 562324 990218 562376 990224
rect 560944 990140 560996 990146
rect 560944 990082 560996 990088
rect 565096 985998 565124 1002458
rect 566476 986134 566504 1004634
rect 567384 1003944 567436 1003950
rect 567384 1003886 567436 1003892
rect 567396 997082 567424 1003886
rect 567856 1001894 567884 1006130
rect 568580 1003672 568632 1003678
rect 568580 1003614 568632 1003620
rect 567764 1001866 567884 1001894
rect 567568 997348 567620 997354
rect 567568 997290 567620 997296
rect 567384 997076 567436 997082
rect 567384 997018 567436 997024
rect 567580 995110 567608 997290
rect 567568 995104 567620 995110
rect 567568 995046 567620 995052
rect 567764 994566 567792 1001866
rect 567936 999116 567988 999122
rect 567936 999058 567988 999064
rect 567948 994838 567976 999058
rect 568592 997422 568620 1003614
rect 568580 997416 568632 997422
rect 568580 997358 568632 997364
rect 569236 996946 569264 1006878
rect 571984 1006052 572036 1006058
rect 571984 1005994 572036 1006000
rect 570604 1005440 570656 1005446
rect 570604 1005382 570656 1005388
rect 570144 997212 570196 997218
rect 570144 997154 570196 997160
rect 569224 996940 569276 996946
rect 569224 996882 569276 996888
rect 567936 994832 567988 994838
rect 567936 994774 567988 994780
rect 567752 994560 567804 994566
rect 567752 994502 567804 994508
rect 570156 994430 570184 997154
rect 570616 996130 570644 1005382
rect 570788 998436 570840 998442
rect 570788 998378 570840 998384
rect 570604 996124 570656 996130
rect 570604 996066 570656 996072
rect 570800 994809 570828 998378
rect 571996 997694 572024 1005994
rect 573364 1005576 573416 1005582
rect 573364 1005518 573416 1005524
rect 571984 997688 572036 997694
rect 571984 997630 572036 997636
rect 573376 997218 573404 1005518
rect 574744 1005304 574796 1005310
rect 574744 1005246 574796 1005252
rect 574100 1001224 574152 1001230
rect 574100 1001166 574152 1001172
rect 573364 997212 573416 997218
rect 573364 997154 573416 997160
rect 570786 994800 570842 994809
rect 570786 994735 570842 994744
rect 570144 994424 570196 994430
rect 570144 994366 570196 994372
rect 574112 994090 574140 1001166
rect 574100 994084 574152 994090
rect 574100 994026 574152 994032
rect 574756 993954 574784 1005246
rect 618168 999184 618220 999190
rect 618168 999126 618220 999132
rect 625528 999184 625580 999190
rect 625528 999126 625580 999132
rect 590568 997688 590620 997694
rect 590568 997630 590620 997636
rect 590384 997416 590436 997422
rect 590384 997358 590436 997364
rect 590396 996690 590424 997358
rect 590580 997098 590608 997630
rect 618180 997354 618208 999126
rect 591304 997348 591356 997354
rect 591304 997290 591356 997296
rect 618168 997348 618220 997354
rect 618168 997290 618220 997296
rect 590580 997070 590792 997098
rect 590566 996976 590622 996985
rect 590566 996911 590568 996920
rect 590620 996911 590622 996920
rect 590568 996882 590620 996888
rect 590566 996704 590622 996713
rect 590396 996662 590566 996690
rect 590566 996639 590622 996648
rect 590764 996441 590792 997070
rect 590750 996432 590806 996441
rect 590750 996367 590806 996376
rect 590566 995072 590622 995081
rect 590566 995007 590622 995016
rect 590580 994702 590608 995007
rect 590568 994696 590620 994702
rect 590568 994638 590620 994644
rect 591316 994430 591344 997290
rect 622400 997212 622452 997218
rect 622400 997154 622452 997160
rect 620284 997076 620336 997082
rect 620284 997018 620336 997024
rect 620296 995489 620324 997018
rect 622412 996033 622440 997154
rect 622398 996024 622454 996033
rect 622398 995959 622454 995968
rect 620282 995480 620338 995489
rect 620282 995415 620338 995424
rect 625540 994430 625568 999126
rect 625712 997824 625764 997830
rect 625712 997766 625764 997772
rect 625724 994838 625752 997766
rect 625896 995988 625948 995994
rect 625896 995930 625948 995936
rect 625908 995518 625936 995930
rect 642088 995920 642140 995926
rect 642088 995862 642140 995868
rect 642100 995761 642128 995862
rect 626630 995752 626686 995761
rect 627182 995752 627238 995761
rect 626686 995710 626888 995738
rect 626630 995687 626686 995696
rect 627918 995752 627974 995761
rect 627238 995710 627532 995738
rect 627182 995687 627238 995696
rect 633990 995752 634046 995761
rect 627974 995710 628176 995738
rect 627918 995687 627974 995696
rect 635830 995752 635886 995761
rect 634046 995710 634340 995738
rect 635536 995710 635830 995738
rect 633990 995687 634046 995696
rect 635830 995687 635886 995696
rect 642086 995752 642142 995761
rect 642086 995687 642142 995696
rect 625896 995512 625948 995518
rect 625896 995454 625948 995460
rect 629668 995512 629720 995518
rect 631506 995480 631562 995489
rect 629720 995460 630016 995466
rect 629668 995454 630016 995460
rect 629680 995438 630016 995454
rect 630232 995438 630568 995466
rect 630876 995438 631212 995466
rect 625712 994832 625764 994838
rect 625712 994774 625764 994780
rect 630232 994430 630260 995438
rect 630876 994838 630904 995438
rect 631562 995438 631856 995466
rect 634556 995438 634892 995466
rect 635844 995438 636180 995466
rect 637040 995438 637376 995466
rect 638572 995438 638908 995466
rect 631506 995415 631562 995424
rect 630864 994832 630916 994838
rect 634556 994809 634584 995438
rect 630864 994774 630916 994780
rect 634542 994800 634598 994809
rect 634542 994735 634598 994744
rect 591304 994424 591356 994430
rect 591304 994366 591356 994372
rect 625528 994424 625580 994430
rect 625528 994366 625580 994372
rect 630220 994424 630272 994430
rect 630220 994366 630272 994372
rect 574744 993948 574796 993954
rect 574744 993890 574796 993896
rect 635844 993546 635872 995438
rect 637040 995110 637068 995438
rect 637028 995104 637080 995110
rect 637028 995046 637080 995052
rect 635832 993540 635884 993546
rect 635832 993482 635884 993488
rect 608600 993064 608652 993070
rect 608600 993006 608652 993012
rect 576306 990992 576362 991001
rect 576306 990927 576362 990936
rect 566464 986128 566516 986134
rect 566464 986070 566516 986076
rect 560116 985992 560168 985998
rect 560116 985934 560168 985940
rect 565084 985992 565136 985998
rect 565084 985934 565136 985940
rect 560128 983620 560156 985934
rect 576320 983620 576348 990927
rect 592500 986128 592552 986134
rect 592500 986070 592552 986076
rect 592512 983620 592540 986070
rect 608612 983634 608640 993006
rect 638880 992322 638908 995438
rect 639064 995438 639216 995466
rect 639524 995438 639860 995466
rect 640720 995438 641056 995466
rect 639064 994566 639092 995438
rect 639524 994702 639552 995438
rect 639512 994696 639564 994702
rect 639512 994638 639564 994644
rect 639052 994560 639104 994566
rect 639052 994502 639104 994508
rect 640720 993410 640748 995438
rect 660578 995072 660634 995081
rect 660578 995007 660580 995016
rect 660632 995007 660634 995016
rect 660580 994977 660632 994983
rect 660764 994628 660816 994634
rect 660764 994570 660816 994576
rect 660776 993818 660804 994570
rect 660948 994560 661000 994566
rect 660948 994502 661000 994508
rect 660764 993812 660816 993818
rect 660764 993754 660816 993760
rect 660960 993682 660988 994502
rect 660948 993676 661000 993682
rect 660948 993618 661000 993624
rect 640708 993404 640760 993410
rect 640708 993346 640760 993352
rect 667204 992928 667256 992934
rect 667204 992870 667256 992876
rect 638868 992316 638920 992322
rect 638868 992258 638920 992264
rect 640800 992316 640852 992322
rect 640800 992258 640852 992264
rect 624976 985992 625028 985998
rect 624976 985934 625028 985940
rect 608612 983606 608810 983634
rect 624988 983620 625016 985934
rect 640812 983634 640840 992258
rect 658924 991500 658976 991506
rect 658924 991442 658976 991448
rect 640812 983606 641194 983634
rect 62118 976032 62174 976041
rect 62118 975967 62174 975976
rect 62132 975730 62160 975967
rect 651654 975896 651710 975905
rect 651654 975831 651710 975840
rect 651668 975730 651696 975831
rect 62120 975724 62172 975730
rect 62120 975666 62172 975672
rect 651656 975724 651708 975730
rect 651656 975666 651708 975672
rect 62118 962976 62174 962985
rect 62118 962911 62174 962920
rect 62132 961926 62160 962911
rect 651470 962568 651526 962577
rect 651470 962503 651526 962512
rect 651484 961926 651512 962503
rect 62120 961920 62172 961926
rect 62120 961862 62172 961868
rect 651472 961920 651524 961926
rect 651472 961862 651524 961868
rect 62118 949920 62174 949929
rect 62118 949855 62174 949864
rect 62132 946014 62160 949855
rect 652206 949376 652262 949385
rect 652206 949311 652262 949320
rect 652220 948122 652248 949311
rect 652208 948116 652260 948122
rect 652208 948058 652260 948064
rect 62120 946008 62172 946014
rect 62120 945950 62172 945956
rect 651472 937032 651524 937038
rect 651472 936974 651524 936980
rect 651484 936193 651512 936974
rect 651470 936184 651526 936193
rect 651470 936119 651526 936128
rect 658936 936057 658964 991442
rect 665824 961920 665876 961926
rect 665824 961862 665876 961868
rect 661682 957808 661738 957817
rect 661682 957743 661738 957752
rect 660304 948116 660356 948122
rect 660304 948058 660356 948064
rect 660316 941769 660344 948058
rect 660302 941760 660358 941769
rect 660302 941695 660358 941704
rect 661696 937038 661724 957743
rect 665836 939865 665864 961862
rect 665822 939856 665878 939865
rect 665822 939791 665878 939800
rect 667216 937145 667244 992870
rect 669964 990276 670016 990282
rect 669964 990218 670016 990224
rect 668584 990140 668636 990146
rect 668584 990082 668636 990088
rect 668596 937689 668624 990082
rect 669976 938505 670004 990218
rect 672724 975724 672776 975730
rect 672724 975666 672776 975672
rect 672538 952232 672594 952241
rect 672538 952167 672594 952176
rect 669962 938496 670018 938505
rect 669962 938431 670018 938440
rect 668582 937680 668638 937689
rect 668582 937615 668638 937624
rect 667202 937136 667258 937145
rect 667202 937071 667258 937080
rect 661684 937032 661736 937038
rect 661684 936974 661736 936980
rect 670974 936456 671030 936465
rect 670974 936391 671030 936400
rect 658922 936048 658978 936057
rect 658922 935983 658978 935992
rect 669226 929520 669282 929529
rect 669226 929455 669282 929464
rect 62118 923808 62174 923817
rect 62118 923743 62174 923752
rect 62132 923302 62160 923743
rect 62120 923296 62172 923302
rect 62120 923238 62172 923244
rect 651470 922720 651526 922729
rect 651470 922655 651526 922664
rect 651484 921874 651512 922655
rect 651472 921868 651524 921874
rect 651472 921810 651524 921816
rect 663064 921868 663116 921874
rect 663064 921810 663116 921816
rect 62118 910752 62174 910761
rect 62118 910687 62174 910696
rect 62132 909498 62160 910687
rect 652390 909528 652446 909537
rect 62120 909492 62172 909498
rect 652390 909463 652392 909472
rect 62120 909434 62172 909440
rect 652444 909463 652446 909472
rect 652392 909434 652444 909440
rect 62118 897832 62174 897841
rect 62118 897767 62174 897776
rect 62132 897054 62160 897767
rect 62120 897048 62172 897054
rect 62120 896990 62172 896996
rect 651470 896200 651526 896209
rect 651470 896135 651526 896144
rect 651484 895694 651512 896135
rect 651472 895688 651524 895694
rect 651472 895630 651524 895636
rect 55862 892800 55918 892809
rect 55862 892735 55918 892744
rect 54482 892528 54538 892537
rect 54482 892463 54538 892472
rect 53286 892256 53342 892265
rect 53286 892191 53342 892200
rect 651654 882872 651710 882881
rect 651654 882807 651710 882816
rect 651668 881890 651696 882807
rect 651656 881884 651708 881890
rect 651656 881826 651708 881832
rect 62118 871720 62174 871729
rect 62118 871655 62174 871664
rect 62132 870874 62160 871655
rect 62120 870868 62172 870874
rect 62120 870810 62172 870816
rect 651470 869680 651526 869689
rect 651470 869615 651526 869624
rect 651484 869446 651512 869615
rect 651472 869440 651524 869446
rect 651472 869382 651524 869388
rect 658924 869440 658976 869446
rect 658924 869382 658976 869388
rect 62118 858664 62174 858673
rect 62118 858599 62174 858608
rect 62132 858430 62160 858599
rect 62120 858424 62172 858430
rect 62120 858366 62172 858372
rect 651470 856352 651526 856361
rect 651470 856287 651526 856296
rect 651484 852174 651512 856287
rect 651472 852168 651524 852174
rect 651472 852110 651524 852116
rect 62118 845608 62174 845617
rect 62118 845543 62174 845552
rect 62132 844626 62160 845543
rect 54484 844620 54536 844626
rect 54484 844562 54536 844568
rect 62120 844620 62172 844626
rect 62120 844562 62172 844568
rect 53102 799096 53158 799105
rect 53102 799031 53158 799040
rect 54496 774353 54524 844562
rect 651838 843024 651894 843033
rect 651838 842959 651894 842968
rect 651852 841838 651880 842959
rect 651840 841832 651892 841838
rect 651840 841774 651892 841780
rect 62762 832552 62818 832561
rect 62762 832487 62818 832496
rect 62118 819496 62174 819505
rect 62118 819431 62174 819440
rect 62132 818378 62160 819431
rect 62120 818372 62172 818378
rect 62120 818314 62172 818320
rect 62118 806576 62174 806585
rect 62118 806511 62174 806520
rect 62132 806002 62160 806511
rect 62120 805996 62172 806002
rect 62120 805938 62172 805944
rect 62118 793656 62174 793665
rect 55864 793620 55916 793626
rect 62118 793591 62120 793600
rect 55864 793562 55916 793568
rect 62172 793591 62174 793600
rect 62120 793562 62172 793568
rect 54482 774344 54538 774353
rect 54482 774279 54538 774288
rect 51722 773528 51778 773537
rect 51722 773463 51778 773472
rect 51724 753568 51776 753574
rect 51724 753510 51776 753516
rect 50342 730552 50398 730561
rect 50342 730487 50398 730496
rect 50344 714876 50396 714882
rect 50344 714818 50396 714824
rect 48962 669352 49018 669361
rect 48962 669287 49018 669296
rect 47584 662448 47636 662454
rect 47584 662390 47636 662396
rect 47306 637936 47362 637945
rect 47306 637871 47362 637880
rect 47122 637664 47178 637673
rect 47122 637599 47178 637608
rect 47136 618633 47164 637599
rect 47122 618624 47178 618633
rect 47122 618559 47178 618568
rect 47320 615641 47348 637871
rect 47306 615632 47362 615641
rect 47306 615567 47362 615576
rect 46940 612740 46992 612746
rect 46940 612682 46992 612688
rect 46110 598088 46166 598097
rect 46110 598023 46166 598032
rect 47596 582457 47624 662390
rect 47766 636984 47822 636993
rect 47766 636919 47822 636928
rect 47780 618361 47808 636919
rect 50356 626657 50384 714818
rect 51736 691393 51764 753510
rect 54484 741124 54536 741130
rect 54484 741066 54536 741072
rect 51722 691384 51778 691393
rect 51722 691319 51778 691328
rect 53104 688696 53156 688702
rect 53104 688638 53156 688644
rect 51724 674892 51776 674898
rect 51724 674834 51776 674840
rect 51736 646649 51764 674834
rect 51722 646640 51778 646649
rect 51722 646575 51778 646584
rect 53116 644745 53144 688638
rect 54496 688129 54524 741066
rect 55876 730153 55904 793562
rect 62776 788633 62804 832487
rect 651470 829832 651526 829841
rect 651470 829767 651526 829776
rect 651484 829462 651512 829767
rect 651472 829456 651524 829462
rect 651472 829398 651524 829404
rect 651470 816504 651526 816513
rect 651470 816439 651526 816448
rect 651484 815658 651512 816439
rect 651472 815652 651524 815658
rect 651472 815594 651524 815600
rect 651470 803312 651526 803321
rect 651470 803247 651472 803256
rect 651524 803247 651526 803256
rect 651472 803218 651524 803224
rect 651470 789984 651526 789993
rect 651470 789919 651526 789928
rect 651484 789410 651512 789919
rect 651472 789404 651524 789410
rect 651472 789346 651524 789352
rect 62762 788624 62818 788633
rect 62762 788559 62818 788568
rect 62762 780464 62818 780473
rect 62762 780399 62818 780408
rect 62118 767408 62174 767417
rect 62118 767343 62120 767352
rect 62172 767343 62174 767352
rect 62120 767314 62172 767320
rect 62118 754352 62174 754361
rect 62118 754287 62174 754296
rect 62132 753574 62160 754287
rect 62120 753568 62172 753574
rect 62120 753510 62172 753516
rect 62776 743073 62804 780399
rect 652390 776656 652446 776665
rect 652390 776591 652446 776600
rect 652404 775606 652432 776591
rect 652392 775600 652444 775606
rect 652392 775542 652444 775548
rect 651470 763328 651526 763337
rect 651470 763263 651472 763272
rect 651524 763263 651526 763272
rect 651472 763234 651524 763240
rect 651470 750136 651526 750145
rect 651470 750071 651526 750080
rect 651484 749426 651512 750071
rect 651472 749420 651524 749426
rect 651472 749362 651524 749368
rect 62762 743064 62818 743073
rect 62762 742999 62818 743008
rect 62118 741296 62174 741305
rect 62118 741231 62174 741240
rect 62132 741130 62160 741231
rect 62120 741124 62172 741130
rect 62120 741066 62172 741072
rect 651838 736808 651894 736817
rect 651838 736743 651894 736752
rect 651852 735622 651880 736743
rect 651840 735616 651892 735622
rect 651840 735558 651892 735564
rect 55862 730144 55918 730153
rect 55862 730079 55918 730088
rect 62762 728240 62818 728249
rect 62762 728175 62818 728184
rect 62118 715320 62174 715329
rect 62118 715255 62174 715264
rect 62132 714882 62160 715255
rect 62120 714876 62172 714882
rect 62120 714818 62172 714824
rect 62118 702264 62174 702273
rect 62118 702199 62174 702208
rect 62132 701078 62160 702199
rect 55864 701072 55916 701078
rect 55864 701014 55916 701020
rect 62120 701072 62172 701078
rect 62120 701014 62172 701020
rect 54482 688120 54538 688129
rect 54482 688055 54538 688064
rect 54484 647896 54536 647902
rect 54484 647838 54536 647844
rect 53102 644736 53158 644745
rect 53102 644671 53158 644680
rect 51724 636268 51776 636274
rect 51724 636210 51776 636216
rect 50342 626648 50398 626657
rect 50342 626583 50398 626592
rect 48964 623824 49016 623830
rect 48964 623766 49016 623772
rect 47766 618352 47822 618361
rect 47766 618287 47822 618296
rect 48976 601361 49004 623766
rect 51736 601769 51764 636210
rect 51722 601760 51778 601769
rect 51722 601695 51778 601704
rect 48962 601352 49018 601361
rect 48962 601287 49018 601296
rect 54496 600953 54524 647838
rect 55876 643249 55904 701014
rect 62776 689489 62804 728175
rect 651470 723480 651526 723489
rect 651470 723415 651526 723424
rect 651484 723178 651512 723415
rect 651472 723172 651524 723178
rect 651472 723114 651524 723120
rect 658936 716009 658964 869382
rect 660304 829456 660356 829462
rect 660304 829398 660356 829404
rect 660316 778977 660344 829398
rect 661684 815652 661736 815658
rect 661684 815594 661736 815600
rect 660302 778968 660358 778977
rect 660302 778903 660358 778912
rect 660304 763224 660356 763230
rect 660304 763166 660356 763172
rect 658922 716000 658978 716009
rect 658922 715935 658978 715944
rect 652574 710288 652630 710297
rect 652574 710223 652630 710232
rect 652588 709374 652616 710223
rect 652576 709368 652628 709374
rect 652576 709310 652628 709316
rect 652392 696992 652444 696998
rect 652390 696960 652392 696969
rect 652444 696960 652446 696969
rect 652390 696895 652446 696904
rect 62762 689480 62818 689489
rect 62762 689415 62818 689424
rect 62118 689208 62174 689217
rect 62118 689143 62174 689152
rect 62132 688702 62160 689143
rect 62120 688696 62172 688702
rect 62120 688638 62172 688644
rect 651838 683632 651894 683641
rect 651838 683567 651894 683576
rect 651852 683194 651880 683567
rect 651840 683188 651892 683194
rect 651840 683130 651892 683136
rect 658924 683188 658976 683194
rect 658924 683130 658976 683136
rect 62118 676152 62174 676161
rect 62118 676087 62174 676096
rect 62132 674898 62160 676087
rect 62120 674892 62172 674898
rect 62120 674834 62172 674840
rect 652390 670440 652446 670449
rect 652390 670375 652446 670384
rect 652404 669390 652432 670375
rect 652392 669384 652444 669390
rect 652392 669326 652444 669332
rect 62118 663096 62174 663105
rect 62118 663031 62174 663040
rect 62132 662454 62160 663031
rect 62120 662448 62172 662454
rect 62120 662390 62172 662396
rect 651654 657112 651710 657121
rect 651654 657047 651710 657056
rect 651668 656946 651696 657047
rect 651656 656940 651708 656946
rect 651656 656882 651708 656888
rect 62118 650040 62174 650049
rect 62118 649975 62174 649984
rect 62132 647902 62160 649975
rect 62120 647896 62172 647902
rect 62120 647838 62172 647844
rect 651470 643784 651526 643793
rect 651470 643719 651526 643728
rect 55862 643240 55918 643249
rect 55862 643175 55918 643184
rect 651484 643142 651512 643719
rect 651472 643136 651524 643142
rect 651472 643078 651524 643084
rect 62118 637120 62174 637129
rect 62118 637055 62174 637064
rect 62132 636274 62160 637055
rect 62120 636268 62172 636274
rect 62120 636210 62172 636216
rect 651562 630592 651618 630601
rect 651562 630527 651618 630536
rect 651576 628590 651604 630527
rect 651564 628584 651616 628590
rect 651564 628526 651616 628532
rect 62118 624064 62174 624073
rect 62118 623999 62174 624008
rect 62132 623830 62160 623999
rect 62120 623824 62172 623830
rect 62120 623766 62172 623772
rect 651470 617264 651526 617273
rect 651470 617199 651526 617208
rect 651484 616894 651512 617199
rect 651472 616888 651524 616894
rect 651472 616830 651524 616836
rect 62118 611008 62174 611017
rect 62118 610943 62174 610952
rect 62132 608666 62160 610943
rect 56048 608660 56100 608666
rect 56048 608602 56100 608608
rect 62120 608660 62172 608666
rect 62120 608602 62172 608608
rect 54482 600944 54538 600953
rect 54482 600879 54538 600888
rect 48964 597576 49016 597582
rect 48964 597518 49016 597524
rect 47582 582448 47638 582457
rect 47582 582383 47638 582392
rect 48976 557841 49004 597518
rect 50344 583772 50396 583778
rect 50344 583714 50396 583720
rect 48962 557832 49018 557841
rect 48962 557767 49018 557776
rect 50356 557569 50384 583714
rect 55864 558136 55916 558142
rect 55864 558078 55916 558084
rect 50342 557560 50398 557569
rect 50342 557495 50398 557504
rect 45650 556880 45706 556889
rect 45650 556815 45706 556824
rect 45006 555656 45062 555665
rect 45006 555591 45062 555600
rect 44638 555248 44694 555257
rect 44638 555183 44694 555192
rect 44270 554432 44326 554441
rect 44270 554367 44326 554376
rect 43810 548176 43866 548185
rect 43810 548111 43866 548120
rect 43824 355337 43852 548111
rect 43994 547088 44050 547097
rect 43994 547023 44050 547032
rect 44008 355722 44036 547023
rect 44284 427281 44312 554367
rect 44454 552392 44510 552401
rect 44454 552327 44510 552336
rect 44468 534313 44496 552327
rect 44454 534304 44510 534313
rect 44454 534239 44510 534248
rect 44652 428097 44680 555183
rect 44914 551168 44970 551177
rect 44914 551103 44970 551112
rect 44928 549386 44956 551103
rect 45098 549536 45154 549545
rect 45098 549471 45154 549480
rect 44928 549358 45048 549386
rect 44822 548720 44878 548729
rect 44822 548655 44878 548664
rect 44836 536897 44864 548655
rect 44822 536888 44878 536897
rect 44822 536823 44878 536832
rect 45020 532681 45048 549358
rect 45112 547874 45140 549471
rect 45282 549128 45338 549137
rect 45282 549063 45338 549072
rect 45112 547846 45232 547874
rect 45204 534074 45232 547846
rect 45296 543734 45324 549063
rect 45296 543706 45416 543734
rect 45388 537441 45416 543706
rect 45374 537432 45430 537441
rect 45374 537367 45430 537376
rect 45204 534046 45324 534074
rect 45296 533361 45324 534046
rect 45282 533352 45338 533361
rect 45282 533287 45338 533296
rect 45006 532672 45062 532681
rect 45006 532607 45062 532616
rect 45664 429729 45692 556815
rect 46018 556064 46074 556073
rect 46018 555999 46074 556008
rect 45650 429720 45706 429729
rect 45650 429655 45706 429664
rect 45834 429312 45890 429321
rect 45834 429247 45890 429256
rect 45650 428496 45706 428505
rect 45650 428431 45706 428440
rect 44638 428088 44694 428097
rect 44638 428023 44694 428032
rect 44730 427680 44786 427689
rect 44730 427615 44786 427624
rect 44270 427272 44326 427281
rect 44270 427207 44326 427216
rect 44270 426864 44326 426873
rect 44270 426799 44326 426808
rect 44284 384033 44312 426799
rect 44454 423192 44510 423201
rect 44454 423127 44510 423136
rect 44468 402937 44496 423127
rect 44454 402928 44510 402937
rect 44454 402863 44510 402872
rect 44744 384849 44772 427615
rect 45098 423600 45154 423609
rect 45098 423535 45154 423544
rect 44914 422376 44970 422385
rect 44914 422311 44970 422320
rect 44928 405657 44956 422311
rect 44914 405648 44970 405657
rect 44914 405583 44970 405592
rect 45112 402529 45140 423535
rect 45466 421560 45522 421569
rect 45466 421495 45522 421504
rect 45282 421152 45338 421161
rect 45282 421087 45338 421096
rect 45296 407833 45324 421087
rect 45282 407824 45338 407833
rect 45282 407759 45338 407768
rect 45480 406745 45508 421495
rect 45466 406736 45522 406745
rect 45466 406671 45522 406680
rect 45098 402520 45154 402529
rect 45098 402455 45154 402464
rect 45282 386064 45338 386073
rect 45282 385999 45338 386008
rect 45098 385248 45154 385257
rect 45098 385183 45154 385192
rect 44730 384840 44786 384849
rect 44730 384775 44786 384784
rect 44270 384024 44326 384033
rect 44270 383959 44326 383968
rect 44546 379944 44602 379953
rect 44546 379879 44602 379888
rect 44178 377496 44234 377505
rect 44178 377431 44234 377440
rect 44192 356697 44220 377431
rect 44362 376272 44418 376281
rect 44362 376207 44418 376216
rect 44376 360194 44404 376207
rect 44560 360194 44588 379879
rect 44914 379536 44970 379545
rect 44914 379471 44970 379480
rect 44730 379128 44786 379137
rect 44730 379063 44786 379072
rect 44744 369854 44772 379063
rect 44928 369854 44956 379471
rect 45112 369854 45140 385183
rect 45296 379514 45324 385999
rect 45664 385665 45692 428431
rect 45848 387297 45876 429247
rect 46032 428913 46060 555999
rect 47584 545148 47636 545154
rect 47584 545090 47636 545096
rect 46204 506524 46256 506530
rect 46204 506466 46256 506472
rect 46018 428904 46074 428913
rect 46018 428839 46074 428848
rect 45834 387288 45890 387297
rect 45834 387223 45890 387232
rect 45650 385656 45706 385665
rect 45650 385591 45706 385600
rect 45834 384432 45890 384441
rect 45834 384367 45890 384376
rect 45650 383616 45706 383625
rect 45650 383551 45706 383560
rect 45296 379486 45508 379514
rect 44652 369826 44772 369854
rect 44836 369826 44956 369854
rect 45020 369826 45140 369854
rect 44652 364290 44680 369826
rect 44836 365809 44864 369826
rect 44822 365800 44878 365809
rect 44822 365735 44878 365744
rect 44822 364304 44878 364313
rect 44652 364262 44822 364290
rect 44822 364239 44878 364248
rect 44376 360166 44496 360194
rect 44560 360166 44680 360194
rect 44178 356688 44234 356697
rect 44178 356623 44234 356632
rect 44468 356289 44496 360166
rect 44652 359961 44680 360166
rect 44638 359952 44694 359961
rect 44638 359887 44694 359896
rect 44454 356280 44510 356289
rect 44454 356215 44510 356224
rect 44008 355694 44312 355722
rect 43810 355328 43866 355337
rect 43810 355263 43866 355272
rect 44284 355008 44312 355694
rect 44638 355600 44694 355609
rect 44638 355535 44694 355544
rect 44652 355026 44680 355535
rect 44822 355328 44878 355337
rect 44822 355263 44878 355272
rect 44640 355020 44692 355026
rect 44284 354980 44496 355008
rect 44468 354634 44496 354980
rect 44640 354962 44692 354968
rect 44468 354606 44726 354634
rect 44836 354618 44864 355263
rect 44575 354544 44627 354550
rect 44468 354504 44575 354532
rect 44468 354362 44496 354504
rect 44575 354486 44627 354492
rect 43640 354334 44496 354362
rect 44698 354362 44726 354606
rect 44824 354612 44876 354618
rect 44824 354554 44876 354560
rect 44811 354482 44956 354498
rect 44799 354476 44956 354482
rect 44851 354470 44956 354476
rect 44799 354418 44851 354424
rect 44698 354346 44839 354362
rect 44698 354340 44851 354346
rect 44698 354334 44799 354340
rect 44799 354282 44851 354288
rect 44928 354226 44956 354470
rect 43548 354198 44956 354226
rect 43258 353696 43314 353705
rect 43258 353631 43314 353640
rect 28538 351248 28594 351257
rect 28538 351183 28594 351192
rect 8588 345100 8616 345236
rect 9048 345100 9076 345236
rect 9508 345100 9536 345236
rect 9968 345100 9996 345236
rect 10428 345100 10456 345236
rect 10888 345100 10916 345236
rect 11348 345100 11376 345236
rect 11808 345100 11836 345236
rect 12268 345100 12296 345236
rect 12728 345100 12756 345236
rect 13188 345100 13216 345236
rect 13648 345100 13676 345236
rect 14108 345100 14136 345236
rect 28552 343913 28580 351183
rect 45020 350534 45048 369826
rect 45190 356688 45246 356697
rect 45246 356646 45416 356674
rect 45190 356623 45246 356632
rect 45190 356280 45246 356289
rect 45190 356215 45246 356224
rect 45204 353870 45232 356215
rect 45192 353864 45244 353870
rect 45192 353806 45244 353812
rect 45146 353728 45198 353734
rect 45144 353696 45146 353705
rect 45198 353696 45200 353705
rect 45144 353631 45200 353640
rect 45388 353546 45416 356646
rect 45371 353518 45416 353546
rect 45371 353326 45399 353518
rect 45359 353320 45411 353326
rect 45359 353262 45411 353268
rect 44836 350506 45048 350534
rect 40222 345536 40278 345545
rect 40222 345471 40278 345480
rect 28538 343904 28594 343913
rect 28538 343839 28594 343848
rect 35806 343904 35862 343913
rect 35806 343839 35862 343848
rect 35820 343670 35848 343839
rect 40236 343670 40264 345471
rect 35808 343664 35860 343670
rect 35808 343606 35860 343612
rect 40224 343664 40276 343670
rect 40224 343606 40276 343612
rect 44836 342553 44864 350506
rect 45480 343369 45508 379486
rect 45466 343360 45522 343369
rect 45466 343295 45522 343304
rect 44822 342544 44878 342553
rect 44822 342479 44878 342488
rect 45466 341320 45522 341329
rect 45466 341255 45522 341264
rect 35806 339824 35862 339833
rect 35806 339759 35862 339768
rect 35820 339522 35848 339759
rect 35808 339516 35860 339522
rect 35808 339458 35860 339464
rect 37556 339516 37608 339522
rect 37556 339458 37608 339464
rect 35162 339008 35218 339017
rect 35162 338943 35218 338952
rect 33782 338192 33838 338201
rect 33782 338127 33838 338136
rect 33796 327729 33824 338127
rect 35176 329089 35204 338943
rect 37568 336569 37596 339458
rect 37554 336560 37610 336569
rect 37554 336495 37610 336504
rect 42798 334656 42854 334665
rect 42798 334591 42854 334600
rect 43166 334656 43222 334665
rect 43166 334591 43222 334600
rect 44178 334656 44234 334665
rect 44178 334591 44234 334600
rect 44362 334656 44418 334665
rect 44362 334591 44418 334600
rect 35162 329080 35218 329089
rect 35162 329015 35218 329024
rect 33782 327720 33838 327729
rect 33782 327655 33838 327664
rect 42168 326210 42196 326264
rect 42168 326182 42288 326210
rect 41786 325408 41842 325417
rect 41786 325343 41842 325352
rect 41800 325040 41828 325343
rect 41878 324728 41934 324737
rect 41878 324663 41934 324672
rect 41892 324428 41920 324663
rect 42260 324329 42288 326182
rect 42246 324320 42302 324329
rect 42246 324255 42302 324264
rect 42182 323734 42472 323762
rect 42246 323640 42302 323649
rect 42246 323575 42302 323584
rect 42062 322824 42118 322833
rect 42062 322759 42118 322768
rect 42076 322592 42104 322759
rect 42260 321382 42288 323575
rect 42444 321473 42472 323734
rect 42430 321464 42486 321473
rect 42430 321399 42486 321408
rect 42182 321354 42288 321382
rect 42430 321192 42486 321201
rect 42430 321127 42486 321136
rect 42444 320739 42472 321127
rect 42182 320711 42472 320739
rect 42430 320104 42486 320113
rect 42182 320062 42430 320090
rect 42430 320039 42486 320048
rect 41786 319968 41842 319977
rect 41786 319903 41842 319912
rect 41800 319532 41828 319903
rect 42812 318794 42840 334591
rect 42982 334384 43038 334393
rect 42982 334319 43038 334328
rect 42996 323649 43024 334319
rect 42982 323640 43038 323649
rect 42982 323575 43038 323584
rect 43180 322833 43208 334591
rect 43626 322960 43682 322969
rect 43626 322895 43682 322904
rect 43166 322824 43222 322833
rect 43166 322759 43222 322768
rect 42812 318766 43024 318794
rect 42996 317098 43024 318766
rect 42536 317070 43024 317098
rect 42536 317059 42564 317070
rect 42182 317031 42564 317059
rect 41786 316840 41842 316849
rect 41786 316775 41842 316784
rect 41800 316404 41828 316775
rect 42154 316024 42210 316033
rect 42154 315959 42210 315968
rect 42168 315757 42196 315959
rect 41786 315616 41842 315625
rect 41786 315551 41842 315560
rect 41800 315180 41828 315551
rect 42154 313712 42210 313721
rect 42154 313647 42210 313656
rect 42168 313344 42196 313647
rect 42430 312760 42486 312769
rect 42182 312718 42430 312746
rect 42430 312695 42486 312704
rect 41970 312624 42026 312633
rect 41970 312559 42026 312568
rect 41984 312052 42012 312559
rect 41786 303104 41842 303113
rect 41786 303039 41842 303048
rect 8588 301988 8616 302124
rect 9048 301988 9076 302124
rect 9508 301988 9536 302124
rect 9968 301988 9996 302124
rect 10428 301988 10456 302124
rect 10888 301988 10916 302124
rect 11348 301988 11376 302124
rect 11808 301988 11836 302124
rect 12268 301988 12296 302124
rect 12728 301988 12756 302124
rect 13188 301988 13216 302124
rect 13648 301988 13676 302124
rect 14108 301988 14136 302124
rect 41800 300937 41828 303039
rect 41786 300928 41842 300937
rect 41786 300863 41842 300872
rect 42798 297256 42854 297265
rect 42798 297191 42854 297200
rect 41786 296848 41842 296857
rect 41786 296783 41842 296792
rect 41326 296032 41382 296041
rect 41326 295967 41382 295976
rect 39302 294808 39358 294817
rect 39302 294743 39358 294752
rect 39316 284782 39344 294743
rect 41340 292074 41368 295967
rect 41800 292913 41828 296783
rect 41786 292904 41842 292913
rect 41786 292839 41842 292848
rect 41786 292224 41842 292233
rect 41524 292182 41786 292210
rect 41524 292074 41552 292182
rect 41786 292159 41842 292168
rect 41340 292046 41552 292074
rect 41326 290320 41382 290329
rect 41326 290255 41382 290264
rect 41340 284986 41368 290255
rect 41328 284980 41380 284986
rect 41328 284922 41380 284928
rect 41696 284980 41748 284986
rect 41748 284940 42380 284968
rect 41696 284922 41748 284928
rect 39304 284776 39356 284782
rect 39304 284718 39356 284724
rect 41696 284776 41748 284782
rect 41748 284724 42288 284730
rect 41696 284718 42288 284724
rect 41708 284702 42288 284718
rect 42260 283059 42288 284702
rect 42182 283031 42288 283059
rect 42352 281874 42380 284940
rect 42182 281846 42380 281874
rect 41970 281480 42026 281489
rect 41970 281415 42026 281424
rect 41984 281180 42012 281415
rect 42182 280554 42472 280582
rect 42154 279848 42210 279857
rect 42154 279783 42210 279792
rect 42168 279344 42196 279783
rect 42444 278769 42472 280554
rect 42430 278760 42486 278769
rect 42430 278695 42486 278704
rect 42430 278216 42486 278225
rect 42168 278066 42196 278188
rect 42260 278174 42430 278202
rect 42260 278066 42288 278174
rect 42430 278151 42486 278160
rect 42168 278038 42288 278066
rect 41786 277944 41842 277953
rect 41786 277879 41842 277888
rect 41800 277508 41828 277879
rect 42246 277672 42302 277681
rect 42246 277607 42302 277616
rect 42062 277128 42118 277137
rect 42062 277063 42118 277072
rect 42076 276896 42104 277063
rect 42062 276720 42118 276729
rect 42062 276655 42118 276664
rect 42076 276352 42104 276655
rect 41786 274272 41842 274281
rect 41786 274207 41842 274216
rect 41800 273836 41828 274207
rect 42076 273057 42104 273224
rect 42062 273048 42118 273057
rect 42062 272983 42118 272992
rect 42062 272776 42118 272785
rect 42062 272711 42118 272720
rect 42076 272544 42104 272711
rect 42260 272014 42288 277607
rect 42182 271986 42288 272014
rect 41786 270464 41842 270473
rect 41786 270399 41842 270408
rect 41800 270164 41828 270399
rect 42182 269507 42472 269535
rect 41786 269104 41842 269113
rect 41786 269039 41842 269048
rect 41800 268872 41828 269039
rect 42444 267753 42472 269507
rect 42430 267744 42486 267753
rect 42812 267734 42840 297191
rect 42982 295216 43038 295225
rect 42982 295151 43038 295160
rect 42996 276729 43024 295151
rect 43166 293176 43222 293185
rect 43166 293111 43222 293120
rect 43180 279857 43208 293111
rect 43442 291136 43498 291145
rect 43442 291071 43498 291080
rect 43166 279848 43222 279857
rect 43166 279783 43222 279792
rect 42982 276720 43038 276729
rect 42982 276655 43038 276664
rect 42812 267706 43024 267734
rect 42430 267679 42486 267688
rect 35806 259992 35862 260001
rect 35806 259927 35862 259936
rect 8588 258740 8616 258876
rect 9048 258740 9076 258876
rect 9508 258740 9536 258876
rect 9968 258740 9996 258876
rect 10428 258740 10456 258876
rect 10888 258740 10916 258876
rect 11348 258740 11376 258876
rect 11808 258740 11836 258876
rect 12268 258740 12296 258876
rect 12728 258740 12756 258876
rect 13188 258740 13216 258876
rect 13648 258740 13676 258876
rect 14108 258740 14136 258876
rect 35820 258369 35848 259927
rect 35806 258360 35862 258369
rect 35806 258295 35862 258304
rect 42798 254824 42854 254833
rect 42798 254759 42854 254768
rect 35622 253464 35678 253473
rect 35622 253399 35678 253408
rect 35636 252618 35664 253399
rect 35806 253056 35862 253065
rect 35806 252991 35862 253000
rect 35820 252754 35848 252991
rect 35808 252748 35860 252754
rect 35808 252690 35860 252696
rect 41696 252748 41748 252754
rect 41696 252690 41748 252696
rect 35624 252612 35676 252618
rect 35624 252554 35676 252560
rect 40684 252612 40736 252618
rect 40684 252554 40736 252560
rect 35806 252240 35862 252249
rect 35806 252175 35862 252184
rect 35820 251258 35848 252175
rect 35808 251252 35860 251258
rect 35808 251194 35860 251200
rect 37924 251252 37976 251258
rect 37924 251194 37976 251200
rect 34426 246936 34482 246945
rect 34426 246871 34482 246880
rect 34440 242214 34468 246871
rect 37936 242894 37964 251194
rect 37924 242888 37976 242894
rect 37924 242830 37976 242836
rect 34428 242208 34480 242214
rect 34428 242150 34480 242156
rect 40696 241505 40724 252554
rect 41708 248414 41736 252690
rect 41708 248386 42288 248414
rect 42260 244274 42288 248386
rect 42260 244246 42656 244274
rect 41696 242888 41748 242894
rect 41694 242856 41696 242865
rect 41748 242856 41750 242865
rect 41694 242791 41750 242800
rect 42430 242856 42486 242865
rect 42430 242791 42486 242800
rect 41696 242208 41748 242214
rect 41748 242156 42380 242162
rect 41696 242150 42380 242156
rect 41708 242134 42380 242150
rect 40682 241496 40738 241505
rect 40682 241431 40738 241440
rect 41786 240136 41842 240145
rect 41786 240071 41842 240080
rect 41800 239836 41828 240071
rect 42352 238663 42380 242134
rect 42182 238635 42380 238663
rect 42444 238105 42472 242791
rect 42430 238096 42486 238105
rect 42430 238031 42486 238040
rect 42182 237986 42288 238014
rect 42260 237946 42288 237986
rect 42628 237946 42656 244246
rect 42260 237918 42656 237946
rect 41800 235929 41828 236164
rect 41786 235920 41842 235929
rect 41786 235855 41842 235864
rect 42430 235920 42486 235929
rect 42430 235855 42486 235864
rect 42444 234983 42472 235855
rect 42182 234955 42472 234983
rect 42182 234314 42472 234342
rect 42246 234152 42302 234161
rect 42246 234087 42302 234096
rect 42260 233695 42288 234087
rect 42182 233667 42288 233695
rect 42444 233695 42472 234314
rect 42444 233667 42656 233695
rect 42168 233158 42288 233186
rect 42168 233104 42196 233158
rect 42260 233118 42288 233158
rect 42260 233090 42472 233118
rect 42444 232257 42472 233090
rect 42628 232529 42656 233667
rect 42614 232520 42670 232529
rect 42614 232455 42670 232464
rect 42430 232248 42486 232257
rect 42430 232183 42486 232192
rect 42430 231840 42486 231849
rect 42430 231775 42486 231784
rect 42444 230670 42472 231775
rect 42182 230642 42472 230670
rect 42154 230480 42210 230489
rect 42154 230415 42210 230424
rect 42168 229976 42196 230415
rect 42182 229350 42288 229378
rect 41970 228984 42026 228993
rect 41970 228919 42026 228928
rect 41984 228820 42012 228919
rect 42260 227361 42288 229350
rect 42430 227624 42486 227633
rect 42430 227559 42486 227568
rect 42246 227352 42302 227361
rect 42246 227287 42302 227296
rect 42444 226998 42472 227559
rect 42168 226930 42196 226984
rect 42260 226970 42472 226998
rect 42260 226930 42288 226970
rect 42168 226902 42288 226930
rect 42168 226358 42288 226386
rect 42168 226304 42196 226358
rect 42260 226318 42288 226358
rect 42260 226290 42656 226318
rect 42430 226128 42486 226137
rect 42430 226063 42486 226072
rect 42444 225706 42472 226063
rect 42182 225678 42472 225706
rect 42246 225584 42302 225593
rect 42246 225519 42302 225528
rect 28538 222864 28594 222873
rect 28538 222799 28594 222808
rect 8588 215492 8616 215628
rect 9048 215492 9076 215628
rect 9508 215492 9536 215628
rect 9968 215492 9996 215628
rect 10428 215492 10456 215628
rect 10888 215492 10916 215628
rect 11348 215492 11376 215628
rect 11808 215492 11836 215628
rect 12268 215492 12296 215628
rect 12728 215492 12756 215628
rect 13188 215492 13216 215628
rect 13648 215492 13676 215628
rect 14108 215492 14136 215628
rect 28552 214305 28580 222799
rect 42260 219434 42288 225519
rect 42628 224913 42656 226290
rect 42614 224904 42670 224913
rect 42614 224839 42670 224848
rect 41708 219406 42288 219434
rect 28538 214296 28594 214305
rect 28538 214231 28594 214240
rect 41326 214296 41382 214305
rect 41326 214231 41382 214240
rect 41340 213994 41368 214231
rect 41708 213994 41736 219406
rect 41328 213988 41380 213994
rect 41328 213930 41380 213936
rect 41696 213988 41748 213994
rect 41696 213930 41748 213936
rect 41142 212256 41198 212265
rect 41142 212191 41198 212200
rect 41156 211206 41184 212191
rect 42812 212129 42840 254759
rect 42996 254425 43024 267706
rect 43258 256456 43314 256465
rect 43258 256391 43314 256400
rect 43272 256306 43300 256391
rect 43272 256278 43392 256306
rect 43166 255640 43222 255649
rect 43166 255575 43222 255584
rect 42982 254416 43038 254425
rect 42982 254351 43038 254360
rect 43180 234614 43208 255575
rect 43364 234614 43392 256278
rect 42996 234586 43208 234614
rect 43272 234586 43392 234614
rect 42996 212945 43024 234586
rect 43272 213761 43300 234586
rect 43258 213752 43314 213761
rect 43258 213687 43314 213696
rect 42982 212936 43038 212945
rect 42982 212871 43038 212880
rect 42798 212120 42854 212129
rect 42798 212055 42854 212064
rect 41326 211848 41382 211857
rect 41326 211783 41382 211792
rect 41340 211342 41368 211783
rect 41328 211336 41380 211342
rect 41328 211278 41380 211284
rect 41696 211336 41748 211342
rect 41696 211278 41748 211284
rect 41144 211200 41196 211206
rect 41144 211142 41196 211148
rect 41512 211200 41564 211206
rect 41512 211142 41564 211148
rect 41326 210216 41382 210225
rect 41326 210151 41382 210160
rect 41142 209808 41198 209817
rect 41142 209743 41198 209752
rect 41156 207369 41184 209743
rect 41340 209409 41368 210151
rect 41326 209400 41382 209409
rect 41326 209335 41382 209344
rect 41326 208992 41382 209001
rect 41326 208927 41382 208936
rect 41142 207360 41198 207369
rect 41142 207295 41198 207304
rect 40958 206952 41014 206961
rect 40958 206887 41014 206896
rect 35806 204096 35862 204105
rect 35806 204031 35862 204040
rect 35820 202201 35848 204031
rect 40972 203289 41000 206887
rect 41340 204513 41368 208927
rect 41326 204504 41382 204513
rect 41326 204439 41382 204448
rect 40958 203280 41014 203289
rect 40958 203215 41014 203224
rect 35806 202192 35862 202201
rect 35806 202127 35862 202136
rect 41524 200705 41552 211142
rect 41708 208593 41736 211278
rect 41694 208584 41750 208593
rect 41694 208519 41750 208528
rect 42798 207632 42854 207641
rect 42798 207567 42854 207576
rect 41510 200696 41566 200705
rect 41510 200631 41566 200640
rect 41786 197160 41842 197169
rect 41786 197095 41842 197104
rect 41800 196656 41828 197095
rect 42154 195800 42210 195809
rect 42154 195735 42210 195744
rect 42168 195432 42196 195735
rect 41878 195256 41934 195265
rect 41878 195191 41934 195200
rect 41892 194820 41920 195191
rect 42430 193216 42486 193225
rect 42430 193151 42486 193160
rect 42444 192998 42472 193151
rect 42168 192930 42196 192984
rect 42260 192970 42472 192998
rect 42260 192930 42288 192970
rect 42168 192902 42288 192930
rect 42168 191706 42196 191760
rect 42338 191720 42394 191729
rect 42168 191678 42338 191706
rect 42338 191655 42394 191664
rect 42430 191176 42486 191185
rect 42168 191026 42196 191148
rect 42260 191134 42430 191162
rect 42260 191026 42288 191134
rect 42430 191111 42486 191120
rect 42168 190998 42288 191026
rect 42430 190496 42486 190505
rect 42182 190454 42430 190482
rect 42430 190431 42486 190440
rect 42430 189952 42486 189961
rect 42182 189910 42430 189938
rect 42430 189887 42486 189896
rect 42430 187640 42486 187649
rect 42430 187575 42486 187584
rect 42444 187459 42472 187575
rect 42182 187431 42472 187459
rect 42430 186824 42486 186833
rect 42182 186782 42430 186810
rect 42430 186759 42486 186768
rect 42812 186266 42840 207567
rect 42982 206408 43038 206417
rect 42982 206343 43038 206352
rect 42996 191185 43024 206343
rect 43258 203280 43314 203289
rect 43258 203215 43314 203224
rect 42982 191176 43038 191185
rect 42982 191111 43038 191120
rect 43272 186833 43300 203215
rect 43258 186824 43314 186833
rect 43258 186759 43314 186768
rect 42536 186238 42840 186266
rect 42536 186198 42564 186238
rect 42168 186130 42196 186184
rect 42260 186170 42564 186198
rect 42260 186130 42288 186170
rect 42168 186102 42288 186130
rect 41786 185872 41842 185881
rect 41786 185807 41842 185816
rect 41800 185605 41828 185807
rect 41786 184104 41842 184113
rect 41786 184039 41842 184048
rect 41800 183765 41828 184039
rect 42430 183152 42486 183161
rect 42182 183110 42430 183138
rect 42430 183087 42486 183096
rect 42182 182463 42472 182491
rect 42444 180713 42472 182463
rect 42430 180704 42486 180713
rect 42430 180639 42486 180648
rect 43456 51785 43484 291071
rect 43640 257689 43668 322895
rect 44192 321201 44220 334591
rect 44178 321192 44234 321201
rect 44178 321127 44234 321136
rect 44376 320113 44404 334591
rect 44362 320104 44418 320113
rect 44362 320039 44418 320048
rect 44546 311400 44602 311409
rect 44546 311335 44602 311344
rect 44362 311128 44418 311137
rect 44362 311063 44418 311072
rect 44376 300121 44404 311063
rect 44362 300112 44418 300121
rect 44362 300047 44418 300056
rect 44178 299704 44234 299713
rect 44178 299639 44234 299648
rect 43994 293584 44050 293593
rect 43994 293519 44050 293528
rect 43810 291544 43866 291553
rect 43810 291479 43866 291488
rect 43824 278225 43852 291479
rect 43810 278216 43866 278225
rect 43810 278151 43866 278160
rect 44008 273057 44036 293519
rect 43994 273048 44050 273057
rect 43994 272983 44050 272992
rect 43626 257680 43682 257689
rect 43626 257615 43682 257624
rect 44192 256873 44220 299639
rect 44560 299305 44588 311335
rect 44546 299296 44602 299305
rect 44546 299231 44602 299240
rect 45190 298888 45246 298897
rect 45190 298823 45246 298832
rect 44362 298072 44418 298081
rect 44362 298007 44418 298016
rect 44178 256864 44234 256873
rect 44178 256799 44234 256808
rect 44376 255241 44404 298007
rect 44822 294672 44878 294681
rect 44822 294607 44878 294616
rect 44638 293992 44694 294001
rect 44638 293927 44694 293936
rect 44652 273254 44680 293927
rect 44468 273226 44680 273254
rect 44468 272898 44496 273226
rect 44468 272870 44588 272898
rect 44560 272785 44588 272870
rect 44546 272776 44602 272785
rect 44546 272711 44602 272720
rect 44362 255232 44418 255241
rect 44362 255167 44418 255176
rect 44178 254008 44234 254017
rect 44178 253943 44234 253952
rect 43626 249112 43682 249121
rect 43626 249047 43682 249056
rect 43640 231849 43668 249047
rect 43810 241496 43866 241505
rect 43810 241431 43866 241440
rect 43626 231840 43682 231849
rect 43626 231775 43682 231784
rect 43824 227633 43852 241431
rect 43810 227624 43866 227633
rect 43810 227559 43866 227568
rect 44192 211313 44220 253943
rect 44362 250336 44418 250345
rect 44362 250271 44418 250280
rect 44376 230489 44404 250271
rect 44546 248704 44602 248713
rect 44546 248639 44602 248648
rect 44560 234161 44588 248639
rect 44546 234152 44602 234161
rect 44546 234087 44602 234096
rect 44362 230480 44418 230489
rect 44362 230415 44418 230424
rect 44836 214985 44864 294607
rect 45006 291816 45062 291825
rect 45006 291751 45062 291760
rect 45020 277137 45048 291751
rect 45006 277128 45062 277137
rect 45006 277063 45062 277072
rect 45204 273254 45232 298823
rect 45480 298489 45508 341255
rect 45664 340921 45692 383551
rect 45848 341737 45876 384367
rect 46216 367033 46244 506466
rect 47596 430137 47624 545090
rect 50344 532772 50396 532778
rect 50344 532714 50396 532720
rect 48964 491972 49016 491978
rect 48964 491914 49016 491920
rect 47582 430128 47638 430137
rect 47582 430063 47638 430072
rect 46938 426456 46994 426465
rect 46938 426391 46994 426400
rect 46952 399809 46980 426391
rect 46938 399800 46994 399809
rect 46938 399735 46994 399744
rect 47768 389292 47820 389298
rect 47768 389234 47820 389240
rect 46938 380760 46994 380769
rect 46938 380695 46994 380704
rect 46202 367024 46258 367033
rect 46202 366959 46258 366968
rect 46952 356017 46980 380695
rect 47122 380352 47178 380361
rect 47122 380287 47178 380296
rect 47136 357377 47164 380287
rect 47122 357368 47178 357377
rect 47122 357303 47178 357312
rect 46938 356008 46994 356017
rect 46938 355943 46994 355952
rect 46204 347064 46256 347070
rect 46204 347006 46256 347012
rect 45834 341728 45890 341737
rect 45834 341663 45890 341672
rect 45650 340912 45706 340921
rect 45650 340847 45706 340856
rect 45742 340096 45798 340105
rect 45742 340031 45798 340040
rect 45756 313721 45784 340031
rect 45926 338056 45982 338065
rect 45926 337991 45982 338000
rect 45940 324329 45968 337991
rect 45926 324320 45982 324329
rect 45926 324255 45982 324264
rect 45742 313712 45798 313721
rect 45742 313647 45798 313656
rect 45466 298480 45522 298489
rect 45466 298415 45522 298424
rect 45468 298172 45520 298178
rect 45468 298114 45520 298120
rect 45480 294681 45508 298114
rect 45466 294672 45522 294681
rect 45466 294607 45522 294616
rect 45558 294400 45614 294409
rect 45558 294335 45614 294344
rect 45112 273226 45232 273254
rect 45112 256057 45140 273226
rect 45572 267753 45600 294335
rect 45558 267744 45614 267753
rect 45558 267679 45614 267688
rect 46216 257281 46244 347006
rect 47582 333160 47638 333169
rect 47582 333095 47638 333104
rect 46202 257272 46258 257281
rect 46202 257207 46258 257216
rect 45098 256048 45154 256057
rect 45098 255983 45154 255992
rect 45558 252784 45614 252793
rect 45558 252719 45614 252728
rect 45006 248296 45062 248305
rect 45006 248231 45062 248240
rect 45020 235929 45048 248231
rect 45006 235920 45062 235929
rect 45006 235855 45062 235864
rect 45572 226137 45600 252719
rect 47030 251968 47086 251977
rect 47030 251903 47086 251912
rect 45834 251152 45890 251161
rect 45834 251087 45890 251096
rect 45558 226128 45614 226137
rect 45558 226063 45614 226072
rect 45848 224913 45876 251087
rect 46018 249520 46074 249529
rect 46018 249455 46074 249464
rect 46032 232529 46060 249455
rect 46202 247888 46258 247897
rect 46202 247823 46258 247832
rect 46018 232520 46074 232529
rect 46018 232455 46074 232464
rect 45834 224904 45890 224913
rect 45834 224839 45890 224848
rect 44822 214976 44878 214985
rect 44822 214911 44878 214920
rect 44178 211304 44234 211313
rect 44178 211239 44234 211248
rect 44178 208040 44234 208049
rect 44178 207975 44234 207984
rect 43810 205592 43866 205601
rect 43810 205527 43866 205536
rect 43626 202192 43682 202201
rect 43626 202127 43682 202136
rect 43442 51776 43498 51785
rect 43442 51711 43498 51720
rect 43640 42838 43668 202127
rect 43824 190505 43852 205527
rect 43994 205184 44050 205193
rect 43994 205119 44050 205128
rect 44008 191729 44036 205119
rect 43994 191720 44050 191729
rect 43994 191655 44050 191664
rect 43810 190496 43866 190505
rect 43810 190431 43866 190440
rect 44192 183161 44220 207975
rect 44362 206816 44418 206825
rect 44362 206751 44418 206760
rect 44376 193225 44404 206751
rect 44638 206000 44694 206009
rect 44638 205935 44694 205944
rect 44652 204626 44680 205935
rect 44822 204776 44878 204785
rect 44822 204711 44878 204720
rect 44652 204598 44772 204626
rect 44546 203960 44602 203969
rect 44546 203895 44602 203904
rect 44560 195809 44588 203895
rect 44546 195800 44602 195809
rect 44546 195735 44602 195744
rect 44362 193216 44418 193225
rect 44362 193151 44418 193160
rect 44744 190454 44772 204598
rect 44652 190426 44772 190454
rect 44652 187649 44680 190426
rect 44638 187640 44694 187649
rect 44638 187575 44694 187584
rect 44178 183152 44234 183161
rect 44178 183087 44234 183096
rect 44836 74534 44864 204711
rect 44836 74506 45508 74534
rect 45480 49162 45508 74506
rect 46216 50386 46244 247823
rect 47044 232257 47072 251903
rect 47214 250744 47270 250753
rect 47214 250679 47270 250688
rect 47030 232248 47086 232257
rect 47030 232183 47086 232192
rect 47228 227361 47256 250679
rect 47214 227352 47270 227361
rect 47214 227287 47270 227296
rect 46938 209672 46994 209681
rect 46938 209607 46994 209616
rect 46386 203552 46442 203561
rect 46386 203487 46442 203496
rect 46204 50380 46256 50386
rect 46204 50322 46256 50328
rect 45468 49156 45520 49162
rect 45468 49098 45520 49104
rect 46400 49026 46428 203487
rect 46952 180713 46980 209607
rect 47122 208856 47178 208865
rect 47122 208791 47178 208800
rect 47136 189961 47164 208791
rect 47122 189952 47178 189961
rect 47122 189887 47178 189896
rect 46938 180704 46994 180713
rect 46938 180639 46994 180648
rect 47596 51746 47624 333095
rect 47780 300529 47808 389234
rect 48976 387025 49004 491914
rect 50356 430953 50384 532714
rect 54484 518968 54536 518974
rect 54484 518910 54536 518916
rect 51724 480276 51776 480282
rect 51724 480218 51776 480224
rect 50528 440292 50580 440298
rect 50528 440234 50580 440240
rect 50342 430944 50398 430953
rect 50342 430879 50398 430888
rect 48962 387016 49018 387025
rect 48962 386951 49018 386960
rect 50344 362976 50396 362982
rect 50344 362918 50396 362924
rect 48962 334112 49018 334121
rect 48962 334047 49018 334056
rect 47766 300520 47822 300529
rect 47766 300455 47822 300464
rect 47766 247480 47822 247489
rect 47766 247415 47822 247424
rect 47584 51740 47636 51746
rect 47584 51682 47636 51688
rect 47780 50522 47808 247415
rect 47950 213344 48006 213353
rect 47950 213279 48006 213288
rect 47964 190505 47992 213279
rect 48134 210896 48190 210905
rect 48134 210831 48190 210840
rect 48148 194449 48176 210831
rect 48134 194440 48190 194449
rect 48134 194375 48190 194384
rect 47950 190496 48006 190505
rect 47950 190431 48006 190440
rect 47768 50516 47820 50522
rect 47768 50458 47820 50464
rect 48976 49298 49004 334047
rect 50356 303113 50384 362918
rect 50540 351257 50568 440234
rect 51736 386753 51764 480218
rect 51908 466472 51960 466478
rect 51908 466414 51960 466420
rect 51722 386744 51778 386753
rect 51722 386679 51778 386688
rect 51920 386481 51948 466414
rect 53104 454096 53156 454102
rect 53104 454038 53156 454044
rect 51906 386472 51962 386481
rect 51906 386407 51962 386416
rect 51908 375420 51960 375426
rect 51908 375362 51960 375368
rect 50526 351248 50582 351257
rect 50526 351183 50582 351192
rect 51724 310548 51776 310554
rect 51724 310490 51776 310496
rect 50342 303104 50398 303113
rect 50342 303039 50398 303048
rect 50342 290728 50398 290737
rect 50342 290663 50398 290672
rect 49146 289912 49202 289921
rect 49146 289847 49202 289856
rect 49160 51882 49188 289847
rect 49330 208584 49386 208593
rect 49330 208519 49386 208528
rect 49344 196489 49372 208519
rect 49514 200696 49570 200705
rect 49514 200631 49570 200640
rect 49330 196480 49386 196489
rect 49330 196415 49386 196424
rect 49528 192409 49556 200631
rect 49514 192400 49570 192409
rect 49514 192335 49570 192344
rect 50356 52018 50384 290663
rect 50526 246528 50582 246537
rect 50526 246463 50582 246472
rect 50344 52012 50396 52018
rect 50344 51954 50396 51960
rect 49148 51876 49200 51882
rect 49148 51818 49200 51824
rect 50540 50658 50568 246463
rect 51736 222873 51764 310490
rect 51920 301345 51948 375362
rect 53116 321473 53144 454038
rect 54496 430545 54524 518910
rect 54482 430536 54538 430545
rect 54482 430471 54538 430480
rect 54484 427848 54536 427854
rect 54484 427790 54536 427796
rect 54496 344321 54524 427790
rect 55876 408513 55904 558078
rect 56060 540297 56088 608602
rect 651470 603936 651526 603945
rect 651470 603871 651526 603880
rect 651484 603158 651512 603871
rect 651472 603152 651524 603158
rect 651472 603094 651524 603100
rect 62118 597952 62174 597961
rect 62118 597887 62174 597896
rect 62132 597582 62160 597887
rect 62120 597576 62172 597582
rect 62120 597518 62172 597524
rect 652390 590744 652446 590753
rect 652390 590679 652392 590688
rect 652444 590679 652446 590688
rect 652392 590650 652444 590656
rect 62118 584896 62174 584905
rect 62118 584831 62174 584840
rect 62132 583778 62160 584831
rect 62120 583772 62172 583778
rect 62120 583714 62172 583720
rect 658936 579737 658964 683130
rect 660316 625297 660344 763166
rect 661696 670721 661724 815594
rect 663076 760481 663104 921810
rect 665824 909492 665876 909498
rect 665824 909434 665876 909440
rect 664444 881884 664496 881890
rect 664444 881826 664496 881832
rect 664456 868737 664484 881826
rect 664442 868728 664498 868737
rect 664442 868663 664498 868672
rect 664444 852168 664496 852174
rect 664444 852110 664496 852116
rect 663062 760472 663118 760481
rect 663062 760407 663118 760416
rect 661868 735616 661920 735622
rect 661868 735558 661920 735564
rect 661682 670712 661738 670721
rect 661682 670647 661738 670656
rect 661880 628561 661908 735558
rect 663064 723172 663116 723178
rect 663064 723114 663116 723120
rect 663076 689353 663104 723114
rect 664456 716553 664484 852110
rect 665836 761569 665864 909434
rect 666466 879200 666522 879209
rect 666466 879135 666522 879144
rect 666282 778424 666338 778433
rect 666282 778359 666338 778368
rect 665822 761560 665878 761569
rect 665822 761495 665878 761504
rect 665824 749420 665876 749426
rect 665824 749362 665876 749368
rect 664442 716544 664498 716553
rect 664442 716479 664498 716488
rect 664444 709368 664496 709374
rect 664444 709310 664496 709316
rect 663062 689344 663118 689353
rect 663062 689279 663118 689288
rect 663064 656940 663116 656946
rect 663064 656882 663116 656888
rect 661866 628552 661922 628561
rect 661866 628487 661922 628496
rect 660302 625288 660358 625297
rect 660302 625223 660358 625232
rect 660304 616888 660356 616894
rect 660304 616830 660356 616836
rect 660316 599593 660344 616830
rect 661684 603152 661736 603158
rect 661684 603094 661736 603100
rect 660302 599584 660358 599593
rect 660302 599519 660358 599528
rect 658922 579728 658978 579737
rect 658922 579663 658978 579672
rect 651470 577416 651526 577425
rect 651470 577351 651526 577360
rect 651484 576910 651512 577351
rect 651472 576904 651524 576910
rect 651472 576846 651524 576852
rect 62118 571840 62174 571849
rect 62118 571775 62174 571784
rect 62132 569265 62160 571775
rect 62118 569256 62174 569265
rect 62118 569191 62174 569200
rect 651654 564088 651710 564097
rect 651654 564023 651710 564032
rect 651668 563106 651696 564023
rect 651656 563100 651708 563106
rect 651656 563042 651708 563048
rect 658924 563100 658976 563106
rect 658924 563042 658976 563048
rect 62118 558784 62174 558793
rect 62118 558719 62174 558728
rect 62132 558142 62160 558719
rect 62120 558136 62172 558142
rect 62120 558078 62172 558084
rect 658936 554033 658964 563042
rect 658922 554024 658978 554033
rect 658922 553959 658978 553968
rect 651470 550896 651526 550905
rect 651470 550831 651526 550840
rect 651484 550662 651512 550831
rect 651472 550656 651524 550662
rect 651472 550598 651524 550604
rect 660304 550656 660356 550662
rect 660304 550598 660356 550604
rect 62118 545864 62174 545873
rect 62118 545799 62174 545808
rect 62132 545154 62160 545799
rect 62120 545148 62172 545154
rect 62120 545090 62172 545096
rect 56046 540288 56102 540297
rect 56046 540223 56102 540232
rect 651470 537568 651526 537577
rect 651470 537503 651526 537512
rect 651484 536858 651512 537503
rect 651472 536852 651524 536858
rect 651472 536794 651524 536800
rect 62118 532808 62174 532817
rect 62118 532743 62120 532752
rect 62172 532743 62174 532752
rect 62120 532714 62172 532720
rect 651838 524240 651894 524249
rect 651838 524175 651894 524184
rect 651852 523054 651880 524175
rect 651840 523048 651892 523054
rect 651840 522990 651892 522996
rect 62118 519752 62174 519761
rect 62118 519687 62174 519696
rect 62132 518974 62160 519687
rect 62120 518968 62172 518974
rect 62120 518910 62172 518916
rect 651470 511048 651526 511057
rect 651470 510983 651526 510992
rect 651484 510678 651512 510983
rect 651472 510672 651524 510678
rect 651472 510614 651524 510620
rect 659108 510672 659160 510678
rect 659108 510614 659160 510620
rect 62118 506696 62174 506705
rect 62118 506631 62174 506640
rect 62132 506530 62160 506631
rect 62120 506524 62172 506530
rect 62120 506466 62172 506472
rect 652574 497720 652630 497729
rect 652574 497655 652630 497664
rect 652588 494766 652616 497655
rect 652576 494760 652628 494766
rect 652576 494702 652628 494708
rect 62118 493640 62174 493649
rect 62118 493575 62174 493584
rect 62132 491978 62160 493575
rect 62120 491972 62172 491978
rect 62120 491914 62172 491920
rect 651470 484528 651526 484537
rect 651470 484463 651472 484472
rect 651524 484463 651526 484472
rect 651472 484434 651524 484440
rect 62118 480584 62174 480593
rect 62118 480519 62174 480528
rect 62132 480282 62160 480519
rect 62120 480276 62172 480282
rect 62120 480218 62172 480224
rect 651470 471200 651526 471209
rect 651470 471135 651526 471144
rect 651484 470626 651512 471135
rect 651472 470620 651524 470626
rect 651472 470562 651524 470568
rect 62118 467528 62174 467537
rect 62118 467463 62174 467472
rect 62132 466478 62160 467463
rect 62120 466472 62172 466478
rect 62120 466414 62172 466420
rect 652390 457872 652446 457881
rect 652390 457807 652446 457816
rect 652404 456822 652432 457807
rect 652392 456816 652444 456822
rect 652392 456758 652444 456764
rect 62118 454608 62174 454617
rect 62118 454543 62174 454552
rect 62132 454102 62160 454543
rect 62120 454096 62172 454102
rect 62120 454038 62172 454044
rect 651470 444544 651526 444553
rect 651470 444479 651472 444488
rect 651524 444479 651526 444488
rect 651472 444450 651524 444456
rect 62118 441552 62174 441561
rect 62118 441487 62174 441496
rect 62132 440298 62160 441487
rect 62120 440292 62172 440298
rect 62120 440234 62172 440240
rect 651470 431352 651526 431361
rect 651470 431287 651526 431296
rect 651484 430642 651512 431287
rect 651472 430636 651524 430642
rect 651472 430578 651524 430584
rect 62118 428496 62174 428505
rect 62118 428431 62174 428440
rect 62132 427854 62160 428431
rect 62120 427848 62172 427854
rect 62120 427790 62172 427796
rect 651838 418024 651894 418033
rect 651838 417959 651894 417968
rect 651852 416838 651880 417959
rect 651840 416832 651892 416838
rect 651840 416774 651892 416780
rect 62762 415440 62818 415449
rect 62762 415375 62818 415384
rect 55862 408504 55918 408513
rect 55862 408439 55918 408448
rect 62118 402384 62174 402393
rect 62118 402319 62174 402328
rect 62132 401674 62160 402319
rect 55864 401668 55916 401674
rect 55864 401610 55916 401616
rect 62120 401668 62172 401674
rect 62120 401610 62172 401616
rect 54482 344312 54538 344321
rect 54482 344247 54538 344256
rect 54484 336796 54536 336802
rect 54484 336738 54536 336744
rect 53102 321464 53158 321473
rect 53102 321399 53158 321408
rect 51906 301336 51962 301345
rect 51906 301271 51962 301280
rect 54496 260001 54524 336738
rect 55876 278769 55904 401610
rect 62118 389328 62174 389337
rect 62118 389263 62120 389272
rect 62172 389263 62174 389272
rect 62120 389234 62172 389240
rect 62118 376272 62174 376281
rect 62118 376207 62174 376216
rect 62132 375426 62160 376207
rect 62120 375420 62172 375426
rect 62120 375362 62172 375368
rect 62118 363352 62174 363361
rect 62118 363287 62174 363296
rect 62132 362982 62160 363287
rect 62120 362976 62172 362982
rect 62120 362918 62172 362924
rect 62118 350296 62174 350305
rect 62118 350231 62174 350240
rect 62132 347070 62160 350231
rect 62120 347064 62172 347070
rect 62120 347006 62172 347012
rect 62776 345681 62804 415375
rect 651470 404696 651526 404705
rect 651470 404631 651526 404640
rect 651484 404394 651512 404631
rect 651472 404388 651524 404394
rect 651472 404330 651524 404336
rect 652574 391504 652630 391513
rect 652574 391439 652630 391448
rect 652588 390590 652616 391439
rect 652576 390584 652628 390590
rect 652576 390526 652628 390532
rect 658924 390584 658976 390590
rect 658924 390526 658976 390532
rect 652392 378208 652444 378214
rect 652390 378176 652392 378185
rect 652444 378176 652446 378185
rect 652390 378111 652446 378120
rect 651838 364848 651894 364857
rect 651838 364783 651894 364792
rect 651852 364410 651880 364783
rect 651840 364404 651892 364410
rect 651840 364346 651892 364352
rect 652390 351656 652446 351665
rect 652390 351591 652446 351600
rect 652404 350606 652432 351591
rect 652392 350600 652444 350606
rect 652392 350542 652444 350548
rect 62762 345672 62818 345681
rect 62762 345607 62818 345616
rect 652022 338328 652078 338337
rect 652022 338263 652078 338272
rect 62118 337240 62174 337249
rect 62118 337175 62174 337184
rect 62132 336802 62160 337175
rect 62120 336796 62172 336802
rect 62120 336738 62172 336744
rect 651470 325000 651526 325009
rect 651470 324935 651526 324944
rect 651484 324358 651512 324935
rect 651472 324352 651524 324358
rect 651472 324294 651524 324300
rect 651470 311808 651526 311817
rect 651470 311743 651526 311752
rect 62118 311128 62174 311137
rect 62118 311063 62174 311072
rect 62132 310554 62160 311063
rect 651484 310554 651512 311743
rect 62120 310548 62172 310554
rect 62120 310490 62172 310496
rect 651472 310548 651524 310554
rect 651472 310490 651524 310496
rect 62118 298208 62174 298217
rect 62118 298143 62120 298152
rect 62172 298143 62174 298152
rect 62120 298114 62172 298120
rect 651470 285288 651526 285297
rect 651470 285223 651526 285232
rect 62762 285152 62818 285161
rect 62762 285087 62818 285096
rect 55862 278760 55918 278769
rect 55862 278695 55918 278704
rect 54482 259992 54538 260001
rect 54482 259927 54538 259936
rect 57244 228404 57296 228410
rect 57244 228346 57296 228352
rect 56508 227044 56560 227050
rect 56508 226986 56560 226992
rect 51722 222864 51778 222873
rect 51722 222799 51778 222808
rect 56520 218210 56548 226986
rect 55956 218204 56008 218210
rect 55956 218146 56008 218152
rect 56508 218204 56560 218210
rect 56508 218146 56560 218152
rect 55968 217002 55996 218146
rect 57256 218074 57284 228346
rect 60004 225752 60056 225758
rect 60004 225694 60056 225700
rect 59266 224224 59322 224233
rect 59266 224159 59322 224168
rect 57612 218340 57664 218346
rect 57612 218282 57664 218288
rect 56508 218068 56560 218074
rect 56508 218010 56560 218016
rect 57244 218068 57296 218074
rect 57244 218010 57296 218016
rect 56520 217002 56548 218010
rect 57624 217002 57652 218282
rect 58440 218068 58492 218074
rect 58440 218010 58492 218016
rect 58452 217002 58480 218010
rect 59280 217002 59308 224159
rect 59820 218748 59872 218754
rect 59820 218690 59872 218696
rect 59832 217002 59860 218690
rect 60016 218074 60044 225694
rect 61844 225616 61896 225622
rect 62776 225593 62804 285087
rect 651484 284374 651512 285223
rect 651472 284368 651524 284374
rect 651472 284310 651524 284316
rect 65904 272542 65932 277780
rect 67022 277766 67588 277794
rect 65892 272536 65944 272542
rect 65892 272478 65944 272484
rect 67560 270094 67588 277766
rect 68204 271318 68232 277780
rect 68192 271312 68244 271318
rect 68192 271254 68244 271260
rect 67548 270088 67600 270094
rect 67548 270030 67600 270036
rect 69400 269822 69428 277780
rect 70596 275330 70624 277780
rect 70584 275324 70636 275330
rect 70584 275266 70636 275272
rect 71792 274718 71820 277780
rect 71780 274712 71832 274718
rect 71780 274654 71832 274660
rect 72988 271182 73016 277780
rect 74092 274718 74120 277780
rect 73804 274712 73856 274718
rect 73804 274654 73856 274660
rect 74080 274712 74132 274718
rect 74080 274654 74132 274660
rect 72976 271176 73028 271182
rect 72976 271118 73028 271124
rect 69388 269816 69440 269822
rect 69388 269758 69440 269764
rect 73816 267034 73844 274654
rect 75288 273970 75316 277780
rect 76484 275466 76512 277780
rect 76472 275460 76524 275466
rect 76472 275402 76524 275408
rect 77208 274712 77260 274718
rect 77208 274654 77260 274660
rect 75276 273964 75328 273970
rect 75276 273906 75328 273912
rect 75920 270088 75972 270094
rect 75920 270030 75972 270036
rect 75932 267073 75960 270030
rect 77220 269958 77248 274654
rect 77680 274106 77708 277780
rect 77668 274100 77720 274106
rect 77668 274042 77720 274048
rect 78876 270366 78904 277780
rect 78864 270360 78916 270366
rect 78864 270302 78916 270308
rect 80072 270094 80100 277780
rect 81268 274990 81296 277780
rect 81256 274984 81308 274990
rect 81256 274926 81308 274932
rect 82372 272678 82400 277780
rect 82360 272672 82412 272678
rect 82360 272614 82412 272620
rect 83568 271046 83596 277780
rect 84778 277766 85528 277794
rect 83556 271040 83608 271046
rect 83556 270982 83608 270988
rect 85500 270230 85528 277766
rect 85960 275602 85988 277780
rect 85948 275596 86000 275602
rect 85948 275538 86000 275544
rect 86224 274984 86276 274990
rect 86224 274926 86276 274932
rect 85488 270224 85540 270230
rect 85488 270166 85540 270172
rect 80060 270088 80112 270094
rect 80060 270030 80112 270036
rect 77208 269952 77260 269958
rect 77208 269894 77260 269900
rect 86236 267170 86264 274926
rect 87156 268394 87184 277780
rect 88352 275874 88380 277780
rect 88340 275868 88392 275874
rect 88340 275810 88392 275816
rect 89548 271454 89576 277780
rect 90666 277766 91048 277794
rect 91862 277766 92428 277794
rect 89536 271448 89588 271454
rect 89536 271390 89588 271396
rect 91020 268666 91048 277766
rect 91008 268660 91060 268666
rect 91008 268602 91060 268608
rect 92400 268530 92428 277766
rect 93044 274378 93072 277780
rect 93032 274372 93084 274378
rect 93032 274314 93084 274320
rect 94240 272814 94268 277780
rect 95436 274242 95464 277780
rect 96632 275738 96660 277780
rect 96620 275732 96672 275738
rect 96620 275674 96672 275680
rect 97736 274378 97764 277780
rect 98946 277766 99328 277794
rect 100142 277766 100708 277794
rect 101338 277766 102088 277794
rect 95884 274372 95936 274378
rect 95884 274314 95936 274320
rect 97724 274372 97776 274378
rect 97724 274314 97776 274320
rect 95424 274236 95476 274242
rect 95424 274178 95476 274184
rect 94228 272808 94280 272814
rect 94228 272750 94280 272756
rect 92388 268524 92440 268530
rect 92388 268466 92440 268472
rect 87144 268388 87196 268394
rect 87144 268330 87196 268336
rect 95896 267306 95924 274314
rect 99300 268802 99328 277766
rect 100680 270502 100708 277766
rect 100668 270496 100720 270502
rect 100668 270438 100720 270444
rect 102060 269793 102088 277766
rect 102520 272950 102548 277780
rect 103716 276010 103744 277780
rect 103704 276004 103756 276010
rect 103704 275946 103756 275952
rect 102508 272944 102560 272950
rect 102508 272886 102560 272892
rect 104912 271726 104940 277780
rect 104900 271720 104952 271726
rect 104900 271662 104952 271668
rect 106016 271590 106044 277780
rect 107226 277766 107608 277794
rect 108422 277766 108988 277794
rect 109618 277766 110276 277794
rect 106004 271584 106056 271590
rect 106004 271526 106056 271532
rect 102046 269784 102102 269793
rect 102046 269719 102102 269728
rect 99288 268796 99340 268802
rect 99288 268738 99340 268744
rect 99288 268660 99340 268666
rect 99288 268602 99340 268608
rect 99300 267578 99328 268602
rect 107580 267734 107608 277766
rect 108960 268938 108988 277766
rect 108948 268932 109000 268938
rect 108948 268874 109000 268880
rect 110248 268802 110276 277766
rect 110800 275194 110828 277780
rect 110788 275188 110840 275194
rect 110788 275130 110840 275136
rect 111996 273086 112024 277780
rect 111984 273080 112036 273086
rect 111984 273022 112036 273028
rect 113192 270774 113220 277780
rect 114296 274514 114324 277780
rect 115506 277766 115888 277794
rect 114284 274508 114336 274514
rect 114284 274450 114336 274456
rect 113180 270768 113232 270774
rect 113180 270710 113232 270716
rect 115860 269074 115888 277766
rect 116688 272270 116716 277780
rect 117898 277766 118648 277794
rect 116676 272264 116728 272270
rect 116676 272206 116728 272212
rect 115848 269068 115900 269074
rect 115848 269010 115900 269016
rect 110236 268796 110288 268802
rect 110236 268738 110288 268744
rect 118620 268258 118648 277766
rect 119080 269686 119108 277780
rect 120276 274650 120304 277780
rect 120264 274644 120316 274650
rect 120264 274586 120316 274592
rect 121380 271862 121408 277780
rect 122590 277766 122788 277794
rect 121368 271856 121420 271862
rect 121368 271798 121420 271804
rect 122760 270502 122788 277766
rect 123772 271046 123800 277780
rect 124968 273698 124996 277780
rect 126178 277766 126928 277794
rect 124956 273692 125008 273698
rect 124956 273634 125008 273640
rect 123484 271040 123536 271046
rect 123484 270982 123536 270988
rect 123760 271040 123812 271046
rect 123760 270982 123812 270988
rect 119804 270496 119856 270502
rect 119804 270438 119856 270444
rect 122748 270496 122800 270502
rect 122748 270438 122800 270444
rect 119068 269680 119120 269686
rect 119068 269622 119120 269628
rect 118608 268252 118660 268258
rect 118608 268194 118660 268200
rect 107580 267706 107700 267734
rect 99288 267572 99340 267578
rect 99288 267514 99340 267520
rect 107672 267442 107700 267706
rect 107660 267436 107712 267442
rect 107660 267378 107712 267384
rect 95884 267300 95936 267306
rect 95884 267242 95936 267248
rect 86224 267164 86276 267170
rect 86224 267106 86276 267112
rect 75918 267064 75974 267073
rect 73804 267028 73856 267034
rect 75918 266999 75974 267008
rect 73804 266970 73856 266976
rect 119816 266898 119844 270438
rect 119804 266892 119856 266898
rect 119804 266834 119856 266840
rect 123496 266626 123524 270982
rect 126900 269550 126928 277766
rect 127360 273222 127388 277780
rect 127348 273216 127400 273222
rect 127348 273158 127400 273164
rect 128556 272406 128584 277780
rect 129660 274922 129688 277780
rect 129648 274916 129700 274922
rect 129648 274858 129700 274864
rect 130856 273834 130884 277780
rect 132066 277766 132448 277794
rect 133262 277766 133828 277794
rect 130844 273828 130896 273834
rect 130844 273770 130896 273776
rect 128544 272400 128596 272406
rect 128544 272342 128596 272348
rect 126888 269544 126940 269550
rect 126888 269486 126940 269492
rect 132420 267714 132448 277766
rect 133800 270366 133828 277766
rect 134444 270910 134472 277780
rect 135640 275058 135668 277780
rect 136850 277766 137048 277794
rect 135628 275052 135680 275058
rect 135628 274994 135680 275000
rect 136088 274916 136140 274922
rect 136088 274858 136140 274864
rect 134432 270904 134484 270910
rect 134432 270846 134484 270852
rect 132592 270360 132644 270366
rect 132592 270302 132644 270308
rect 133788 270360 133840 270366
rect 133788 270302 133840 270308
rect 132408 267708 132460 267714
rect 132408 267650 132460 267656
rect 132604 266762 132632 270302
rect 136100 269414 136128 274858
rect 136824 272536 136876 272542
rect 136824 272478 136876 272484
rect 136088 269408 136140 269414
rect 136088 269350 136140 269356
rect 132592 266756 132644 266762
rect 132592 266698 132644 266704
rect 123484 266620 123536 266626
rect 123484 266562 123536 266568
rect 136836 264330 136864 272478
rect 137020 268122 137048 277766
rect 137940 272542 137968 277780
rect 137928 272536 137980 272542
rect 137928 272478 137980 272484
rect 139136 271318 139164 277780
rect 140346 277766 140728 277794
rect 141542 277766 141832 277794
rect 140136 275324 140188 275330
rect 140136 275266 140188 275272
rect 138480 271312 138532 271318
rect 138480 271254 138532 271260
rect 139124 271312 139176 271318
rect 139124 271254 139176 271260
rect 137008 268116 137060 268122
rect 137008 268058 137060 268064
rect 138110 267064 138166 267073
rect 138110 266999 138166 267008
rect 136836 264302 137310 264330
rect 138124 264316 138152 266999
rect 138492 264330 138520 271254
rect 139768 269816 139820 269822
rect 139768 269758 139820 269764
rect 138492 264302 138966 264330
rect 139780 264316 139808 269758
rect 140148 264330 140176 275266
rect 140700 269822 140728 277766
rect 141804 271318 141832 277766
rect 142724 274922 142752 277780
rect 143934 277766 144132 277794
rect 145038 277766 145328 277794
rect 143264 275460 143316 275466
rect 143264 275402 143316 275408
rect 142712 274916 142764 274922
rect 142712 274858 142764 274864
rect 142160 273964 142212 273970
rect 142160 273906 142212 273912
rect 141608 271312 141660 271318
rect 141608 271254 141660 271260
rect 141792 271312 141844 271318
rect 141792 271254 141844 271260
rect 140688 269816 140740 269822
rect 140688 269758 140740 269764
rect 141424 267028 141476 267034
rect 141424 266970 141476 266976
rect 140148 264302 140622 264330
rect 141436 264316 141464 266970
rect 141620 266490 141648 271254
rect 141608 266484 141660 266490
rect 141608 266426 141660 266432
rect 142172 265946 142200 273906
rect 143276 271182 143304 275402
rect 142344 271176 142396 271182
rect 142344 271118 142396 271124
rect 143264 271176 143316 271182
rect 143264 271118 143316 271124
rect 142160 265940 142212 265946
rect 142160 265882 142212 265888
rect 142356 265826 142384 271118
rect 144104 269958 144132 277766
rect 145300 274106 145328 277766
rect 146220 274786 146248 277780
rect 146944 275868 146996 275874
rect 146944 275810 146996 275816
rect 146208 274780 146260 274786
rect 146208 274722 146260 274728
rect 145104 274100 145156 274106
rect 145104 274042 145156 274048
rect 145288 274100 145340 274106
rect 145288 274042 145340 274048
rect 144368 271176 144420 271182
rect 144368 271118 144420 271124
rect 143908 269952 143960 269958
rect 143908 269894 143960 269900
rect 144092 269952 144144 269958
rect 144092 269894 144144 269900
rect 142804 265940 142856 265946
rect 142804 265882 142856 265888
rect 142264 265798 142384 265826
rect 142264 264316 142292 265798
rect 142816 264330 142844 265882
rect 142816 264302 143106 264330
rect 143920 264316 143948 269894
rect 144380 264330 144408 271118
rect 145116 264330 145144 274042
rect 146392 270088 146444 270094
rect 146392 270030 146444 270036
rect 144380 264302 144762 264330
rect 145116 264302 145590 264330
rect 146404 264316 146432 270030
rect 146956 269210 146984 275810
rect 147416 273970 147444 277780
rect 148612 275466 148640 277780
rect 149808 275874 149836 277780
rect 149796 275868 149848 275874
rect 149796 275810 149848 275816
rect 150808 275596 150860 275602
rect 150808 275538 150860 275544
rect 148600 275460 148652 275466
rect 148600 275402 148652 275408
rect 149704 274780 149756 274786
rect 149704 274722 149756 274728
rect 147404 273964 147456 273970
rect 147404 273906 147456 273912
rect 148416 273692 148468 273698
rect 148416 273634 148468 273640
rect 148232 272672 148284 272678
rect 148232 272614 148284 272620
rect 146944 269204 146996 269210
rect 146944 269146 146996 269152
rect 148244 267734 148272 272614
rect 148428 267734 148456 273634
rect 149428 270224 149480 270230
rect 149428 270166 149480 270172
rect 148244 267706 148364 267734
rect 148428 267706 148548 267734
rect 148048 267164 148100 267170
rect 148048 267106 148100 267112
rect 146944 267028 146996 267034
rect 146944 266970 146996 266976
rect 146956 266490 146984 266970
rect 147220 266756 147272 266762
rect 147220 266698 147272 266704
rect 146944 266484 146996 266490
rect 146944 266426 146996 266432
rect 147232 264316 147260 266698
rect 148060 264316 148088 267106
rect 148336 264330 148364 267706
rect 148520 266762 148548 267706
rect 148508 266756 148560 266762
rect 148508 266698 148560 266704
rect 149440 264330 149468 270166
rect 149716 267170 149744 274722
rect 150820 267734 150848 275538
rect 151004 274786 151032 277780
rect 150992 274780 151044 274786
rect 150992 274722 151044 274728
rect 152200 272134 152228 277780
rect 152740 274780 152792 274786
rect 152740 274722 152792 274728
rect 152188 272128 152240 272134
rect 152188 272070 152240 272076
rect 152372 271448 152424 271454
rect 152372 271390 152424 271396
rect 152188 268388 152240 268394
rect 152188 268330 152240 268336
rect 150820 267706 151032 267734
rect 149704 267164 149756 267170
rect 149704 267106 149756 267112
rect 150532 266620 150584 266626
rect 150532 266562 150584 266568
rect 148336 264302 148902 264330
rect 149440 264302 149730 264330
rect 150544 264316 150572 266562
rect 151004 264330 151032 267706
rect 151004 264302 151386 264330
rect 152200 264316 152228 268330
rect 152384 267734 152412 271390
rect 152752 268394 152780 274722
rect 153304 270230 153332 277780
rect 154316 277766 154514 277794
rect 154316 271182 154344 277766
rect 155696 273698 155724 277780
rect 156604 275732 156656 275738
rect 156604 275674 156656 275680
rect 155684 273692 155736 273698
rect 155684 273634 155736 273640
rect 155960 272808 156012 272814
rect 155960 272750 156012 272756
rect 154304 271176 154356 271182
rect 154304 271118 154356 271124
rect 154028 270768 154080 270774
rect 154028 270710 154080 270716
rect 153292 270224 153344 270230
rect 153292 270166 153344 270172
rect 153844 269204 153896 269210
rect 153844 269146 153896 269152
rect 152740 268388 152792 268394
rect 152740 268330 152792 268336
rect 152384 267706 152688 267734
rect 152660 264330 152688 267706
rect 152660 264302 153042 264330
rect 153856 264316 153884 269146
rect 154040 266626 154068 270710
rect 155500 268524 155552 268530
rect 155500 268466 155552 268472
rect 154672 267572 154724 267578
rect 154672 267514 154724 267520
rect 154028 266620 154080 266626
rect 154028 266562 154080 266568
rect 154684 264316 154712 267514
rect 155512 264316 155540 268466
rect 155972 264330 156000 272750
rect 156616 266422 156644 275674
rect 156892 275330 156920 277780
rect 158102 277766 158668 277794
rect 159298 277766 160048 277794
rect 156880 275324 156932 275330
rect 156880 275266 156932 275272
rect 157616 274236 157668 274242
rect 157616 274178 157668 274184
rect 157156 267300 157208 267306
rect 157156 267242 157208 267248
rect 156604 266416 156656 266422
rect 156604 266358 156656 266364
rect 155972 264302 156354 264330
rect 157168 264316 157196 267242
rect 157628 264330 157656 274178
rect 158640 270094 158668 277766
rect 158812 274372 158864 274378
rect 158812 274314 158864 274320
rect 158628 270088 158680 270094
rect 158628 270030 158680 270036
rect 157628 264302 158010 264330
rect 158824 264316 158852 274314
rect 160020 268530 160048 277766
rect 160480 275602 160508 277780
rect 160744 276004 160796 276010
rect 160744 275946 160796 275952
rect 160468 275596 160520 275602
rect 160468 275538 160520 275544
rect 160468 268660 160520 268666
rect 160468 268602 160520 268608
rect 160008 268524 160060 268530
rect 160008 268466 160060 268472
rect 159640 266416 159692 266422
rect 159640 266358 159692 266364
rect 159652 264316 159680 266358
rect 160480 264316 160508 268602
rect 160756 267578 160784 275946
rect 161584 272678 161612 277780
rect 162124 272944 162176 272950
rect 162124 272886 162176 272892
rect 161572 272672 161624 272678
rect 161572 272614 161624 272620
rect 161294 269784 161350 269793
rect 161294 269719 161350 269728
rect 160744 267572 160796 267578
rect 160744 267514 160796 267520
rect 161308 264316 161336 269719
rect 161756 266892 161808 266898
rect 161756 266834 161808 266840
rect 161768 264330 161796 266834
rect 162136 266422 162164 272886
rect 162780 271454 162808 277780
rect 163976 274786 164004 277780
rect 165186 277766 165568 277794
rect 165540 276026 165568 277766
rect 165540 275998 165660 276026
rect 166368 276010 166396 277780
rect 164148 275460 164200 275466
rect 164148 275402 164200 275408
rect 163964 274780 164016 274786
rect 163964 274722 164016 274728
rect 164160 271726 164188 275402
rect 164976 275188 165028 275194
rect 164976 275130 165028 275136
rect 163320 271720 163372 271726
rect 163320 271662 163372 271668
rect 164148 271720 164200 271726
rect 164148 271662 164200 271668
rect 162768 271448 162820 271454
rect 162768 271390 162820 271396
rect 162124 266416 162176 266422
rect 162124 266358 162176 266364
rect 162952 266416 163004 266422
rect 162952 266358 163004 266364
rect 161768 264302 162150 264330
rect 162964 264316 162992 266358
rect 163332 264330 163360 271662
rect 164792 271584 164844 271590
rect 164792 271526 164844 271532
rect 164804 267734 164832 271526
rect 164988 267734 165016 275130
rect 165632 274242 165660 275998
rect 166356 276004 166408 276010
rect 166356 275946 166408 275952
rect 167564 275466 167592 277780
rect 167552 275460 167604 275466
rect 167552 275402 167604 275408
rect 167644 275052 167696 275058
rect 167644 274994 167696 275000
rect 166264 274916 166316 274922
rect 166264 274858 166316 274864
rect 165620 274236 165672 274242
rect 165620 274178 165672 274184
rect 166276 272270 166304 274858
rect 166080 272264 166132 272270
rect 166080 272206 166132 272212
rect 166264 272264 166316 272270
rect 166264 272206 166316 272212
rect 166092 270042 166120 272206
rect 166092 270014 166488 270042
rect 166264 268932 166316 268938
rect 166264 268874 166316 268880
rect 164804 267706 164924 267734
rect 164988 267706 165108 267734
rect 164608 267572 164660 267578
rect 164608 267514 164660 267520
rect 163332 264302 163806 264330
rect 164620 264316 164648 267514
rect 164896 264330 164924 267706
rect 165080 266422 165108 267706
rect 165068 266416 165120 266422
rect 165068 266358 165120 266364
rect 164896 264302 165462 264330
rect 166276 264316 166304 268874
rect 166460 267578 166488 270014
rect 166448 267572 166500 267578
rect 166448 267514 166500 267520
rect 167656 267442 167684 274994
rect 168380 273080 168432 273086
rect 168380 273022 168432 273028
rect 167920 268796 167972 268802
rect 167920 268738 167972 268744
rect 167092 267436 167144 267442
rect 167092 267378 167144 267384
rect 167644 267436 167696 267442
rect 167644 267378 167696 267384
rect 167104 264316 167132 267378
rect 167932 264316 167960 268738
rect 168392 264330 168420 273022
rect 168668 268666 168696 277780
rect 169878 277766 170076 277794
rect 170048 270230 170076 277766
rect 171060 275194 171088 277780
rect 171048 275188 171100 275194
rect 171048 275130 171100 275136
rect 172256 274786 172284 277780
rect 173466 277766 173848 277794
rect 172428 275596 172480 275602
rect 172428 275538 172480 275544
rect 170404 274780 170456 274786
rect 170404 274722 170456 274728
rect 172244 274780 172296 274786
rect 172244 274722 172296 274728
rect 169852 270224 169904 270230
rect 169852 270166 169904 270172
rect 170036 270224 170088 270230
rect 170036 270166 170088 270172
rect 168656 268660 168708 268666
rect 168656 268602 168708 268608
rect 169864 266898 169892 270166
rect 170416 267306 170444 274722
rect 171600 274508 171652 274514
rect 171600 274450 171652 274456
rect 171232 269068 171284 269074
rect 171232 269010 171284 269016
rect 170404 267300 170456 267306
rect 170404 267242 170456 267248
rect 169852 266892 169904 266898
rect 169852 266834 169904 266840
rect 170404 266620 170456 266626
rect 170404 266562 170456 266568
rect 169576 266416 169628 266422
rect 169576 266358 169628 266364
rect 168392 264302 168774 264330
rect 169588 264316 169616 266358
rect 170416 264316 170444 266562
rect 171244 264316 171272 269010
rect 171612 264330 171640 274450
rect 172440 268938 172468 275538
rect 173348 269680 173400 269686
rect 173348 269622 173400 269628
rect 172428 268932 172480 268938
rect 172428 268874 172480 268880
rect 172888 267572 172940 267578
rect 172888 267514 172940 267520
rect 171612 264302 172086 264330
rect 172900 264316 172928 267514
rect 173360 264330 173388 269622
rect 173820 268802 173848 277766
rect 174648 275738 174676 277780
rect 174636 275732 174688 275738
rect 174636 275674 174688 275680
rect 174360 274780 174412 274786
rect 174360 274722 174412 274728
rect 174372 269686 174400 274722
rect 175280 274644 175332 274650
rect 175280 274586 175332 274592
rect 174360 269680 174412 269686
rect 174360 269622 174412 269628
rect 173808 268796 173860 268802
rect 173808 268738 173860 268744
rect 174544 268252 174596 268258
rect 174544 268194 174596 268200
rect 173360 264302 173742 264330
rect 174556 264316 174584 268194
rect 175292 264330 175320 274586
rect 175844 270774 175872 277780
rect 176752 271856 176804 271862
rect 176752 271798 176804 271804
rect 175832 270768 175884 270774
rect 175832 270710 175884 270716
rect 176200 270496 176252 270502
rect 176200 270438 176252 270444
rect 175292 264302 175398 264330
rect 176212 264316 176240 270438
rect 176764 264330 176792 271798
rect 176948 270502 176976 277780
rect 178144 271590 178172 277780
rect 179340 274514 179368 277780
rect 179328 274508 179380 274514
rect 179328 274450 179380 274456
rect 180536 274378 180564 277780
rect 181732 275602 181760 277780
rect 182942 277766 183508 277794
rect 184138 277766 184520 277794
rect 182088 276004 182140 276010
rect 182088 275946 182140 275952
rect 181720 275596 181772 275602
rect 181720 275538 181772 275544
rect 180524 274372 180576 274378
rect 180524 274314 180576 274320
rect 181444 273828 181496 273834
rect 181444 273770 181496 273776
rect 179880 273216 179932 273222
rect 179880 273158 179932 273164
rect 178132 271584 178184 271590
rect 178132 271526 178184 271532
rect 177488 271040 177540 271046
rect 177488 270982 177540 270988
rect 176936 270496 176988 270502
rect 176936 270438 176988 270444
rect 177500 264330 177528 270982
rect 178684 269544 178736 269550
rect 178684 269486 178736 269492
rect 176764 264302 177054 264330
rect 177500 264302 177882 264330
rect 178696 264316 178724 269486
rect 179512 266756 179564 266762
rect 179512 266698 179564 266704
rect 179524 264316 179552 266698
rect 179892 264330 179920 273158
rect 181260 272400 181312 272406
rect 181260 272342 181312 272348
rect 180892 269408 180944 269414
rect 180892 269350 180944 269356
rect 180904 264330 180932 269350
rect 181272 267734 181300 272342
rect 181456 267734 181484 273770
rect 182100 273086 182128 275946
rect 182088 273080 182140 273086
rect 182088 273022 182140 273028
rect 183480 269550 183508 277766
rect 184492 271590 184520 277766
rect 185228 271862 185256 277780
rect 185216 271856 185268 271862
rect 185216 271798 185268 271804
rect 184204 271584 184256 271590
rect 184204 271526 184256 271532
rect 184480 271584 184532 271590
rect 184480 271526 184532 271532
rect 183652 270360 183704 270366
rect 183652 270302 183704 270308
rect 183468 269544 183520 269550
rect 183468 269486 183520 269492
rect 183008 268116 183060 268122
rect 183008 268058 183060 268064
rect 181272 267706 181392 267734
rect 181456 267706 181576 267734
rect 181364 264466 181392 267706
rect 181548 266422 181576 267706
rect 183020 266422 183048 268058
rect 181536 266416 181588 266422
rect 181536 266358 181588 266364
rect 182824 266416 182876 266422
rect 182824 266358 182876 266364
rect 183008 266416 183060 266422
rect 183008 266358 183060 266364
rect 181364 264438 181576 264466
rect 181548 264330 181576 264438
rect 179892 264302 180366 264330
rect 180904 264302 181194 264330
rect 181548 264302 182022 264330
rect 182836 264316 182864 266358
rect 183664 264316 183692 270302
rect 184216 267714 184244 271526
rect 184940 270904 184992 270910
rect 184940 270846 184992 270852
rect 184204 267708 184256 267714
rect 184204 267650 184256 267656
rect 184480 267572 184532 267578
rect 184480 267514 184532 267520
rect 184492 264316 184520 267514
rect 184952 264330 184980 270846
rect 186424 270366 186452 277780
rect 187620 272814 187648 277780
rect 188816 276010 188844 277780
rect 188804 276004 188856 276010
rect 188804 275946 188856 275952
rect 187884 275868 187936 275874
rect 187884 275810 187936 275816
rect 187608 272808 187660 272814
rect 187608 272750 187660 272756
rect 187700 272536 187752 272542
rect 187700 272478 187752 272484
rect 186964 271856 187016 271862
rect 186964 271798 187016 271804
rect 186412 270360 186464 270366
rect 186412 270302 186464 270308
rect 186976 267578 187004 271798
rect 186964 267572 187016 267578
rect 186964 267514 187016 267520
rect 186964 267436 187016 267442
rect 186964 267378 187016 267384
rect 186136 266416 186188 266422
rect 186136 266358 186188 266364
rect 184952 264302 185334 264330
rect 186148 264316 186176 266358
rect 186976 264316 187004 267378
rect 187712 264330 187740 272478
rect 187896 271862 187924 275810
rect 189816 274100 189868 274106
rect 189816 274042 189868 274048
rect 187884 271856 187936 271862
rect 187884 271798 187936 271804
rect 189632 271312 189684 271318
rect 189632 271254 189684 271260
rect 188620 269816 188672 269822
rect 188620 269758 188672 269764
rect 187712 264302 187818 264330
rect 188632 264316 188660 269758
rect 189644 267734 189672 271254
rect 189828 267734 189856 274042
rect 190012 272950 190040 277780
rect 191012 275188 191064 275194
rect 191012 275130 191064 275136
rect 190000 272944 190052 272950
rect 190000 272886 190052 272892
rect 190828 269952 190880 269958
rect 190828 269894 190880 269900
rect 189644 267706 189764 267734
rect 189828 267706 189948 267734
rect 189448 267028 189500 267034
rect 189448 266970 189500 266976
rect 189460 264316 189488 266970
rect 189736 264330 189764 267706
rect 189920 267442 189948 267706
rect 189908 267436 189960 267442
rect 189908 267378 189960 267384
rect 190840 264330 190868 269894
rect 191024 267034 191052 275130
rect 191208 274106 191236 277780
rect 191196 274100 191248 274106
rect 191196 274042 191248 274048
rect 192312 272542 192340 277780
rect 193508 273970 193536 277780
rect 194704 277394 194732 277780
rect 194612 277366 194732 277394
rect 195716 277766 195914 277794
rect 193312 273964 193364 273970
rect 193312 273906 193364 273912
rect 193496 273964 193548 273970
rect 193496 273906 193548 273912
rect 192300 272536 192352 272542
rect 192300 272478 192352 272484
rect 191840 272264 191892 272270
rect 191840 272206 191892 272212
rect 191012 267028 191064 267034
rect 191012 266970 191064 266976
rect 191852 264330 191880 272206
rect 192484 272128 192536 272134
rect 192484 272070 192536 272076
rect 192496 266422 192524 272070
rect 193128 267844 193180 267850
rect 193128 267786 193180 267792
rect 193140 267714 193168 267786
rect 193128 267708 193180 267714
rect 193128 267650 193180 267656
rect 192760 267436 192812 267442
rect 192760 267378 192812 267384
rect 192484 266416 192536 266422
rect 192484 266358 192536 266364
rect 189736 264302 190302 264330
rect 190840 264302 191130 264330
rect 191852 264302 191958 264330
rect 192772 264316 192800 267378
rect 193324 264330 193352 273906
rect 194612 269822 194640 277366
rect 194784 271720 194836 271726
rect 194784 271662 194836 271668
rect 194600 269816 194652 269822
rect 194600 269758 194652 269764
rect 194416 267164 194468 267170
rect 194416 267106 194468 267112
rect 193324 264302 193614 264330
rect 194428 264316 194456 267106
rect 194796 264330 194824 271662
rect 195716 271318 195744 277766
rect 196440 271856 196492 271862
rect 196440 271798 196492 271804
rect 195704 271312 195756 271318
rect 195704 271254 195756 271260
rect 196072 268388 196124 268394
rect 196072 268330 196124 268336
rect 194796 264302 195270 264330
rect 196084 264316 196112 268330
rect 196452 264330 196480 271798
rect 197096 271726 197124 277780
rect 198096 273692 198148 273698
rect 198096 273634 198148 273640
rect 197084 271720 197136 271726
rect 197084 271662 197136 271668
rect 197912 271176 197964 271182
rect 197912 271118 197964 271124
rect 197924 267734 197952 271118
rect 198108 267734 198136 273634
rect 198292 271182 198320 277780
rect 199292 275324 199344 275330
rect 199292 275266 199344 275272
rect 198280 271176 198332 271182
rect 198280 271118 198332 271124
rect 197924 267706 198044 267734
rect 198108 267706 198228 267734
rect 197728 266416 197780 266422
rect 197728 266358 197780 266364
rect 196452 264302 196926 264330
rect 197740 264316 197768 266358
rect 198016 264330 198044 267706
rect 198200 267170 198228 267706
rect 198188 267164 198240 267170
rect 198188 267106 198240 267112
rect 199304 266898 199332 275266
rect 199488 274854 199516 277780
rect 199476 274848 199528 274854
rect 199476 274790 199528 274796
rect 200396 268524 200448 268530
rect 200396 268466 200448 268472
rect 200212 267164 200264 267170
rect 200212 267106 200264 267112
rect 199108 266892 199160 266898
rect 199108 266834 199160 266840
rect 199292 266892 199344 266898
rect 199292 266834 199344 266840
rect 199120 264330 199148 266834
rect 198016 264302 198582 264330
rect 199120 264302 199410 264330
rect 200224 264316 200252 267106
rect 200408 266422 200436 268466
rect 200592 268394 200620 277780
rect 201592 270360 201644 270366
rect 201592 270302 201644 270308
rect 201040 270088 201092 270094
rect 201040 270030 201092 270036
rect 200580 268388 200632 268394
rect 200580 268330 200632 268336
rect 200396 266416 200448 266422
rect 200396 266358 200448 266364
rect 201052 264316 201080 270030
rect 201604 266762 201632 270302
rect 201788 269958 201816 277780
rect 202998 277766 203288 277794
rect 202236 274848 202288 274854
rect 202236 274790 202288 274796
rect 202248 270094 202276 274790
rect 203260 272678 203288 277766
rect 203064 272672 203116 272678
rect 203064 272614 203116 272620
rect 203248 272672 203300 272678
rect 203248 272614 203300 272620
rect 202236 270088 202288 270094
rect 202236 270030 202288 270036
rect 201776 269952 201828 269958
rect 201776 269894 201828 269900
rect 201868 266892 201920 266898
rect 201868 266834 201920 266840
rect 201592 266756 201644 266762
rect 201592 266698 201644 266704
rect 201880 264316 201908 266834
rect 202696 266416 202748 266422
rect 202696 266358 202748 266364
rect 202708 264316 202736 266358
rect 203076 264330 203104 272614
rect 204180 270366 204208 277780
rect 205376 271454 205404 277780
rect 206572 274242 206600 277780
rect 207782 277766 208256 277794
rect 205732 274236 205784 274242
rect 205732 274178 205784 274184
rect 206560 274236 206612 274242
rect 206560 274178 206612 274184
rect 204720 271448 204772 271454
rect 204720 271390 204772 271396
rect 205364 271448 205416 271454
rect 205364 271390 205416 271396
rect 204168 270360 204220 270366
rect 204168 270302 204220 270308
rect 204168 269544 204220 269550
rect 204168 269486 204220 269492
rect 204180 267714 204208 269486
rect 204352 268932 204404 268938
rect 204352 268874 204404 268880
rect 204168 267708 204220 267714
rect 204168 267650 204220 267656
rect 203076 264302 203550 264330
rect 204364 264316 204392 268874
rect 204732 264330 204760 271390
rect 205744 264330 205772 274178
rect 207296 273080 207348 273086
rect 207296 273022 207348 273028
rect 206284 270768 206336 270774
rect 206284 270710 206336 270716
rect 206296 267306 206324 270710
rect 206284 267300 206336 267306
rect 206284 267242 206336 267248
rect 206836 267164 206888 267170
rect 206836 267106 206888 267112
rect 207020 267164 207072 267170
rect 207020 267106 207072 267112
rect 204732 264302 205206 264330
rect 205744 264302 206034 264330
rect 206848 264316 206876 267106
rect 207032 266762 207060 267106
rect 207020 266756 207072 266762
rect 207020 266698 207072 266704
rect 207308 264330 207336 273022
rect 208228 268530 208256 277766
rect 208400 275732 208452 275738
rect 208400 275674 208452 275680
rect 208412 268938 208440 275674
rect 208872 274854 208900 277780
rect 209044 275460 209096 275466
rect 209044 275402 209096 275408
rect 208860 274848 208912 274854
rect 208860 274790 208912 274796
rect 208400 268932 208452 268938
rect 208400 268874 208452 268880
rect 208492 268660 208544 268666
rect 208492 268602 208544 268608
rect 208216 268524 208268 268530
rect 208216 268466 208268 268472
rect 207308 264302 207690 264330
rect 208504 264316 208532 268602
rect 209056 264330 209084 275402
rect 210068 274718 210096 277780
rect 211264 275330 211292 277780
rect 212460 275738 212488 277780
rect 212448 275732 212500 275738
rect 212448 275674 212500 275680
rect 211252 275324 211304 275330
rect 211252 275266 211304 275272
rect 211068 274848 211120 274854
rect 211068 274790 211120 274796
rect 210056 274712 210108 274718
rect 210056 274654 210108 274660
rect 211080 270230 211108 274790
rect 212264 274712 212316 274718
rect 212264 274654 212316 274660
rect 210148 270224 210200 270230
rect 210148 270166 210200 270172
rect 211068 270224 211120 270230
rect 211068 270166 211120 270172
rect 209056 264302 209346 264330
rect 210160 264316 210188 270166
rect 210976 269680 211028 269686
rect 210976 269622 211028 269628
rect 210988 264316 211016 269622
rect 212276 268666 212304 274654
rect 213656 274514 213684 277780
rect 214866 277766 215248 277794
rect 215970 277766 216352 277794
rect 213184 274508 213236 274514
rect 213184 274450 213236 274456
rect 213644 274508 213696 274514
rect 213644 274450 213696 274456
rect 212540 272808 212592 272814
rect 212540 272750 212592 272756
rect 212552 272406 212580 272750
rect 212540 272400 212592 272406
rect 212540 272342 212592 272348
rect 212632 268796 212684 268802
rect 212632 268738 212684 268744
rect 212264 268660 212316 268666
rect 212264 268602 212316 268608
rect 211804 267028 211856 267034
rect 211804 266970 211856 266976
rect 211816 264316 211844 266970
rect 212644 264316 212672 268738
rect 213196 266422 213224 274450
rect 214748 270496 214800 270502
rect 214748 270438 214800 270444
rect 214288 268932 214340 268938
rect 214288 268874 214340 268880
rect 213460 267300 213512 267306
rect 213460 267242 213512 267248
rect 213184 266416 213236 266422
rect 213184 266358 213236 266364
rect 213472 264316 213500 267242
rect 214300 264316 214328 268874
rect 214760 264330 214788 270438
rect 215220 268802 215248 277766
rect 216324 271590 216352 277766
rect 216956 274372 217008 274378
rect 216956 274314 217008 274320
rect 215944 271584 215996 271590
rect 215944 271526 215996 271532
rect 216312 271584 216364 271590
rect 216312 271526 216364 271532
rect 215208 268796 215260 268802
rect 215208 268738 215260 268744
rect 215956 267306 215984 271526
rect 216968 267734 216996 274314
rect 217152 272950 217180 277780
rect 218348 275466 218376 277780
rect 218612 275596 218664 275602
rect 218612 275538 218664 275544
rect 218336 275460 218388 275466
rect 218336 275402 218388 275408
rect 217140 272944 217192 272950
rect 217140 272886 217192 272892
rect 217416 272808 217468 272814
rect 217416 272750 217468 272756
rect 216968 267706 217272 267734
rect 216772 267572 216824 267578
rect 216772 267514 216824 267520
rect 215944 267300 215996 267306
rect 215944 267242 215996 267248
rect 215944 266416 215996 266422
rect 215944 266358 215996 266364
rect 214760 264302 215142 264330
rect 215956 264316 215984 266358
rect 216784 264316 216812 267514
rect 217244 264330 217272 267706
rect 217428 267578 217456 272750
rect 218428 267708 218480 267714
rect 218428 267650 218480 267656
rect 217416 267572 217468 267578
rect 217416 267514 217468 267520
rect 217244 264302 217626 264330
rect 218440 264316 218468 267650
rect 218624 264330 218652 275538
rect 218796 272400 218848 272406
rect 218796 272342 218848 272348
rect 218808 267714 218836 272342
rect 219544 270502 219572 277780
rect 220740 275806 220768 277780
rect 221936 277394 221964 277780
rect 221936 277366 222056 277394
rect 221464 276004 221516 276010
rect 221464 275946 221516 275952
rect 220728 275800 220780 275806
rect 220728 275742 220780 275748
rect 219900 275732 219952 275738
rect 219900 275674 219952 275680
rect 219912 272814 219940 275674
rect 219900 272808 219952 272814
rect 219900 272750 219952 272756
rect 219532 270496 219584 270502
rect 219532 270438 219584 270444
rect 220268 270360 220320 270366
rect 220268 270302 220320 270308
rect 218796 267708 218848 267714
rect 218796 267650 218848 267656
rect 220280 267306 220308 270302
rect 220084 267300 220136 267306
rect 220084 267242 220136 267248
rect 220268 267300 220320 267306
rect 220268 267242 220320 267248
rect 218624 264302 219282 264330
rect 220096 264316 220124 267242
rect 220912 267164 220964 267170
rect 220912 267106 220964 267112
rect 220924 264316 220952 267106
rect 221476 266422 221504 275946
rect 221740 267436 221792 267442
rect 221740 267378 221792 267384
rect 221464 266416 221516 266422
rect 221464 266358 221516 266364
rect 221752 264316 221780 267378
rect 222028 267034 222056 277366
rect 223132 273970 223160 277780
rect 224250 277766 224632 277794
rect 222844 273964 222896 273970
rect 222844 273906 222896 273912
rect 223120 273964 223172 273970
rect 223120 273906 223172 273912
rect 222568 267708 222620 267714
rect 222568 267650 222620 267656
rect 222016 267028 222068 267034
rect 222016 266970 222068 266976
rect 222580 264316 222608 267650
rect 222856 266558 222884 273906
rect 224604 271726 224632 277766
rect 224960 275800 225012 275806
rect 224960 275742 225012 275748
rect 224972 274106 225000 275742
rect 225432 275602 225460 277780
rect 225420 275596 225472 275602
rect 225420 275538 225472 275544
rect 224776 274100 224828 274106
rect 224776 274042 224828 274048
rect 224960 274100 225012 274106
rect 224960 274042 225012 274048
rect 224788 273986 224816 274042
rect 224788 273958 225000 273986
rect 224224 271720 224276 271726
rect 224224 271662 224276 271668
rect 224592 271720 224644 271726
rect 224592 271662 224644 271668
rect 223488 268796 223540 268802
rect 223488 268738 223540 268744
rect 223028 267572 223080 267578
rect 223028 267514 223080 267520
rect 222844 266552 222896 266558
rect 222844 266494 222896 266500
rect 223040 264330 223068 267514
rect 223500 267170 223528 268738
rect 224236 267578 224264 271662
rect 224224 267572 224276 267578
rect 224224 267514 224276 267520
rect 223488 267164 223540 267170
rect 223488 267106 223540 267112
rect 224224 266416 224276 266422
rect 224224 266358 224276 266364
rect 223040 264302 223422 264330
rect 224236 264316 224264 266358
rect 224972 264330 225000 273958
rect 225512 272536 225564 272542
rect 225512 272478 225564 272484
rect 225524 264330 225552 272478
rect 226628 269686 226656 277780
rect 227824 277394 227852 277780
rect 227732 277366 227852 277394
rect 228836 277766 229034 277794
rect 230230 277766 230428 277794
rect 227260 269816 227312 269822
rect 227260 269758 227312 269764
rect 226616 269680 226668 269686
rect 226616 269622 226668 269628
rect 226708 266552 226760 266558
rect 226708 266494 226760 266500
rect 224972 264302 225078 264330
rect 225524 264302 225906 264330
rect 226720 264316 226748 266494
rect 227272 264330 227300 269758
rect 227732 268802 227760 277366
rect 228836 271318 228864 277766
rect 227904 271312 227956 271318
rect 227904 271254 227956 271260
rect 228824 271312 228876 271318
rect 228824 271254 228876 271260
rect 227720 268796 227772 268802
rect 227720 268738 227772 268744
rect 227916 264330 227944 271254
rect 229560 271176 229612 271182
rect 229560 271118 229612 271124
rect 229192 267572 229244 267578
rect 229192 267514 229244 267520
rect 227272 264302 227562 264330
rect 227916 264302 228390 264330
rect 229204 264316 229232 267514
rect 229572 264330 229600 271118
rect 230400 270502 230428 277766
rect 231412 271182 231440 277780
rect 232516 275738 232544 277780
rect 232504 275732 232556 275738
rect 232504 275674 232556 275680
rect 232688 275324 232740 275330
rect 232688 275266 232740 275272
rect 231400 271176 231452 271182
rect 231400 271118 231452 271124
rect 230388 270496 230440 270502
rect 230388 270438 230440 270444
rect 230848 270088 230900 270094
rect 230848 270030 230900 270036
rect 229572 264302 230046 264330
rect 230860 264316 230888 270030
rect 232504 269952 232556 269958
rect 232504 269894 232556 269900
rect 231676 268388 231728 268394
rect 231676 268330 231728 268336
rect 231688 264316 231716 268330
rect 232516 264316 232544 269894
rect 232700 267442 232728 275266
rect 233240 272672 233292 272678
rect 233240 272614 233292 272620
rect 232688 267436 232740 267442
rect 232688 267378 232740 267384
rect 233252 264330 233280 272614
rect 233712 270094 233740 277780
rect 234908 277394 234936 277780
rect 234816 277366 234936 277394
rect 234620 274236 234672 274242
rect 234620 274178 234672 274184
rect 233700 270088 233752 270094
rect 233700 270030 233752 270036
rect 234160 267300 234212 267306
rect 234160 267242 234212 267248
rect 233252 264302 233358 264330
rect 234172 264316 234200 267242
rect 234632 265946 234660 274178
rect 234816 269958 234844 277366
rect 236104 272542 236132 277780
rect 236092 272536 236144 272542
rect 236092 272478 236144 272484
rect 234988 271448 235040 271454
rect 234988 271390 235040 271396
rect 234804 269952 234856 269958
rect 234804 269894 234856 269900
rect 234620 265940 234672 265946
rect 234620 265882 234672 265888
rect 235000 264316 235028 271390
rect 237300 271318 237328 277780
rect 238510 277766 238708 277794
rect 236828 271312 236880 271318
rect 236828 271254 236880 271260
rect 237288 271312 237340 271318
rect 237288 271254 237340 271260
rect 236644 268524 236696 268530
rect 236644 268466 236696 268472
rect 235540 265940 235592 265946
rect 235540 265882 235592 265888
rect 235552 264330 235580 265882
rect 235552 264302 235842 264330
rect 236656 264316 236684 268466
rect 236840 267306 236868 271254
rect 237472 270224 237524 270230
rect 237472 270166 237524 270172
rect 236828 267300 236880 267306
rect 236828 267242 236880 267248
rect 237484 264316 237512 270166
rect 238300 268660 238352 268666
rect 238300 268602 238352 268608
rect 238312 264316 238340 268602
rect 238680 268394 238708 277766
rect 239404 275460 239456 275466
rect 239404 275402 239456 275408
rect 239220 272808 239272 272814
rect 239220 272750 239272 272756
rect 238668 268388 238720 268394
rect 238668 268330 238720 268336
rect 239232 267734 239260 272750
rect 239416 267734 239444 275402
rect 239600 272678 239628 277780
rect 240810 277766 241468 277794
rect 240416 274508 240468 274514
rect 240416 274450 240468 274456
rect 239588 272672 239640 272678
rect 239588 272614 239640 272620
rect 239232 267706 239352 267734
rect 239416 267706 239536 267734
rect 239128 267436 239180 267442
rect 239128 267378 239180 267384
rect 239140 264316 239168 267378
rect 239324 264466 239352 267706
rect 239508 266422 239536 267706
rect 239496 266416 239548 266422
rect 239496 266358 239548 266364
rect 239324 264438 239536 264466
rect 239508 264330 239536 264438
rect 240428 264330 240456 274450
rect 241440 268530 241468 277766
rect 241992 277394 242020 277780
rect 241900 277366 242020 277394
rect 241900 271454 241928 277366
rect 243188 274718 243216 277780
rect 244384 275602 244412 277780
rect 245580 277394 245608 277780
rect 245488 277366 245608 277394
rect 243544 275596 243596 275602
rect 243544 275538 243596 275544
rect 244372 275596 244424 275602
rect 244372 275538 244424 275544
rect 243176 274712 243228 274718
rect 243176 274654 243228 274660
rect 242992 272944 243044 272950
rect 242992 272886 243044 272892
rect 242072 271584 242124 271590
rect 242072 271526 242124 271532
rect 241888 271448 241940 271454
rect 241888 271390 241940 271396
rect 241428 268524 241480 268530
rect 241428 268466 241480 268472
rect 241612 267164 241664 267170
rect 241612 267106 241664 267112
rect 239508 264302 239982 264330
rect 240428 264302 240810 264330
rect 241624 264316 241652 267106
rect 242084 264330 242112 271526
rect 242716 270088 242768 270094
rect 242716 270030 242768 270036
rect 242728 267170 242756 270030
rect 242716 267164 242768 267170
rect 242716 267106 242768 267112
rect 243004 264330 243032 272886
rect 243556 266898 243584 275538
rect 244924 270360 244976 270366
rect 244924 270302 244976 270308
rect 243544 266892 243596 266898
rect 243544 266834 243596 266840
rect 244096 266416 244148 266422
rect 244096 266358 244148 266364
rect 242084 264302 242466 264330
rect 243004 264302 243294 264330
rect 244108 264316 244136 266358
rect 244936 264316 244964 270302
rect 245488 270094 245516 277366
rect 245660 275732 245712 275738
rect 245660 275674 245712 275680
rect 245672 274242 245700 275674
rect 246776 275330 246804 277780
rect 247894 277766 248368 277794
rect 247040 275596 247092 275602
rect 247040 275538 247092 275544
rect 246764 275324 246816 275330
rect 246764 275266 246816 275272
rect 245660 274236 245712 274242
rect 245660 274178 245712 274184
rect 245752 274100 245804 274106
rect 245752 274042 245804 274048
rect 245476 270088 245528 270094
rect 245476 270030 245528 270036
rect 245764 264316 245792 274042
rect 247052 273970 247080 275538
rect 248340 274666 248368 277766
rect 249076 275806 249104 277780
rect 249064 275800 249116 275806
rect 249064 275742 249116 275748
rect 249064 274712 249116 274718
rect 248340 274638 248460 274666
rect 249064 274654 249116 274660
rect 247040 273964 247092 273970
rect 247040 273906 247092 273912
rect 247040 273828 247092 273834
rect 247040 273770 247092 273776
rect 246580 267028 246632 267034
rect 246580 266970 246632 266976
rect 246592 264316 246620 266970
rect 247052 264330 247080 273770
rect 247776 271720 247828 271726
rect 247776 271662 247828 271668
rect 247788 264330 247816 271662
rect 248432 271590 248460 274638
rect 248420 271584 248472 271590
rect 248420 271526 248472 271532
rect 249076 267034 249104 274654
rect 250272 269822 250300 277780
rect 249892 269816 249944 269822
rect 249892 269758 249944 269764
rect 250260 269816 250312 269822
rect 250260 269758 250312 269764
rect 249064 267028 249116 267034
rect 249064 266970 249116 266976
rect 249064 266892 249116 266898
rect 249064 266834 249116 266840
rect 247052 264302 247434 264330
rect 247788 264302 248262 264330
rect 249076 264316 249104 266834
rect 249904 264316 249932 269758
rect 251468 269278 251496 277780
rect 252664 272814 252692 277780
rect 253676 277766 253874 277794
rect 253480 275800 253532 275806
rect 253480 275742 253532 275748
rect 253492 274106 253520 275742
rect 253676 275466 253704 277766
rect 253664 275460 253716 275466
rect 253664 275402 253716 275408
rect 254032 274236 254084 274242
rect 254032 274178 254084 274184
rect 253480 274100 253532 274106
rect 253480 274042 253532 274048
rect 252652 272808 252704 272814
rect 252652 272750 252704 272756
rect 253204 272536 253256 272542
rect 253204 272478 253256 272484
rect 252744 271176 252796 271182
rect 252744 271118 252796 271124
rect 252100 270496 252152 270502
rect 252100 270438 252152 270444
rect 251456 269272 251508 269278
rect 251456 269214 251508 269220
rect 250720 268796 250772 268802
rect 250720 268738 250772 268744
rect 250732 264316 250760 268738
rect 251548 267300 251600 267306
rect 251548 267242 251600 267248
rect 251560 264316 251588 267242
rect 252112 264330 252140 270438
rect 252756 264330 252784 271118
rect 253216 266558 253244 272478
rect 253204 266552 253256 266558
rect 253204 266494 253256 266500
rect 252112 264302 252402 264330
rect 252756 264302 253230 264330
rect 254044 264316 254072 274178
rect 254584 272672 254636 272678
rect 254584 272614 254636 272620
rect 254596 266898 254624 272614
rect 255056 272542 255084 277780
rect 256174 277766 256556 277794
rect 255044 272536 255096 272542
rect 255044 272478 255096 272484
rect 255688 269952 255740 269958
rect 255688 269894 255740 269900
rect 254860 267164 254912 267170
rect 254860 267106 254912 267112
rect 254584 266892 254636 266898
rect 254584 266834 254636 266840
rect 254872 264316 254900 267106
rect 255700 264316 255728 269894
rect 256528 268394 256556 277766
rect 256700 275324 256752 275330
rect 256700 275266 256752 275272
rect 256712 268666 256740 275266
rect 257356 274854 257384 277780
rect 257344 274848 257396 274854
rect 257344 274790 257396 274796
rect 256976 271312 257028 271318
rect 256976 271254 257028 271260
rect 256700 268660 256752 268666
rect 256700 268602 256752 268608
rect 256700 268524 256752 268530
rect 256700 268466 256752 268472
rect 256148 268388 256200 268394
rect 256148 268330 256200 268336
rect 256516 268388 256568 268394
rect 256516 268330 256568 268336
rect 256160 266422 256188 268330
rect 256712 266558 256740 268466
rect 256516 266552 256568 266558
rect 256516 266494 256568 266500
rect 256700 266552 256752 266558
rect 256700 266494 256752 266500
rect 256148 266416 256200 266422
rect 256148 266358 256200 266364
rect 256528 264316 256556 266494
rect 256988 264330 257016 271254
rect 258552 270230 258580 277780
rect 259748 275670 259776 277780
rect 259736 275664 259788 275670
rect 259736 275606 259788 275612
rect 260944 275330 260972 277780
rect 262140 277394 262168 277780
rect 262048 277366 262168 277394
rect 261484 275460 261536 275466
rect 261484 275402 261536 275408
rect 260932 275324 260984 275330
rect 260932 275266 260984 275272
rect 259920 274848 259972 274854
rect 259920 274790 259972 274796
rect 259932 271318 259960 274790
rect 260288 271448 260340 271454
rect 260288 271390 260340 271396
rect 259920 271312 259972 271318
rect 259920 271254 259972 271260
rect 258540 270224 258592 270230
rect 258540 270166 258592 270172
rect 258080 269272 258132 269278
rect 258080 269214 258132 269220
rect 258092 266694 258120 269214
rect 259000 266892 259052 266898
rect 259000 266834 259052 266840
rect 258080 266688 258132 266694
rect 258080 266630 258132 266636
rect 258172 266416 258224 266422
rect 258172 266358 258224 266364
rect 256988 264302 257370 264330
rect 258184 264316 258212 266358
rect 259012 264316 259040 266834
rect 259828 266552 259880 266558
rect 259828 266494 259880 266500
rect 259840 264316 259868 266494
rect 260300 264330 260328 271390
rect 261496 267442 261524 275402
rect 262048 269958 262076 277366
rect 262220 273964 262272 273970
rect 262220 273906 262272 273912
rect 262036 269952 262088 269958
rect 262036 269894 262088 269900
rect 261484 267436 261536 267442
rect 261484 267378 261536 267384
rect 261484 267028 261536 267034
rect 261484 266970 261536 266976
rect 260300 264302 260682 264330
rect 261496 264316 261524 266970
rect 262232 264330 262260 273906
rect 263244 271182 263272 277780
rect 264454 277766 264836 277794
rect 264336 271584 264388 271590
rect 264336 271526 264388 271532
rect 263232 271176 263284 271182
rect 263232 271118 263284 271124
rect 263140 270088 263192 270094
rect 263140 270030 263192 270036
rect 262232 264302 262338 264330
rect 263152 264316 263180 270030
rect 263968 268660 264020 268666
rect 263968 268602 264020 268608
rect 263980 264316 264008 268602
rect 264348 264330 264376 271526
rect 264808 267734 264836 277766
rect 265256 274100 265308 274106
rect 265256 274042 265308 274048
rect 264808 267706 265020 267734
rect 264992 267034 265020 267706
rect 264980 267028 265032 267034
rect 264980 266970 265032 266976
rect 265268 264330 265296 274042
rect 265636 273970 265664 277780
rect 265624 273964 265676 273970
rect 265624 273906 265676 273912
rect 266832 270094 266860 277780
rect 268042 277766 268240 277794
rect 267004 275664 267056 275670
rect 267004 275606 267056 275612
rect 266820 270088 266872 270094
rect 266820 270030 266872 270036
rect 266452 269816 266504 269822
rect 266452 269758 266504 269764
rect 264348 264302 264822 264330
rect 265268 264302 265650 264330
rect 266464 264316 266492 269758
rect 267016 267170 267044 275606
rect 267832 272808 267884 272814
rect 267832 272750 267884 272756
rect 267004 267164 267056 267170
rect 267004 267106 267056 267112
rect 267280 266688 267332 266694
rect 267280 266630 267332 266636
rect 267292 264316 267320 266630
rect 267844 264330 267872 272750
rect 268016 270224 268068 270230
rect 268016 270166 268068 270172
rect 268028 266422 268056 270166
rect 268212 269822 268240 277766
rect 269224 277394 269252 277780
rect 269132 277366 269252 277394
rect 270236 277766 270434 277794
rect 268200 269816 268252 269822
rect 268200 269758 268252 269764
rect 269132 268530 269160 277366
rect 270236 272542 270264 277766
rect 269304 272536 269356 272542
rect 269304 272478 269356 272484
rect 270224 272536 270276 272542
rect 270224 272478 270276 272484
rect 269120 268524 269172 268530
rect 269120 268466 269172 268472
rect 268936 267436 268988 267442
rect 268936 267378 268988 267384
rect 268016 266416 268068 266422
rect 268016 266358 268068 266364
rect 267844 264302 268134 264330
rect 268948 264316 268976 267378
rect 269316 264330 269344 272478
rect 271524 271318 271552 277780
rect 272734 277766 273116 277794
rect 270960 271312 271012 271318
rect 270960 271254 271012 271260
rect 271512 271312 271564 271318
rect 271512 271254 271564 271260
rect 270592 268388 270644 268394
rect 270592 268330 270644 268336
rect 269316 264302 269790 264330
rect 270604 264316 270632 268330
rect 270972 264330 271000 271254
rect 273088 269958 273116 277766
rect 273916 275330 273944 277780
rect 273536 275324 273588 275330
rect 273536 275266 273588 275272
rect 273904 275324 273956 275330
rect 273904 275266 273956 275272
rect 272524 269952 272576 269958
rect 272524 269894 272576 269900
rect 273076 269952 273128 269958
rect 273076 269894 273128 269900
rect 272536 266422 272564 269894
rect 273076 267164 273128 267170
rect 273076 267106 273128 267112
rect 272248 266416 272300 266422
rect 272248 266358 272300 266364
rect 272524 266416 272576 266422
rect 272524 266358 272576 266364
rect 270972 264302 271446 264330
rect 272260 264316 272288 266358
rect 273088 264316 273116 267106
rect 273548 264330 273576 275266
rect 275112 270502 275140 277780
rect 276308 271862 276336 277780
rect 277504 275806 277532 277780
rect 277492 275800 277544 275806
rect 277492 275742 277544 275748
rect 276848 273964 276900 273970
rect 276848 273906 276900 273912
rect 276296 271856 276348 271862
rect 276296 271798 276348 271804
rect 275284 271176 275336 271182
rect 275284 271118 275336 271124
rect 275100 270496 275152 270502
rect 275100 270438 275152 270444
rect 274640 270088 274692 270094
rect 274640 270030 274692 270036
rect 274652 266898 274680 270030
rect 274640 266892 274692 266898
rect 274640 266834 274692 266840
rect 274732 266416 274784 266422
rect 274732 266358 274784 266364
rect 273548 264302 273930 264330
rect 274744 264316 274772 266358
rect 275296 264330 275324 271118
rect 276020 270496 276072 270502
rect 276020 270438 276072 270444
rect 276032 267170 276060 270438
rect 276020 267164 276072 267170
rect 276020 267106 276072 267112
rect 276388 267028 276440 267034
rect 276388 266970 276440 266976
rect 275296 264302 275586 264330
rect 276400 264316 276428 266970
rect 276860 264330 276888 273906
rect 278044 271856 278096 271862
rect 278044 271798 278096 271804
rect 278056 267034 278084 271798
rect 278700 270502 278728 277780
rect 279804 271182 279832 277780
rect 281000 272678 281028 277780
rect 282210 277766 282868 277794
rect 280988 272672 281040 272678
rect 280988 272614 281040 272620
rect 280344 272536 280396 272542
rect 280344 272478 280396 272484
rect 279792 271176 279844 271182
rect 279792 271118 279844 271124
rect 278688 270496 278740 270502
rect 278688 270438 278740 270444
rect 278872 269816 278924 269822
rect 278872 269758 278924 269764
rect 278044 267028 278096 267034
rect 278044 266970 278096 266976
rect 278044 266892 278096 266898
rect 278044 266834 278096 266840
rect 276860 264302 277242 264330
rect 278056 264316 278084 266834
rect 278884 264316 278912 269758
rect 279700 268524 279752 268530
rect 279700 268466 279752 268472
rect 279712 264316 279740 268466
rect 280356 264330 280384 272478
rect 280896 271312 280948 271318
rect 280896 271254 280948 271260
rect 280908 264330 280936 271254
rect 282184 269952 282236 269958
rect 282184 269894 282236 269900
rect 280356 264302 280554 264330
rect 280908 264302 281382 264330
rect 282196 264316 282224 269894
rect 282840 269142 282868 277766
rect 283392 275602 283420 277780
rect 283380 275596 283432 275602
rect 283380 275538 283432 275544
rect 284588 275466 284616 277780
rect 285128 275800 285180 275806
rect 285128 275742 285180 275748
rect 284576 275460 284628 275466
rect 284576 275402 284628 275408
rect 283288 275324 283340 275330
rect 283288 275266 283340 275272
rect 282828 269136 282880 269142
rect 282828 269078 282880 269084
rect 283300 264330 283328 275266
rect 283840 267164 283892 267170
rect 283840 267106 283892 267112
rect 283038 264302 283328 264330
rect 283852 264316 283880 267106
rect 284668 267028 284720 267034
rect 284668 266970 284720 266976
rect 284680 264316 284708 266970
rect 285140 264330 285168 275742
rect 285784 269958 285812 277780
rect 286888 272950 286916 277780
rect 286876 272944 286928 272950
rect 286876 272886 286928 272892
rect 287704 272944 287756 272950
rect 287704 272886 287756 272892
rect 286324 272672 286376 272678
rect 286324 272614 286376 272620
rect 285956 270496 286008 270502
rect 285956 270438 286008 270444
rect 285772 269952 285824 269958
rect 285772 269894 285824 269900
rect 285968 264330 285996 270438
rect 286336 267306 286364 272614
rect 287152 271176 287204 271182
rect 287152 271118 287204 271124
rect 286324 267300 286376 267306
rect 286324 267242 286376 267248
rect 285140 264302 285522 264330
rect 285968 264302 286350 264330
rect 287164 264316 287192 271118
rect 287716 266422 287744 272886
rect 288084 271862 288112 277780
rect 289084 275596 289136 275602
rect 289084 275538 289136 275544
rect 288072 271856 288124 271862
rect 288072 271798 288124 271804
rect 288808 269136 288860 269142
rect 288808 269078 288860 269084
rect 287980 267300 288032 267306
rect 287980 267242 288032 267248
rect 287704 266416 287756 266422
rect 287704 266358 287756 266364
rect 287992 264316 288020 267242
rect 288820 264316 288848 269078
rect 289096 267734 289124 275538
rect 289280 274718 289308 277780
rect 290096 275460 290148 275466
rect 290096 275402 290148 275408
rect 289268 274712 289320 274718
rect 289268 274654 289320 274660
rect 289096 267706 289216 267734
rect 289188 264330 289216 267706
rect 290108 264330 290136 275402
rect 290476 275058 290504 277780
rect 290464 275052 290516 275058
rect 290464 274994 290516 275000
rect 291672 270502 291700 277780
rect 292882 277766 293264 277794
rect 292764 274712 292816 274718
rect 292764 274654 292816 274660
rect 291660 270496 291712 270502
rect 291660 270438 291712 270444
rect 291292 269952 291344 269958
rect 291292 269894 291344 269900
rect 289188 264302 289662 264330
rect 290108 264302 290490 264330
rect 291304 264316 291332 269894
rect 292120 266416 292172 266422
rect 292120 266358 292172 266364
rect 292132 264316 292160 266358
rect 292776 265946 292804 274654
rect 293236 271862 293264 277766
rect 292948 271856 293000 271862
rect 292948 271798 293000 271804
rect 293224 271856 293276 271862
rect 293224 271798 293276 271804
rect 292764 265940 292816 265946
rect 292764 265882 292816 265888
rect 292960 264316 292988 271798
rect 294064 269278 294092 277780
rect 294328 275052 294380 275058
rect 294328 274994 294380 275000
rect 294052 269272 294104 269278
rect 294052 269214 294104 269220
rect 293500 265940 293552 265946
rect 293500 265882 293552 265888
rect 293512 264330 293540 265882
rect 294340 264330 294368 274994
rect 295168 274666 295196 277780
rect 296364 274718 296392 277780
rect 297574 277766 297956 277794
rect 296352 274712 296404 274718
rect 295168 274638 295380 274666
rect 296352 274654 296404 274660
rect 295352 269142 295380 274638
rect 295800 271856 295852 271862
rect 295800 271798 295852 271804
rect 295524 270496 295576 270502
rect 295524 270438 295576 270444
rect 295340 269136 295392 269142
rect 295340 269078 295392 269084
rect 295536 267734 295564 270438
rect 295444 267706 295564 267734
rect 293512 264302 293802 264330
rect 294340 264302 294630 264330
rect 295444 264316 295472 267706
rect 295812 264330 295840 271798
rect 297928 270502 297956 277766
rect 298756 274718 298784 277780
rect 298376 274712 298428 274718
rect 298376 274654 298428 274660
rect 298744 274712 298796 274718
rect 298744 274654 298796 274660
rect 297916 270496 297968 270502
rect 297916 270438 297968 270444
rect 297088 269272 297140 269278
rect 297088 269214 297140 269220
rect 295812 264302 296286 264330
rect 297100 264316 297128 269214
rect 297916 269136 297968 269142
rect 297916 269078 297968 269084
rect 297928 264316 297956 269078
rect 298388 264330 298416 274654
rect 299952 270502 299980 277780
rect 301148 277394 301176 277780
rect 301056 277366 301176 277394
rect 302344 277394 302372 277780
rect 302344 277366 302464 277394
rect 300124 274712 300176 274718
rect 300124 274654 300176 274660
rect 299572 270496 299624 270502
rect 299572 270438 299624 270444
rect 299940 270496 299992 270502
rect 299940 270438 299992 270444
rect 298388 264302 298770 264330
rect 299584 264316 299612 270438
rect 300136 264330 300164 274654
rect 300860 270496 300912 270502
rect 300860 270438 300912 270444
rect 300872 264330 300900 270438
rect 301056 266422 301084 277366
rect 301044 266416 301096 266422
rect 301044 266358 301096 266364
rect 302056 266416 302108 266422
rect 302056 266358 302108 266364
rect 300136 264302 300426 264330
rect 300872 264302 301254 264330
rect 302068 264316 302096 266358
rect 302436 264330 302464 277366
rect 303448 270450 303476 277780
rect 304092 277766 304658 277794
rect 305012 277766 305854 277794
rect 306392 277766 307050 277794
rect 307772 277766 308246 277794
rect 303448 270422 303660 270450
rect 303632 264330 303660 270422
rect 304092 264330 304120 277766
rect 305012 264330 305040 277766
rect 306392 266370 306420 277766
rect 307772 267734 307800 277766
rect 309428 277394 309456 277780
rect 310546 277766 310928 277794
rect 309428 277366 309548 277394
rect 306208 266342 306420 266370
rect 307496 267706 307800 267734
rect 302436 264302 302910 264330
rect 303632 264302 303738 264330
rect 304092 264302 304566 264330
rect 305012 264302 305394 264330
rect 306208 264316 306236 266342
rect 307496 264330 307524 267706
rect 308680 266552 308732 266558
rect 308680 266494 308732 266500
rect 307852 266416 307904 266422
rect 307852 266358 307904 266364
rect 307050 264302 307524 264330
rect 307864 264316 307892 266358
rect 308692 264316 308720 266494
rect 309520 266422 309548 277366
rect 309784 270156 309836 270162
rect 309784 270098 309836 270104
rect 309508 266416 309560 266422
rect 309508 266358 309560 266364
rect 309796 264330 309824 270098
rect 310900 266558 310928 277766
rect 311360 277766 311742 277794
rect 311912 277766 312938 277794
rect 313292 277766 314134 277794
rect 314672 277766 315330 277794
rect 311360 270162 311388 277766
rect 311348 270156 311400 270162
rect 311348 270098 311400 270104
rect 310888 266552 310940 266558
rect 310888 266494 310940 266500
rect 311164 266552 311216 266558
rect 311164 266494 311216 266500
rect 310336 266416 310388 266422
rect 310336 266358 310388 266364
rect 309534 264302 309824 264330
rect 310348 264316 310376 266358
rect 311176 264316 311204 266494
rect 311912 266422 311940 277766
rect 312820 266688 312872 266694
rect 312820 266630 312872 266636
rect 311900 266416 311952 266422
rect 311900 266358 311952 266364
rect 312360 266416 312412 266422
rect 312360 266358 312412 266364
rect 312372 264330 312400 266358
rect 312018 264302 312400 264330
rect 312832 264316 312860 266630
rect 313292 266558 313320 277766
rect 314476 269816 314528 269822
rect 314476 269758 314528 269764
rect 313648 267300 313700 267306
rect 313648 267242 313700 267248
rect 313280 266552 313332 266558
rect 313280 266494 313332 266500
rect 313660 264316 313688 267242
rect 314488 264316 314516 269758
rect 314672 266422 314700 277766
rect 316512 277394 316540 277780
rect 316420 277366 316540 277394
rect 317432 277766 317722 277794
rect 318826 277766 319024 277794
rect 315764 271312 315816 271318
rect 315764 271254 315816 271260
rect 314660 266416 314712 266422
rect 314660 266358 314712 266364
rect 315776 264330 315804 271254
rect 316420 266694 316448 277366
rect 316960 270088 317012 270094
rect 316960 270030 317012 270036
rect 316408 266688 316460 266694
rect 316408 266630 316460 266636
rect 316132 266416 316184 266422
rect 316132 266358 316184 266364
rect 315330 264302 315804 264330
rect 316144 264316 316172 266358
rect 316972 264316 317000 270030
rect 317432 267306 317460 277766
rect 318616 271788 318668 271794
rect 318616 271730 318668 271736
rect 317420 267300 317472 267306
rect 317420 267242 317472 267248
rect 317788 266892 317840 266898
rect 317788 266834 317840 266840
rect 317800 264316 317828 266834
rect 318628 264316 318656 271730
rect 318996 269822 319024 277766
rect 320008 271318 320036 277780
rect 320560 277766 321218 277794
rect 321572 277766 322414 277794
rect 322952 277766 323610 277794
rect 319996 271312 320048 271318
rect 319996 271254 320048 271260
rect 318984 269816 319036 269822
rect 318984 269758 319036 269764
rect 319444 269136 319496 269142
rect 319444 269078 319496 269084
rect 319456 264316 319484 269078
rect 320272 266552 320324 266558
rect 320272 266494 320324 266500
rect 320284 264316 320312 266494
rect 320560 266422 320588 277766
rect 321100 270224 321152 270230
rect 321100 270166 321152 270172
rect 320548 266416 320600 266422
rect 320548 266358 320600 266364
rect 321112 264316 321140 270166
rect 321572 270094 321600 277766
rect 322756 273964 322808 273970
rect 322756 273906 322808 273912
rect 321560 270088 321612 270094
rect 321560 270030 321612 270036
rect 321928 266756 321980 266762
rect 321928 266698 321980 266704
rect 321940 264316 321968 266698
rect 322768 264316 322796 273906
rect 322952 266898 322980 277766
rect 324792 271794 324820 277780
rect 325712 277766 326002 277794
rect 324964 274712 325016 274718
rect 324964 274654 325016 274660
rect 324780 271788 324832 271794
rect 324780 271730 324832 271736
rect 323584 270088 323636 270094
rect 323584 270030 323636 270036
rect 322940 266892 322992 266898
rect 322940 266834 322992 266840
rect 323596 264316 323624 270030
rect 324412 267164 324464 267170
rect 324412 267106 324464 267112
rect 324424 264316 324452 267106
rect 324976 266558 325004 274654
rect 325516 271176 325568 271182
rect 325516 271118 325568 271124
rect 324964 266552 325016 266558
rect 324964 266494 325016 266500
rect 325528 264330 325556 271118
rect 325712 269142 325740 277766
rect 327092 274718 327120 277780
rect 327460 277766 328302 277794
rect 328472 277766 329498 277794
rect 327080 274712 327132 274718
rect 327080 274654 327132 274660
rect 327080 270496 327132 270502
rect 327080 270438 327132 270444
rect 326896 269816 326948 269822
rect 326896 269758 326948 269764
rect 325700 269136 325752 269142
rect 325700 269078 325752 269084
rect 326068 268660 326120 268666
rect 326068 268602 326120 268608
rect 325266 264302 325556 264330
rect 326080 264316 326108 268602
rect 326908 264316 326936 269758
rect 327092 266762 327120 270438
rect 327460 270230 327488 277766
rect 328276 275324 328328 275330
rect 328276 275266 328328 275272
rect 327448 270224 327500 270230
rect 327448 270166 327500 270172
rect 328288 268666 328316 275266
rect 328472 270502 328500 277766
rect 330680 273970 330708 277780
rect 331232 277766 331890 277794
rect 330668 273964 330720 273970
rect 330668 273906 330720 273912
rect 330484 273284 330536 273290
rect 330484 273226 330536 273232
rect 329748 271312 329800 271318
rect 329748 271254 329800 271260
rect 328460 270496 328512 270502
rect 328460 270438 328512 270444
rect 329380 269952 329432 269958
rect 329380 269894 329432 269900
rect 328276 268660 328328 268666
rect 328276 268602 328328 268608
rect 327724 268388 327776 268394
rect 327724 268330 327776 268336
rect 327080 266756 327132 266762
rect 327080 266698 327132 266704
rect 327736 264316 327764 268330
rect 328552 266416 328604 266422
rect 328552 266358 328604 266364
rect 328564 264316 328592 266358
rect 329392 264316 329420 269894
rect 329760 266422 329788 271254
rect 330496 267170 330524 273226
rect 331036 272536 331088 272542
rect 331036 272478 331088 272484
rect 330484 267164 330536 267170
rect 330484 267106 330536 267112
rect 330208 266552 330260 266558
rect 330208 266494 330260 266500
rect 329748 266416 329800 266422
rect 329748 266358 329800 266364
rect 330220 264316 330248 266494
rect 331048 264316 331076 272478
rect 331232 270094 331260 277766
rect 333072 273290 333100 277780
rect 333796 273964 333848 273970
rect 333796 273906 333848 273912
rect 333060 273284 333112 273290
rect 333060 273226 333112 273232
rect 331220 270088 331272 270094
rect 331220 270030 331272 270036
rect 331864 269136 331916 269142
rect 331864 269078 331916 269084
rect 331876 264316 331904 269078
rect 333520 267028 333572 267034
rect 333520 266970 333572 266976
rect 332692 266416 332744 266422
rect 332692 266358 332744 266364
rect 332704 264316 332732 266358
rect 333532 264316 333560 266970
rect 333808 266422 333836 273906
rect 334176 271182 334204 277780
rect 335372 275330 335400 277780
rect 335556 277766 336582 277794
rect 336752 277766 337778 277794
rect 335360 275324 335412 275330
rect 335360 275266 335412 275272
rect 334624 271448 334676 271454
rect 334624 271390 334676 271396
rect 334164 271176 334216 271182
rect 334164 271118 334216 271124
rect 334348 267164 334400 267170
rect 334348 267106 334400 267112
rect 333796 266416 333848 266422
rect 333796 266358 333848 266364
rect 334360 264316 334388 267106
rect 334636 266558 334664 271390
rect 335556 269822 335584 277766
rect 336004 270360 336056 270366
rect 336004 270302 336056 270308
rect 335544 269816 335596 269822
rect 335544 269758 335596 269764
rect 335176 267300 335228 267306
rect 335176 267242 335228 267248
rect 334624 266552 334676 266558
rect 334624 266494 334676 266500
rect 335188 264316 335216 267242
rect 336016 264316 336044 270302
rect 336752 268394 336780 277766
rect 338028 274712 338080 274718
rect 338028 274654 338080 274660
rect 336924 269816 336976 269822
rect 336924 269758 336976 269764
rect 336740 268388 336792 268394
rect 336740 268330 336792 268336
rect 336936 267734 336964 269758
rect 338040 269142 338068 274654
rect 338960 271318 338988 277780
rect 339512 277766 340170 277794
rect 339132 274100 339184 274106
rect 339132 274042 339184 274048
rect 338948 271312 339000 271318
rect 338948 271254 339000 271260
rect 338028 269136 338080 269142
rect 338028 269078 338080 269084
rect 337660 268388 337712 268394
rect 337660 268330 337712 268336
rect 336844 267706 336964 267734
rect 336844 264316 336872 267706
rect 337672 264316 337700 268330
rect 339144 267734 339172 274042
rect 339316 271176 339368 271182
rect 339316 271118 339368 271124
rect 338960 267706 339172 267734
rect 338960 264330 338988 267706
rect 338514 264302 338988 264330
rect 339328 264316 339356 271118
rect 339512 269958 339540 277766
rect 340604 271584 340656 271590
rect 340604 271526 340656 271532
rect 339500 269952 339552 269958
rect 339500 269894 339552 269900
rect 340616 264330 340644 271526
rect 341352 271454 341380 277780
rect 342456 272542 342484 277780
rect 343652 274718 343680 277780
rect 343640 274712 343692 274718
rect 343640 274654 343692 274660
rect 344284 274712 344336 274718
rect 344284 274654 344336 274660
rect 343548 272808 343600 272814
rect 343548 272750 343600 272756
rect 342444 272536 342496 272542
rect 342444 272478 342496 272484
rect 341340 271448 341392 271454
rect 341340 271390 341392 271396
rect 341524 271312 341576 271318
rect 341524 271254 341576 271260
rect 340972 267436 341024 267442
rect 340972 267378 341024 267384
rect 340170 264302 340644 264330
rect 340984 264316 341012 267378
rect 341536 267306 341564 271254
rect 341800 269952 341852 269958
rect 341800 269894 341852 269900
rect 341524 267300 341576 267306
rect 341524 267242 341576 267248
rect 341812 264316 341840 269894
rect 342260 269136 342312 269142
rect 342260 269078 342312 269084
rect 342272 267034 342300 269078
rect 343364 268524 343416 268530
rect 343364 268466 343416 268472
rect 342260 267028 342312 267034
rect 342260 266970 342312 266976
rect 342628 266416 342680 266422
rect 342628 266358 342680 266364
rect 342640 264316 342668 266358
rect 343376 264330 343404 268466
rect 343560 266422 343588 272750
rect 344296 267170 344324 274654
rect 344848 273970 344876 277780
rect 345124 277766 346058 277794
rect 344836 273964 344888 273970
rect 344836 273906 344888 273912
rect 344652 273828 344704 273834
rect 344652 273770 344704 273776
rect 344284 267164 344336 267170
rect 344284 267106 344336 267112
rect 343548 266416 343600 266422
rect 343548 266358 343600 266364
rect 344664 264330 344692 273770
rect 345124 269142 345152 277766
rect 347044 275324 347096 275330
rect 347044 275266 347096 275272
rect 345940 270224 345992 270230
rect 345940 270166 345992 270172
rect 345112 269136 345164 269142
rect 345112 269078 345164 269084
rect 345112 266552 345164 266558
rect 345112 266494 345164 266500
rect 343376 264302 343482 264330
rect 344310 264302 344692 264330
rect 345124 264316 345152 266494
rect 345952 264316 345980 270166
rect 346768 270088 346820 270094
rect 346768 270030 346820 270036
rect 346780 264316 346808 270030
rect 347056 267442 347084 275266
rect 347240 274718 347268 277780
rect 347228 274712 347280 274718
rect 347228 274654 347280 274660
rect 347412 274712 347464 274718
rect 347412 274654 347464 274660
rect 347424 270366 347452 274654
rect 348436 271318 348464 277780
rect 349632 274718 349660 277780
rect 350552 277766 350750 277794
rect 351946 277766 352144 277794
rect 349804 275460 349856 275466
rect 349804 275402 349856 275408
rect 349620 274712 349672 274718
rect 349620 274654 349672 274660
rect 349816 273834 349844 275402
rect 349804 273828 349856 273834
rect 349804 273770 349856 273776
rect 350356 273828 350408 273834
rect 350356 273770 350408 273776
rect 349804 272672 349856 272678
rect 349804 272614 349856 272620
rect 348884 271448 348936 271454
rect 348884 271390 348936 271396
rect 348424 271312 348476 271318
rect 348424 271254 348476 271260
rect 347412 270360 347464 270366
rect 347412 270302 347464 270308
rect 347044 267436 347096 267442
rect 347044 267378 347096 267384
rect 347596 266416 347648 266422
rect 347596 266358 347648 266364
rect 347608 264316 347636 266358
rect 348896 264330 348924 271390
rect 349252 266892 349304 266898
rect 349252 266834 349304 266840
rect 348450 264302 348924 264330
rect 349264 264316 349292 266834
rect 349816 266422 349844 272614
rect 349804 266416 349856 266422
rect 349804 266358 349856 266364
rect 350368 264330 350396 273770
rect 350552 269822 350580 277766
rect 351184 274236 351236 274242
rect 351184 274178 351236 274184
rect 350540 269816 350592 269822
rect 350540 269758 350592 269764
rect 350908 267436 350960 267442
rect 350908 267378 350960 267384
rect 350106 264302 350396 264330
rect 350920 264316 350948 267378
rect 351196 266558 351224 274178
rect 351736 269816 351788 269822
rect 351736 269758 351788 269764
rect 351184 266552 351236 266558
rect 351184 266494 351236 266500
rect 351748 264316 351776 269758
rect 352116 268394 352144 277766
rect 353128 274106 353156 277780
rect 353116 274100 353168 274106
rect 353116 274042 353168 274048
rect 354324 271182 354352 277780
rect 355152 277766 355534 277794
rect 355152 271590 355180 277766
rect 356716 275330 356744 277780
rect 357452 277766 357926 277794
rect 356704 275324 356756 275330
rect 356704 275266 356756 275272
rect 357256 274848 357308 274854
rect 357256 274790 357308 274796
rect 356888 272536 356940 272542
rect 356888 272478 356940 272484
rect 355140 271584 355192 271590
rect 355140 271526 355192 271532
rect 355324 271584 355376 271590
rect 355324 271526 355376 271532
rect 354588 271312 354640 271318
rect 354588 271254 354640 271260
rect 354312 271176 354364 271182
rect 354312 271118 354364 271124
rect 352104 268388 352156 268394
rect 352104 268330 352156 268336
rect 352564 268388 352616 268394
rect 352564 268330 352616 268336
rect 352576 264316 352604 268330
rect 353392 267164 353444 267170
rect 353392 267106 353444 267112
rect 353404 264316 353432 267106
rect 354600 264330 354628 271254
rect 355336 266898 355364 271526
rect 355876 268660 355928 268666
rect 355876 268602 355928 268608
rect 355324 266892 355376 266898
rect 355324 266834 355376 266840
rect 355048 266416 355100 266422
rect 355048 266358 355100 266364
rect 354246 264302 354628 264330
rect 355060 264316 355088 266358
rect 355888 264316 355916 268602
rect 356704 266892 356756 266898
rect 356704 266834 356756 266840
rect 356716 264316 356744 266834
rect 356900 266422 356928 272478
rect 357268 268530 357296 274790
rect 357452 269958 357480 277766
rect 359016 272814 359044 277780
rect 359464 275324 359516 275330
rect 359464 275266 359516 275272
rect 359004 272808 359056 272814
rect 359004 272750 359056 272756
rect 359188 270360 359240 270366
rect 359188 270302 359240 270308
rect 357440 269952 357492 269958
rect 357440 269894 357492 269900
rect 357256 268524 357308 268530
rect 357256 268466 357308 268472
rect 357532 268524 357584 268530
rect 357532 268466 357584 268472
rect 356888 266416 356940 266422
rect 356888 266358 356940 266364
rect 357544 264316 357572 268466
rect 358360 266416 358412 266422
rect 358360 266358 358412 266364
rect 358372 264316 358400 266358
rect 359200 264316 359228 270302
rect 359476 267442 359504 275266
rect 360212 274854 360240 277780
rect 361408 275466 361436 277780
rect 361396 275460 361448 275466
rect 361396 275402 361448 275408
rect 360200 274848 360252 274854
rect 360200 274790 360252 274796
rect 360200 274712 360252 274718
rect 360200 274654 360252 274660
rect 360212 270502 360240 274654
rect 362604 274242 362632 277780
rect 362960 275460 363012 275466
rect 362960 275402 363012 275408
rect 362592 274236 362644 274242
rect 362592 274178 362644 274184
rect 362776 274100 362828 274106
rect 362776 274042 362828 274048
rect 360844 272808 360896 272814
rect 360844 272750 360896 272756
rect 360200 270496 360252 270502
rect 360200 270438 360252 270444
rect 360200 270224 360252 270230
rect 360200 270166 360252 270172
rect 360212 267734 360240 270166
rect 360028 267706 360240 267734
rect 359464 267436 359516 267442
rect 359464 267378 359516 267384
rect 360028 264316 360056 267706
rect 360856 266422 360884 272750
rect 362788 271266 362816 274042
rect 362972 271454 363000 275402
rect 363800 274718 363828 277780
rect 364352 277766 365010 277794
rect 363788 274712 363840 274718
rect 363788 274654 363840 274660
rect 363604 271720 363656 271726
rect 363604 271662 363656 271668
rect 362960 271448 363012 271454
rect 362960 271390 363012 271396
rect 362788 271238 362908 271266
rect 362684 271176 362736 271182
rect 362684 271118 362736 271124
rect 361120 267436 361172 267442
rect 361120 267378 361172 267384
rect 360844 266416 360896 266422
rect 360844 266358 360896 266364
rect 361132 264330 361160 267378
rect 361672 266416 361724 266422
rect 361672 266358 361724 266364
rect 360870 264302 361160 264330
rect 361684 264316 361712 266358
rect 362696 264330 362724 271118
rect 362880 266422 362908 271238
rect 363328 267300 363380 267306
rect 363328 267242 363380 267248
rect 362868 266416 362920 266422
rect 362868 266358 362920 266364
rect 362526 264302 362724 264330
rect 363340 264316 363368 267242
rect 363616 267170 363644 271662
rect 364352 270094 364380 277766
rect 366100 272678 366128 277780
rect 367296 275466 367324 277780
rect 367836 275596 367888 275602
rect 367836 275538 367888 275544
rect 367284 275460 367336 275466
rect 367284 275402 367336 275408
rect 366364 275052 366416 275058
rect 366364 274994 366416 275000
rect 366376 273970 366404 274994
rect 366364 273964 366416 273970
rect 366364 273906 366416 273912
rect 367008 273964 367060 273970
rect 367008 273906 367060 273912
rect 366088 272672 366140 272678
rect 366088 272614 366140 272620
rect 366364 271448 366416 271454
rect 366364 271390 366416 271396
rect 364340 270088 364392 270094
rect 364340 270030 364392 270036
rect 364984 270088 365036 270094
rect 364984 270030 365036 270036
rect 364156 269952 364208 269958
rect 364156 269894 364208 269900
rect 363604 267164 363656 267170
rect 363604 267106 363656 267112
rect 364168 264316 364196 269894
rect 364996 264316 365024 270030
rect 365812 267164 365864 267170
rect 365812 267106 365864 267112
rect 365824 264316 365852 267106
rect 366376 266898 366404 271390
rect 366364 266892 366416 266898
rect 366364 266834 366416 266840
rect 367020 264330 367048 273906
rect 367848 268666 367876 275538
rect 368296 274372 368348 274378
rect 368296 274314 368348 274320
rect 367836 268660 367888 268666
rect 367836 268602 367888 268608
rect 368112 267028 368164 267034
rect 368112 266970 368164 266976
rect 367468 266416 367520 266422
rect 367468 266358 367520 266364
rect 366666 264302 367048 264330
rect 367480 264316 367508 266358
rect 368124 264330 368152 266970
rect 368308 266422 368336 274314
rect 368492 271590 368520 277780
rect 368848 275868 368900 275874
rect 368848 275810 368900 275816
rect 368480 271584 368532 271590
rect 368480 271526 368532 271532
rect 368860 268394 368888 275810
rect 369688 275058 369716 277780
rect 370884 275330 370912 277780
rect 371252 277766 372094 277794
rect 370872 275324 370924 275330
rect 370872 275266 370924 275272
rect 369676 275052 369728 275058
rect 369676 274994 369728 275000
rect 369860 274848 369912 274854
rect 369860 274790 369912 274796
rect 369492 271584 369544 271590
rect 369492 271526 369544 271532
rect 368848 268388 368900 268394
rect 368848 268330 368900 268336
rect 368296 266416 368348 266422
rect 368296 266358 368348 266364
rect 369504 264330 369532 271526
rect 369872 271318 369900 274790
rect 370964 272672 371016 272678
rect 370964 272614 371016 272620
rect 369860 271312 369912 271318
rect 369860 271254 369912 271260
rect 369952 268388 370004 268394
rect 369952 268330 370004 268336
rect 368124 264302 368322 264330
rect 369150 264302 369532 264330
rect 369964 264316 369992 268330
rect 370976 264330 371004 272614
rect 371252 269822 371280 277766
rect 373276 275874 373304 277780
rect 373264 275868 373316 275874
rect 373264 275810 373316 275816
rect 373264 275732 373316 275738
rect 373264 275674 373316 275680
rect 372528 271312 372580 271318
rect 372528 271254 372580 271260
rect 371240 269816 371292 269822
rect 371240 269758 371292 269764
rect 372344 268796 372396 268802
rect 372344 268738 372396 268744
rect 371608 266416 371660 266422
rect 371608 266358 371660 266364
rect 370806 264302 371004 264330
rect 371620 264316 371648 266358
rect 372356 264330 372384 268738
rect 372540 266422 372568 271254
rect 373276 267734 373304 275674
rect 374380 271726 374408 277780
rect 375576 274854 375604 277780
rect 376772 277394 376800 277780
rect 376772 277366 376892 277394
rect 376668 275460 376720 275466
rect 376668 275402 376720 275408
rect 375564 274848 375616 274854
rect 375564 274790 375616 274796
rect 376680 273970 376708 275402
rect 376668 273964 376720 273970
rect 376668 273906 376720 273912
rect 376576 273828 376628 273834
rect 376576 273770 376628 273776
rect 375288 271856 375340 271862
rect 375288 271798 375340 271804
rect 374368 271720 374420 271726
rect 374368 271662 374420 271668
rect 374920 269816 374972 269822
rect 374920 269758 374972 269764
rect 373092 267706 373304 267734
rect 373092 267442 373120 267706
rect 373264 267572 373316 267578
rect 373264 267514 373316 267520
rect 373080 267436 373132 267442
rect 373080 267378 373132 267384
rect 372528 266416 372580 266422
rect 372528 266358 372580 266364
rect 372356 264302 372462 264330
rect 373276 264316 373304 267514
rect 374092 266416 374144 266422
rect 374092 266358 374144 266364
rect 374104 264316 374132 266358
rect 374932 264316 374960 269758
rect 375300 266422 375328 271798
rect 375748 267436 375800 267442
rect 375748 267378 375800 267384
rect 375288 266416 375340 266422
rect 375288 266358 375340 266364
rect 375760 264316 375788 267378
rect 376588 264316 376616 273770
rect 376864 272542 376892 277366
rect 377968 275602 377996 277780
rect 377956 275596 378008 275602
rect 377956 275538 378008 275544
rect 377404 275324 377456 275330
rect 377404 275266 377456 275272
rect 376852 272536 376904 272542
rect 376852 272478 376904 272484
rect 377416 271590 377444 275266
rect 378784 274508 378836 274514
rect 378784 274450 378836 274456
rect 377404 271584 377456 271590
rect 377404 271526 377456 271532
rect 377036 270496 377088 270502
rect 377036 270438 377088 270444
rect 377048 267306 377076 270438
rect 377772 267708 377824 267714
rect 377772 267650 377824 267656
rect 377036 267300 377088 267306
rect 377036 267242 377088 267248
rect 377784 267034 377812 267650
rect 377772 267028 377824 267034
rect 377772 266970 377824 266976
rect 378796 266422 378824 274450
rect 379164 271454 379192 277780
rect 379532 277766 380374 277794
rect 379336 271584 379388 271590
rect 379336 271526 379388 271532
rect 379152 271448 379204 271454
rect 379152 271390 379204 271396
rect 378968 267028 379020 267034
rect 378968 266970 379020 266976
rect 377404 266416 377456 266422
rect 377404 266358 377456 266364
rect 378784 266416 378836 266422
rect 378784 266358 378836 266364
rect 377416 264316 377444 266358
rect 378980 264466 379008 266970
rect 378704 264438 379008 264466
rect 378704 264330 378732 264438
rect 379348 264330 379376 271526
rect 379532 268530 379560 277766
rect 381556 272814 381584 277780
rect 382292 277766 382674 277794
rect 383672 277766 383870 277794
rect 382004 273080 382056 273086
rect 382004 273022 382056 273028
rect 381544 272808 381596 272814
rect 381544 272750 381596 272756
rect 380808 272536 380860 272542
rect 380808 272478 380860 272484
rect 379520 268524 379572 268530
rect 379520 268466 379572 268472
rect 380624 266892 380676 266898
rect 380624 266834 380676 266840
rect 379888 266416 379940 266422
rect 379888 266358 379940 266364
rect 378258 264302 378732 264330
rect 379086 264302 379376 264330
rect 379900 264316 379928 266358
rect 380636 264330 380664 266834
rect 380820 266422 380848 272478
rect 380808 266416 380860 266422
rect 380808 266358 380860 266364
rect 382016 264330 382044 273022
rect 382292 270366 382320 277766
rect 382464 275596 382516 275602
rect 382464 275538 382516 275544
rect 382476 271318 382504 275538
rect 382464 271312 382516 271318
rect 382464 271254 382516 271260
rect 383384 271312 383436 271318
rect 383384 271254 383436 271260
rect 382280 270360 382332 270366
rect 382280 270302 382332 270308
rect 382372 268660 382424 268666
rect 382372 268602 382424 268608
rect 380636 264302 380742 264330
rect 381570 264302 382044 264330
rect 382384 264316 382412 268602
rect 383396 264330 383424 271254
rect 383672 270230 383700 277766
rect 385052 275738 385080 277780
rect 385040 275732 385092 275738
rect 385040 275674 385092 275680
rect 384948 274644 385000 274650
rect 384948 274586 385000 274592
rect 384764 271720 384816 271726
rect 384764 271662 384816 271668
rect 383660 270224 383712 270230
rect 383660 270166 383712 270172
rect 383660 269544 383712 269550
rect 383660 269486 383712 269492
rect 383672 266762 383700 269486
rect 383660 266756 383712 266762
rect 383660 266698 383712 266704
rect 384028 266416 384080 266422
rect 384028 266358 384080 266364
rect 383226 264302 383424 264330
rect 384040 264316 384068 266358
rect 384776 264330 384804 271662
rect 384960 266422 384988 274586
rect 386248 274242 386276 277780
rect 387168 277766 387458 277794
rect 387904 277766 388654 277794
rect 389192 277766 389758 277794
rect 390572 277766 390954 277794
rect 391952 277766 392150 277794
rect 386236 274236 386288 274242
rect 386236 274178 386288 274184
rect 385684 274100 385736 274106
rect 385684 274042 385736 274048
rect 385696 267714 385724 274042
rect 387168 271182 387196 277766
rect 387708 274780 387760 274786
rect 387708 274722 387760 274728
rect 387720 274378 387748 274722
rect 387708 274372 387760 274378
rect 387708 274314 387760 274320
rect 387616 271448 387668 271454
rect 387616 271390 387668 271396
rect 387156 271176 387208 271182
rect 387156 271118 387208 271124
rect 387432 269680 387484 269686
rect 387432 269622 387484 269628
rect 385684 267708 385736 267714
rect 385684 267650 385736 267656
rect 387248 267708 387300 267714
rect 387248 267650 387300 267656
rect 385684 267164 385736 267170
rect 385684 267106 385736 267112
rect 384948 266416 385000 266422
rect 384948 266358 385000 266364
rect 384776 264302 384882 264330
rect 385696 264316 385724 267106
rect 386512 266416 386564 266422
rect 386512 266358 386564 266364
rect 386524 264316 386552 266358
rect 387260 264330 387288 267650
rect 387444 267578 387472 269622
rect 387432 267572 387484 267578
rect 387432 267514 387484 267520
rect 387628 266422 387656 271390
rect 387904 270502 387932 277766
rect 388812 272944 388864 272950
rect 388812 272886 388864 272892
rect 387892 270496 387944 270502
rect 387892 270438 387944 270444
rect 388168 270224 388220 270230
rect 388168 270166 388220 270172
rect 387616 266416 387668 266422
rect 387616 266358 387668 266364
rect 387260 264302 387366 264330
rect 388180 264316 388208 270166
rect 388824 264330 388852 272886
rect 389192 269958 389220 277766
rect 390376 270360 390428 270366
rect 390376 270302 390428 270308
rect 389180 269952 389232 269958
rect 389180 269894 389232 269900
rect 390192 269952 390244 269958
rect 390192 269894 390244 269900
rect 390204 266898 390232 269894
rect 390388 267442 390416 270302
rect 390572 270094 390600 277766
rect 391756 271176 391808 271182
rect 391756 271118 391808 271124
rect 390560 270088 390612 270094
rect 390560 270030 390612 270036
rect 390376 267436 390428 267442
rect 390376 267378 390428 267384
rect 390652 267436 390704 267442
rect 390652 267378 390704 267384
rect 390192 266892 390244 266898
rect 390192 266834 390244 266840
rect 389824 266688 389876 266694
rect 389824 266630 389876 266636
rect 388824 264302 389022 264330
rect 389836 264316 389864 266630
rect 390664 264316 390692 267378
rect 391768 264330 391796 271118
rect 391952 269550 391980 277766
rect 393332 275466 393360 277780
rect 393780 275868 393832 275874
rect 393780 275810 393832 275816
rect 393320 275460 393372 275466
rect 393320 275402 393372 275408
rect 393792 271590 393820 275810
rect 394528 274786 394556 277780
rect 395172 277766 395738 277794
rect 394516 274780 394568 274786
rect 394516 274722 394568 274728
rect 395172 274106 395200 277766
rect 395436 275460 395488 275466
rect 395436 275402 395488 275408
rect 395160 274100 395212 274106
rect 395160 274042 395212 274048
rect 394332 272808 394384 272814
rect 394332 272750 394384 272756
rect 393780 271584 393832 271590
rect 393780 271526 393832 271532
rect 391940 269544 391992 269550
rect 391940 269486 391992 269492
rect 392124 269544 392176 269550
rect 392124 269486 392176 269492
rect 392136 267034 392164 269486
rect 393136 268524 393188 268530
rect 393136 268466 393188 268472
rect 392124 267028 392176 267034
rect 392124 266970 392176 266976
rect 392308 267028 392360 267034
rect 392308 266970 392360 266976
rect 391506 264302 391796 264330
rect 392320 264316 392348 266970
rect 393148 264316 393176 268466
rect 394344 264330 394372 272750
rect 395448 271862 395476 275402
rect 396920 275330 396948 277780
rect 397472 277766 398038 277794
rect 396908 275324 396960 275330
rect 396908 275266 396960 275272
rect 397092 274780 397144 274786
rect 397092 274722 397144 274728
rect 395620 274100 395672 274106
rect 395620 274042 395672 274048
rect 395436 271856 395488 271862
rect 395436 271798 395488 271804
rect 395632 271674 395660 274042
rect 395356 271646 395660 271674
rect 394792 267300 394844 267306
rect 394792 267242 394844 267248
rect 393990 264302 394372 264330
rect 394804 264316 394832 267242
rect 395356 266694 395384 271646
rect 395528 271584 395580 271590
rect 395528 271526 395580 271532
rect 395540 267442 395568 271526
rect 397104 268802 397132 274722
rect 397276 274372 397328 274378
rect 397276 274314 397328 274320
rect 397092 268796 397144 268802
rect 397092 268738 397144 268744
rect 395528 267436 395580 267442
rect 395528 267378 395580 267384
rect 397092 267436 397144 267442
rect 397092 267378 397144 267384
rect 395344 266688 395396 266694
rect 395344 266630 395396 266636
rect 395620 266552 395672 266558
rect 395620 266494 395672 266500
rect 395632 264316 395660 266494
rect 396448 266416 396500 266422
rect 396448 266358 396500 266364
rect 396460 264316 396488 266358
rect 397104 264330 397132 267378
rect 397288 266422 397316 274314
rect 397472 268394 397500 277766
rect 399220 272678 399248 277780
rect 400220 275732 400272 275738
rect 400220 275674 400272 275680
rect 400232 274650 400260 275674
rect 400416 275602 400444 277780
rect 400404 275596 400456 275602
rect 400404 275538 400456 275544
rect 400404 275324 400456 275330
rect 400404 275266 400456 275272
rect 400220 274644 400272 274650
rect 400220 274586 400272 274592
rect 400128 274508 400180 274514
rect 400128 274450 400180 274456
rect 399208 272672 399260 272678
rect 399208 272614 399260 272620
rect 398748 268796 398800 268802
rect 398748 268738 398800 268744
rect 397460 268388 397512 268394
rect 397460 268330 397512 268336
rect 398760 267714 398788 268738
rect 399760 268388 399812 268394
rect 399760 268330 399812 268336
rect 398748 267708 398800 267714
rect 398748 267650 398800 267656
rect 398104 266756 398156 266762
rect 398104 266698 398156 266704
rect 397276 266416 397328 266422
rect 397276 266358 397328 266364
rect 397104 264302 397302 264330
rect 398116 264316 398144 266698
rect 398932 266416 398984 266422
rect 398932 266358 398984 266364
rect 398944 264316 398972 266358
rect 399772 264316 399800 268330
rect 400140 266422 400168 274450
rect 400416 272950 400444 275266
rect 401612 274802 401640 277780
rect 401980 277766 402822 277794
rect 401980 277394 402008 277766
rect 401520 274786 401640 274802
rect 401508 274780 401640 274786
rect 401560 274774 401640 274780
rect 401704 277366 402008 277394
rect 401508 274722 401560 274728
rect 401508 273216 401560 273222
rect 401508 273158 401560 273164
rect 400404 272944 400456 272950
rect 400404 272886 400456 272892
rect 400588 270496 400640 270502
rect 400588 270438 400640 270444
rect 400128 266416 400180 266422
rect 400128 266358 400180 266364
rect 400600 264316 400628 270438
rect 401520 267734 401548 273158
rect 401704 269686 401732 277366
rect 403440 275596 403492 275602
rect 403440 275538 403492 275544
rect 403452 271182 403480 275538
rect 404004 275466 404032 277780
rect 404372 277766 405214 277794
rect 405752 277766 406318 277794
rect 403992 275460 404044 275466
rect 403992 275402 404044 275408
rect 403992 274644 404044 274650
rect 403992 274586 404044 274592
rect 403440 271176 403492 271182
rect 403440 271118 403492 271124
rect 401692 269680 401744 269686
rect 401692 269622 401744 269628
rect 401876 269680 401928 269686
rect 401876 269622 401928 269628
rect 401428 267706 401548 267734
rect 401428 264316 401456 267706
rect 401888 267170 401916 269622
rect 404004 267734 404032 274586
rect 404176 270768 404228 270774
rect 404176 270710 404228 270716
rect 403912 267706 404032 267734
rect 402244 267572 402296 267578
rect 402244 267514 402296 267520
rect 401876 267164 401928 267170
rect 401876 267106 401928 267112
rect 402256 264316 402284 267514
rect 403072 266416 403124 266422
rect 403072 266358 403124 266364
rect 403084 264316 403112 266358
rect 403912 264316 403940 267706
rect 404188 266422 404216 270710
rect 404372 269822 404400 277766
rect 405004 271176 405056 271182
rect 405004 271118 405056 271124
rect 404360 269816 404412 269822
rect 404360 269758 404412 269764
rect 404728 267708 404780 267714
rect 404728 267650 404780 267656
rect 404176 266416 404228 266422
rect 404176 266358 404228 266364
rect 404740 264316 404768 267650
rect 405016 266558 405044 271118
rect 405752 270366 405780 277766
rect 407500 273970 407528 277780
rect 407764 275460 407816 275466
rect 407764 275402 407816 275408
rect 407488 273964 407540 273970
rect 407488 273906 407540 273912
rect 406844 272944 406896 272950
rect 406844 272886 406896 272892
rect 405740 270360 405792 270366
rect 405740 270302 405792 270308
rect 405556 266892 405608 266898
rect 405556 266834 405608 266840
rect 405004 266552 405056 266558
rect 405004 266494 405056 266500
rect 405568 264316 405596 266834
rect 406856 264330 406884 272886
rect 407776 272814 407804 275402
rect 408696 274242 408724 277780
rect 408684 274236 408736 274242
rect 408684 274178 408736 274184
rect 409236 273964 409288 273970
rect 409236 273906 409288 273912
rect 407764 272808 407816 272814
rect 407764 272750 407816 272756
rect 408408 272808 408460 272814
rect 408408 272750 408460 272756
rect 407212 270360 407264 270366
rect 407212 270302 407264 270308
rect 406410 264302 406884 264330
rect 407224 264316 407252 270302
rect 408420 264330 408448 272750
rect 409248 264330 409276 273906
rect 409696 270088 409748 270094
rect 409696 270030 409748 270036
rect 408066 264302 408448 264330
rect 408894 264302 409276 264330
rect 409708 264316 409736 270030
rect 409892 269550 409920 277780
rect 410064 276004 410116 276010
rect 410064 275946 410116 275952
rect 410076 270230 410104 275946
rect 411088 275874 411116 277780
rect 412008 277766 412298 277794
rect 412652 277766 413402 277794
rect 411076 275868 411128 275874
rect 411076 275810 411128 275816
rect 412008 272542 412036 277766
rect 412272 272672 412324 272678
rect 412272 272614 412324 272620
rect 411996 272536 412048 272542
rect 411996 272478 412048 272484
rect 410064 270224 410116 270230
rect 410064 270166 410116 270172
rect 410800 270224 410852 270230
rect 410800 270166 410852 270172
rect 409880 269544 409932 269550
rect 409880 269486 409932 269492
rect 410812 264330 410840 270166
rect 412284 266422 412312 272614
rect 412652 269958 412680 277766
rect 414584 273086 414612 277780
rect 415412 277766 415794 277794
rect 415216 274780 415268 274786
rect 415216 274722 415268 274728
rect 414572 273080 414624 273086
rect 414572 273022 414624 273028
rect 413928 272536 413980 272542
rect 413928 272478 413980 272484
rect 412640 269952 412692 269958
rect 412640 269894 412692 269900
rect 412456 269816 412508 269822
rect 412456 269758 412508 269764
rect 411352 266416 411404 266422
rect 411352 266358 411404 266364
rect 412272 266416 412324 266422
rect 412272 266358 412324 266364
rect 410550 264302 410840 264330
rect 411364 264316 411392 266358
rect 412468 264330 412496 269758
rect 413008 269068 413060 269074
rect 413008 269010 413060 269016
rect 412206 264302 412496 264330
rect 413020 264316 413048 269010
rect 413940 267734 413968 272478
rect 415228 271726 415256 274722
rect 415216 271720 415268 271726
rect 415216 271662 415268 271668
rect 414480 270632 414532 270638
rect 414480 270574 414532 270580
rect 413848 267706 413968 267734
rect 413848 264316 413876 267706
rect 414492 266762 414520 270574
rect 414664 269952 414716 269958
rect 414664 269894 414716 269900
rect 414480 266756 414532 266762
rect 414480 266698 414532 266704
rect 414676 264316 414704 269894
rect 415412 268666 415440 277766
rect 416976 271318 417004 277780
rect 418172 275738 418200 277780
rect 418160 275732 418212 275738
rect 418160 275674 418212 275680
rect 418344 275732 418396 275738
rect 418344 275674 418396 275680
rect 418356 274378 418384 275674
rect 419368 274786 419396 277780
rect 419736 277766 420578 277794
rect 419540 276004 419592 276010
rect 419540 275946 419592 275952
rect 419356 274780 419408 274786
rect 419356 274722 419408 274728
rect 419552 274514 419580 275946
rect 419540 274508 419592 274514
rect 419540 274450 419592 274456
rect 418344 274372 418396 274378
rect 418344 274314 418396 274320
rect 419172 274372 419224 274378
rect 419172 274314 419224 274320
rect 418804 271720 418856 271726
rect 418804 271662 418856 271668
rect 416964 271312 417016 271318
rect 416964 271254 417016 271260
rect 418068 270904 418120 270910
rect 418068 270846 418120 270852
rect 415400 268660 415452 268666
rect 415400 268602 415452 268608
rect 416688 268660 416740 268666
rect 416688 268602 416740 268608
rect 416700 267306 416728 268602
rect 418080 267734 418108 270846
rect 417988 267706 418108 267734
rect 416688 267300 416740 267306
rect 416688 267242 416740 267248
rect 415492 267164 415544 267170
rect 415492 267106 415544 267112
rect 415504 264316 415532 267106
rect 416320 266620 416372 266626
rect 416320 266562 416372 266568
rect 416332 264316 416360 266562
rect 417148 266416 417200 266422
rect 417148 266358 417200 266364
rect 417160 264316 417188 266358
rect 417988 264316 418016 267706
rect 418816 267034 418844 271662
rect 418804 267028 418856 267034
rect 418804 266970 418856 266976
rect 419184 264330 419212 274314
rect 419736 269686 419764 277766
rect 420736 274508 420788 274514
rect 420736 274450 420788 274456
rect 419724 269680 419776 269686
rect 419724 269622 419776 269628
rect 419816 269408 419868 269414
rect 419816 269350 419868 269356
rect 419632 267300 419684 267306
rect 419632 267242 419684 267248
rect 418830 264302 419212 264330
rect 419644 264316 419672 267242
rect 419828 266422 419856 269350
rect 419816 266416 419868 266422
rect 419816 266358 419868 266364
rect 420748 264330 420776 274450
rect 421668 271454 421696 277780
rect 422312 277766 422878 277794
rect 421656 271448 421708 271454
rect 421656 271390 421708 271396
rect 421564 271312 421616 271318
rect 421564 271254 421616 271260
rect 421576 267442 421604 271254
rect 422116 269680 422168 269686
rect 422116 269622 422168 269628
rect 421564 267436 421616 267442
rect 421564 267378 421616 267384
rect 421288 266484 421340 266490
rect 421288 266426 421340 266432
rect 420486 264302 420776 264330
rect 421300 264316 421328 266426
rect 422128 264316 422156 269622
rect 422312 268802 422340 277766
rect 424060 275874 424088 277780
rect 424048 275868 424100 275874
rect 424048 275810 424100 275816
rect 425256 275330 425284 277780
rect 425244 275324 425296 275330
rect 425244 275266 425296 275272
rect 426256 275052 426308 275058
rect 426256 274994 426308 275000
rect 424968 272264 425020 272270
rect 424968 272206 425020 272212
rect 424600 269544 424652 269550
rect 424600 269486 424652 269492
rect 422300 268796 422352 268802
rect 422300 268738 422352 268744
rect 422300 268116 422352 268122
rect 422300 268058 422352 268064
rect 422312 267578 422340 268058
rect 422300 267572 422352 267578
rect 422300 267514 422352 267520
rect 422944 267028 422996 267034
rect 422944 266970 422996 266976
rect 422956 264316 422984 266970
rect 423772 266756 423824 266762
rect 423772 266698 423824 266704
rect 423784 264316 423812 266698
rect 424612 264316 424640 269486
rect 424980 266762 425008 272206
rect 425704 271448 425756 271454
rect 425704 271390 425756 271396
rect 425716 266898 425744 271390
rect 425704 266892 425756 266898
rect 425704 266834 425756 266840
rect 426072 266892 426124 266898
rect 426072 266834 426124 266840
rect 424968 266756 425020 266762
rect 424968 266698 425020 266704
rect 425428 266756 425480 266762
rect 425428 266698 425480 266704
rect 425440 264316 425468 266698
rect 426084 264330 426112 266834
rect 426268 266762 426296 274994
rect 426452 274106 426480 277780
rect 427452 274236 427504 274242
rect 427452 274178 427504 274184
rect 426440 274100 426492 274106
rect 426440 274042 426492 274048
rect 426256 266756 426308 266762
rect 426256 266698 426308 266704
rect 427464 264330 427492 274178
rect 427648 271590 427676 277780
rect 428844 275602 428872 277780
rect 429672 277766 429962 277794
rect 430592 277766 431158 277794
rect 428832 275596 428884 275602
rect 428832 275538 428884 275544
rect 427820 275324 427872 275330
rect 427820 275266 427872 275272
rect 427832 273222 427860 275266
rect 428924 275188 428976 275194
rect 428924 275130 428976 275136
rect 427820 273216 427872 273222
rect 427820 273158 427872 273164
rect 427636 271584 427688 271590
rect 427636 271526 427688 271532
rect 428740 268932 428792 268938
rect 428740 268874 428792 268880
rect 427912 266756 427964 266762
rect 427912 266698 427964 266704
rect 426084 264302 426282 264330
rect 427110 264302 427492 264330
rect 427924 264316 427952 266698
rect 428752 264316 428780 268874
rect 428936 266762 428964 275130
rect 429672 271726 429700 277766
rect 429844 273080 429896 273086
rect 429844 273022 429896 273028
rect 429660 271720 429712 271726
rect 429660 271662 429712 271668
rect 429568 268252 429620 268258
rect 429568 268194 429620 268200
rect 428924 266756 428976 266762
rect 428924 266698 428976 266704
rect 429580 264316 429608 268194
rect 429856 267714 429884 273022
rect 430592 268530 430620 277766
rect 432340 275466 432368 277780
rect 433352 277766 433550 277794
rect 432788 275868 432840 275874
rect 432788 275810 432840 275816
rect 432328 275460 432380 275466
rect 432328 275402 432380 275408
rect 431684 273828 431736 273834
rect 431684 273770 431736 273776
rect 430580 268524 430632 268530
rect 430580 268466 430632 268472
rect 429844 267708 429896 267714
rect 429844 267650 429896 267656
rect 430396 267572 430448 267578
rect 430396 267514 430448 267520
rect 430408 264316 430436 267514
rect 431696 264330 431724 273770
rect 432052 266416 432104 266422
rect 432052 266358 432104 266364
rect 431250 264302 431724 264330
rect 432064 264316 432092 266358
rect 432800 264330 432828 275810
rect 432972 271448 433024 271454
rect 432972 271390 433024 271396
rect 432984 270638 433012 271390
rect 432972 270632 433024 270638
rect 432972 270574 433024 270580
rect 433156 270632 433208 270638
rect 433156 270574 433208 270580
rect 433168 266422 433196 270574
rect 433352 268666 433380 277766
rect 434444 271856 434496 271862
rect 434444 271798 434496 271804
rect 433708 268796 433760 268802
rect 433708 268738 433760 268744
rect 433340 268660 433392 268666
rect 433340 268602 433392 268608
rect 433156 266416 433208 266422
rect 433156 266358 433208 266364
rect 432800 264302 432906 264330
rect 433720 264316 433748 268738
rect 434456 264330 434484 271798
rect 434732 271046 434760 277780
rect 435928 275738 435956 277780
rect 435916 275732 435968 275738
rect 435916 275674 435968 275680
rect 435732 275596 435784 275602
rect 435732 275538 435784 275544
rect 434720 271040 434772 271046
rect 434720 270982 434772 270988
rect 434904 271040 434956 271046
rect 434904 270982 434956 270988
rect 434916 270638 434944 270982
rect 434904 270632 434956 270638
rect 434904 270574 434956 270580
rect 435744 264330 435772 275538
rect 437032 271318 437060 277780
rect 437952 277766 438242 277794
rect 437204 271720 437256 271726
rect 437204 271662 437256 271668
rect 437020 271312 437072 271318
rect 437020 271254 437072 271260
rect 436192 268660 436244 268666
rect 436192 268602 436244 268608
rect 434456 264302 434562 264330
rect 435390 264302 435772 264330
rect 436204 264316 436232 268602
rect 436744 267708 436796 267714
rect 436744 267650 436796 267656
rect 436560 267436 436612 267442
rect 436560 267378 436612 267384
rect 436572 266898 436600 267378
rect 436756 267170 436784 267650
rect 436744 267164 436796 267170
rect 436744 267106 436796 267112
rect 436560 266892 436612 266898
rect 436560 266834 436612 266840
rect 437216 264330 437244 271662
rect 437952 271454 437980 277766
rect 439424 276010 439452 277780
rect 440252 277766 440634 277794
rect 441632 277766 441830 277794
rect 439412 276004 439464 276010
rect 439412 275946 439464 275952
rect 438860 275460 438912 275466
rect 438860 275402 438912 275408
rect 438872 274650 438900 275402
rect 438860 274644 438912 274650
rect 438860 274586 438912 274592
rect 439320 273556 439372 273562
rect 439320 273498 439372 273504
rect 438124 273216 438176 273222
rect 438124 273158 438176 273164
rect 437940 271448 437992 271454
rect 437940 271390 437992 271396
rect 437848 266756 437900 266762
rect 437848 266698 437900 266704
rect 437046 264302 437244 264330
rect 437860 264316 437888 266698
rect 438136 266626 438164 273158
rect 438676 266892 438728 266898
rect 438676 266834 438728 266840
rect 438124 266620 438176 266626
rect 438124 266562 438176 266568
rect 438688 264316 438716 266834
rect 439332 266422 439360 273498
rect 439964 271448 440016 271454
rect 439964 271390 440016 271396
rect 439320 266416 439372 266422
rect 439320 266358 439372 266364
rect 439976 264330 440004 271390
rect 440252 268394 440280 277766
rect 441344 275596 441396 275602
rect 441344 275538 441396 275544
rect 441160 268524 441212 268530
rect 441160 268466 441212 268472
rect 440240 268388 440292 268394
rect 440240 268330 440292 268336
rect 440332 266416 440384 266422
rect 440332 266358 440384 266364
rect 439530 264302 440004 264330
rect 440344 264316 440372 266358
rect 441172 264316 441200 268466
rect 441356 266422 441384 275538
rect 441632 270502 441660 277766
rect 443012 275330 443040 277780
rect 443288 277766 444222 277794
rect 443000 275324 443052 275330
rect 443000 275266 443052 275272
rect 442908 271584 442960 271590
rect 442908 271526 442960 271532
rect 441620 270496 441672 270502
rect 441620 270438 441672 270444
rect 441620 269272 441672 269278
rect 441620 269214 441672 269220
rect 441632 267714 441660 269214
rect 441620 267708 441672 267714
rect 441620 267650 441672 267656
rect 442724 267708 442776 267714
rect 442724 267650 442776 267656
rect 441344 266416 441396 266422
rect 441344 266358 441396 266364
rect 441988 266416 442040 266422
rect 441988 266358 442040 266364
rect 442000 264316 442028 266358
rect 442736 264330 442764 267650
rect 442920 266422 442948 271526
rect 443288 268122 443316 277766
rect 445024 274644 445076 274650
rect 445024 274586 445076 274592
rect 443644 268388 443696 268394
rect 443644 268330 443696 268336
rect 443276 268116 443328 268122
rect 443276 268058 443328 268064
rect 442908 266416 442960 266422
rect 442908 266358 442960 266364
rect 442736 264302 442842 264330
rect 443656 264316 443684 268330
rect 445036 267442 445064 274586
rect 445312 270774 445340 277780
rect 446508 275466 446536 277780
rect 446496 275460 446548 275466
rect 446496 275402 446548 275408
rect 446404 274780 446456 274786
rect 446404 274722 446456 274728
rect 446416 273970 446444 274722
rect 446588 274100 446640 274106
rect 446588 274042 446640 274048
rect 446404 273964 446456 273970
rect 446404 273906 446456 273912
rect 445668 271312 445720 271318
rect 445668 271254 445720 271260
rect 445300 270768 445352 270774
rect 445300 270710 445352 270716
rect 445024 267436 445076 267442
rect 445024 267378 445076 267384
rect 445300 267164 445352 267170
rect 445300 267106 445352 267112
rect 444472 266416 444524 266422
rect 444472 266358 444524 266364
rect 444484 264316 444512 266358
rect 445312 264316 445340 267106
rect 445680 266422 445708 271254
rect 446600 267306 446628 274042
rect 447704 273086 447732 277780
rect 447692 273080 447744 273086
rect 447692 273022 447744 273028
rect 447784 272128 447836 272134
rect 447784 272070 447836 272076
rect 446588 267300 446640 267306
rect 446588 267242 446640 267248
rect 446956 266620 447008 266626
rect 446956 266562 447008 266568
rect 445668 266416 445720 266422
rect 445668 266358 445720 266364
rect 446128 266416 446180 266422
rect 446128 266358 446180 266364
rect 446140 264316 446168 266358
rect 446968 264316 446996 266562
rect 447796 266422 447824 272070
rect 448900 271182 448928 277780
rect 450096 272950 450124 277780
rect 451306 277766 451504 277794
rect 450544 275460 450596 275466
rect 450544 275402 450596 275408
rect 450084 272944 450136 272950
rect 450084 272886 450136 272892
rect 448888 271176 448940 271182
rect 448888 271118 448940 271124
rect 449808 271176 449860 271182
rect 449808 271118 449860 271124
rect 448612 267844 448664 267850
rect 448612 267786 448664 267792
rect 447784 266416 447836 266422
rect 447784 266358 447836 266364
rect 448152 266416 448204 266422
rect 448152 266358 448204 266364
rect 448164 264330 448192 266358
rect 447810 264302 448192 264330
rect 448624 264316 448652 267786
rect 449820 264330 449848 271118
rect 450268 267436 450320 267442
rect 450268 267378 450320 267384
rect 449466 264302 449848 264330
rect 450280 264316 450308 267378
rect 450556 266422 450584 275402
rect 451096 273080 451148 273086
rect 451096 273022 451148 273028
rect 450728 267164 450780 267170
rect 450728 267106 450780 267112
rect 450740 266490 450768 267106
rect 450728 266484 450780 266490
rect 450728 266426 450780 266432
rect 450544 266416 450596 266422
rect 450544 266358 450596 266364
rect 451108 264316 451136 273022
rect 451476 270366 451504 277766
rect 452120 277766 452502 277794
rect 452120 272814 452148 277766
rect 453592 274786 453620 277780
rect 454052 277766 454802 277794
rect 455432 277766 455998 277794
rect 453764 275324 453816 275330
rect 453764 275266 453816 275272
rect 453580 274780 453632 274786
rect 453580 274722 453632 274728
rect 452108 272808 452160 272814
rect 452108 272750 452160 272756
rect 452292 272808 452344 272814
rect 452292 272750 452344 272756
rect 451464 270360 451516 270366
rect 451464 270302 451516 270308
rect 452304 264330 452332 272750
rect 453776 270586 453804 275266
rect 453684 270558 453804 270586
rect 452568 267164 452620 267170
rect 452568 267106 452620 267112
rect 452580 266626 452608 267106
rect 453684 266626 453712 270558
rect 453856 270496 453908 270502
rect 453856 270438 453908 270444
rect 452568 266620 452620 266626
rect 452568 266562 452620 266568
rect 452752 266620 452804 266626
rect 452752 266562 452804 266568
rect 453672 266620 453724 266626
rect 453672 266562 453724 266568
rect 451950 264302 452332 264330
rect 452764 264316 452792 266562
rect 453868 264330 453896 270438
rect 454052 270094 454080 277766
rect 455432 270230 455460 277766
rect 456064 276004 456116 276010
rect 456064 275946 456116 275952
rect 456076 270910 456104 275946
rect 457180 272678 457208 277780
rect 458192 277766 458390 277794
rect 459586 277766 459784 277794
rect 457444 273692 457496 273698
rect 457444 273634 457496 273640
rect 457168 272672 457220 272678
rect 457168 272614 457220 272620
rect 456064 270904 456116 270910
rect 456064 270846 456116 270852
rect 456064 270632 456116 270638
rect 456064 270574 456116 270580
rect 455420 270224 455472 270230
rect 455420 270166 455472 270172
rect 454040 270088 454092 270094
rect 454040 270030 454092 270036
rect 455052 270088 455104 270094
rect 455052 270030 455104 270036
rect 455064 267034 455092 270030
rect 455236 267300 455288 267306
rect 455236 267242 455288 267248
rect 455052 267028 455104 267034
rect 455052 266970 455104 266976
rect 454408 266620 454460 266626
rect 454408 266562 454460 266568
rect 453606 264302 453896 264330
rect 454420 264316 454448 266562
rect 455248 264316 455276 267242
rect 456076 267170 456104 270574
rect 456432 270360 456484 270366
rect 456432 270302 456484 270308
rect 456064 267164 456116 267170
rect 456064 267106 456116 267112
rect 455420 267028 455472 267034
rect 455420 266970 455472 266976
rect 455432 266626 455460 266970
rect 455420 266620 455472 266626
rect 455420 266562 455472 266568
rect 456444 264330 456472 270302
rect 457456 267578 457484 273634
rect 457996 272944 458048 272950
rect 457996 272886 458048 272892
rect 457812 272400 457864 272406
rect 457812 272342 457864 272348
rect 457824 267734 457852 272342
rect 457732 267706 457852 267734
rect 457444 267572 457496 267578
rect 457444 267514 457496 267520
rect 456892 266620 456944 266626
rect 456892 266562 456944 266568
rect 456090 264302 456472 264330
rect 456904 264316 456932 266562
rect 457732 264316 457760 267706
rect 458008 266626 458036 272886
rect 458192 269822 458220 277766
rect 459192 270768 459244 270774
rect 459192 270710 459244 270716
rect 458180 269816 458232 269822
rect 458180 269758 458232 269764
rect 458548 269816 458600 269822
rect 458548 269758 458600 269764
rect 457996 266620 458048 266626
rect 457996 266562 458048 266568
rect 458560 264316 458588 269758
rect 459204 264330 459232 270710
rect 459756 269074 459784 277766
rect 460676 272542 460704 277780
rect 460952 277766 461886 277794
rect 462332 277766 463082 277794
rect 460664 272536 460716 272542
rect 460664 272478 460716 272484
rect 460952 269958 460980 277766
rect 461952 272672 462004 272678
rect 461952 272614 462004 272620
rect 461400 270224 461452 270230
rect 461400 270166 461452 270172
rect 460940 269952 460992 269958
rect 460940 269894 460992 269900
rect 459744 269068 459796 269074
rect 459744 269010 459796 269016
rect 459560 268116 459612 268122
rect 459560 268058 459612 268064
rect 459572 267034 459600 268058
rect 459560 267028 459612 267034
rect 459560 266970 459612 266976
rect 460204 266620 460256 266626
rect 460204 266562 460256 266568
rect 459204 264302 459402 264330
rect 460216 264316 460244 266562
rect 461412 264330 461440 270166
rect 461964 267734 461992 272614
rect 462332 269278 462360 277766
rect 464264 273222 464292 277780
rect 465092 277766 465474 277794
rect 464804 273420 464856 273426
rect 464804 273362 464856 273368
rect 464252 273216 464304 273222
rect 464252 273158 464304 273164
rect 463516 269952 463568 269958
rect 463516 269894 463568 269900
rect 462320 269272 462372 269278
rect 462320 269214 462372 269220
rect 461058 264302 461440 264330
rect 461872 267706 461992 267734
rect 461872 264316 461900 267706
rect 462688 267572 462740 267578
rect 462688 267514 462740 267520
rect 462700 264316 462728 267514
rect 463528 264316 463556 269894
rect 464816 264330 464844 273362
rect 465092 269414 465120 277766
rect 466656 276010 466684 277780
rect 466644 276004 466696 276010
rect 466644 275946 466696 275952
rect 466828 276004 466880 276010
rect 466828 275946 466880 275952
rect 466840 272406 466868 275946
rect 467852 274378 467880 277780
rect 467840 274372 467892 274378
rect 467840 274314 467892 274320
rect 468956 274106 468984 277780
rect 469404 274916 469456 274922
rect 469404 274858 469456 274864
rect 468944 274100 468996 274106
rect 468944 274042 468996 274048
rect 469128 274100 469180 274106
rect 469128 274042 469180 274048
rect 468484 273964 468536 273970
rect 468484 273906 468536 273912
rect 467748 272536 467800 272542
rect 467748 272478 467800 272484
rect 466828 272400 466880 272406
rect 466828 272342 466880 272348
rect 465080 269408 465132 269414
rect 465080 269350 465132 269356
rect 466000 269272 466052 269278
rect 466000 269214 466052 269220
rect 465172 266892 465224 266898
rect 465172 266834 465224 266840
rect 464370 264302 464844 264330
rect 465184 264316 465212 266834
rect 466012 264316 466040 269214
rect 467562 267064 467618 267073
rect 467562 266999 467618 267008
rect 466828 266756 466880 266762
rect 466828 266698 466880 266704
rect 466840 264316 466868 266698
rect 467576 264330 467604 266999
rect 467760 266762 467788 272478
rect 468496 267034 468524 273906
rect 469140 273426 469168 274042
rect 469128 273420 469180 273426
rect 469128 273362 469180 273368
rect 468758 269784 468814 269793
rect 468758 269719 468814 269728
rect 468484 267028 468536 267034
rect 468484 266970 468536 266976
rect 467748 266756 467800 266762
rect 467748 266698 467800 266704
rect 468772 264330 468800 269719
rect 469220 269068 469272 269074
rect 469220 269010 469272 269016
rect 468944 267572 468996 267578
rect 468944 267514 468996 267520
rect 468956 267034 468984 267514
rect 469232 267322 469260 269010
rect 469416 268258 469444 274858
rect 470152 274514 470180 277780
rect 470140 274508 470192 274514
rect 470140 274450 470192 274456
rect 471348 273562 471376 277780
rect 472176 277766 472558 277794
rect 473372 277766 473754 277794
rect 471980 274236 472032 274242
rect 471980 274178 472032 274184
rect 471992 273970 472020 274178
rect 471980 273964 472032 273970
rect 471980 273906 472032 273912
rect 471336 273556 471388 273562
rect 471336 273498 471388 273504
rect 471612 273216 471664 273222
rect 471612 273158 471664 273164
rect 470508 272400 470560 272406
rect 470508 272342 470560 272348
rect 469404 268252 469456 268258
rect 469404 268194 469456 268200
rect 469140 267294 469260 267322
rect 469140 267170 469168 267294
rect 470520 267170 470548 272342
rect 470966 269240 471022 269249
rect 470966 269175 471022 269184
rect 469128 267164 469180 267170
rect 469128 267106 469180 267112
rect 469312 267164 469364 267170
rect 469312 267106 469364 267112
rect 470508 267164 470560 267170
rect 470508 267106 470560 267112
rect 468944 267028 468996 267034
rect 468944 266970 468996 266976
rect 467576 264302 467682 264330
rect 468510 264302 468800 264330
rect 469324 264316 469352 267106
rect 470140 266892 470192 266898
rect 470140 266834 470192 266840
rect 470152 264316 470180 266834
rect 470980 264316 471008 269175
rect 471624 264330 471652 273158
rect 472176 269686 472204 277766
rect 473084 273556 473136 273562
rect 473084 273498 473136 273504
rect 472164 269680 472216 269686
rect 472164 269622 472216 269628
rect 473096 264330 473124 273498
rect 473372 270094 473400 277766
rect 474372 274508 474424 274514
rect 474372 274450 474424 274456
rect 473360 270088 473412 270094
rect 473360 270030 473412 270036
rect 473268 267164 473320 267170
rect 473268 267106 473320 267112
rect 473280 266762 473308 267106
rect 474384 266762 474412 274450
rect 474936 272270 474964 277780
rect 475568 274100 475620 274106
rect 475568 274042 475620 274048
rect 475580 273562 475608 274042
rect 475568 273556 475620 273562
rect 475568 273498 475620 273504
rect 475936 273420 475988 273426
rect 475936 273362 475988 273368
rect 474924 272264 474976 272270
rect 474924 272206 474976 272212
rect 474648 269680 474700 269686
rect 474648 269622 474700 269628
rect 473268 266756 473320 266762
rect 473268 266698 473320 266704
rect 473452 266756 473504 266762
rect 473452 266698 473504 266704
rect 474372 266756 474424 266762
rect 474372 266698 474424 266704
rect 471624 264302 471822 264330
rect 472650 264302 473124 264330
rect 473464 264316 473492 266698
rect 474660 264330 474688 269622
rect 475108 267572 475160 267578
rect 475108 267514 475160 267520
rect 474306 264302 474688 264330
rect 475120 264316 475148 267514
rect 475948 264316 475976 273362
rect 476132 269550 476160 277780
rect 477236 275058 477264 277780
rect 477224 275052 477276 275058
rect 477224 274994 477276 275000
rect 478432 274650 478460 277780
rect 479352 277766 479642 277794
rect 478972 274712 479024 274718
rect 478972 274654 479024 274660
rect 478420 274644 478472 274650
rect 478420 274586 478472 274592
rect 478788 273556 478840 273562
rect 478788 273498 478840 273504
rect 478602 271416 478658 271425
rect 478602 271351 478658 271360
rect 476120 269544 476172 269550
rect 476120 269486 476172 269492
rect 476764 269544 476816 269550
rect 476764 269486 476816 269492
rect 476776 264316 476804 269486
rect 478616 266762 478644 271351
rect 477592 266756 477644 266762
rect 477592 266698 477644 266704
rect 478604 266756 478656 266762
rect 478604 266698 478656 266704
rect 477604 264316 477632 266698
rect 478800 264330 478828 273498
rect 478984 268938 479012 274654
rect 479352 274378 479380 277766
rect 480824 275058 480852 277780
rect 481548 275188 481600 275194
rect 481548 275130 481600 275136
rect 480812 275052 480864 275058
rect 480812 274994 480864 275000
rect 481560 274378 481588 275130
rect 482020 274718 482048 277780
rect 482836 276684 482888 276690
rect 482836 276626 482888 276632
rect 482008 274712 482060 274718
rect 482008 274654 482060 274660
rect 482192 274644 482244 274650
rect 482192 274586 482244 274592
rect 479340 274372 479392 274378
rect 479340 274314 479392 274320
rect 479524 274372 479576 274378
rect 479524 274314 479576 274320
rect 481548 274372 481600 274378
rect 481548 274314 481600 274320
rect 479536 274106 479564 274314
rect 482204 274242 482232 274586
rect 481364 274236 481416 274242
rect 481364 274178 481416 274184
rect 482192 274236 482244 274242
rect 482192 274178 482244 274184
rect 479524 274100 479576 274106
rect 479524 274042 479576 274048
rect 479708 272264 479760 272270
rect 479708 272206 479760 272212
rect 478972 268932 479024 268938
rect 478972 268874 479024 268880
rect 479720 267578 479748 272206
rect 479708 267572 479760 267578
rect 479708 267514 479760 267520
rect 480076 266348 480128 266354
rect 480076 266290 480128 266296
rect 479248 265396 479300 265402
rect 479248 265338 479300 265344
rect 478446 264302 478828 264330
rect 479260 264316 479288 265338
rect 480088 264316 480116 266290
rect 481376 264330 481404 274178
rect 481732 265532 481784 265538
rect 481732 265474 481784 265480
rect 480930 264302 481404 264330
rect 481744 264316 481772 265474
rect 482848 264330 482876 276626
rect 483216 274922 483244 277780
rect 483204 274916 483256 274922
rect 483204 274858 483256 274864
rect 483664 274780 483716 274786
rect 483664 274722 483716 274728
rect 483676 267714 483704 274722
rect 484320 273698 484348 277780
rect 485516 273834 485544 277780
rect 485504 273828 485556 273834
rect 485504 273770 485556 273776
rect 484308 273692 484360 273698
rect 484308 273634 484360 273640
rect 484492 273692 484544 273698
rect 484492 273634 484544 273640
rect 484504 273578 484532 273634
rect 484320 273550 484532 273578
rect 483664 267708 483716 267714
rect 483664 267650 483716 267656
rect 483848 267708 483900 267714
rect 483848 267650 483900 267656
rect 483388 266756 483440 266762
rect 483388 266698 483440 266704
rect 482586 264302 482876 264330
rect 483400 264316 483428 266698
rect 483860 264330 483888 267650
rect 484032 267572 484084 267578
rect 484032 267514 484084 267520
rect 484044 267034 484072 267514
rect 484032 267028 484084 267034
rect 484032 266970 484084 266976
rect 484320 266762 484348 273550
rect 486712 271046 486740 277780
rect 487908 275874 487936 277780
rect 488552 277766 489118 277794
rect 487896 275868 487948 275874
rect 487896 275810 487948 275816
rect 487804 275052 487856 275058
rect 487804 274994 487856 275000
rect 487068 274372 487120 274378
rect 487068 274314 487120 274320
rect 486700 271040 486752 271046
rect 486700 270982 486752 270988
rect 487080 266762 487108 274314
rect 487816 267578 487844 274994
rect 488356 273828 488408 273834
rect 488356 273770 488408 273776
rect 487804 267572 487856 267578
rect 487804 267514 487856 267520
rect 487528 266892 487580 266898
rect 487528 266834 487580 266840
rect 484308 266756 484360 266762
rect 484308 266698 484360 266704
rect 485872 266756 485924 266762
rect 485872 266698 485924 266704
rect 487068 266756 487120 266762
rect 487068 266698 487120 266704
rect 485044 266212 485096 266218
rect 485044 266154 485096 266160
rect 483860 264302 484242 264330
rect 485056 264316 485084 266154
rect 485884 264316 485912 266698
rect 486700 266076 486752 266082
rect 486700 266018 486752 266024
rect 486712 264316 486740 266018
rect 487540 264316 487568 266834
rect 488368 264316 488396 273770
rect 488552 268802 488580 277766
rect 490300 271862 490328 277780
rect 491496 275738 491524 277780
rect 491864 277766 492614 277794
rect 491484 275732 491536 275738
rect 491484 275674 491536 275680
rect 490564 274916 490616 274922
rect 490564 274858 490616 274864
rect 490288 271856 490340 271862
rect 490288 271798 490340 271804
rect 488540 268796 488592 268802
rect 488540 268738 488592 268744
rect 489184 267980 489236 267986
rect 489184 267922 489236 267928
rect 489196 264316 489224 267922
rect 490012 267708 490064 267714
rect 490012 267650 490064 267656
rect 490024 264316 490052 267650
rect 490576 266626 490604 274858
rect 491864 268666 491892 277766
rect 493796 277394 493824 277780
rect 493704 277366 493824 277394
rect 493704 271726 493732 277366
rect 493876 275732 493928 275738
rect 493876 275674 493928 275680
rect 493888 274786 493916 275674
rect 493876 274780 493928 274786
rect 493876 274722 493928 274728
rect 494992 274106 495020 277780
rect 495452 277766 496202 277794
rect 497016 277766 497398 277794
rect 494980 274100 495032 274106
rect 494980 274042 495032 274048
rect 493692 271720 493744 271726
rect 493692 271662 493744 271668
rect 495256 271040 495308 271046
rect 495256 270982 495308 270988
rect 492588 270904 492640 270910
rect 492588 270846 492640 270852
rect 491852 268660 491904 268666
rect 491852 268602 491904 268608
rect 492220 268524 492272 268530
rect 492220 268466 492272 268472
rect 492232 268410 492260 268466
rect 492140 268382 492260 268410
rect 492140 268258 492168 268382
rect 492128 268252 492180 268258
rect 492128 268194 492180 268200
rect 492312 268252 492364 268258
rect 492312 268194 492364 268200
rect 492324 267986 492352 268194
rect 490840 267980 490892 267986
rect 490840 267922 490892 267928
rect 492312 267980 492364 267986
rect 492312 267922 492364 267928
rect 490564 266620 490616 266626
rect 490564 266562 490616 266568
rect 490852 264316 490880 267922
rect 492600 266626 492628 270846
rect 493324 267980 493376 267986
rect 493324 267922 493376 267928
rect 491668 266620 491720 266626
rect 491668 266562 491720 266568
rect 492588 266620 492640 266626
rect 492588 266562 492640 266568
rect 491680 264316 491708 266562
rect 492496 265940 492548 265946
rect 492496 265882 492548 265888
rect 492508 264316 492536 265882
rect 493336 264316 493364 267922
rect 494980 266756 495032 266762
rect 494980 266698 495032 266704
rect 494152 266620 494204 266626
rect 494152 266562 494204 266568
rect 494164 264316 494192 266562
rect 494992 264316 495020 266698
rect 495268 266626 495296 270982
rect 495452 269074 495480 277766
rect 496544 271856 496596 271862
rect 496544 271798 496596 271804
rect 495440 269068 495492 269074
rect 495440 269010 495492 269016
rect 495808 269068 495860 269074
rect 495808 269010 495860 269016
rect 495256 266620 495308 266626
rect 495256 266562 495308 266568
rect 495820 264316 495848 269010
rect 496556 264330 496584 271798
rect 497016 271454 497044 277766
rect 498580 275602 498608 277780
rect 498568 275596 498620 275602
rect 498568 275538 498620 275544
rect 499776 274786 499804 277780
rect 500512 277766 500894 277794
rect 498476 274780 498528 274786
rect 498476 274722 498528 274728
rect 499764 274780 499816 274786
rect 499764 274722 499816 274728
rect 497004 271448 497056 271454
rect 497004 271390 497056 271396
rect 497278 269512 497334 269521
rect 497278 269447 497334 269456
rect 497292 267714 497320 269447
rect 498292 268932 498344 268938
rect 498292 268874 498344 268880
rect 497280 267708 497332 267714
rect 497280 267650 497332 267656
rect 497464 266620 497516 266626
rect 497464 266562 497516 266568
rect 496556 264302 496662 264330
rect 497476 264316 497504 266562
rect 498304 264316 498332 268874
rect 498488 268666 498516 274722
rect 499488 271720 499540 271726
rect 499488 271662 499540 271668
rect 498476 268660 498528 268666
rect 498476 268602 498528 268608
rect 499500 264330 499528 271662
rect 500512 271590 500540 277766
rect 502076 275738 502104 277780
rect 502352 277766 503286 277794
rect 502064 275732 502116 275738
rect 502064 275674 502116 275680
rect 501604 274780 501656 274786
rect 501604 274722 501656 274728
rect 500868 274236 500920 274242
rect 500868 274178 500920 274184
rect 500500 271584 500552 271590
rect 500500 271526 500552 271532
rect 500684 268796 500736 268802
rect 500684 268738 500736 268744
rect 499672 267708 499724 267714
rect 499672 267650 499724 267656
rect 499684 266762 499712 267650
rect 499672 266756 499724 266762
rect 499672 266698 499724 266704
rect 499856 266756 499908 266762
rect 499856 266698 499908 266704
rect 499868 266642 499896 266698
rect 499776 266614 499896 266642
rect 499776 266490 499804 266614
rect 499764 266484 499816 266490
rect 499764 266426 499816 266432
rect 499948 266484 500000 266490
rect 499948 266426 500000 266432
rect 499146 264302 499528 264330
rect 499960 264316 499988 266426
rect 500696 264330 500724 268738
rect 500880 266490 500908 274178
rect 501616 266762 501644 274722
rect 501972 271584 502024 271590
rect 501972 271526 502024 271532
rect 501604 266756 501656 266762
rect 501604 266698 501656 266704
rect 500868 266484 500920 266490
rect 500868 266426 500920 266432
rect 501984 264330 502012 271526
rect 502352 268394 502380 277766
rect 504468 271318 504496 277780
rect 504732 275868 504784 275874
rect 504732 275810 504784 275816
rect 504456 271312 504508 271318
rect 504456 271254 504508 271260
rect 503260 268660 503312 268666
rect 503260 268602 503312 268608
rect 502340 268388 502392 268394
rect 502340 268330 502392 268336
rect 502432 266756 502484 266762
rect 502432 266698 502484 266704
rect 500696 264302 500802 264330
rect 501630 264302 502012 264330
rect 502444 264316 502472 266698
rect 503272 264316 503300 268602
rect 504088 266484 504140 266490
rect 504088 266426 504140 266432
rect 504100 264316 504128 266426
rect 504744 264330 504772 275810
rect 505664 274786 505692 277780
rect 505836 275732 505888 275738
rect 505836 275674 505888 275680
rect 505652 274780 505704 274786
rect 505652 274722 505704 274728
rect 504916 271448 504968 271454
rect 504916 271390 504968 271396
rect 504928 266490 504956 271390
rect 505848 267442 505876 275674
rect 506480 274780 506532 274786
rect 506480 274722 506532 274728
rect 506110 268424 506166 268433
rect 506110 268359 506166 268368
rect 505836 267436 505888 267442
rect 505836 267378 505888 267384
rect 504916 266484 504968 266490
rect 504916 266426 504968 266432
rect 506124 264330 506152 268359
rect 506492 267850 506520 274722
rect 506860 272134 506888 277780
rect 506848 272128 506900 272134
rect 506848 272070 506900 272076
rect 507674 271144 507730 271153
rect 507674 271079 507730 271088
rect 506480 267844 506532 267850
rect 506480 267786 506532 267792
rect 507400 267436 507452 267442
rect 507400 267378 507452 267384
rect 506572 266484 506624 266490
rect 506572 266426 506624 266432
rect 504744 264302 504942 264330
rect 505770 264302 506152 264330
rect 506584 264316 506612 266426
rect 507412 264316 507440 267378
rect 507688 266490 507716 271079
rect 507964 270638 507992 277780
rect 509160 275466 509188 277780
rect 510068 275596 510120 275602
rect 510068 275538 510120 275544
rect 509148 275460 509200 275466
rect 509148 275402 509200 275408
rect 509148 271312 509200 271318
rect 509148 271254 509200 271260
rect 507952 270632 508004 270638
rect 507952 270574 508004 270580
rect 507860 269408 507912 269414
rect 507860 269350 507912 269356
rect 507872 267578 507900 269350
rect 509160 267734 509188 271254
rect 509700 270632 509752 270638
rect 509700 270574 509752 270580
rect 509068 267706 509188 267734
rect 507860 267572 507912 267578
rect 507860 267514 507912 267520
rect 508228 267572 508280 267578
rect 508228 267514 508280 267520
rect 507860 267300 507912 267306
rect 507860 267242 507912 267248
rect 507872 266490 507900 267242
rect 507676 266484 507728 266490
rect 507676 266426 507728 266432
rect 507860 266484 507912 266490
rect 507860 266426 507912 266432
rect 508240 264316 508268 267514
rect 509068 264316 509096 267706
rect 509712 267073 509740 270574
rect 509884 267300 509936 267306
rect 509884 267242 509936 267248
rect 509698 267064 509754 267073
rect 509698 266999 509754 267008
rect 509896 264316 509924 267242
rect 510080 266490 510108 275538
rect 510356 274786 510384 277780
rect 510344 274780 510396 274786
rect 510344 274722 510396 274728
rect 510528 274780 510580 274786
rect 510528 274722 510580 274728
rect 510540 270638 510568 274722
rect 511552 271182 511580 277780
rect 512748 275738 512776 277780
rect 512736 275732 512788 275738
rect 512736 275674 512788 275680
rect 512184 275460 512236 275466
rect 512184 275402 512236 275408
rect 511540 271176 511592 271182
rect 511540 271118 511592 271124
rect 511908 271176 511960 271182
rect 511908 271118 511960 271124
rect 510528 270632 510580 270638
rect 510528 270574 510580 270580
rect 510712 268524 510764 268530
rect 510712 268466 510764 268472
rect 510068 266484 510120 266490
rect 510068 266426 510120 266432
rect 510724 264316 510752 268466
rect 511920 264330 511948 271118
rect 512196 267170 512224 275402
rect 513194 273864 513250 273873
rect 513194 273799 513250 273808
rect 512184 267164 512236 267170
rect 512184 267106 512236 267112
rect 512368 267164 512420 267170
rect 512368 267106 512420 267112
rect 511566 264302 511948 264330
rect 512380 264316 512408 267106
rect 513208 264316 513236 273799
rect 513944 273086 513972 277780
rect 513932 273080 513984 273086
rect 513932 273022 513984 273028
rect 515140 272814 515168 277780
rect 516244 275330 516272 277780
rect 516612 277766 517454 277794
rect 517900 277766 518650 277794
rect 516416 275732 516468 275738
rect 516416 275674 516468 275680
rect 516232 275324 516284 275330
rect 516232 275266 516284 275272
rect 515128 272808 515180 272814
rect 515128 272750 515180 272756
rect 514024 272128 514076 272134
rect 514024 272070 514076 272076
rect 514036 266898 514064 272070
rect 516428 271946 516456 275674
rect 516060 271918 516456 271946
rect 514024 266892 514076 266898
rect 514024 266834 514076 266840
rect 514392 266892 514444 266898
rect 514392 266834 514444 266840
rect 514404 264330 514432 266834
rect 516060 266490 516088 271918
rect 516612 270502 516640 277766
rect 517336 272808 517388 272814
rect 517336 272750 517388 272756
rect 516600 270496 516652 270502
rect 516600 270438 516652 270444
rect 517150 267336 517206 267345
rect 517150 267271 517206 267280
rect 514852 266484 514904 266490
rect 514852 266426 514904 266432
rect 516048 266484 516100 266490
rect 516048 266426 516100 266432
rect 516508 266484 516560 266490
rect 516508 266426 516560 266432
rect 514050 264302 514432 264330
rect 514864 264316 514892 266426
rect 515680 265804 515732 265810
rect 515680 265746 515732 265752
rect 515692 264316 515720 265746
rect 516520 264316 516548 266426
rect 517164 264330 517192 267271
rect 517348 266490 517376 272750
rect 517704 270496 517756 270502
rect 517704 270438 517756 270444
rect 517716 267306 517744 270438
rect 517900 268394 517928 277766
rect 519832 275602 519860 277780
rect 520292 277766 521042 277794
rect 519820 275596 519872 275602
rect 519820 275538 519872 275544
rect 520096 273080 520148 273086
rect 520096 273022 520148 273028
rect 517888 268388 517940 268394
rect 517888 268330 517940 268336
rect 519818 267608 519874 267617
rect 519818 267543 519874 267552
rect 517704 267300 517756 267306
rect 517704 267242 517756 267248
rect 517520 266892 517572 266898
rect 517520 266834 517572 266840
rect 518992 266892 519044 266898
rect 518992 266834 519044 266840
rect 517532 266490 517560 266834
rect 517336 266484 517388 266490
rect 517336 266426 517388 266432
rect 517520 266484 517572 266490
rect 517520 266426 517572 266432
rect 518164 265668 518216 265674
rect 518164 265610 518216 265616
rect 517164 264302 517362 264330
rect 518176 264316 518204 265610
rect 519004 264316 519032 266834
rect 519832 264316 519860 267543
rect 520108 266898 520136 273022
rect 520292 270366 520320 277766
rect 522224 272950 522252 277780
rect 523420 276010 523448 277780
rect 524524 277394 524552 277780
rect 525720 277394 525748 277780
rect 524432 277366 524552 277394
rect 525628 277366 525748 277394
rect 523408 276004 523460 276010
rect 523408 275946 523460 275952
rect 523040 275596 523092 275602
rect 523040 275538 523092 275544
rect 522394 274136 522450 274145
rect 522394 274071 522450 274080
rect 522212 272944 522264 272950
rect 522212 272886 522264 272892
rect 521566 272776 521622 272785
rect 521566 272711 521622 272720
rect 520280 270360 520332 270366
rect 520280 270302 520332 270308
rect 521580 267734 521608 272711
rect 521488 267706 521608 267734
rect 520648 267164 520700 267170
rect 520648 267106 520700 267112
rect 520096 266892 520148 266898
rect 520096 266834 520148 266840
rect 520660 264316 520688 267106
rect 521488 264316 521516 267706
rect 522408 267578 522436 274071
rect 523052 270774 523080 275538
rect 523684 275324 523736 275330
rect 523684 275266 523736 275272
rect 523696 274514 523724 275266
rect 523684 274508 523736 274514
rect 523684 274450 523736 274456
rect 524052 272944 524104 272950
rect 524052 272886 524104 272892
rect 523040 270768 523092 270774
rect 523040 270710 523092 270716
rect 523132 270360 523184 270366
rect 523132 270302 523184 270308
rect 522396 267572 522448 267578
rect 522396 267514 522448 267520
rect 522304 266892 522356 266898
rect 522304 266834 522356 266840
rect 522316 264316 522344 266834
rect 523144 264316 523172 270302
rect 524064 267734 524092 272886
rect 524432 269822 524460 277366
rect 525154 275632 525210 275641
rect 525628 275602 525656 277366
rect 525800 276004 525852 276010
rect 525800 275946 525852 275952
rect 525154 275567 525210 275576
rect 525616 275596 525668 275602
rect 524420 269816 524472 269822
rect 524420 269758 524472 269764
rect 523972 267706 524092 267734
rect 523684 267572 523736 267578
rect 523684 267514 523736 267520
rect 523696 267034 523724 267514
rect 523684 267028 523736 267034
rect 523684 266970 523736 266976
rect 523972 264316 524000 267706
rect 524236 267164 524288 267170
rect 524236 267106 524288 267112
rect 524248 266898 524276 267106
rect 524236 266892 524288 266898
rect 524236 266834 524288 266840
rect 525168 264330 525196 275567
rect 525616 275538 525668 275544
rect 525812 272814 525840 275946
rect 525982 275632 526038 275641
rect 525982 275567 525984 275576
rect 526036 275567 526038 275576
rect 525984 275538 526036 275544
rect 526916 274922 526944 277780
rect 527192 277766 528126 277794
rect 526904 274916 526956 274922
rect 526904 274858 526956 274864
rect 525800 272808 525852 272814
rect 525800 272750 525852 272756
rect 526812 272808 526864 272814
rect 526812 272750 526864 272756
rect 526444 270768 526496 270774
rect 526444 270710 526496 270716
rect 525616 270088 525668 270094
rect 525616 270030 525668 270036
rect 524814 264302 525196 264330
rect 525628 264316 525656 270030
rect 526456 267714 526484 270710
rect 526444 267708 526496 267714
rect 526444 267650 526496 267656
rect 526824 264330 526852 272750
rect 527192 270230 527220 277766
rect 529308 272678 529336 277780
rect 529570 275224 529626 275233
rect 529570 275159 529626 275168
rect 529296 272672 529348 272678
rect 529296 272614 529348 272620
rect 527180 270224 527232 270230
rect 527180 270166 527232 270172
rect 528100 270224 528152 270230
rect 528100 270166 528152 270172
rect 527272 267708 527324 267714
rect 527272 267650 527324 267656
rect 526470 264302 526852 264330
rect 527284 264316 527312 267650
rect 528112 264316 528140 270166
rect 528928 266892 528980 266898
rect 528928 266834 528980 266840
rect 528940 264316 528968 266834
rect 529584 264330 529612 275159
rect 530504 275058 530532 277780
rect 531332 277766 531622 277794
rect 530492 275052 530544 275058
rect 530492 274994 530544 275000
rect 530676 275052 530728 275058
rect 530676 274994 530728 275000
rect 529756 272672 529808 272678
rect 529756 272614 529808 272620
rect 529768 266898 529796 272614
rect 530688 267578 530716 274994
rect 530950 270328 531006 270337
rect 530950 270263 531006 270272
rect 530676 267572 530728 267578
rect 530676 267514 530728 267520
rect 529756 266892 529808 266898
rect 529756 266834 529808 266840
rect 530964 264330 530992 270263
rect 531332 269958 531360 277766
rect 532804 273970 532832 277780
rect 534000 275466 534028 277780
rect 534184 277766 535210 277794
rect 533988 275460 534040 275466
rect 533988 275402 534040 275408
rect 533436 274100 533488 274106
rect 533436 274042 533488 274048
rect 532792 273964 532844 273970
rect 532792 273906 532844 273912
rect 531320 269952 531372 269958
rect 531320 269894 531372 269900
rect 531688 269952 531740 269958
rect 531688 269894 531740 269900
rect 531700 264330 531728 269894
rect 532240 267572 532292 267578
rect 532240 267514 532292 267520
rect 529584 264302 529782 264330
rect 530610 264302 530992 264330
rect 531438 264302 531728 264330
rect 532252 264316 532280 267514
rect 533448 264330 533476 274042
rect 533894 272504 533950 272513
rect 533894 272439 533950 272448
rect 533094 264302 533476 264330
rect 533908 264316 533936 272439
rect 534184 269278 534212 277766
rect 535736 275460 535788 275466
rect 535736 275402 535788 275408
rect 535552 269816 535604 269822
rect 535552 269758 535604 269764
rect 534172 269272 534224 269278
rect 534172 269214 534224 269220
rect 534724 268388 534776 268394
rect 534724 268330 534776 268336
rect 534736 264316 534764 268330
rect 535564 264316 535592 269758
rect 535748 268394 535776 275402
rect 536392 272542 536420 277780
rect 537312 277766 537602 277794
rect 537312 274786 537340 277766
rect 538784 274786 538812 277780
rect 537300 274780 537352 274786
rect 537300 274722 537352 274728
rect 537668 274780 537720 274786
rect 537668 274722 537720 274728
rect 538772 274780 538824 274786
rect 538772 274722 538824 274728
rect 539508 274780 539560 274786
rect 539508 274722 539560 274728
rect 537484 274508 537536 274514
rect 537484 274450 537536 274456
rect 536380 272536 536432 272542
rect 536380 272478 536432 272484
rect 535736 268388 535788 268394
rect 535736 268330 535788 268336
rect 536380 268388 536432 268394
rect 536380 268330 536432 268336
rect 536392 264316 536420 268330
rect 537208 267028 537260 267034
rect 537208 266970 537260 266976
rect 537220 264316 537248 266970
rect 537496 266898 537524 274450
rect 537680 269793 537708 274722
rect 539324 272536 539376 272542
rect 539324 272478 539376 272484
rect 538034 270056 538090 270065
rect 538034 269991 538090 270000
rect 537666 269784 537722 269793
rect 537666 269719 537722 269728
rect 537484 266892 537536 266898
rect 537484 266834 537536 266840
rect 538048 264316 538076 269991
rect 539336 264330 539364 272478
rect 539520 269249 539548 274722
rect 539888 272406 539916 277780
rect 541084 275058 541112 277780
rect 542096 277766 542294 277794
rect 541072 275052 541124 275058
rect 541072 274994 541124 275000
rect 542096 274786 542124 277766
rect 542268 275052 542320 275058
rect 542268 274994 542320 275000
rect 542084 274780 542136 274786
rect 542084 274722 542136 274728
rect 542084 273964 542136 273970
rect 542084 273906 542136 273912
rect 539876 272400 539928 272406
rect 539876 272342 539928 272348
rect 541624 272400 541676 272406
rect 541624 272342 541676 272348
rect 540518 269784 540574 269793
rect 540518 269719 540574 269728
rect 539506 269240 539562 269249
rect 539506 269175 539562 269184
rect 539690 267064 539746 267073
rect 539690 266999 539746 267008
rect 538890 264302 539364 264330
rect 539704 264316 539732 266999
rect 540532 264316 540560 269719
rect 541636 266898 541664 272342
rect 540980 266892 541032 266898
rect 540980 266834 541032 266840
rect 541624 266892 541676 266898
rect 541624 266834 541676 266840
rect 541900 266892 541952 266898
rect 541900 266834 541952 266840
rect 540992 266490 541020 266834
rect 540980 266484 541032 266490
rect 540980 266426 541032 266432
rect 541348 266484 541400 266490
rect 541348 266426 541400 266432
rect 541360 264316 541388 266426
rect 541912 264194 541940 266834
rect 542096 266490 542124 273906
rect 542280 273426 542308 274994
rect 543280 274916 543332 274922
rect 543280 274858 543332 274864
rect 542268 273420 542320 273426
rect 542268 273362 542320 273368
rect 542084 266484 542136 266490
rect 542084 266426 542136 266432
rect 543292 264330 543320 274858
rect 543476 273222 543504 277780
rect 544672 275194 544700 277780
rect 545868 275330 545896 277780
rect 546512 277766 547078 277794
rect 545856 275324 545908 275330
rect 545856 275266 545908 275272
rect 546040 275324 546092 275330
rect 546040 275266 546092 275272
rect 544660 275188 544712 275194
rect 544660 275130 544712 275136
rect 546052 273562 546080 275266
rect 546040 273556 546092 273562
rect 546040 273498 546092 273504
rect 543464 273216 543516 273222
rect 543464 273158 543516 273164
rect 546512 269686 546540 277766
rect 548168 272270 548196 277780
rect 549364 275058 549392 277780
rect 549916 277766 550574 277794
rect 549352 275052 549404 275058
rect 549352 274994 549404 275000
rect 548156 272264 548208 272270
rect 548156 272206 548208 272212
rect 546500 269680 546552 269686
rect 546500 269622 546552 269628
rect 549916 269550 549944 277766
rect 551560 275052 551612 275058
rect 551560 274994 551612 275000
rect 549904 269544 549956 269550
rect 549904 269486 549956 269492
rect 551572 267986 551600 274994
rect 551756 271425 551784 277780
rect 552952 275330 552980 277780
rect 553412 277766 554162 277794
rect 554792 277766 555266 277794
rect 552940 275324 552992 275330
rect 552940 275266 552992 275272
rect 553124 275324 553176 275330
rect 553124 275266 553176 275272
rect 552664 275188 552716 275194
rect 552664 275130 552716 275136
rect 552676 273698 552704 275130
rect 553136 275058 553164 275266
rect 553124 275052 553176 275058
rect 553124 274994 553176 275000
rect 552664 273692 552716 273698
rect 552664 273634 552716 273640
rect 552664 273556 552716 273562
rect 552664 273498 552716 273504
rect 551742 271416 551798 271425
rect 551742 271351 551798 271360
rect 551560 267980 551612 267986
rect 551560 267922 551612 267928
rect 552676 266626 552704 273498
rect 552664 266620 552716 266626
rect 552664 266562 552716 266568
rect 553412 265402 553440 277766
rect 554792 266354 554820 277766
rect 556448 274650 556476 277780
rect 557644 277394 557672 277780
rect 557552 277366 557672 277394
rect 556436 274644 556488 274650
rect 556436 274586 556488 274592
rect 554780 266348 554832 266354
rect 554780 266290 554832 266296
rect 557552 265538 557580 277366
rect 558840 276690 558868 277780
rect 558828 276684 558880 276690
rect 558828 276626 558880 276632
rect 560036 275194 560064 277780
rect 560312 277766 561246 277794
rect 561692 277766 562442 277794
rect 560024 275188 560076 275194
rect 560024 275130 560076 275136
rect 559564 275052 559616 275058
rect 559564 274994 559616 275000
rect 559576 273834 559604 274994
rect 559748 274644 559800 274650
rect 559748 274586 559800 274592
rect 559564 273828 559616 273834
rect 559564 273770 559616 273776
rect 559760 266762 559788 274586
rect 560312 269414 560340 277766
rect 560300 269408 560352 269414
rect 560300 269350 560352 269356
rect 559748 266756 559800 266762
rect 559748 266698 559800 266704
rect 561692 266218 561720 277766
rect 563532 274378 563560 277780
rect 564452 277766 564742 277794
rect 563520 274372 563572 274378
rect 563520 274314 563572 274320
rect 563704 274372 563756 274378
rect 563704 274314 563756 274320
rect 563716 267617 563744 274314
rect 563702 267608 563758 267617
rect 563702 267543 563758 267552
rect 561680 266212 561732 266218
rect 561680 266154 561732 266160
rect 564452 266082 564480 277766
rect 565924 272134 565952 277780
rect 567120 275058 567148 277780
rect 567396 277766 568330 277794
rect 568592 277766 569526 277794
rect 569972 277766 570722 277794
rect 567108 275052 567160 275058
rect 567108 274994 567160 275000
rect 565912 272128 565964 272134
rect 565912 272070 565964 272076
rect 567396 268122 567424 277766
rect 568592 269521 568620 277766
rect 568578 269512 568634 269521
rect 568578 269447 568634 269456
rect 569972 268258 570000 277766
rect 571812 270910 571840 277780
rect 572732 277766 573022 277794
rect 571800 270904 571852 270910
rect 571800 270846 571852 270852
rect 569960 268252 570012 268258
rect 569960 268194 570012 268200
rect 567384 268116 567436 268122
rect 567384 268058 567436 268064
rect 564440 266076 564492 266082
rect 564440 266018 564492 266024
rect 572732 265946 572760 277766
rect 574204 275330 574232 277780
rect 574192 275324 574244 275330
rect 574192 275266 574244 275272
rect 575400 271046 575428 277780
rect 575388 271040 575440 271046
rect 575388 270982 575440 270988
rect 576124 271040 576176 271046
rect 576124 270982 576176 270988
rect 576136 267442 576164 270982
rect 576596 270774 576624 277780
rect 576872 277766 577806 277794
rect 576584 270768 576636 270774
rect 576584 270710 576636 270716
rect 576872 269074 576900 277766
rect 578896 271862 578924 277780
rect 580092 273562 580120 277780
rect 581012 277766 581302 277794
rect 580080 273556 580132 273562
rect 580080 273498 580132 273504
rect 578884 271856 578936 271862
rect 578884 271798 578936 271804
rect 576860 269068 576912 269074
rect 576860 269010 576912 269016
rect 581012 268938 581040 277766
rect 582484 271726 582512 277780
rect 583680 274242 583708 277780
rect 584140 277766 584890 277794
rect 585612 277766 586086 277794
rect 583668 274236 583720 274242
rect 583668 274178 583720 274184
rect 582472 271720 582524 271726
rect 582472 271662 582524 271668
rect 581000 268932 581052 268938
rect 581000 268874 581052 268880
rect 582196 268932 582248 268938
rect 582196 268874 582248 268880
rect 576124 267436 576176 267442
rect 576124 267378 576176 267384
rect 582208 267306 582236 268874
rect 584140 268802 584168 277766
rect 585612 271590 585640 277766
rect 587176 274650 587204 277780
rect 587912 277766 588386 277794
rect 587164 274644 587216 274650
rect 587164 274586 587216 274592
rect 585600 271584 585652 271590
rect 585600 271526 585652 271532
rect 585784 271584 585836 271590
rect 585784 271526 585836 271532
rect 584128 268796 584180 268802
rect 584128 268738 584180 268744
rect 585796 267345 585824 271526
rect 587912 268666 587940 277766
rect 589568 271454 589596 277780
rect 590764 275874 590792 277780
rect 591040 277766 591974 277794
rect 590752 275868 590804 275874
rect 590752 275810 590804 275816
rect 589556 271448 589608 271454
rect 589556 271390 589608 271396
rect 587900 268660 587952 268666
rect 587900 268602 587952 268608
rect 591040 268433 591068 277766
rect 592684 271448 592736 271454
rect 592684 271390 592736 271396
rect 591026 268424 591082 268433
rect 591026 268359 591082 268368
rect 592696 267714 592724 271390
rect 593156 271153 593184 277780
rect 593142 271144 593198 271153
rect 593142 271079 593198 271088
rect 594352 271046 594380 277780
rect 595456 274145 595484 277780
rect 595442 274136 595498 274145
rect 595442 274071 595498 274080
rect 596652 271318 596680 277780
rect 597572 277766 597862 277794
rect 596640 271312 596692 271318
rect 596640 271254 596692 271260
rect 596824 271312 596876 271318
rect 596824 271254 596876 271260
rect 594340 271040 594392 271046
rect 594340 270982 594392 270988
rect 592684 267708 592736 267714
rect 592684 267650 592736 267656
rect 596836 267578 596864 271254
rect 597572 270502 597600 277766
rect 599044 277394 599072 277780
rect 598952 277366 599072 277394
rect 597560 270496 597612 270502
rect 597560 270438 597612 270444
rect 598952 268530 598980 277366
rect 600240 271182 600268 277780
rect 600424 277766 601450 277794
rect 600228 271176 600280 271182
rect 600228 271118 600280 271124
rect 600424 268938 600452 277766
rect 602540 273873 602568 277780
rect 602526 273864 602582 273873
rect 602526 273799 602582 273808
rect 603736 272406 603764 277780
rect 604932 275738 604960 277780
rect 605852 277766 606142 277794
rect 604920 275732 604972 275738
rect 604920 275674 604972 275680
rect 605104 275732 605156 275738
rect 605104 275674 605156 275680
rect 603724 272400 603776 272406
rect 603724 272342 603776 272348
rect 602344 271176 602396 271182
rect 602344 271118 602396 271124
rect 600412 268932 600464 268938
rect 600412 268874 600464 268880
rect 598940 268524 598992 268530
rect 598940 268466 598992 268472
rect 596824 267572 596876 267578
rect 596824 267514 596876 267520
rect 585782 267336 585838 267345
rect 582196 267300 582248 267306
rect 585782 267271 585838 267280
rect 582196 267242 582248 267248
rect 602356 266898 602384 271118
rect 605116 270366 605144 275674
rect 605104 270360 605156 270366
rect 605104 270302 605156 270308
rect 602344 266892 602396 266898
rect 602344 266834 602396 266840
rect 572720 265940 572772 265946
rect 572720 265882 572772 265888
rect 605852 265810 605880 277766
rect 607324 276010 607352 277780
rect 607312 276004 607364 276010
rect 607312 275946 607364 275952
rect 608520 271590 608548 277780
rect 608704 277766 609730 277794
rect 608508 271584 608560 271590
rect 608508 271526 608560 271532
rect 605840 265804 605892 265810
rect 605840 265746 605892 265752
rect 608704 265674 608732 277766
rect 610820 273086 610848 277780
rect 612016 274378 612044 277780
rect 613212 274514 613240 277780
rect 613200 274508 613252 274514
rect 613200 274450 613252 274456
rect 612004 274372 612056 274378
rect 612004 274314 612056 274320
rect 610808 273080 610860 273086
rect 610808 273022 610860 273028
rect 614408 272785 614436 277780
rect 615604 277394 615632 277780
rect 615512 277366 615632 277394
rect 614394 272776 614450 272785
rect 614394 272711 614450 272720
rect 615512 267170 615540 277366
rect 616800 275738 616828 277780
rect 616788 275732 616840 275738
rect 616788 275674 616840 275680
rect 617996 272950 618024 277780
rect 619100 275602 619128 277780
rect 619652 277766 620310 277794
rect 619088 275596 619140 275602
rect 619088 275538 619140 275544
rect 619180 274712 619232 274718
rect 619180 274654 619232 274660
rect 617984 272944 618036 272950
rect 617984 272886 618036 272892
rect 619192 270230 619220 274654
rect 619180 270224 619232 270230
rect 619180 270166 619232 270172
rect 619652 270094 619680 277766
rect 621492 272814 621520 277780
rect 621480 272808 621532 272814
rect 621480 272750 621532 272756
rect 622688 271454 622716 277780
rect 623884 274718 623912 277780
rect 623872 274712 623924 274718
rect 623872 274654 623924 274660
rect 625080 272678 625108 277780
rect 625804 275596 625856 275602
rect 625804 275538 625856 275544
rect 625068 272672 625120 272678
rect 625068 272614 625120 272620
rect 622676 271448 622728 271454
rect 622676 271390 622728 271396
rect 619640 270088 619692 270094
rect 619640 270030 619692 270036
rect 615500 267164 615552 267170
rect 615500 267106 615552 267112
rect 625816 267073 625844 275538
rect 626184 275233 626212 277780
rect 626552 277766 627394 277794
rect 627932 277766 628590 277794
rect 626170 275224 626226 275233
rect 626170 275159 626226 275168
rect 626552 270337 626580 277766
rect 626538 270328 626594 270337
rect 626538 270263 626594 270272
rect 627932 269958 627960 277766
rect 629772 271318 629800 277780
rect 630968 274106 630996 277780
rect 630956 274100 631008 274106
rect 630956 274042 631008 274048
rect 632164 272513 632192 277780
rect 633360 275466 633388 277780
rect 633544 277766 634478 277794
rect 634832 277766 635674 277794
rect 636212 277766 636870 277794
rect 637592 277766 638066 277794
rect 633348 275460 633400 275466
rect 633348 275402 633400 275408
rect 632150 272504 632206 272513
rect 632150 272439 632206 272448
rect 629760 271312 629812 271318
rect 629760 271254 629812 271260
rect 627920 269952 627972 269958
rect 627920 269894 627972 269900
rect 633544 269822 633572 277766
rect 633532 269816 633584 269822
rect 633532 269758 633584 269764
rect 634832 268394 634860 277766
rect 634820 268388 634872 268394
rect 634820 268330 634872 268336
rect 625802 267064 625858 267073
rect 636212 267034 636240 277766
rect 637592 270065 637620 277766
rect 639248 272542 639276 277780
rect 640444 275602 640472 277780
rect 640720 277766 641654 277794
rect 640432 275596 640484 275602
rect 640432 275538 640484 275544
rect 639236 272536 639288 272542
rect 639236 272478 639288 272484
rect 637578 270056 637634 270065
rect 637578 269991 637634 270000
rect 640720 269793 640748 277766
rect 642744 273970 642772 277780
rect 642732 273964 642784 273970
rect 642732 273906 642784 273912
rect 643940 271182 643968 277780
rect 645136 274922 645164 277780
rect 645872 277766 646346 277794
rect 647252 277766 647542 277794
rect 645124 274916 645176 274922
rect 645124 274858 645176 274864
rect 643928 271176 643980 271182
rect 643928 271118 643980 271124
rect 640706 269784 640762 269793
rect 640706 269719 640762 269728
rect 625802 266999 625858 267008
rect 636200 267028 636252 267034
rect 636200 266970 636252 266976
rect 608692 265668 608744 265674
rect 608692 265610 608744 265616
rect 557540 265532 557592 265538
rect 557540 265474 557592 265480
rect 553400 265396 553452 265402
rect 553400 265338 553452 265344
rect 543030 264302 543320 264330
rect 541912 264166 542202 264194
rect 554410 262168 554466 262177
rect 554410 262103 554466 262112
rect 554424 260914 554452 262103
rect 577504 261656 577556 261662
rect 577504 261598 577556 261604
rect 570604 261520 570656 261526
rect 570604 261462 570656 261468
rect 554412 260908 554464 260914
rect 554412 260850 554464 260856
rect 568580 260908 568632 260914
rect 568580 260850 568632 260856
rect 554318 259992 554374 260001
rect 554318 259927 554374 259936
rect 554332 259486 554360 259927
rect 554320 259480 554372 259486
rect 554320 259422 554372 259428
rect 560944 259480 560996 259486
rect 560944 259422 560996 259428
rect 553950 257816 554006 257825
rect 553950 257751 554006 257760
rect 553964 256766 553992 257751
rect 553952 256760 554004 256766
rect 553952 256702 554004 256708
rect 559564 256760 559616 256766
rect 559564 256702 559616 256708
rect 553490 255640 553546 255649
rect 553490 255575 553546 255584
rect 553504 249082 553532 255575
rect 554410 253464 554466 253473
rect 554410 253399 554466 253408
rect 554424 252618 554452 253399
rect 554412 252612 554464 252618
rect 554412 252554 554464 252560
rect 554134 251288 554190 251297
rect 554134 251223 554136 251232
rect 554188 251223 554190 251232
rect 556804 251252 556856 251258
rect 554136 251194 554188 251200
rect 556804 251194 556856 251200
rect 553858 249112 553914 249121
rect 553492 249076 553544 249082
rect 553858 249047 553914 249056
rect 553492 249018 553544 249024
rect 553872 246362 553900 249047
rect 554410 246936 554466 246945
rect 554410 246871 554466 246880
rect 553860 246356 553912 246362
rect 553860 246298 553912 246304
rect 554424 245682 554452 246871
rect 554412 245676 554464 245682
rect 554412 245618 554464 245624
rect 553398 244760 553454 244769
rect 553398 244695 553454 244704
rect 553412 244322 553440 244695
rect 553400 244316 553452 244322
rect 553400 244258 553452 244264
rect 555424 244316 555476 244322
rect 555424 244258 555476 244264
rect 553950 242584 554006 242593
rect 553950 242519 554006 242528
rect 553964 241534 553992 242519
rect 553952 241528 554004 241534
rect 553952 241470 554004 241476
rect 554042 240408 554098 240417
rect 554042 240343 554098 240352
rect 129648 230920 129700 230926
rect 129648 230862 129700 230868
rect 104808 230784 104860 230790
rect 104808 230726 104860 230732
rect 97908 230648 97960 230654
rect 97908 230590 97960 230596
rect 91008 230512 91060 230518
rect 91008 230454 91060 230460
rect 71042 230072 71098 230081
rect 71042 230007 71098 230016
rect 86224 230036 86276 230042
rect 65522 229800 65578 229809
rect 65522 229735 65578 229744
rect 64142 228576 64198 228585
rect 64142 228511 64198 228520
rect 63408 226296 63460 226302
rect 63408 226238 63460 226244
rect 61844 225558 61896 225564
rect 62762 225584 62818 225593
rect 60648 221740 60700 221746
rect 60648 221682 60700 221688
rect 60004 218068 60056 218074
rect 60004 218010 60056 218016
rect 60660 217002 60688 221682
rect 61856 217002 61884 225558
rect 62762 225519 62818 225528
rect 63224 224256 63276 224262
rect 63224 224198 63276 224204
rect 63236 218074 63264 224198
rect 62580 218068 62632 218074
rect 62580 218010 62632 218016
rect 63224 218068 63276 218074
rect 63224 218010 63276 218016
rect 62592 217002 62620 218010
rect 63420 217002 63448 226238
rect 64156 218346 64184 228511
rect 64786 222864 64842 222873
rect 64786 222799 64842 222808
rect 64144 218340 64196 218346
rect 64144 218282 64196 218288
rect 64236 218204 64288 218210
rect 64236 218146 64288 218152
rect 64248 217002 64276 218146
rect 64800 217002 64828 222799
rect 65536 218210 65564 229735
rect 68192 227180 68244 227186
rect 68192 227122 68244 227128
rect 66902 224496 66958 224505
rect 66902 224431 66958 224440
rect 66720 220652 66772 220658
rect 66720 220594 66772 220600
rect 65524 218204 65576 218210
rect 65524 218146 65576 218152
rect 65892 218068 65944 218074
rect 65892 218010 65944 218016
rect 65904 217002 65932 218010
rect 66732 217002 66760 220594
rect 66916 218074 66944 224431
rect 68204 218754 68232 227122
rect 70124 225888 70176 225894
rect 70124 225830 70176 225836
rect 68928 222896 68980 222902
rect 68928 222838 68980 222844
rect 68192 218748 68244 218754
rect 68192 218690 68244 218696
rect 68744 218340 68796 218346
rect 68744 218282 68796 218288
rect 67548 218204 67600 218210
rect 67548 218146 67600 218152
rect 66904 218068 66956 218074
rect 66904 218010 66956 218016
rect 67560 217002 67588 218146
rect 68376 218068 68428 218074
rect 68376 218010 68428 218016
rect 68388 217002 68416 218010
rect 55660 216974 55996 217002
rect 56488 216974 56548 217002
rect 57316 216974 57652 217002
rect 58144 216974 58480 217002
rect 58972 216974 59308 217002
rect 59800 216974 59860 217002
rect 60628 216974 60688 217002
rect 61456 216974 61884 217002
rect 62284 216974 62620 217002
rect 63112 216974 63448 217002
rect 63940 216974 64276 217002
rect 64768 216974 64828 217002
rect 65596 216974 65932 217002
rect 66424 216974 66760 217002
rect 67252 216974 67588 217002
rect 68080 216974 68416 217002
rect 68756 217002 68784 218282
rect 68940 218074 68968 222838
rect 68928 218068 68980 218074
rect 68928 218010 68980 218016
rect 70136 217002 70164 225830
rect 70858 218648 70914 218657
rect 70858 218583 70914 218592
rect 70872 217002 70900 218583
rect 71056 218210 71084 230007
rect 86224 229978 86276 229984
rect 73802 228304 73858 228313
rect 73802 228239 73858 228248
rect 72422 224768 72478 224777
rect 72422 224703 72478 224712
rect 71686 223136 71742 223145
rect 71686 223071 71742 223080
rect 71044 218204 71096 218210
rect 71044 218146 71096 218152
rect 71700 217002 71728 223071
rect 72436 218346 72464 224703
rect 73068 220108 73120 220114
rect 73068 220050 73120 220056
rect 72424 218340 72476 218346
rect 72424 218282 72476 218288
rect 72516 218068 72568 218074
rect 72516 218010 72568 218016
rect 72528 217002 72556 218010
rect 73080 217002 73108 220050
rect 73816 218074 73844 228239
rect 81348 227316 81400 227322
rect 81348 227258 81400 227264
rect 79966 226944 80022 226953
rect 79966 226879 80022 226888
rect 76564 224392 76616 224398
rect 76564 224334 76616 224340
rect 75828 223032 75880 223038
rect 75828 222974 75880 222980
rect 74172 221604 74224 221610
rect 74172 221546 74224 221552
rect 73804 218068 73856 218074
rect 73804 218010 73856 218016
rect 74184 217002 74212 221546
rect 75644 218204 75696 218210
rect 75644 218146 75696 218152
rect 75000 218068 75052 218074
rect 75000 218010 75052 218016
rect 75012 217002 75040 218010
rect 75656 217002 75684 218146
rect 75840 218074 75868 222974
rect 76380 220244 76432 220250
rect 76380 220186 76432 220192
rect 75828 218068 75880 218074
rect 75828 218010 75880 218016
rect 76392 217002 76420 220186
rect 76576 218210 76604 224334
rect 78404 223304 78456 223310
rect 78404 223246 78456 223252
rect 77206 218920 77262 218929
rect 77206 218855 77262 218864
rect 76564 218204 76616 218210
rect 76564 218146 76616 218152
rect 77220 217002 77248 218855
rect 78416 217002 78444 223246
rect 79784 220380 79836 220386
rect 79784 220322 79836 220328
rect 79048 218068 79100 218074
rect 79048 218010 79100 218016
rect 79060 217002 79088 218010
rect 79796 217002 79824 220322
rect 79980 218074 80008 226879
rect 81164 223168 81216 223174
rect 81164 223110 81216 223116
rect 79968 218068 80020 218074
rect 79968 218010 80020 218016
rect 80796 218068 80848 218074
rect 80796 218010 80848 218016
rect 80808 217002 80836 218010
rect 68756 216974 68908 217002
rect 69736 216974 70164 217002
rect 70564 216974 70900 217002
rect 71392 216974 71728 217002
rect 72220 216974 72556 217002
rect 73048 216974 73108 217002
rect 73876 216974 74212 217002
rect 74704 216974 75040 217002
rect 75532 216974 75684 217002
rect 76360 216974 76420 217002
rect 77188 216974 77248 217002
rect 78016 216974 78444 217002
rect 78844 216974 79088 217002
rect 79672 216974 79824 217002
rect 80500 216974 80836 217002
rect 81176 217002 81204 223110
rect 81360 218074 81388 227258
rect 84108 226024 84160 226030
rect 84108 225966 84160 225972
rect 82542 225584 82598 225593
rect 82542 225519 82598 225528
rect 81348 218068 81400 218074
rect 81348 218010 81400 218016
rect 82556 217002 82584 225519
rect 83924 218748 83976 218754
rect 83924 218690 83976 218696
rect 83280 218068 83332 218074
rect 83280 218010 83332 218016
rect 83292 217002 83320 218010
rect 83936 217002 83964 218690
rect 84120 218074 84148 225966
rect 85488 224528 85540 224534
rect 85488 224470 85540 224476
rect 84936 221468 84988 221474
rect 84936 221410 84988 221416
rect 84108 218068 84160 218074
rect 84108 218010 84160 218016
rect 84948 217002 84976 221410
rect 85500 217002 85528 224470
rect 86236 221610 86264 229978
rect 89626 227216 89682 227225
rect 89626 227151 89682 227160
rect 89166 225856 89222 225865
rect 89166 225791 89222 225800
rect 88248 223440 88300 223446
rect 88248 223382 88300 223388
rect 86224 221604 86276 221610
rect 86224 221546 86276 221552
rect 86592 220516 86644 220522
rect 86592 220458 86644 220464
rect 86604 217002 86632 220458
rect 87420 219020 87472 219026
rect 87420 218962 87472 218968
rect 87432 217002 87460 218962
rect 88260 217002 88288 223382
rect 89180 217002 89208 225791
rect 89640 217002 89668 227151
rect 91020 219434 91048 230454
rect 95240 229628 95292 229634
rect 95240 229570 95292 229576
rect 94504 229220 94556 229226
rect 94504 229162 94556 229168
rect 93768 228540 93820 228546
rect 93768 228482 93820 228488
rect 92386 223408 92442 223417
rect 92386 223343 92442 223352
rect 91560 221604 91612 221610
rect 91560 221546 91612 221552
rect 90836 219406 91048 219434
rect 90836 217002 90864 219406
rect 91572 217002 91600 221546
rect 92400 217002 92428 223343
rect 93584 219156 93636 219162
rect 93584 219098 93636 219104
rect 93216 218068 93268 218074
rect 93216 218010 93268 218016
rect 93228 217002 93256 218010
rect 81176 216974 81328 217002
rect 82156 216974 82584 217002
rect 82984 216974 83320 217002
rect 83812 216974 83964 217002
rect 84640 216974 84976 217002
rect 85468 216974 85528 217002
rect 86296 216974 86632 217002
rect 87124 216974 87460 217002
rect 87952 216974 88288 217002
rect 88780 216974 89208 217002
rect 89608 216974 89668 217002
rect 90436 216974 90864 217002
rect 91264 216974 91600 217002
rect 92092 216974 92428 217002
rect 92920 216974 93256 217002
rect 93596 217002 93624 219098
rect 93780 218074 93808 228482
rect 94516 221746 94544 229162
rect 95252 227322 95280 229570
rect 95240 227316 95292 227322
rect 95240 227258 95292 227264
rect 96528 227316 96580 227322
rect 96528 227258 96580 227264
rect 94504 221740 94556 221746
rect 94504 221682 94556 221688
rect 94872 221740 94924 221746
rect 94872 221682 94924 221688
rect 93768 218068 93820 218074
rect 93768 218010 93820 218016
rect 94884 217002 94912 221682
rect 95698 221504 95754 221513
rect 95698 221439 95754 221448
rect 95712 217002 95740 221439
rect 96540 217002 96568 227258
rect 97722 221776 97778 221785
rect 97722 221711 97778 221720
rect 97356 218068 97408 218074
rect 97356 218010 97408 218016
rect 97368 217002 97396 218010
rect 93596 216974 93748 217002
rect 94576 216974 94912 217002
rect 95404 216974 95740 217002
rect 96232 216974 96568 217002
rect 97060 216974 97396 217002
rect 97736 217002 97764 221711
rect 97920 218074 97948 230590
rect 100668 228812 100720 228818
rect 100668 228754 100720 228760
rect 99104 226160 99156 226166
rect 99104 226102 99156 226108
rect 97908 218068 97960 218074
rect 97908 218010 97960 218016
rect 99116 217002 99144 226102
rect 100484 218884 100536 218890
rect 100484 218826 100536 218832
rect 99840 218068 99892 218074
rect 99840 218010 99892 218016
rect 99852 217002 99880 218010
rect 100496 217002 100524 218826
rect 100680 218074 100708 228754
rect 103244 227452 103296 227458
rect 103244 227394 103296 227400
rect 102048 223576 102100 223582
rect 102048 223518 102100 223524
rect 101496 221876 101548 221882
rect 101496 221818 101548 221824
rect 100668 218068 100720 218074
rect 100668 218010 100720 218016
rect 101508 217002 101536 221818
rect 102060 217002 102088 223518
rect 103256 217002 103284 227394
rect 104624 222012 104676 222018
rect 104624 221954 104676 221960
rect 103980 218068 104032 218074
rect 103980 218010 104032 218016
rect 103992 217002 104020 218010
rect 104636 217002 104664 221954
rect 104820 218074 104848 230726
rect 106922 230344 106978 230353
rect 106922 230279 106978 230288
rect 106188 228676 106240 228682
rect 106188 228618 106240 228624
rect 105728 224664 105780 224670
rect 105728 224606 105780 224612
rect 104808 218068 104860 218074
rect 104808 218010 104860 218016
rect 105740 217002 105768 224606
rect 106200 217002 106228 228618
rect 106936 219026 106964 230279
rect 126888 230172 126940 230178
rect 126888 230114 126940 230120
rect 117228 229900 117280 229906
rect 117228 229842 117280 229848
rect 110328 229764 110380 229770
rect 110328 229706 110380 229712
rect 109868 227588 109920 227594
rect 109868 227530 109920 227536
rect 108946 222048 109002 222057
rect 108946 221983 109002 221992
rect 108120 220788 108172 220794
rect 108120 220730 108172 220736
rect 106924 219020 106976 219026
rect 106924 218962 106976 218968
rect 107292 219020 107344 219026
rect 107292 218962 107344 218968
rect 107304 217002 107332 218962
rect 108132 217002 108160 220730
rect 108304 219428 108356 219434
rect 108304 219370 108356 219376
rect 108316 218890 108344 219370
rect 108304 218884 108356 218890
rect 108304 218826 108356 218832
rect 108960 217002 108988 221983
rect 109880 217002 109908 227530
rect 110340 217002 110368 229706
rect 113086 228848 113142 228857
rect 113086 228783 113142 228792
rect 112904 224800 112956 224806
rect 112904 224742 112956 224748
rect 111432 222148 111484 222154
rect 111432 222090 111484 222096
rect 111444 217002 111472 222090
rect 112916 218074 112944 224742
rect 112260 218068 112312 218074
rect 112260 218010 112312 218016
rect 112904 218068 112956 218074
rect 112904 218010 112956 218016
rect 112272 217002 112300 218010
rect 113100 217002 113128 228783
rect 117044 227724 117096 227730
rect 117044 227666 117096 227672
rect 115664 224120 115716 224126
rect 115664 224062 115716 224068
rect 114468 219972 114520 219978
rect 114468 219914 114520 219920
rect 113916 219020 113968 219026
rect 113916 218962 113968 218968
rect 113928 217002 113956 218962
rect 114480 217002 114508 219914
rect 115676 217002 115704 224062
rect 117056 218074 117084 227666
rect 116400 218068 116452 218074
rect 116400 218010 116452 218016
rect 117044 218068 117096 218074
rect 117044 218010 117096 218016
rect 116412 217002 116440 218010
rect 117240 217002 117268 229842
rect 126428 229084 126480 229090
rect 126428 229026 126480 229032
rect 119804 228948 119856 228954
rect 119804 228890 119856 228896
rect 118608 224936 118660 224942
rect 118608 224878 118660 224884
rect 118054 220144 118110 220153
rect 118054 220079 118110 220088
rect 118068 217002 118096 220079
rect 118620 217002 118648 224878
rect 119816 217002 119844 228890
rect 122748 226908 122800 226914
rect 122748 226850 122800 226856
rect 122288 223984 122340 223990
rect 122288 223926 122340 223932
rect 121368 221332 121420 221338
rect 121368 221274 121420 221280
rect 120540 218612 120592 218618
rect 120540 218554 120592 218560
rect 120552 217002 120580 218554
rect 121380 217002 121408 221274
rect 122300 217002 122328 223926
rect 122760 217002 122788 226850
rect 125506 226128 125562 226137
rect 125506 226063 125562 226072
rect 124678 220416 124734 220425
rect 124678 220351 124734 220360
rect 123852 219156 123904 219162
rect 123852 219098 123904 219104
rect 123864 217002 123892 219098
rect 124692 217002 124720 220351
rect 125520 217002 125548 226063
rect 126440 217002 126468 229026
rect 126900 217002 126928 230114
rect 129464 226772 129516 226778
rect 129464 226714 129516 226720
rect 127992 219836 128044 219842
rect 127992 219778 128044 219784
rect 128004 217002 128032 219778
rect 128636 218068 128688 218074
rect 128636 218010 128688 218016
rect 128648 217002 128676 218010
rect 129476 217002 129504 226714
rect 129660 218074 129688 230862
rect 133696 230308 133748 230314
rect 133696 230250 133748 230256
rect 133708 229094 133736 230250
rect 133880 229356 133932 229362
rect 133880 229298 133932 229304
rect 133892 229094 133920 229298
rect 133708 229066 133828 229094
rect 133892 229066 134012 229094
rect 133604 228268 133656 228274
rect 133604 228210 133656 228216
rect 132224 225480 132276 225486
rect 132224 225422 132276 225428
rect 131028 222760 131080 222766
rect 131028 222702 131080 222708
rect 130476 218204 130528 218210
rect 130476 218146 130528 218152
rect 129648 218068 129700 218074
rect 129648 218010 129700 218016
rect 130488 217002 130516 218146
rect 131040 217002 131068 222702
rect 132236 217002 132264 225422
rect 133616 218074 133644 228210
rect 132960 218068 133012 218074
rect 132960 218010 133012 218016
rect 133604 218068 133656 218074
rect 133604 218010 133656 218016
rect 132972 217002 133000 218010
rect 133800 217002 133828 229066
rect 133984 226302 134012 229066
rect 141160 228410 141188 231676
rect 141148 228404 141200 228410
rect 141148 228346 141200 228352
rect 139308 228132 139360 228138
rect 139308 228074 139360 228080
rect 136362 227488 136418 227497
rect 136362 227423 136418 227432
rect 133972 226296 134024 226302
rect 133972 226238 134024 226244
rect 135168 226296 135220 226302
rect 135168 226238 135220 226244
rect 134708 222488 134760 222494
rect 134708 222430 134760 222436
rect 134720 217002 134748 222430
rect 135180 217002 135208 226238
rect 136376 217002 136404 227423
rect 138848 225344 138900 225350
rect 138848 225286 138900 225292
rect 137928 219700 137980 219706
rect 137928 219642 137980 219648
rect 137100 218476 137152 218482
rect 137100 218418 137152 218424
rect 137112 217002 137140 218418
rect 137940 217002 137968 219642
rect 138860 217002 138888 225286
rect 139320 217002 139348 228074
rect 140504 227996 140556 228002
rect 140504 227938 140556 227944
rect 140044 223848 140096 223854
rect 140044 223790 140096 223796
rect 140056 219298 140084 223790
rect 140044 219292 140096 219298
rect 140044 219234 140096 219240
rect 140516 217002 140544 227938
rect 141804 225758 141832 231676
rect 142448 227050 142476 231676
rect 143092 228585 143120 231676
rect 143078 228576 143134 228585
rect 143078 228511 143134 228520
rect 143172 227860 143224 227866
rect 143172 227802 143224 227808
rect 142436 227044 142488 227050
rect 142436 226986 142488 226992
rect 141792 225752 141844 225758
rect 141792 225694 141844 225700
rect 142068 225752 142120 225758
rect 142068 225694 142120 225700
rect 141240 221060 141292 221066
rect 141240 221002 141292 221008
rect 141252 217002 141280 221002
rect 142080 217002 142108 225694
rect 142896 218068 142948 218074
rect 142896 218010 142948 218016
rect 142908 217002 142936 218010
rect 97736 216974 97888 217002
rect 98716 216974 99144 217002
rect 99544 216974 99880 217002
rect 100372 216974 100524 217002
rect 101200 216974 101536 217002
rect 102028 216974 102088 217002
rect 102856 216974 103284 217002
rect 103684 216974 104020 217002
rect 104512 216974 104664 217002
rect 105340 216974 105768 217002
rect 106168 216974 106228 217002
rect 106996 216974 107332 217002
rect 107824 216974 108160 217002
rect 108652 216974 108988 217002
rect 109480 216974 109908 217002
rect 110308 216974 110368 217002
rect 111136 216974 111472 217002
rect 111964 216974 112300 217002
rect 112792 216974 113128 217002
rect 113620 216974 113956 217002
rect 114448 216974 114508 217002
rect 115276 216974 115704 217002
rect 116104 216974 116440 217002
rect 116932 216974 117268 217002
rect 117760 216974 118096 217002
rect 118588 216974 118648 217002
rect 119416 216974 119844 217002
rect 120244 216974 120580 217002
rect 121072 216974 121408 217002
rect 121900 216974 122328 217002
rect 122728 216974 122788 217002
rect 123556 216974 123892 217002
rect 124384 216974 124720 217002
rect 125212 216974 125548 217002
rect 126040 216974 126468 217002
rect 126868 216974 126928 217002
rect 127696 216974 128032 217002
rect 128524 216974 128676 217002
rect 129352 216974 129504 217002
rect 130180 216974 130516 217002
rect 131008 216974 131068 217002
rect 131836 216974 132264 217002
rect 132664 216974 133000 217002
rect 133492 216974 133828 217002
rect 134320 216974 134748 217002
rect 135148 216974 135208 217002
rect 135976 216974 136404 217002
rect 136804 216974 137140 217002
rect 137632 216974 137968 217002
rect 138460 216974 138888 217002
rect 139288 216974 139348 217002
rect 140116 216974 140544 217002
rect 140944 216974 141280 217002
rect 141772 216974 142108 217002
rect 142600 216974 142936 217002
rect 143184 217002 143212 227802
rect 143736 227186 143764 231676
rect 144184 229492 144236 229498
rect 144184 229434 144236 229440
rect 143724 227180 143776 227186
rect 143724 227122 143776 227128
rect 143356 227044 143408 227050
rect 143356 226986 143408 226992
rect 143368 218074 143396 226986
rect 144196 220658 144224 229434
rect 144380 225622 144408 231676
rect 144368 225616 144420 225622
rect 144368 225558 144420 225564
rect 145024 224233 145052 231676
rect 145668 229226 145696 231676
rect 146312 229362 146340 231676
rect 146680 231662 146970 231690
rect 146300 229356 146352 229362
rect 146300 229298 146352 229304
rect 145656 229220 145708 229226
rect 145656 229162 145708 229168
rect 146208 229220 146260 229226
rect 146208 229162 146260 229168
rect 146024 228404 146076 228410
rect 146024 228346 146076 228352
rect 145010 224224 145066 224233
rect 145010 224159 145066 224168
rect 146036 223938 146064 228346
rect 146220 228002 146248 229162
rect 146208 227996 146260 228002
rect 146208 227938 146260 227944
rect 146036 223910 146248 223938
rect 146024 222624 146076 222630
rect 146024 222566 146076 222572
rect 144184 220652 144236 220658
rect 144184 220594 144236 220600
rect 144552 220652 144604 220658
rect 144552 220594 144604 220600
rect 143356 218068 143408 218074
rect 143356 218010 143408 218016
rect 144564 217002 144592 220594
rect 146036 218074 146064 222566
rect 145380 218068 145432 218074
rect 145380 218010 145432 218016
rect 146024 218068 146076 218074
rect 146024 218010 146076 218016
rect 145392 217002 145420 218010
rect 146220 217002 146248 223910
rect 146680 222873 146708 231662
rect 147600 224262 147628 231676
rect 148244 229809 148272 231676
rect 148230 229800 148286 229809
rect 148230 229735 148286 229744
rect 148888 229498 148916 231676
rect 148876 229492 148928 229498
rect 148876 229434 148928 229440
rect 148692 229356 148744 229362
rect 148692 229298 148744 229304
rect 148704 227866 148732 229298
rect 148692 227860 148744 227866
rect 148692 227802 148744 227808
rect 147588 224256 147640 224262
rect 147588 224198 147640 224204
rect 146850 223952 146906 223961
rect 146850 223887 146906 223896
rect 146666 222864 146722 222873
rect 146666 222799 146722 222808
rect 146864 219434 146892 223887
rect 149532 222902 149560 231676
rect 149808 231662 150190 231690
rect 149808 224505 149836 231662
rect 150820 230081 150848 231676
rect 150806 230072 150862 230081
rect 150806 230007 150862 230016
rect 150440 229492 150492 229498
rect 150440 229434 150492 229440
rect 150072 226636 150124 226642
rect 150072 226578 150124 226584
rect 149794 224496 149850 224505
rect 149794 224431 149850 224440
rect 149520 222896 149572 222902
rect 149520 222838 149572 222844
rect 148692 221196 148744 221202
rect 148692 221138 148744 221144
rect 147586 220688 147642 220697
rect 147586 220623 147642 220632
rect 146852 219428 146904 219434
rect 146852 219370 146904 219376
rect 147036 219292 147088 219298
rect 147036 219234 147088 219240
rect 147048 217002 147076 219234
rect 147600 217002 147628 220623
rect 148704 217002 148732 221138
rect 150084 218074 150112 226578
rect 150452 223530 150480 229434
rect 151464 225894 151492 231676
rect 151452 225888 151504 225894
rect 151452 225830 151504 225836
rect 151728 224256 151780 224262
rect 151728 224198 151780 224204
rect 150268 223502 150480 223530
rect 149520 218068 149572 218074
rect 149520 218010 149572 218016
rect 150072 218068 150124 218074
rect 150072 218010 150124 218016
rect 149532 217002 149560 218010
rect 150268 217002 150296 223502
rect 151266 222864 151322 222873
rect 151266 222799 151322 222808
rect 151280 217002 151308 222799
rect 151740 217002 151768 224198
rect 152108 223145 152136 231676
rect 152752 224777 152780 231676
rect 153410 231662 153608 231690
rect 153580 229094 153608 231662
rect 153488 229066 153608 229094
rect 153764 231662 154054 231690
rect 152924 227996 152976 228002
rect 152924 227938 152976 227944
rect 152738 224768 152794 224777
rect 152738 224703 152794 224712
rect 152094 223136 152150 223145
rect 152094 223071 152150 223080
rect 152936 217002 152964 227938
rect 153488 218657 153516 229066
rect 153764 220114 153792 231662
rect 154304 223168 154356 223174
rect 154304 223110 154356 223116
rect 154316 222358 154344 223110
rect 154684 223038 154712 231676
rect 155328 228313 155356 231676
rect 155972 230042 156000 231676
rect 156156 231662 156630 231690
rect 155960 230036 156012 230042
rect 155960 229978 156012 229984
rect 155314 228304 155370 228313
rect 155314 228239 155370 228248
rect 155776 225888 155828 225894
rect 155776 225830 155828 225836
rect 155592 225208 155644 225214
rect 155592 225150 155644 225156
rect 154672 223032 154724 223038
rect 154672 222974 154724 222980
rect 154488 222896 154540 222902
rect 154488 222838 154540 222844
rect 154304 222352 154356 222358
rect 154304 222294 154356 222300
rect 153752 220108 153804 220114
rect 153752 220050 153804 220056
rect 153660 219428 153712 219434
rect 153660 219370 153712 219376
rect 153474 218648 153530 218657
rect 153474 218583 153530 218592
rect 153672 217002 153700 219370
rect 154500 217002 154528 222838
rect 155316 218068 155368 218074
rect 155316 218010 155368 218016
rect 155328 217002 155356 218010
rect 143184 216974 143428 217002
rect 144256 216974 144592 217002
rect 145084 216974 145420 217002
rect 145912 216974 146248 217002
rect 146740 216974 147076 217002
rect 147568 216974 147628 217002
rect 148396 216974 148732 217002
rect 149224 216974 149560 217002
rect 150052 216974 150296 217002
rect 150880 216974 151308 217002
rect 151708 216974 151768 217002
rect 152536 216974 152964 217002
rect 153364 216974 153700 217002
rect 154192 216974 154528 217002
rect 155020 216974 155356 217002
rect 155604 217002 155632 225150
rect 155788 218074 155816 225830
rect 156156 220250 156184 231662
rect 156604 227180 156656 227186
rect 156604 227122 156656 227128
rect 156616 226642 156644 227122
rect 156604 226636 156656 226642
rect 156604 226578 156656 226584
rect 157064 223304 157116 223310
rect 157064 223246 157116 223252
rect 156144 220244 156196 220250
rect 156144 220186 156196 220192
rect 155776 218068 155828 218074
rect 155776 218010 155828 218016
rect 157076 217002 157104 223246
rect 157260 223174 157288 231676
rect 157904 229094 157932 231676
rect 158180 231662 158562 231690
rect 158916 231662 159206 231690
rect 158180 229094 158208 231662
rect 157812 229066 157932 229094
rect 157996 229066 158208 229094
rect 157812 224398 157840 229066
rect 157800 224392 157852 224398
rect 157800 224334 157852 224340
rect 157996 223394 158024 229066
rect 158444 225616 158496 225622
rect 158444 225558 158496 225564
rect 157536 223366 158024 223394
rect 157248 223168 157300 223174
rect 157248 223110 157300 223116
rect 157536 218929 157564 223366
rect 157800 220108 157852 220114
rect 157800 220050 157852 220056
rect 157522 218920 157578 218929
rect 157522 218855 157578 218864
rect 157812 217002 157840 220050
rect 158456 217002 158484 225558
rect 158916 220386 158944 231662
rect 159272 223168 159324 223174
rect 159272 223110 159324 223116
rect 158904 220380 158956 220386
rect 158904 220322 158956 220328
rect 159284 218890 159312 223110
rect 159836 222358 159864 231676
rect 160192 230036 160244 230042
rect 160192 229978 160244 229984
rect 160008 226636 160060 226642
rect 160008 226578 160060 226584
rect 159824 222352 159876 222358
rect 159824 222294 159876 222300
rect 159272 218884 159324 218890
rect 159272 218826 159324 218832
rect 159824 218340 159876 218346
rect 159824 218282 159876 218288
rect 159456 218068 159508 218074
rect 159456 218010 159508 218016
rect 159468 217002 159496 218010
rect 155604 216974 155848 217002
rect 156676 216974 157104 217002
rect 157504 216974 157840 217002
rect 158332 216974 158484 217002
rect 159160 216974 159496 217002
rect 159836 217002 159864 218282
rect 160020 218074 160048 226578
rect 160204 223310 160232 229978
rect 160480 226953 160508 231676
rect 161124 229634 161152 231676
rect 161112 229628 161164 229634
rect 161112 229570 161164 229576
rect 161296 229628 161348 229634
rect 161296 229570 161348 229576
rect 160466 226944 160522 226953
rect 160466 226879 160522 226888
rect 160192 223304 160244 223310
rect 160192 223246 160244 223252
rect 161308 219434 161336 229570
rect 161768 226030 161796 231676
rect 162044 231662 162426 231690
rect 161756 226024 161808 226030
rect 161756 225966 161808 225972
rect 161480 221740 161532 221746
rect 161480 221682 161532 221688
rect 161492 220930 161520 221682
rect 162044 221610 162072 231662
rect 163056 225593 163084 231676
rect 163240 231662 163714 231690
rect 163042 225584 163098 225593
rect 163042 225519 163098 225528
rect 162032 221604 162084 221610
rect 162032 221546 162084 221552
rect 161940 221468 161992 221474
rect 161940 221410 161992 221416
rect 161480 220924 161532 220930
rect 161480 220866 161532 220872
rect 161480 220244 161532 220250
rect 161480 220186 161532 220192
rect 160744 219428 161336 219434
rect 160796 219406 161336 219428
rect 160744 219370 160796 219376
rect 160192 218748 160244 218754
rect 160192 218690 160244 218696
rect 160204 218074 160232 218690
rect 161492 218090 161520 220186
rect 160008 218068 160060 218074
rect 160008 218010 160060 218016
rect 160192 218068 160244 218074
rect 160192 218010 160244 218016
rect 161216 218062 161520 218090
rect 161216 217002 161244 218062
rect 161952 217002 161980 221410
rect 162768 218748 162820 218754
rect 162768 218690 162820 218696
rect 162780 217002 162808 218690
rect 163240 218074 163268 231662
rect 164056 223032 164108 223038
rect 164056 222974 164108 222980
rect 163596 219428 163648 219434
rect 163596 219370 163648 219376
rect 163228 218068 163280 218074
rect 163228 218010 163280 218016
rect 163608 217002 163636 219370
rect 159836 216974 159988 217002
rect 160816 216974 161244 217002
rect 161644 216974 161980 217002
rect 162472 216974 162808 217002
rect 163300 216974 163636 217002
rect 164068 217002 164096 222974
rect 164344 220522 164372 231676
rect 164988 223446 165016 231676
rect 165632 224534 165660 231676
rect 166276 230353 166304 231676
rect 166262 230344 166318 230353
rect 166262 230279 166318 230288
rect 166920 227225 166948 231676
rect 167288 231662 167578 231690
rect 166906 227216 166962 227225
rect 166906 227151 166962 227160
rect 166080 225072 166132 225078
rect 166080 225014 166132 225020
rect 165620 224528 165672 224534
rect 165620 224470 165672 224476
rect 165344 224392 165396 224398
rect 165344 224334 165396 224340
rect 164976 223440 165028 223446
rect 164976 223382 165028 223388
rect 164332 220516 164384 220522
rect 164332 220458 164384 220464
rect 165356 217002 165384 224334
rect 166092 219026 166120 225014
rect 166448 223440 166500 223446
rect 166448 223382 166500 223388
rect 166080 219020 166132 219026
rect 166080 218962 166132 218968
rect 166460 218618 166488 223382
rect 167288 221746 167316 231662
rect 168208 225865 168236 231676
rect 168852 230518 168880 231676
rect 168840 230512 168892 230518
rect 168840 230454 168892 230460
rect 169496 228546 169524 231676
rect 169772 231662 170154 231690
rect 169484 228540 169536 228546
rect 169484 228482 169536 228488
rect 169022 228304 169078 228313
rect 169022 228239 169078 228248
rect 168194 225856 168250 225865
rect 168194 225791 168250 225800
rect 167550 224224 167606 224233
rect 167550 224159 167606 224168
rect 167276 221740 167328 221746
rect 167276 221682 167328 221688
rect 166632 219020 166684 219026
rect 166632 218962 166684 218968
rect 166448 218612 166500 218618
rect 166448 218554 166500 218560
rect 166644 218074 166672 218962
rect 166906 218648 166962 218657
rect 166906 218583 166962 218592
rect 166080 218068 166132 218074
rect 166080 218010 166132 218016
rect 166632 218068 166684 218074
rect 166632 218010 166684 218016
rect 166092 217002 166120 218010
rect 166920 217002 166948 218583
rect 167564 218210 167592 224159
rect 168288 223168 168340 223174
rect 168288 223110 168340 223116
rect 167552 218204 167604 218210
rect 167552 218146 167604 218152
rect 168104 218204 168156 218210
rect 168104 218146 168156 218152
rect 167736 218068 167788 218074
rect 167736 218010 167788 218016
rect 167748 217002 167776 218010
rect 164068 216974 164128 217002
rect 164956 216974 165384 217002
rect 165784 216974 166120 217002
rect 166612 216974 166948 217002
rect 167440 216974 167776 217002
rect 168116 217002 168144 218146
rect 168300 218074 168328 223110
rect 169036 218754 169064 228239
rect 169484 227860 169536 227866
rect 169484 227802 169536 227808
rect 169024 218748 169076 218754
rect 169024 218690 169076 218696
rect 168288 218068 168340 218074
rect 168288 218010 168340 218016
rect 169496 217002 169524 227802
rect 169772 220930 169800 231662
rect 169944 228540 169996 228546
rect 169944 228482 169996 228488
rect 169956 227866 169984 228482
rect 169944 227860 169996 227866
rect 169944 227802 169996 227808
rect 170784 223417 170812 231676
rect 171428 223854 171456 231676
rect 172072 227322 172100 231676
rect 172060 227316 172112 227322
rect 172060 227258 172112 227264
rect 172336 224528 172388 224534
rect 172336 224470 172388 224476
rect 171416 223848 171468 223854
rect 171416 223790 171468 223796
rect 170770 223408 170826 223417
rect 170770 223343 170826 223352
rect 170586 221232 170642 221241
rect 170586 221167 170642 221176
rect 169760 220924 169812 220930
rect 169760 220866 169812 220872
rect 170220 218612 170272 218618
rect 170220 218554 170272 218560
rect 170232 217002 170260 218554
rect 170600 218210 170628 221167
rect 171048 220380 171100 220386
rect 171048 220322 171100 220328
rect 170588 218204 170640 218210
rect 170588 218146 170640 218152
rect 171060 217002 171088 220322
rect 172152 218204 172204 218210
rect 172152 218146 172204 218152
rect 171876 218068 171928 218074
rect 171876 218010 171928 218016
rect 171888 217002 171916 218010
rect 168116 216974 168268 217002
rect 169096 216974 169524 217002
rect 169924 216974 170260 217002
rect 170752 216974 171088 217002
rect 171580 216974 171916 217002
rect 172164 217002 172192 218146
rect 172348 218074 172376 224470
rect 172716 221785 172744 231676
rect 172992 231662 173374 231690
rect 172702 221776 172758 221785
rect 172702 221711 172758 221720
rect 172992 221513 173020 231662
rect 174004 230654 174032 231676
rect 173992 230648 174044 230654
rect 173992 230590 174044 230596
rect 174648 228818 174676 231676
rect 175306 231662 175504 231690
rect 174636 228812 174688 228818
rect 174636 228754 174688 228760
rect 173164 227316 173216 227322
rect 173164 227258 173216 227264
rect 172978 221504 173034 221513
rect 172978 221439 173034 221448
rect 172520 220924 172572 220930
rect 172520 220866 172572 220872
rect 172532 218890 172560 220866
rect 173176 219026 173204 227258
rect 175188 223848 175240 223854
rect 175188 223790 175240 223796
rect 173164 219020 173216 219026
rect 173164 218962 173216 218968
rect 173532 219020 173584 219026
rect 173532 218962 173584 218968
rect 172520 218884 172572 218890
rect 172520 218826 172572 218832
rect 172336 218068 172388 218074
rect 172336 218010 172388 218016
rect 173544 217002 173572 218962
rect 174912 218884 174964 218890
rect 174912 218826 174964 218832
rect 174360 218748 174412 218754
rect 174360 218690 174412 218696
rect 174372 217002 174400 218690
rect 174924 218482 174952 218826
rect 174912 218476 174964 218482
rect 174912 218418 174964 218424
rect 175200 217002 175228 223790
rect 175476 221882 175504 231662
rect 175936 226166 175964 231676
rect 176304 231662 176594 231690
rect 175924 226160 175976 226166
rect 175924 226102 175976 226108
rect 176304 223961 176332 231662
rect 176476 228812 176528 228818
rect 176476 228754 176528 228760
rect 176290 223952 176346 223961
rect 176290 223887 176346 223896
rect 175464 221876 175516 221882
rect 175464 221818 175516 221824
rect 176292 218476 176344 218482
rect 176292 218418 176344 218424
rect 176016 218068 176068 218074
rect 176016 218010 176068 218016
rect 176028 217002 176056 218010
rect 172164 216974 172408 217002
rect 173236 216974 173572 217002
rect 174064 216974 174400 217002
rect 174892 216974 175228 217002
rect 175720 216974 176056 217002
rect 176304 217002 176332 218418
rect 176488 218074 176516 228754
rect 177224 227458 177252 231676
rect 177408 231662 177882 231690
rect 177408 229094 177436 231662
rect 177408 229066 177528 229094
rect 177212 227452 177264 227458
rect 177212 227394 177264 227400
rect 177304 226500 177356 226506
rect 177304 226442 177356 226448
rect 177316 218210 177344 226442
rect 177500 222018 177528 229066
rect 178512 223582 178540 231676
rect 179156 230790 179184 231676
rect 179144 230784 179196 230790
rect 179144 230726 179196 230732
rect 179800 228682 179828 231676
rect 179984 231662 180458 231690
rect 179788 228676 179840 228682
rect 179788 228618 179840 228624
rect 178500 223576 178552 223582
rect 178500 223518 178552 223524
rect 178684 222352 178736 222358
rect 178684 222294 178736 222300
rect 177488 222012 177540 222018
rect 177488 221954 177540 221960
rect 177672 221740 177724 221746
rect 177672 221682 177724 221688
rect 177304 218204 177356 218210
rect 177304 218146 177356 218152
rect 176476 218068 176528 218074
rect 176476 218010 176528 218016
rect 177684 217002 177712 221682
rect 178500 221604 178552 221610
rect 178500 221546 178552 221552
rect 178512 217002 178540 221546
rect 178696 218890 178724 222294
rect 179984 220794 180012 231662
rect 181088 224670 181116 231676
rect 181076 224664 181128 224670
rect 181076 224606 181128 224612
rect 181732 223310 181760 231676
rect 182376 227594 182404 231676
rect 182560 231662 183034 231690
rect 182364 227588 182416 227594
rect 182364 227530 182416 227536
rect 181904 223712 181956 223718
rect 181904 223654 181956 223660
rect 181720 223304 181772 223310
rect 181720 223246 181772 223252
rect 179972 220788 180024 220794
rect 179972 220730 180024 220736
rect 180708 220516 180760 220522
rect 180708 220458 180760 220464
rect 179512 219564 179564 219570
rect 179512 219506 179564 219512
rect 179328 219020 179380 219026
rect 179328 218962 179380 218968
rect 178684 218884 178736 218890
rect 178684 218826 178736 218832
rect 179340 217002 179368 218962
rect 179524 218754 179552 219506
rect 179512 218748 179564 218754
rect 179512 218690 179564 218696
rect 180156 218748 180208 218754
rect 180156 218690 180208 218696
rect 180168 217002 180196 218690
rect 180720 217002 180748 220458
rect 181916 217002 181944 223654
rect 182560 222154 182588 231662
rect 183468 228676 183520 228682
rect 183468 228618 183520 228624
rect 182824 227588 182876 227594
rect 182824 227530 182876 227536
rect 182548 222148 182600 222154
rect 182548 222090 182600 222096
rect 182836 219026 182864 227530
rect 183100 219156 183152 219162
rect 183100 219098 183152 219104
rect 182824 219020 182876 219026
rect 182824 218962 182876 218968
rect 183112 218482 183140 219098
rect 183100 218476 183152 218482
rect 183100 218418 183152 218424
rect 183284 218476 183336 218482
rect 183284 218418 183336 218424
rect 182640 218068 182692 218074
rect 182640 218010 182692 218016
rect 182652 217002 182680 218010
rect 183296 217002 183324 218418
rect 183480 218074 183508 228618
rect 183664 222057 183692 231676
rect 184308 229770 184336 231676
rect 184296 229764 184348 229770
rect 184296 229706 184348 229712
rect 184480 229764 184532 229770
rect 184480 229706 184532 229712
rect 184020 222148 184072 222154
rect 184020 222090 184072 222096
rect 183650 222048 183706 222057
rect 183650 221983 183706 221992
rect 183468 218068 183520 218074
rect 183468 218010 183520 218016
rect 184032 217002 184060 222090
rect 184492 219434 184520 229706
rect 184952 228857 184980 231676
rect 185136 231662 185610 231690
rect 185872 231662 186254 231690
rect 184938 228848 184994 228857
rect 184938 228783 184994 228792
rect 185136 219978 185164 231662
rect 185400 227452 185452 227458
rect 185400 227394 185452 227400
rect 185412 226914 185440 227394
rect 185584 227316 185636 227322
rect 185584 227258 185636 227264
rect 185596 226914 185624 227258
rect 185400 226908 185452 226914
rect 185400 226850 185452 226856
rect 185584 226908 185636 226914
rect 185584 226850 185636 226856
rect 185584 224936 185636 224942
rect 185584 224878 185636 224884
rect 185596 223718 185624 224878
rect 185872 224806 185900 231662
rect 186044 226024 186096 226030
rect 186044 225966 186096 225972
rect 185860 224800 185912 224806
rect 185860 224742 185912 224748
rect 185768 224664 185820 224670
rect 185768 224606 185820 224612
rect 185584 223712 185636 223718
rect 185584 223654 185636 223660
rect 185124 219972 185176 219978
rect 185124 219914 185176 219920
rect 185780 219434 185808 224606
rect 184204 219428 184520 219434
rect 184256 219406 184520 219428
rect 185596 219406 185808 219434
rect 184204 219370 184256 219376
rect 185596 218074 185624 219406
rect 184848 218068 184900 218074
rect 184848 218010 184900 218016
rect 185584 218068 185636 218074
rect 185584 218010 185636 218016
rect 184860 217002 184888 218010
rect 186056 217002 186084 225966
rect 186884 225078 186912 231676
rect 187528 227730 187556 231676
rect 187896 231662 188186 231690
rect 187516 227724 187568 227730
rect 187516 227666 187568 227672
rect 186872 225072 186924 225078
rect 186872 225014 186924 225020
rect 186320 224664 186372 224670
rect 186320 224606 186372 224612
rect 186332 223582 186360 224606
rect 186320 223576 186372 223582
rect 186320 223518 186372 223524
rect 187608 220788 187660 220794
rect 187608 220730 187660 220736
rect 186780 219020 186832 219026
rect 186780 218962 186832 218968
rect 186792 217002 186820 218962
rect 187620 217002 187648 220730
rect 187896 220153 187924 231662
rect 188816 224126 188844 231676
rect 189460 229906 189488 231676
rect 189448 229900 189500 229906
rect 189448 229842 189500 229848
rect 189724 229900 189776 229906
rect 189724 229842 189776 229848
rect 188988 227316 189040 227322
rect 188988 227258 189040 227264
rect 188804 224120 188856 224126
rect 188804 224062 188856 224068
rect 187882 220144 187938 220153
rect 187882 220079 187938 220088
rect 188436 218068 188488 218074
rect 188436 218010 188488 218016
rect 188448 217002 188476 218010
rect 189000 217002 189028 227258
rect 189448 221876 189500 221882
rect 189448 221818 189500 221824
rect 189460 218074 189488 221818
rect 189736 219162 189764 229842
rect 190104 228954 190132 231676
rect 190656 231662 190762 231690
rect 191024 231662 191406 231690
rect 190092 228948 190144 228954
rect 190092 228890 190144 228896
rect 189908 224120 189960 224126
rect 189908 224062 189960 224068
rect 189920 219298 189948 224062
rect 190656 221338 190684 231662
rect 191024 223718 191052 231662
rect 191472 224936 191524 224942
rect 191472 224878 191524 224884
rect 191012 223712 191064 223718
rect 191012 223654 191064 223660
rect 190644 221332 190696 221338
rect 190644 221274 190696 221280
rect 189908 219292 189960 219298
rect 189908 219234 189960 219240
rect 189724 219156 189776 219162
rect 189724 219098 189776 219104
rect 190092 218204 190144 218210
rect 190092 218146 190144 218152
rect 189448 218068 189500 218074
rect 189448 218010 189500 218016
rect 190104 217002 190132 218146
rect 190920 218068 190972 218074
rect 190920 218010 190972 218016
rect 190932 217002 190960 218010
rect 191484 217002 191512 224878
rect 192036 223446 192064 231676
rect 192680 227458 192708 231676
rect 193128 228948 193180 228954
rect 193128 228890 193180 228896
rect 192668 227452 192720 227458
rect 192668 227394 192720 227400
rect 192024 223440 192076 223446
rect 192024 223382 192076 223388
rect 191656 223304 191708 223310
rect 191656 223246 191708 223252
rect 191668 218074 191696 223246
rect 192944 219428 192996 219434
rect 192944 219370 192996 219376
rect 191656 218068 191708 218074
rect 191656 218010 191708 218016
rect 192576 218068 192628 218074
rect 192576 218010 192628 218016
rect 192588 217002 192616 218010
rect 176304 216974 176548 217002
rect 177376 216974 177712 217002
rect 178204 216974 178540 217002
rect 179032 216974 179368 217002
rect 179860 216974 180196 217002
rect 180688 216974 180748 217002
rect 181516 216974 181944 217002
rect 182344 216974 182680 217002
rect 183172 216974 183324 217002
rect 184000 216974 184060 217002
rect 184828 216974 184888 217002
rect 185656 216974 186084 217002
rect 186484 216974 186820 217002
rect 187312 216974 187648 217002
rect 188140 216974 188476 217002
rect 188968 216974 189028 217002
rect 189796 216974 190132 217002
rect 190624 216974 190960 217002
rect 191452 216974 191512 217002
rect 192280 216974 192616 217002
rect 192956 217002 192984 219370
rect 193140 218074 193168 228890
rect 193324 220425 193352 231676
rect 193968 223990 193996 231676
rect 194626 231662 195008 231690
rect 193956 223984 194008 223990
rect 193956 223926 194008 223932
rect 194324 223576 194376 223582
rect 194324 223518 194376 223524
rect 193310 220416 193366 220425
rect 193310 220351 193366 220360
rect 193128 218068 193180 218074
rect 193128 218010 193180 218016
rect 194336 217002 194364 223518
rect 194980 220930 195008 231662
rect 195256 229090 195284 231676
rect 195624 231662 195914 231690
rect 195244 229084 195296 229090
rect 195244 229026 195296 229032
rect 195152 222012 195204 222018
rect 195152 221954 195204 221960
rect 194968 220924 195020 220930
rect 194968 220866 195020 220872
rect 195164 217002 195192 221954
rect 195624 219842 195652 231662
rect 196072 230444 196124 230450
rect 196072 230386 196124 230392
rect 195888 225072 195940 225078
rect 195888 225014 195940 225020
rect 195612 219836 195664 219842
rect 195612 219778 195664 219784
rect 195900 217002 195928 225014
rect 196084 222766 196112 230386
rect 196544 226137 196572 231676
rect 197188 230178 197216 231676
rect 197176 230172 197228 230178
rect 197176 230114 197228 230120
rect 197452 230172 197504 230178
rect 197452 230114 197504 230120
rect 196530 226128 196586 226137
rect 196530 226063 196586 226072
rect 196808 223984 196860 223990
rect 196808 223926 196860 223932
rect 196072 222760 196124 222766
rect 196072 222702 196124 222708
rect 196820 218346 196848 223926
rect 197268 223440 197320 223446
rect 197268 223382 197320 223388
rect 196808 218340 196860 218346
rect 196808 218282 196860 218288
rect 196716 218068 196768 218074
rect 196716 218010 196768 218016
rect 196728 217002 196756 218010
rect 197280 217002 197308 223382
rect 197464 222494 197492 230114
rect 197832 226778 197860 231676
rect 198476 230450 198504 231676
rect 199120 230926 199148 231676
rect 199108 230920 199160 230926
rect 199108 230862 199160 230868
rect 198464 230444 198516 230450
rect 198464 230386 198516 230392
rect 198464 227452 198516 227458
rect 198464 227394 198516 227400
rect 197820 226772 197872 226778
rect 197820 226714 197872 226720
rect 197452 222488 197504 222494
rect 197452 222430 197504 222436
rect 198476 217002 198504 227394
rect 199764 224233 199792 231676
rect 200408 228274 200436 231676
rect 201052 230178 201080 231676
rect 201040 230172 201092 230178
rect 201040 230114 201092 230120
rect 200396 228268 200448 228274
rect 200396 228210 200448 228216
rect 200672 227860 200724 227866
rect 200672 227802 200724 227808
rect 200028 227724 200080 227730
rect 200028 227666 200080 227672
rect 199750 224224 199806 224233
rect 199750 224159 199806 224168
rect 199844 219156 199896 219162
rect 199844 219098 199896 219104
rect 199200 218340 199252 218346
rect 199200 218282 199252 218288
rect 199212 217002 199240 218282
rect 199856 217002 199884 219098
rect 200040 218346 200068 227666
rect 200684 218618 200712 227802
rect 201696 225486 201724 231676
rect 202340 230314 202368 231676
rect 202328 230308 202380 230314
rect 202328 230250 202380 230256
rect 202144 230172 202196 230178
rect 202144 230114 202196 230120
rect 201684 225480 201736 225486
rect 201684 225422 201736 225428
rect 201408 221332 201460 221338
rect 201408 221274 201460 221280
rect 200856 219972 200908 219978
rect 200856 219914 200908 219920
rect 200672 218612 200724 218618
rect 200672 218554 200724 218560
rect 200028 218340 200080 218346
rect 200028 218282 200080 218288
rect 200868 217002 200896 219914
rect 201420 217002 201448 221274
rect 202156 218482 202184 230114
rect 202984 227497 203012 231676
rect 203168 231662 203642 231690
rect 202970 227488 203026 227497
rect 202970 227423 203026 227432
rect 202604 225480 202656 225486
rect 202604 225422 202656 225428
rect 202144 218476 202196 218482
rect 202144 218418 202196 218424
rect 202616 217002 202644 225422
rect 203168 219706 203196 231662
rect 204272 226302 204300 231676
rect 204260 226296 204312 226302
rect 204260 226238 204312 226244
rect 204168 222488 204220 222494
rect 204168 222430 204220 222436
rect 203156 219700 203208 219706
rect 203156 219642 203208 219648
rect 203340 218476 203392 218482
rect 203340 218418 203392 218424
rect 203352 217002 203380 218418
rect 203892 218340 203944 218346
rect 203892 218282 203944 218288
rect 203904 218074 203932 218282
rect 203892 218068 203944 218074
rect 203892 218010 203944 218016
rect 204180 217002 204208 222430
rect 204916 222358 204944 231676
rect 205272 229084 205324 229090
rect 205272 229026 205324 229032
rect 204904 222352 204956 222358
rect 204904 222294 204956 222300
rect 204996 218068 205048 218074
rect 204996 218010 205048 218016
rect 205008 217002 205036 218010
rect 192956 216974 193108 217002
rect 193936 216974 194364 217002
rect 194764 216974 195192 217002
rect 195592 216974 195928 217002
rect 196420 216974 196756 217002
rect 197248 216974 197308 217002
rect 198076 216974 198504 217002
rect 198904 216974 199240 217002
rect 199732 216974 199884 217002
rect 200560 216974 200896 217002
rect 201388 216974 201448 217002
rect 202216 216974 202644 217002
rect 203044 216974 203380 217002
rect 203872 216974 204208 217002
rect 204700 216974 205036 217002
rect 205284 217002 205312 229026
rect 205560 228138 205588 231676
rect 205836 231662 206218 231690
rect 206388 231662 206862 231690
rect 205548 228132 205600 228138
rect 205548 228074 205600 228080
rect 205456 226160 205508 226166
rect 205456 226102 205508 226108
rect 205468 218074 205496 226102
rect 205836 221066 205864 231662
rect 206388 225350 206416 231662
rect 207492 229226 207520 231676
rect 207664 230444 207716 230450
rect 207664 230386 207716 230392
rect 207480 229220 207532 229226
rect 207480 229162 207532 229168
rect 206376 225344 206428 225350
rect 206376 225286 206428 225292
rect 206560 225344 206612 225350
rect 206560 225286 206612 225292
rect 205824 221060 205876 221066
rect 205824 221002 205876 221008
rect 206572 219434 206600 225286
rect 207480 219836 207532 219842
rect 207480 219778 207532 219784
rect 206296 219406 206600 219434
rect 206296 218657 206324 219406
rect 206282 218648 206338 218657
rect 206282 218583 206338 218592
rect 206652 218612 206704 218618
rect 206652 218554 206704 218560
rect 205456 218068 205508 218074
rect 205456 218010 205508 218016
rect 206664 217002 206692 218554
rect 207492 217002 207520 219778
rect 207676 218346 207704 230386
rect 208136 227050 208164 231676
rect 208596 231662 208794 231690
rect 208124 227044 208176 227050
rect 208124 226986 208176 226992
rect 208124 222760 208176 222766
rect 208124 222702 208176 222708
rect 207664 218340 207716 218346
rect 207664 218282 207716 218288
rect 208136 217002 208164 222702
rect 208596 220658 208624 231662
rect 209424 225758 209452 231676
rect 210068 229362 210096 231676
rect 210056 229356 210108 229362
rect 210056 229298 210108 229304
rect 210424 229356 210476 229362
rect 210424 229298 210476 229304
rect 209412 225752 209464 225758
rect 209412 225694 209464 225700
rect 209596 225752 209648 225758
rect 209596 225694 209648 225700
rect 208584 220652 208636 220658
rect 208584 220594 208636 220600
rect 209608 219434 209636 225694
rect 209240 219406 209636 219434
rect 209240 217002 209268 219406
rect 210436 219298 210464 229298
rect 210712 228410 210740 231676
rect 210700 228404 210752 228410
rect 210700 228346 210752 228352
rect 210884 228268 210936 228274
rect 210884 228210 210936 228216
rect 209688 219292 209740 219298
rect 209688 219234 209740 219240
rect 210424 219292 210476 219298
rect 210424 219234 210476 219240
rect 209700 217002 209728 219234
rect 210896 217002 210924 228210
rect 211356 220697 211384 231676
rect 212000 222630 212028 231676
rect 212356 226908 212408 226914
rect 212356 226850 212408 226856
rect 211988 222624 212040 222630
rect 211988 222566 212040 222572
rect 211342 220688 211398 220697
rect 211342 220623 211398 220632
rect 211620 218068 211672 218074
rect 211620 218010 211672 218016
rect 211632 217002 211660 218010
rect 212368 217002 212396 226850
rect 212644 224126 212672 231676
rect 213092 229220 213144 229226
rect 213092 229162 213144 229168
rect 212632 224120 212684 224126
rect 212632 224062 212684 224068
rect 213104 218482 213132 229162
rect 213288 227186 213316 231676
rect 213276 227180 213328 227186
rect 213276 227122 213328 227128
rect 213932 222873 213960 231676
rect 214116 231662 214590 231690
rect 213918 222864 213974 222873
rect 213918 222799 213974 222808
rect 213828 222624 213880 222630
rect 213828 222566 213880 222572
rect 213092 218476 213144 218482
rect 213092 218418 213144 218424
rect 213276 218340 213328 218346
rect 213276 218282 213328 218288
rect 213288 217002 213316 218282
rect 213840 217002 213868 222566
rect 214116 221202 214144 231662
rect 215220 229498 215248 231676
rect 215208 229492 215260 229498
rect 215208 229434 215260 229440
rect 215024 228404 215076 228410
rect 215024 228346 215076 228352
rect 214104 221196 214156 221202
rect 214104 221138 214156 221144
rect 214380 219292 214432 219298
rect 214380 219234 214432 219240
rect 214392 218618 214420 219234
rect 214564 218884 214616 218890
rect 214564 218826 214616 218832
rect 214380 218612 214432 218618
rect 214380 218554 214432 218560
rect 214576 218482 214604 218826
rect 214748 218612 214800 218618
rect 214748 218554 214800 218560
rect 214564 218476 214616 218482
rect 214564 218418 214616 218424
rect 214760 218346 214788 218554
rect 214748 218340 214800 218346
rect 214748 218282 214800 218288
rect 215036 217002 215064 228346
rect 215864 228002 215892 231676
rect 216232 231662 216522 231690
rect 215852 227996 215904 228002
rect 215852 227938 215904 227944
rect 216232 222902 216260 231662
rect 217152 224262 217180 231676
rect 217796 229634 217824 231676
rect 217784 229628 217836 229634
rect 217784 229570 217836 229576
rect 217324 229492 217376 229498
rect 217324 229434 217376 229440
rect 217140 224256 217192 224262
rect 217140 224198 217192 224204
rect 216588 224120 216640 224126
rect 216588 224062 216640 224068
rect 216220 222896 216272 222902
rect 216220 222838 216272 222844
rect 215208 221196 215260 221202
rect 215208 221138 215260 221144
rect 215220 218074 215248 221138
rect 216404 220652 216456 220658
rect 216404 220594 216456 220600
rect 215208 218068 215260 218074
rect 215208 218010 215260 218016
rect 215760 218068 215812 218074
rect 215760 218010 215812 218016
rect 215772 217002 215800 218010
rect 216416 217002 216444 220594
rect 216600 218074 216628 224062
rect 217336 220658 217364 229434
rect 218440 225214 218468 231676
rect 218624 231662 219098 231690
rect 218428 225208 218480 225214
rect 218428 225150 218480 225156
rect 217784 222896 217836 222902
rect 217784 222838 217836 222844
rect 217324 220652 217376 220658
rect 217324 220594 217376 220600
rect 217508 220652 217560 220658
rect 217508 220594 217560 220600
rect 217520 219434 217548 220594
rect 217152 219406 217548 219434
rect 216588 218068 216640 218074
rect 216588 218010 216640 218016
rect 217152 217002 217180 219406
rect 205284 216974 205528 217002
rect 206356 216974 206692 217002
rect 207184 216974 207520 217002
rect 208012 216974 208164 217002
rect 208840 216974 209268 217002
rect 209668 216974 209728 217002
rect 210496 216974 210924 217002
rect 211324 216974 211660 217002
rect 212152 216974 212396 217002
rect 212980 216974 213316 217002
rect 213808 216974 213868 217002
rect 214636 216974 215064 217002
rect 215464 216974 215800 217002
rect 216292 216974 216444 217002
rect 217120 216974 217180 217002
rect 217796 217002 217824 222838
rect 218624 220114 218652 231662
rect 219164 226296 219216 226302
rect 219164 226238 219216 226244
rect 218612 220108 218664 220114
rect 218612 220050 218664 220056
rect 219176 217002 219204 226238
rect 219728 225894 219756 231676
rect 220372 230042 220400 231676
rect 220360 230036 220412 230042
rect 220360 229978 220412 229984
rect 221016 226642 221044 231676
rect 221292 231662 221674 231690
rect 221004 226636 221056 226642
rect 221004 226578 221056 226584
rect 219716 225888 219768 225894
rect 219716 225830 219768 225836
rect 220636 225888 220688 225894
rect 220636 225830 220688 225836
rect 219900 218340 219952 218346
rect 219900 218282 219952 218288
rect 219912 217002 219940 218282
rect 220648 217002 220676 225830
rect 220820 220244 220872 220250
rect 220820 220186 220872 220192
rect 220832 218482 220860 220186
rect 221292 220114 221320 231662
rect 222016 228132 222068 228138
rect 222016 228074 222068 228080
rect 221280 220108 221332 220114
rect 221280 220050 221332 220056
rect 220820 218476 220872 218482
rect 220820 218418 220872 218424
rect 221556 218068 221608 218074
rect 221556 218010 221608 218016
rect 221568 217002 221596 218010
rect 217796 216974 217948 217002
rect 218776 216974 219204 217002
rect 219604 216974 219940 217002
rect 220432 216974 220676 217002
rect 221260 216974 221596 217002
rect 222028 217002 222056 228074
rect 222304 225622 222332 231676
rect 222292 225616 222344 225622
rect 222292 225558 222344 225564
rect 222948 223990 222976 231676
rect 223592 228313 223620 231676
rect 223578 228304 223634 228313
rect 223578 228239 223634 228248
rect 223304 224256 223356 224262
rect 223304 224198 223356 224204
rect 222936 223984 222988 223990
rect 222936 223926 222988 223932
rect 222568 221060 222620 221066
rect 222568 221002 222620 221008
rect 222580 218074 222608 221002
rect 222568 218068 222620 218074
rect 222568 218010 222620 218016
rect 223316 217002 223344 224198
rect 224236 223038 224264 231676
rect 224420 231662 224894 231690
rect 224224 223032 224276 223038
rect 224224 222974 224276 222980
rect 224420 221474 224448 231662
rect 224960 230036 225012 230042
rect 224960 229978 225012 229984
rect 224776 227180 224828 227186
rect 224776 227122 224828 227128
rect 224592 226772 224644 226778
rect 224592 226714 224644 226720
rect 224408 221468 224460 221474
rect 224408 221410 224460 221416
rect 224604 218074 224632 226714
rect 224040 218068 224092 218074
rect 224040 218010 224092 218016
rect 224592 218068 224644 218074
rect 224592 218010 224644 218016
rect 224052 217002 224080 218010
rect 224788 217002 224816 227122
rect 224972 224262 225000 229978
rect 225524 229770 225552 231676
rect 225512 229764 225564 229770
rect 225512 229706 225564 229712
rect 226168 227050 226196 231676
rect 226156 227044 226208 227050
rect 226156 226986 226208 226992
rect 225512 225208 225564 225214
rect 225512 225150 225564 225156
rect 224960 224256 225012 224262
rect 224960 224198 225012 224204
rect 225524 218210 225552 225150
rect 226156 223984 226208 223990
rect 226156 223926 226208 223932
rect 225972 218476 226024 218482
rect 225972 218418 226024 218424
rect 225512 218204 225564 218210
rect 225512 218146 225564 218152
rect 225696 218068 225748 218074
rect 225696 218010 225748 218016
rect 225708 217002 225736 218010
rect 222028 216974 222088 217002
rect 222916 216974 223344 217002
rect 223744 216974 224080 217002
rect 224572 216974 224816 217002
rect 225400 216974 225736 217002
rect 225984 217002 226012 218418
rect 226168 218074 226196 223926
rect 226812 223174 226840 231676
rect 227456 224398 227484 231676
rect 228100 225350 228128 231676
rect 228744 228546 228772 231676
rect 229112 231662 229402 231690
rect 229572 231662 230046 231690
rect 228732 228540 228784 228546
rect 228732 228482 228784 228488
rect 228732 227044 228784 227050
rect 228732 226986 228784 226992
rect 228088 225344 228140 225350
rect 228088 225286 228140 225292
rect 227444 224392 227496 224398
rect 227444 224334 227496 224340
rect 227444 223712 227496 223718
rect 227444 223654 227496 223660
rect 226800 223168 226852 223174
rect 226800 223110 226852 223116
rect 226156 218068 226208 218074
rect 226156 218010 226208 218016
rect 227456 217002 227484 223654
rect 228180 220924 228232 220930
rect 228180 220866 228232 220872
rect 228192 217002 228220 220866
rect 228744 217002 228772 226986
rect 229112 220386 229140 231662
rect 229572 221241 229600 231662
rect 230480 230172 230532 230178
rect 230480 230114 230532 230120
rect 230492 223530 230520 230114
rect 230676 227866 230704 231676
rect 230664 227860 230716 227866
rect 230664 227802 230716 227808
rect 231320 226506 231348 231676
rect 231964 229094 231992 231676
rect 231964 229066 232084 229094
rect 231308 226500 231360 226506
rect 231308 226442 231360 226448
rect 231584 224256 231636 224262
rect 231584 224198 231636 224204
rect 230400 223502 230520 223530
rect 229558 221232 229614 221241
rect 229558 221167 229614 221176
rect 229100 220380 229152 220386
rect 229100 220322 229152 220328
rect 230204 220108 230256 220114
rect 230204 220050 230256 220056
rect 229836 218068 229888 218074
rect 229836 218010 229888 218016
rect 229848 217002 229876 218010
rect 225984 216974 226228 217002
rect 227056 216974 227484 217002
rect 227884 216974 228220 217002
rect 228712 216974 228772 217002
rect 229540 216974 229876 217002
rect 230216 217002 230244 220050
rect 230400 218074 230428 223502
rect 230388 218068 230440 218074
rect 230388 218010 230440 218016
rect 231596 217002 231624 224198
rect 231860 220516 231912 220522
rect 231860 220458 231912 220464
rect 231872 218754 231900 220458
rect 232056 219570 232084 229066
rect 232608 224534 232636 231676
rect 233266 231662 233464 231690
rect 232596 224528 232648 224534
rect 232596 224470 232648 224476
rect 233148 224528 233200 224534
rect 233148 224470 233200 224476
rect 232044 219564 232096 219570
rect 232044 219506 232096 219512
rect 232964 218884 233016 218890
rect 232964 218826 233016 218832
rect 231860 218748 231912 218754
rect 231860 218690 231912 218696
rect 232320 218068 232372 218074
rect 232320 218010 232372 218016
rect 232332 217002 232360 218010
rect 232976 217002 233004 218826
rect 233160 218074 233188 224470
rect 233436 220250 233464 231662
rect 233896 228818 233924 231676
rect 234172 231662 234554 231690
rect 233884 228812 233936 228818
rect 233884 228754 233936 228760
rect 234172 221746 234200 231662
rect 234528 228812 234580 228818
rect 234528 228754 234580 228760
rect 234160 221740 234212 221746
rect 234160 221682 234212 221688
rect 234344 221468 234396 221474
rect 234344 221410 234396 221416
rect 233424 220244 233476 220250
rect 233424 220186 233476 220192
rect 233884 219428 233936 219434
rect 233884 219370 233936 219376
rect 233896 218754 233924 219370
rect 233884 218748 233936 218754
rect 233884 218690 233936 218696
rect 233148 218068 233200 218074
rect 233148 218010 233200 218016
rect 233976 218068 234028 218074
rect 233976 218010 234028 218016
rect 233988 217002 234016 218010
rect 230216 216974 230368 217002
rect 231196 216974 231624 217002
rect 232024 216974 232360 217002
rect 232852 216974 233004 217002
rect 233680 216974 234016 217002
rect 234356 217002 234384 221410
rect 234540 218074 234568 228754
rect 235184 223854 235212 231676
rect 235828 229906 235856 231676
rect 235816 229900 235868 229906
rect 235816 229842 235868 229848
rect 235724 228540 235776 228546
rect 235724 228482 235776 228488
rect 235172 223848 235224 223854
rect 235172 223790 235224 223796
rect 234528 218068 234580 218074
rect 234528 218010 234580 218016
rect 235736 217002 235764 228482
rect 236472 227594 236500 231676
rect 236656 231662 237130 231690
rect 237392 231662 237774 231690
rect 238036 231662 238418 231690
rect 236460 227588 236512 227594
rect 236460 227530 236512 227536
rect 236656 220386 236684 231662
rect 237392 221610 237420 231662
rect 237380 221604 237432 221610
rect 237380 221546 237432 221552
rect 238036 220522 238064 231662
rect 239048 228682 239076 231676
rect 239232 231662 239706 231690
rect 239036 228676 239088 228682
rect 239036 228618 239088 228624
rect 238668 223032 238720 223038
rect 238668 222974 238720 222980
rect 238024 220516 238076 220522
rect 238024 220458 238076 220464
rect 236644 220380 236696 220386
rect 236644 220322 236696 220328
rect 237288 220244 237340 220250
rect 237288 220186 237340 220192
rect 236460 219700 236512 219706
rect 236460 219642 236512 219648
rect 235908 219564 235960 219570
rect 235908 219506 235960 219512
rect 235920 219026 235948 219506
rect 235908 219020 235960 219026
rect 235908 218962 235960 218968
rect 236472 217002 236500 219642
rect 237300 217002 237328 220186
rect 238116 219020 238168 219026
rect 238116 218962 238168 218968
rect 238128 217002 238156 218962
rect 238680 217002 238708 222974
rect 239232 222154 239260 231662
rect 239404 225616 239456 225622
rect 239404 225558 239456 225564
rect 239220 222148 239272 222154
rect 239220 222090 239272 222096
rect 238852 221604 238904 221610
rect 238852 221546 238904 221552
rect 238864 218754 238892 221546
rect 239416 219026 239444 225558
rect 240336 224670 240364 231676
rect 240980 230314 241008 231676
rect 240968 230308 241020 230314
rect 240968 230250 241020 230256
rect 241624 226030 241652 231676
rect 241808 231662 242282 231690
rect 241612 226024 241664 226030
rect 241612 225966 241664 225972
rect 240324 224664 240376 224670
rect 240324 224606 240376 224612
rect 241244 224392 241296 224398
rect 241244 224334 241296 224340
rect 240600 220380 240652 220386
rect 240600 220322 240652 220328
rect 239404 219020 239456 219026
rect 239404 218962 239456 218968
rect 239772 219020 239824 219026
rect 239772 218962 239824 218968
rect 238852 218748 238904 218754
rect 238852 218690 238904 218696
rect 239784 217002 239812 218962
rect 240612 217002 240640 220322
rect 241256 217002 241284 224334
rect 241808 220794 241836 231662
rect 242532 230308 242584 230314
rect 242532 230250 242584 230256
rect 241796 220788 241848 220794
rect 241796 220730 241848 220736
rect 242256 218068 242308 218074
rect 242256 218010 242308 218016
rect 242268 217002 242296 218010
rect 234356 216974 234508 217002
rect 235336 216974 235764 217002
rect 236164 216974 236500 217002
rect 236992 216974 237328 217002
rect 237820 216974 238156 217002
rect 238648 216974 238708 217002
rect 239476 216974 239812 217002
rect 240304 216974 240640 217002
rect 241132 216974 241284 217002
rect 241960 216974 242296 217002
rect 242544 217002 242572 230250
rect 242716 227588 242768 227594
rect 242716 227530 242768 227536
rect 242728 218074 242756 227530
rect 242912 224806 242940 231676
rect 243096 231662 243570 231690
rect 242900 224800 242952 224806
rect 242900 224742 242952 224748
rect 243096 219570 243124 231662
rect 244200 227322 244228 231676
rect 244188 227316 244240 227322
rect 244188 227258 244240 227264
rect 244844 223310 244872 231676
rect 245120 231662 245502 231690
rect 244832 223304 244884 223310
rect 244832 223246 244884 223252
rect 244004 222352 244056 222358
rect 244004 222294 244056 222300
rect 243084 219564 243136 219570
rect 243084 219506 243136 219512
rect 242716 218068 242768 218074
rect 242716 218010 242768 218016
rect 244016 217002 244044 222294
rect 245120 221882 245148 231662
rect 245568 225344 245620 225350
rect 245568 225286 245620 225292
rect 245108 221876 245160 221882
rect 245108 221818 245160 221824
rect 244740 218748 244792 218754
rect 244740 218690 244792 218696
rect 244752 217002 244780 218690
rect 245580 217002 245608 225286
rect 246132 225214 246160 231676
rect 246776 228954 246804 231676
rect 246764 228948 246816 228954
rect 246764 228890 246816 228896
rect 246304 228676 246356 228682
rect 246304 228618 246356 228624
rect 246120 225208 246172 225214
rect 246120 225150 246172 225156
rect 246316 218754 246344 228618
rect 247420 223582 247448 231676
rect 248064 224942 248092 231676
rect 248616 231662 248722 231690
rect 248052 224936 248104 224942
rect 248052 224878 248104 224884
rect 247408 223576 247460 223582
rect 247408 223518 247460 223524
rect 248144 223168 248196 223174
rect 248144 223110 248196 223116
rect 247132 221740 247184 221746
rect 247132 221682 247184 221688
rect 246948 220516 247000 220522
rect 246948 220458 247000 220464
rect 246488 219020 246540 219026
rect 246488 218962 246540 218968
rect 246500 218754 246528 218962
rect 246304 218748 246356 218754
rect 246304 218690 246356 218696
rect 246488 218748 246540 218754
rect 246488 218690 246540 218696
rect 246396 218204 246448 218210
rect 246396 218146 246448 218152
rect 246408 217002 246436 218146
rect 246960 217002 246988 220458
rect 247144 219162 247172 221682
rect 247132 219156 247184 219162
rect 247132 219098 247184 219104
rect 248156 217002 248184 223110
rect 248616 221610 248644 231662
rect 249352 225078 249380 231676
rect 249340 225072 249392 225078
rect 249340 225014 249392 225020
rect 249616 224664 249668 224670
rect 249616 224606 249668 224612
rect 248604 221604 248656 221610
rect 248604 221546 248656 221552
rect 249248 219020 249300 219026
rect 249248 218962 249300 218968
rect 249260 218210 249288 218962
rect 249248 218204 249300 218210
rect 249248 218146 249300 218152
rect 249432 218204 249484 218210
rect 249432 218146 249484 218152
rect 248880 218068 248932 218074
rect 248880 218010 248932 218016
rect 248892 217002 248920 218010
rect 249444 217002 249472 218146
rect 249628 218074 249656 224606
rect 249996 223446 250024 231676
rect 250180 231662 250654 231690
rect 249984 223440 250036 223446
rect 249984 223382 250036 223388
rect 250180 222018 250208 231662
rect 251284 230450 251312 231676
rect 251272 230444 251324 230450
rect 251272 230386 251324 230392
rect 251732 229628 251784 229634
rect 251732 229570 251784 229576
rect 251744 229094 251772 229570
rect 251928 229094 251956 231676
rect 252586 231662 252784 231690
rect 251744 229066 251864 229094
rect 251928 229066 252048 229094
rect 251088 227316 251140 227322
rect 251088 227258 251140 227264
rect 250168 222012 250220 222018
rect 250168 221954 250220 221960
rect 250536 221604 250588 221610
rect 250536 221546 250588 221552
rect 249616 218068 249668 218074
rect 249616 218010 249668 218016
rect 250548 217002 250576 221546
rect 251100 217002 251128 227258
rect 251836 218210 251864 229066
rect 252020 227730 252048 229066
rect 252284 227996 252336 228002
rect 252284 227938 252336 227944
rect 252008 227724 252060 227730
rect 252008 227666 252060 227672
rect 251824 218204 251876 218210
rect 251824 218146 251876 218152
rect 252296 217002 252324 227938
rect 252756 219978 252784 231662
rect 253216 227458 253244 231676
rect 253400 231662 253874 231690
rect 253204 227452 253256 227458
rect 253204 227394 253256 227400
rect 253400 221746 253428 231662
rect 254504 225486 254532 231676
rect 254780 231662 255162 231690
rect 255424 231662 255806 231690
rect 254492 225480 254544 225486
rect 254492 225422 254544 225428
rect 253756 223576 253808 223582
rect 253756 223518 253808 223524
rect 253388 221740 253440 221746
rect 253388 221682 253440 221688
rect 253572 221740 253624 221746
rect 253572 221682 253624 221688
rect 252744 219972 252796 219978
rect 252744 219914 252796 219920
rect 253020 219428 253072 219434
rect 253020 219370 253072 219376
rect 253032 217002 253060 219370
rect 253584 219298 253612 221682
rect 253572 219292 253624 219298
rect 253572 219234 253624 219240
rect 253768 217002 253796 223518
rect 254780 222494 254808 231662
rect 255136 226024 255188 226030
rect 255136 225966 255188 225972
rect 254952 225480 255004 225486
rect 254952 225422 255004 225428
rect 254768 222488 254820 222494
rect 254768 222430 254820 222436
rect 254676 218068 254728 218074
rect 254676 218010 254728 218016
rect 254688 217002 254716 218010
rect 242544 216974 242788 217002
rect 243616 216974 244044 217002
rect 244444 216974 244780 217002
rect 245272 216974 245608 217002
rect 246100 216974 246436 217002
rect 246928 216974 246988 217002
rect 247756 216974 248184 217002
rect 248584 216974 248920 217002
rect 249412 216974 249472 217002
rect 250240 216974 250576 217002
rect 251068 216974 251128 217002
rect 251896 216974 252324 217002
rect 252724 216974 253060 217002
rect 253552 216974 253796 217002
rect 254380 216974 254716 217002
rect 254964 217002 254992 225422
rect 255148 218074 255176 225966
rect 255424 221338 255452 231662
rect 256436 229226 256464 231676
rect 256608 230444 256660 230450
rect 256608 230386 256660 230392
rect 256424 229220 256476 229226
rect 256424 229162 256476 229168
rect 255412 221332 255464 221338
rect 255412 221274 255464 221280
rect 256620 219434 256648 230386
rect 257080 229090 257108 231676
rect 257264 231662 257738 231690
rect 257264 229094 257292 231662
rect 257068 229084 257120 229090
rect 257264 229066 257384 229094
rect 257068 229026 257120 229032
rect 257160 219972 257212 219978
rect 257160 219914 257212 219920
rect 256436 219406 256648 219434
rect 255136 218068 255188 218074
rect 255136 218010 255188 218016
rect 256436 217002 256464 219406
rect 257172 217002 257200 219914
rect 257356 219842 257384 229066
rect 257804 228948 257856 228954
rect 257804 228890 257856 228896
rect 257344 219836 257396 219842
rect 257344 219778 257396 219784
rect 257816 217002 257844 228890
rect 258368 226166 258396 231676
rect 258644 231662 259026 231690
rect 258356 226160 258408 226166
rect 258356 226102 258408 226108
rect 258080 221876 258132 221882
rect 258080 221818 258132 221824
rect 258092 218346 258120 221818
rect 258644 221746 258672 231662
rect 259368 227452 259420 227458
rect 259368 227394 259420 227400
rect 258632 221740 258684 221746
rect 258632 221682 258684 221688
rect 259184 219292 259236 219298
rect 259184 219234 259236 219240
rect 258080 218340 258132 218346
rect 258080 218282 258132 218288
rect 258816 218068 258868 218074
rect 258816 218010 258868 218016
rect 258828 217002 258856 218010
rect 254964 216974 255208 217002
rect 256036 216974 256464 217002
rect 256864 216974 257200 217002
rect 257692 216974 257844 217002
rect 258520 216974 258856 217002
rect 259196 217002 259224 219234
rect 259380 218074 259408 227394
rect 259656 225758 259684 231676
rect 260300 228274 260328 231676
rect 260288 228268 260340 228274
rect 260288 228210 260340 228216
rect 259644 225752 259696 225758
rect 259644 225694 259696 225700
rect 260104 225004 260156 225010
rect 260104 224946 260156 224952
rect 260116 218618 260144 224946
rect 260944 222766 260972 231676
rect 261312 231662 261602 231690
rect 261312 229362 261340 231662
rect 261300 229356 261352 229362
rect 261300 229298 261352 229304
rect 261484 229356 261536 229362
rect 261484 229298 261536 229304
rect 260932 222760 260984 222766
rect 260932 222702 260984 222708
rect 260472 221740 260524 221746
rect 260472 221682 260524 221688
rect 260104 218612 260156 218618
rect 260104 218554 260156 218560
rect 259368 218068 259420 218074
rect 259368 218010 259420 218016
rect 260484 217002 260512 221682
rect 261300 220788 261352 220794
rect 261300 220730 261352 220736
rect 261312 217002 261340 220730
rect 261496 219706 261524 229298
rect 262232 226914 262260 231676
rect 262220 226908 262272 226914
rect 262220 226850 262272 226856
rect 262128 223304 262180 223310
rect 262128 223246 262180 223252
rect 261484 219700 261536 219706
rect 261484 219642 261536 219648
rect 262140 217002 262168 223246
rect 262876 222630 262904 231676
rect 263152 231662 263534 231690
rect 262864 222624 262916 222630
rect 262864 222566 262916 222572
rect 263152 221202 263180 231662
rect 263416 227724 263468 227730
rect 263416 227666 263468 227672
rect 263140 221196 263192 221202
rect 263140 221138 263192 221144
rect 262956 218612 263008 218618
rect 262956 218554 263008 218560
rect 262968 217002 262996 218554
rect 259196 216974 259348 217002
rect 260176 216974 260512 217002
rect 261004 216974 261340 217002
rect 261832 216974 262168 217002
rect 262660 216974 262996 217002
rect 263428 217002 263456 227666
rect 264164 225010 264192 231676
rect 264440 231662 264822 231690
rect 265084 231662 265466 231690
rect 264152 225004 264204 225010
rect 264152 224946 264204 224952
rect 264440 224126 264468 231662
rect 264704 225752 264756 225758
rect 264704 225694 264756 225700
rect 264428 224120 264480 224126
rect 264428 224062 264480 224068
rect 264716 217002 264744 225694
rect 265084 220658 265112 231662
rect 265624 229084 265676 229090
rect 265624 229026 265676 229032
rect 265072 220652 265124 220658
rect 265072 220594 265124 220600
rect 265636 218482 265664 229026
rect 266096 228410 266124 231676
rect 266740 229498 266768 231676
rect 266728 229492 266780 229498
rect 266728 229434 266780 229440
rect 266084 228404 266136 228410
rect 266084 228346 266136 228352
rect 267384 226302 267412 231676
rect 267372 226296 267424 226302
rect 267372 226238 267424 226244
rect 268028 225894 268056 231676
rect 268016 225888 268068 225894
rect 268016 225830 268068 225836
rect 266268 224936 266320 224942
rect 266268 224878 266320 224884
rect 265624 218476 265676 218482
rect 265624 218418 265676 218424
rect 266084 218476 266136 218482
rect 266084 218418 266136 218424
rect 265440 218068 265492 218074
rect 265440 218010 265492 218016
rect 265452 217002 265480 218010
rect 266096 217002 266124 218418
rect 266280 218074 266308 224878
rect 267372 223440 267424 223446
rect 267372 223382 267424 223388
rect 267096 222148 267148 222154
rect 267096 222090 267148 222096
rect 266268 218068 266320 218074
rect 266268 218010 266320 218016
rect 267108 217002 267136 222090
rect 263428 216974 263488 217002
rect 264316 216974 264744 217002
rect 265144 216974 265480 217002
rect 265972 216974 266124 217002
rect 266800 216974 267136 217002
rect 267384 217002 267412 223382
rect 268672 222902 268700 231676
rect 269224 231662 269330 231690
rect 268844 225888 268896 225894
rect 268844 225830 268896 225836
rect 268660 222896 268712 222902
rect 268660 222838 268712 222844
rect 268856 217002 268884 225830
rect 269224 221882 269252 231662
rect 269960 228138 269988 231676
rect 270132 229764 270184 229770
rect 270132 229706 270184 229712
rect 269948 228132 270000 228138
rect 269948 228074 270000 228080
rect 269948 222012 270000 222018
rect 269948 221954 270000 221960
rect 269212 221876 269264 221882
rect 269212 221818 269264 221824
rect 269580 218068 269632 218074
rect 269580 218010 269632 218016
rect 269592 217002 269620 218010
rect 267384 216974 267628 217002
rect 268456 216974 268884 217002
rect 269284 216974 269620 217002
rect 269960 217002 269988 221954
rect 270144 218074 270172 229706
rect 270604 226778 270632 231676
rect 270880 231662 271262 231690
rect 270592 226772 270644 226778
rect 270592 226714 270644 226720
rect 270880 221066 270908 231662
rect 271892 230042 271920 231676
rect 271880 230036 271932 230042
rect 271880 229978 271932 229984
rect 271788 228404 271840 228410
rect 271788 228346 271840 228352
rect 271328 224800 271380 224806
rect 271328 224742 271380 224748
rect 270868 221060 270920 221066
rect 270868 221002 270920 221008
rect 270132 218068 270184 218074
rect 270132 218010 270184 218016
rect 271340 217002 271368 224742
rect 271800 217002 271828 228346
rect 272536 223990 272564 231676
rect 272524 223984 272576 223990
rect 272524 223926 272576 223932
rect 273180 223718 273208 231676
rect 273824 227186 273852 231676
rect 274468 229090 274496 231676
rect 274456 229084 274508 229090
rect 274456 229026 274508 229032
rect 274640 229084 274692 229090
rect 274640 229026 274692 229032
rect 274652 228970 274680 229026
rect 274284 228942 274680 228970
rect 273812 227180 273864 227186
rect 273812 227122 273864 227128
rect 273168 223712 273220 223718
rect 273168 223654 273220 223660
rect 273076 219564 273128 219570
rect 273076 219506 273128 219512
rect 272524 219428 272576 219434
rect 272524 219370 272576 219376
rect 272536 218482 272564 219370
rect 273088 218890 273116 219506
rect 273076 218884 273128 218890
rect 273076 218826 273128 218832
rect 272524 218476 272576 218482
rect 272524 218418 272576 218424
rect 272892 218476 272944 218482
rect 272892 218418 272944 218424
rect 272904 217002 272932 218418
rect 274284 218074 274312 228942
rect 274456 227180 274508 227186
rect 274456 227122 274508 227128
rect 273720 218068 273772 218074
rect 273720 218010 273772 218016
rect 274272 218068 274324 218074
rect 274272 218010 274324 218016
rect 273732 217002 273760 218010
rect 274468 217002 274496 227122
rect 275112 227050 275140 231676
rect 275296 231662 275770 231690
rect 276124 231662 276414 231690
rect 275100 227044 275152 227050
rect 275100 226986 275152 226992
rect 275296 220114 275324 231662
rect 275468 226908 275520 226914
rect 275468 226850 275520 226856
rect 275284 220108 275336 220114
rect 275284 220050 275336 220056
rect 275480 217002 275508 226850
rect 275836 224120 275888 224126
rect 275836 224062 275888 224068
rect 269960 216974 270112 217002
rect 270940 216974 271368 217002
rect 271768 216974 271828 217002
rect 272596 216974 272932 217002
rect 273424 216974 273760 217002
rect 274252 216974 274496 217002
rect 275080 216974 275508 217002
rect 275848 217002 275876 224062
rect 276124 220930 276152 231662
rect 277044 230178 277072 231676
rect 277032 230172 277084 230178
rect 277032 230114 277084 230120
rect 276664 229492 276716 229498
rect 276664 229434 276716 229440
rect 276112 220924 276164 220930
rect 276112 220866 276164 220872
rect 276676 218618 276704 229434
rect 277688 224534 277716 231676
rect 278332 228818 278360 231676
rect 278320 228812 278372 228818
rect 278320 228754 278372 228760
rect 277676 224528 277728 224534
rect 277676 224470 277728 224476
rect 278976 224262 279004 231676
rect 279252 231662 279634 231690
rect 278964 224256 279016 224262
rect 278964 224198 279016 224204
rect 278412 222896 278464 222902
rect 278412 222838 278464 222844
rect 277860 221876 277912 221882
rect 277860 221818 277912 221824
rect 277032 220652 277084 220658
rect 277032 220594 277084 220600
rect 276664 218612 276716 218618
rect 276664 218554 276716 218560
rect 277044 217002 277072 220594
rect 277872 217002 277900 221818
rect 278424 217002 278452 222838
rect 279252 219570 279280 231662
rect 280264 228546 280292 231676
rect 280540 231662 280922 231690
rect 281566 231662 281764 231690
rect 280252 228540 280304 228546
rect 280252 228482 280304 228488
rect 280540 220250 280568 231662
rect 280804 227860 280856 227866
rect 280804 227802 280856 227808
rect 280528 220244 280580 220250
rect 280528 220186 280580 220192
rect 280068 220108 280120 220114
rect 280068 220050 280120 220056
rect 279240 219564 279292 219570
rect 279240 219506 279292 219512
rect 279516 218612 279568 218618
rect 279516 218554 279568 218560
rect 279528 217002 279556 218554
rect 280080 217002 280108 220050
rect 280816 218754 280844 227802
rect 281264 224256 281316 224262
rect 281264 224198 281316 224204
rect 280804 218748 280856 218754
rect 280804 218690 280856 218696
rect 281276 217002 281304 224198
rect 281736 221474 281764 231662
rect 282196 229362 282224 231676
rect 282184 229356 282236 229362
rect 282184 229298 282236 229304
rect 282552 224528 282604 224534
rect 282552 224470 282604 224476
rect 281724 221468 281776 221474
rect 281724 221410 281776 221416
rect 282564 218074 282592 224470
rect 282840 223038 282868 231676
rect 283116 231662 283498 231690
rect 282828 223032 282880 223038
rect 282828 222974 282880 222980
rect 282828 221332 282880 221338
rect 282828 221274 282880 221280
rect 282000 218068 282052 218074
rect 282000 218010 282052 218016
rect 282552 218068 282604 218074
rect 282552 218010 282604 218016
rect 282012 217002 282040 218010
rect 282840 217002 282868 221274
rect 283116 220386 283144 231662
rect 283564 229900 283616 229906
rect 283564 229842 283616 229848
rect 283576 221338 283604 229842
rect 284128 225622 284156 231676
rect 284772 227866 284800 231676
rect 284760 227860 284812 227866
rect 284760 227802 284812 227808
rect 285416 227594 285444 231676
rect 285588 228812 285640 228818
rect 285588 228754 285640 228760
rect 285404 227588 285456 227594
rect 285404 227530 285456 227536
rect 284944 227044 284996 227050
rect 284944 226986 284996 226992
rect 284116 225616 284168 225622
rect 284116 225558 284168 225564
rect 284024 221468 284076 221474
rect 284024 221410 284076 221416
rect 283564 221332 283616 221338
rect 283564 221274 283616 221280
rect 283104 220380 283156 220386
rect 283104 220322 283156 220328
rect 283656 220244 283708 220250
rect 283656 220186 283708 220192
rect 283668 217002 283696 220186
rect 284036 219026 284064 221410
rect 284024 219020 284076 219026
rect 284024 218962 284076 218968
rect 284956 218074 284984 226986
rect 285600 219434 285628 228754
rect 286060 222358 286088 231676
rect 286704 224398 286732 231676
rect 287348 230314 287376 231676
rect 287336 230308 287388 230314
rect 287336 230250 287388 230256
rect 286968 226296 287020 226302
rect 286968 226238 287020 226244
rect 286692 224392 286744 224398
rect 286692 224334 286744 224340
rect 286048 222352 286100 222358
rect 286048 222294 286100 222300
rect 285416 219406 285628 219434
rect 284208 218068 284260 218074
rect 284208 218010 284260 218016
rect 284944 218068 284996 218074
rect 284944 218010 284996 218016
rect 284220 217002 284248 218010
rect 285416 217002 285444 219406
rect 286140 218884 286192 218890
rect 286140 218826 286192 218832
rect 286152 217002 286180 218826
rect 286980 217002 287008 226238
rect 287992 225350 288020 231676
rect 288544 231662 288650 231690
rect 288348 228540 288400 228546
rect 288348 228482 288400 228488
rect 288164 225616 288216 225622
rect 288164 225558 288216 225564
rect 287980 225344 288032 225350
rect 287980 225286 288032 225292
rect 287796 218068 287848 218074
rect 287796 218010 287848 218016
rect 287808 217002 287836 218010
rect 275848 216974 275908 217002
rect 276736 216974 277072 217002
rect 277564 216974 277900 217002
rect 278392 216974 278452 217002
rect 279220 216974 279556 217002
rect 280048 216974 280108 217002
rect 280876 216974 281304 217002
rect 281704 216974 282040 217002
rect 282532 216974 282868 217002
rect 283360 216974 283696 217002
rect 284188 216974 284248 217002
rect 285016 216974 285444 217002
rect 285844 216974 286180 217002
rect 286672 216974 287008 217002
rect 287500 216974 287836 217002
rect 288176 217002 288204 225558
rect 288360 218074 288388 228482
rect 288544 220522 288572 231662
rect 288716 229356 288768 229362
rect 288716 229298 288768 229304
rect 288728 224126 288756 229298
rect 289280 228682 289308 231676
rect 289268 228676 289320 228682
rect 289268 228618 289320 228624
rect 288716 224120 288768 224126
rect 288716 224062 288768 224068
rect 289084 223916 289136 223922
rect 289084 223858 289136 223864
rect 288532 220516 288584 220522
rect 288532 220458 288584 220464
rect 288532 219836 288584 219842
rect 288532 219778 288584 219784
rect 288544 218482 288572 219778
rect 289096 219026 289124 223858
rect 289924 221474 289952 231676
rect 290568 224670 290596 231676
rect 291226 231662 291424 231690
rect 290556 224664 290608 224670
rect 290556 224606 290608 224612
rect 291108 224392 291160 224398
rect 291108 224334 291160 224340
rect 290924 222760 290976 222766
rect 290924 222702 290976 222708
rect 289912 221468 289964 221474
rect 289912 221410 289964 221416
rect 289084 219020 289136 219026
rect 289084 218962 289136 218968
rect 288532 218476 288584 218482
rect 288532 218418 288584 218424
rect 289452 218204 289504 218210
rect 289452 218146 289504 218152
rect 288348 218068 288400 218074
rect 288348 218010 288400 218016
rect 289464 217002 289492 218146
rect 290936 218074 290964 222702
rect 290280 218068 290332 218074
rect 290280 218010 290332 218016
rect 290924 218068 290976 218074
rect 290924 218010 290976 218016
rect 290292 217002 290320 218010
rect 291120 217002 291148 224334
rect 291396 221610 291424 231662
rect 291856 223174 291884 231676
rect 292500 229634 292528 231676
rect 292488 229628 292540 229634
rect 292488 229570 292540 229576
rect 293144 228002 293172 231676
rect 293512 231662 293802 231690
rect 293132 227996 293184 228002
rect 293132 227938 293184 227944
rect 293512 223582 293540 231662
rect 293684 227588 293736 227594
rect 293684 227530 293736 227536
rect 293500 223576 293552 223582
rect 293500 223518 293552 223524
rect 291844 223168 291896 223174
rect 291844 223110 291896 223116
rect 292488 223032 292540 223038
rect 292488 222974 292540 222980
rect 291384 221604 291436 221610
rect 291384 221546 291436 221552
rect 292304 221468 292356 221474
rect 292304 221410 292356 221416
rect 292316 219298 292344 221410
rect 292304 219292 292356 219298
rect 292304 219234 292356 219240
rect 291936 218748 291988 218754
rect 291936 218690 291988 218696
rect 291948 217002 291976 218690
rect 292500 217002 292528 222974
rect 293696 217002 293724 227530
rect 294432 227322 294460 231676
rect 294800 231662 295090 231690
rect 294604 230172 294656 230178
rect 294604 230114 294656 230120
rect 294420 227316 294472 227322
rect 294420 227258 294472 227264
rect 294420 219020 294472 219026
rect 294420 218962 294472 218968
rect 294432 217002 294460 218962
rect 294616 218210 294644 230114
rect 294800 223922 294828 231662
rect 295720 225486 295748 231676
rect 295996 231662 296378 231690
rect 295708 225480 295760 225486
rect 295708 225422 295760 225428
rect 295156 224664 295208 224670
rect 295156 224606 295208 224612
rect 294788 223916 294840 223922
rect 294788 223858 294840 223864
rect 294604 218204 294656 218210
rect 294604 218146 294656 218152
rect 295168 217002 295196 224606
rect 295996 219978 296024 231662
rect 296628 226160 296680 226166
rect 296628 226102 296680 226108
rect 296444 221604 296496 221610
rect 296444 221546 296496 221552
rect 295984 219972 296036 219978
rect 295984 219914 296036 219920
rect 296076 218068 296128 218074
rect 296076 218010 296128 218016
rect 296088 217002 296116 218010
rect 288176 216974 288328 217002
rect 289156 216974 289492 217002
rect 289984 216974 290320 217002
rect 290812 216974 291148 217002
rect 291640 216974 291976 217002
rect 292468 216974 292528 217002
rect 293296 216974 293724 217002
rect 294124 216974 294460 217002
rect 294952 216974 295196 217002
rect 295780 216974 296116 217002
rect 296456 217002 296484 221546
rect 296640 218074 296668 226102
rect 297008 226030 297036 231676
rect 297652 230450 297680 231676
rect 297640 230444 297692 230450
rect 297640 230386 297692 230392
rect 297364 227860 297416 227866
rect 297364 227802 297416 227808
rect 296996 226024 297048 226030
rect 296996 225966 297048 225972
rect 297376 219434 297404 227802
rect 298296 227458 298324 231676
rect 298572 231662 298954 231690
rect 298572 229094 298600 231662
rect 298480 229066 298600 229094
rect 298284 227452 298336 227458
rect 298284 227394 298336 227400
rect 298480 221898 298508 229066
rect 299584 228954 299612 231676
rect 299768 231662 300242 231690
rect 299572 228948 299624 228954
rect 299572 228890 299624 228896
rect 298388 221870 298508 221898
rect 298388 221746 298416 221870
rect 298376 221740 298428 221746
rect 298376 221682 298428 221688
rect 298560 221740 298612 221746
rect 298560 221682 298612 221688
rect 297364 219428 297416 219434
rect 297364 219370 297416 219376
rect 296628 218068 296680 218074
rect 296628 218010 296680 218016
rect 297732 218068 297784 218074
rect 297732 218010 297784 218016
rect 297744 217002 297772 218010
rect 298572 217002 298600 221682
rect 299768 221474 299796 231662
rect 300124 230036 300176 230042
rect 300124 229978 300176 229984
rect 299756 221468 299808 221474
rect 299756 221410 299808 221416
rect 299204 220380 299256 220386
rect 299204 220322 299256 220328
rect 299216 217002 299244 220322
rect 300136 219434 300164 229978
rect 300872 223310 300900 231676
rect 301516 227730 301544 231676
rect 301792 231662 302174 231690
rect 301504 227724 301556 227730
rect 301504 227666 301556 227672
rect 300860 223304 300912 223310
rect 300860 223246 300912 223252
rect 300768 223168 300820 223174
rect 300768 223110 300820 223116
rect 300044 219406 300164 219434
rect 300044 218074 300072 219406
rect 300584 219156 300636 219162
rect 300584 219098 300636 219104
rect 300032 218068 300084 218074
rect 300032 218010 300084 218016
rect 300216 218068 300268 218074
rect 300216 218010 300268 218016
rect 300228 217002 300256 218010
rect 296456 216974 296608 217002
rect 297436 216974 297772 217002
rect 298264 216974 298600 217002
rect 299092 216974 299244 217002
rect 299920 216974 300256 217002
rect 300596 217002 300624 219098
rect 300780 218074 300808 223110
rect 301792 220794 301820 231662
rect 302804 229498 302832 231676
rect 302792 229492 302844 229498
rect 302792 229434 302844 229440
rect 301964 227452 302016 227458
rect 301964 227394 302016 227400
rect 301780 220788 301832 220794
rect 301780 220730 301832 220736
rect 300768 218068 300820 218074
rect 300768 218010 300820 218016
rect 301976 217002 302004 227394
rect 303252 226024 303304 226030
rect 303252 225966 303304 225972
rect 302700 221468 302752 221474
rect 302700 221410 302752 221416
rect 302712 217002 302740 221410
rect 303264 217002 303292 225966
rect 303448 224942 303476 231676
rect 303816 231662 304106 231690
rect 303436 224936 303488 224942
rect 303436 224878 303488 224884
rect 303816 222154 303844 231662
rect 304736 225758 304764 231676
rect 304908 228676 304960 228682
rect 304908 228618 304960 228624
rect 304724 225752 304776 225758
rect 304724 225694 304776 225700
rect 303804 222148 303856 222154
rect 303804 222090 303856 222096
rect 304920 219434 304948 228618
rect 305380 227866 305408 231676
rect 305644 230308 305696 230314
rect 305644 230250 305696 230256
rect 305368 227860 305420 227866
rect 305368 227802 305420 227808
rect 304828 219406 304948 219434
rect 304356 218068 304408 218074
rect 304356 218010 304408 218016
rect 304368 217002 304396 218010
rect 300596 216974 300748 217002
rect 301576 216974 302004 217002
rect 302404 216974 302740 217002
rect 303232 216974 303292 217002
rect 304060 216974 304396 217002
rect 304828 217002 304856 219406
rect 305656 218074 305684 230250
rect 306024 225894 306052 231676
rect 306576 231662 306682 231690
rect 306012 225888 306064 225894
rect 306012 225830 306064 225836
rect 306104 225752 306156 225758
rect 306104 225694 306156 225700
rect 305644 218068 305696 218074
rect 305644 218010 305696 218016
rect 306116 217002 306144 225694
rect 306576 222018 306604 231662
rect 307024 223576 307076 223582
rect 307024 223518 307076 223524
rect 306564 222012 306616 222018
rect 306564 221954 306616 221960
rect 306840 222012 306892 222018
rect 306840 221954 306892 221960
rect 306852 217002 306880 221954
rect 307036 218482 307064 223518
rect 307312 223446 307340 231676
rect 307956 229770 307984 231676
rect 307944 229764 307996 229770
rect 307944 229706 307996 229712
rect 308600 228410 308628 231676
rect 309244 229090 309272 231676
rect 309232 229084 309284 229090
rect 309232 229026 309284 229032
rect 309692 229084 309744 229090
rect 309692 229026 309744 229032
rect 308588 228404 308640 228410
rect 308588 228346 308640 228352
rect 309048 228404 309100 228410
rect 309048 228346 309100 228352
rect 308864 227316 308916 227322
rect 308864 227258 308916 227264
rect 307300 223440 307352 223446
rect 307300 223382 307352 223388
rect 307668 219292 307720 219298
rect 307668 219234 307720 219240
rect 307024 218476 307076 218482
rect 307024 218418 307076 218424
rect 307680 217002 307708 219234
rect 308496 218068 308548 218074
rect 308496 218010 308548 218016
rect 308508 217002 308536 218010
rect 304828 216974 304888 217002
rect 305716 216974 306144 217002
rect 306544 216974 306880 217002
rect 307372 216974 307708 217002
rect 308200 216974 308536 217002
rect 308876 217002 308904 227258
rect 309060 218074 309088 228346
rect 309704 219434 309732 229026
rect 309888 224806 309916 231676
rect 309876 224800 309928 224806
rect 309876 224742 309928 224748
rect 310152 220516 310204 220522
rect 310152 220458 310204 220464
rect 309704 219406 309824 219434
rect 309796 219026 309824 219406
rect 309784 219020 309836 219026
rect 309784 218962 309836 218968
rect 309048 218068 309100 218074
rect 309048 218010 309100 218016
rect 310164 217002 310192 220458
rect 310532 219842 310560 231676
rect 311176 226914 311204 231676
rect 311452 231662 311834 231690
rect 311164 226908 311216 226914
rect 311164 226850 311216 226856
rect 311452 220658 311480 231662
rect 311900 230444 311952 230450
rect 311900 230386 311952 230392
rect 311912 223802 311940 230386
rect 312464 227186 312492 231676
rect 313108 229362 313136 231676
rect 313096 229356 313148 229362
rect 313096 229298 313148 229304
rect 312912 228948 312964 228954
rect 312912 228890 312964 228896
rect 312452 227180 312504 227186
rect 312452 227122 312504 227128
rect 311820 223774 311940 223802
rect 311440 220652 311492 220658
rect 311440 220594 311492 220600
rect 311624 220652 311676 220658
rect 311624 220594 311676 220600
rect 310520 219836 310572 219842
rect 310520 219778 310572 219784
rect 310980 218068 311032 218074
rect 310980 218010 311032 218016
rect 310992 217002 311020 218010
rect 311636 217002 311664 220594
rect 311820 218074 311848 223774
rect 311808 218068 311860 218074
rect 311808 218010 311860 218016
rect 312636 218068 312688 218074
rect 312636 218010 312688 218016
rect 312648 217002 312676 218010
rect 308876 216974 309028 217002
rect 309856 216974 310192 217002
rect 310684 216974 311020 217002
rect 311512 216974 311664 217002
rect 312340 216974 312676 217002
rect 312924 217002 312952 228890
rect 313096 224800 313148 224806
rect 313096 224742 313148 224748
rect 313108 218074 313136 224742
rect 313752 222902 313780 231676
rect 313936 231662 314410 231690
rect 314856 231662 315054 231690
rect 315408 231662 315698 231690
rect 313740 222896 313792 222902
rect 313740 222838 313792 222844
rect 313936 220946 313964 231662
rect 314856 221882 314884 231662
rect 315408 223582 315436 231662
rect 316328 224534 316356 231676
rect 316604 231662 316986 231690
rect 316316 224528 316368 224534
rect 316316 224470 316368 224476
rect 315396 223576 315448 223582
rect 315396 223518 315448 223524
rect 315672 223304 315724 223310
rect 315672 223246 315724 223252
rect 314844 221876 314896 221882
rect 314844 221818 314896 221824
rect 313752 220918 313964 220946
rect 313752 220114 313780 220918
rect 313924 220788 313976 220794
rect 313924 220730 313976 220736
rect 313740 220108 313792 220114
rect 313740 220050 313792 220056
rect 313936 218890 313964 220730
rect 314292 219020 314344 219026
rect 314292 218962 314344 218968
rect 313924 218884 313976 218890
rect 313924 218826 313976 218832
rect 313096 218068 313148 218074
rect 313096 218010 313148 218016
rect 314304 217002 314332 218962
rect 315684 218074 315712 223246
rect 315856 222896 315908 222902
rect 315856 222838 315908 222844
rect 315120 218068 315172 218074
rect 315120 218010 315172 218016
rect 315672 218068 315724 218074
rect 315672 218010 315724 218016
rect 315132 217002 315160 218010
rect 315868 217002 315896 222838
rect 316604 220250 316632 231662
rect 316868 224528 316920 224534
rect 316868 224470 316920 224476
rect 316592 220244 316644 220250
rect 316592 220186 316644 220192
rect 316880 217002 316908 224470
rect 317616 224262 317644 231676
rect 318260 229906 318288 231676
rect 318248 229900 318300 229906
rect 318248 229842 318300 229848
rect 318064 229764 318116 229770
rect 318064 229706 318116 229712
rect 317604 224256 317656 224262
rect 317604 224198 317656 224204
rect 318076 218074 318104 229706
rect 318904 228818 318932 231676
rect 318892 228812 318944 228818
rect 318892 228754 318944 228760
rect 319548 226302 319576 231676
rect 319812 227180 319864 227186
rect 319812 227122 319864 227128
rect 319536 226296 319588 226302
rect 319536 226238 319588 226244
rect 318432 220108 318484 220114
rect 318432 220050 318484 220056
rect 317328 218068 317380 218074
rect 317328 218010 317380 218016
rect 318064 218068 318116 218074
rect 318064 218010 318116 218016
rect 317340 217002 317368 218010
rect 318444 217002 318472 220050
rect 319260 218068 319312 218074
rect 319260 218010 319312 218016
rect 319272 217002 319300 218010
rect 319824 217002 319852 227122
rect 320192 227050 320220 231676
rect 320376 231662 320850 231690
rect 320180 227044 320232 227050
rect 320180 226986 320232 226992
rect 319996 225888 320048 225894
rect 319996 225830 320048 225836
rect 320008 218074 320036 225830
rect 320376 220794 320404 231662
rect 320824 229084 320876 229090
rect 320824 229026 320876 229032
rect 320836 228818 320864 229026
rect 320824 228812 320876 228818
rect 320824 228754 320876 228760
rect 321480 225622 321508 231676
rect 321848 231662 322138 231690
rect 321468 225616 321520 225622
rect 321468 225558 321520 225564
rect 321468 224936 321520 224942
rect 321468 224878 321520 224884
rect 320364 220788 320416 220794
rect 320364 220730 320416 220736
rect 320916 218612 320968 218618
rect 320916 218554 320968 218560
rect 319996 218068 320048 218074
rect 319996 218010 320048 218016
rect 320928 217002 320956 218554
rect 321480 217002 321508 224878
rect 321848 222766 321876 231662
rect 322768 228546 322796 231676
rect 323412 230178 323440 231676
rect 323400 230172 323452 230178
rect 323400 230114 323452 230120
rect 323584 230172 323636 230178
rect 323584 230114 323636 230120
rect 322756 228540 322808 228546
rect 322756 228482 322808 228488
rect 322572 224256 322624 224262
rect 322572 224198 322624 224204
rect 321836 222760 321888 222766
rect 321836 222702 321888 222708
rect 322584 217002 322612 224198
rect 322848 223440 322900 223446
rect 322848 223382 322900 223388
rect 322860 219162 322888 223382
rect 323400 219428 323452 219434
rect 323400 219370 323452 219376
rect 322848 219156 322900 219162
rect 322848 219098 322900 219104
rect 323412 217002 323440 219370
rect 323596 218754 323624 230114
rect 324056 229094 324084 231676
rect 324700 230178 324728 231676
rect 324688 230172 324740 230178
rect 324688 230114 324740 230120
rect 324964 229900 325016 229906
rect 324964 229842 325016 229848
rect 323872 229066 324084 229094
rect 323872 224398 323900 229066
rect 324044 225616 324096 225622
rect 324044 225558 324096 225564
rect 323860 224392 323912 224398
rect 323860 224334 323912 224340
rect 324056 219434 324084 225558
rect 324976 224954 325004 229842
rect 325344 227594 325372 231676
rect 325332 227588 325384 227594
rect 325332 227530 325384 227536
rect 325516 227044 325568 227050
rect 325516 226986 325568 226992
rect 324884 224926 325004 224954
rect 324884 219434 324912 224926
rect 325528 219434 325556 226986
rect 325988 224670 326016 231676
rect 325976 224664 326028 224670
rect 325976 224606 326028 224612
rect 326632 223038 326660 231676
rect 327276 228818 327304 231676
rect 327552 231662 327934 231690
rect 327264 228812 327316 228818
rect 327264 228754 327316 228760
rect 326804 228540 326856 228546
rect 326804 228482 326856 228488
rect 326620 223032 326672 223038
rect 326620 222974 326672 222980
rect 324044 219428 324096 219434
rect 324044 219370 324096 219376
rect 324228 219428 324280 219434
rect 324228 219370 324280 219376
rect 324872 219428 324924 219434
rect 324872 219370 324924 219376
rect 325056 219428 325108 219434
rect 325056 219370 325108 219376
rect 325516 219428 325568 219434
rect 325516 219370 325568 219376
rect 323584 218748 323636 218754
rect 323584 218690 323636 218696
rect 324240 217002 324268 219370
rect 325068 217002 325096 219370
rect 325608 219156 325660 219162
rect 325608 219098 325660 219104
rect 325620 217002 325648 219098
rect 326816 217002 326844 228482
rect 327552 221610 327580 231662
rect 327724 229084 327776 229090
rect 327724 229026 327776 229032
rect 327540 221604 327592 221610
rect 327540 221546 327592 221552
rect 327736 219434 327764 229026
rect 328564 221746 328592 231676
rect 329208 226166 329236 231676
rect 329852 230042 329880 231676
rect 330128 231662 330510 231690
rect 329840 230036 329892 230042
rect 329840 229978 329892 229984
rect 329196 226160 329248 226166
rect 329196 226102 329248 226108
rect 330128 223174 330156 231662
rect 331140 227458 331168 231676
rect 331416 231662 331798 231690
rect 331128 227452 331180 227458
rect 331128 227394 331180 227400
rect 330484 226160 330536 226166
rect 330484 226102 330536 226108
rect 330116 223168 330168 223174
rect 330116 223110 330168 223116
rect 329748 223032 329800 223038
rect 329748 222974 329800 222980
rect 328552 221740 328604 221746
rect 328552 221682 328604 221688
rect 328368 221604 328420 221610
rect 328368 221546 328420 221552
rect 327724 219428 327776 219434
rect 327724 219370 327776 219376
rect 327540 219292 327592 219298
rect 327540 219234 327592 219240
rect 327552 217002 327580 219234
rect 328380 217002 328408 221546
rect 329196 220244 329248 220250
rect 329196 220186 329248 220192
rect 329208 217002 329236 220186
rect 329760 217002 329788 222974
rect 330496 219162 330524 226102
rect 330852 222148 330904 222154
rect 330852 222090 330904 222096
rect 330484 219156 330536 219162
rect 330484 219098 330536 219104
rect 330864 217002 330892 222090
rect 331416 220386 331444 231662
rect 332428 223446 332456 231676
rect 333072 226030 333100 231676
rect 333716 228682 333744 231676
rect 334084 231662 334374 231690
rect 333704 228676 333756 228682
rect 333704 228618 333756 228624
rect 333888 227452 333940 227458
rect 333888 227394 333940 227400
rect 333060 226024 333112 226030
rect 333060 225966 333112 225972
rect 332416 223440 332468 223446
rect 332416 223382 332468 223388
rect 331680 221740 331732 221746
rect 331680 221682 331732 221688
rect 331404 220380 331456 220386
rect 331404 220322 331456 220328
rect 331692 217002 331720 221682
rect 333704 218748 333756 218754
rect 333704 218690 333756 218696
rect 332508 218204 332560 218210
rect 332508 218146 332560 218152
rect 332520 217002 332548 218146
rect 333336 218068 333388 218074
rect 333336 218010 333388 218016
rect 333348 217002 333376 218010
rect 312924 216974 313168 217002
rect 313996 216974 314332 217002
rect 314824 216974 315160 217002
rect 315652 216974 315896 217002
rect 316480 216974 316908 217002
rect 317308 216974 317368 217002
rect 318136 216974 318472 217002
rect 318964 216974 319300 217002
rect 319792 216974 319852 217002
rect 320620 216974 320956 217002
rect 321448 216974 321508 217002
rect 322276 216974 322612 217002
rect 323104 216974 323440 217002
rect 323932 216974 324268 217002
rect 324760 216974 325096 217002
rect 325588 216974 325648 217002
rect 326416 216974 326844 217002
rect 327244 216974 327580 217002
rect 328072 216974 328408 217002
rect 328900 216974 329236 217002
rect 329728 216974 329788 217002
rect 330556 216974 330892 217002
rect 331384 216974 331720 217002
rect 332212 216974 332548 217002
rect 333040 216974 333376 217002
rect 333716 217002 333744 218690
rect 333900 218074 333928 227394
rect 334084 221474 334112 231662
rect 335004 230314 335032 231676
rect 335464 231662 335662 231690
rect 334992 230308 335044 230314
rect 334992 230250 335044 230256
rect 335084 228812 335136 228818
rect 335084 228754 335136 228760
rect 334072 221468 334124 221474
rect 334072 221410 334124 221416
rect 333888 218068 333940 218074
rect 333888 218010 333940 218016
rect 335096 217002 335124 228754
rect 335464 222018 335492 231662
rect 336292 228410 336320 231676
rect 336280 228404 336332 228410
rect 336280 228346 336332 228352
rect 336648 228404 336700 228410
rect 336648 228346 336700 228352
rect 336464 223168 336516 223174
rect 336464 223110 336516 223116
rect 335452 222012 335504 222018
rect 335452 221954 335504 221960
rect 335268 221468 335320 221474
rect 335268 221410 335320 221416
rect 335280 218210 335308 221410
rect 335268 218204 335320 218210
rect 335268 218146 335320 218152
rect 336476 218074 336504 223110
rect 335820 218068 335872 218074
rect 335820 218010 335872 218016
rect 336464 218068 336516 218074
rect 336464 218010 336516 218016
rect 335832 217002 335860 218010
rect 336660 217002 336688 228346
rect 336936 225758 336964 231676
rect 337580 229090 337608 231676
rect 337844 230036 337896 230042
rect 337844 229978 337896 229984
rect 337568 229084 337620 229090
rect 337568 229026 337620 229032
rect 336924 225752 336976 225758
rect 336924 225694 336976 225700
rect 337856 219434 337884 229978
rect 338224 220522 338252 231676
rect 338592 231662 338882 231690
rect 338592 220658 338620 231662
rect 339512 227322 339540 231676
rect 340156 230450 340184 231676
rect 340144 230444 340196 230450
rect 340144 230386 340196 230392
rect 340800 228954 340828 231676
rect 340788 228948 340840 228954
rect 340788 228890 340840 228896
rect 340144 228676 340196 228682
rect 340144 228618 340196 228624
rect 339500 227316 339552 227322
rect 339500 227258 339552 227264
rect 338948 220788 339000 220794
rect 338948 220730 339000 220736
rect 338580 220652 338632 220658
rect 338580 220594 338632 220600
rect 338212 220516 338264 220522
rect 338212 220458 338264 220464
rect 338028 220380 338080 220386
rect 338028 220322 338080 220328
rect 337580 219406 337884 219434
rect 337580 217002 337608 219406
rect 338040 217002 338068 220322
rect 338960 219026 338988 220730
rect 338948 219020 339000 219026
rect 338948 218962 339000 218968
rect 340156 218210 340184 228618
rect 340696 225752 340748 225758
rect 340696 225694 340748 225700
rect 340512 219020 340564 219026
rect 340512 218962 340564 218968
rect 339132 218204 339184 218210
rect 339132 218146 339184 218152
rect 340144 218204 340196 218210
rect 340144 218146 340196 218152
rect 339144 217002 339172 218146
rect 339960 218068 340012 218074
rect 339960 218010 340012 218016
rect 339972 217002 340000 218010
rect 340524 217002 340552 218962
rect 340708 218074 340736 225694
rect 341444 223310 341472 231676
rect 342088 224806 342116 231676
rect 342456 231662 342746 231690
rect 343008 231662 343390 231690
rect 343836 231662 344034 231690
rect 342076 224800 342128 224806
rect 342076 224742 342128 224748
rect 341892 224392 341944 224398
rect 341892 224334 341944 224340
rect 341432 223304 341484 223310
rect 341432 223246 341484 223252
rect 340696 218068 340748 218074
rect 340696 218010 340748 218016
rect 341616 218068 341668 218074
rect 341616 218010 341668 218016
rect 341628 217002 341656 218010
rect 333716 216974 333868 217002
rect 334696 216974 335124 217002
rect 335524 216974 335860 217002
rect 336352 216974 336688 217002
rect 337180 216974 337608 217002
rect 338008 216974 338068 217002
rect 338836 216974 339172 217002
rect 339664 216974 340000 217002
rect 340492 216974 340552 217002
rect 341320 216974 341656 217002
rect 341904 217002 341932 224334
rect 342076 223304 342128 223310
rect 342076 223246 342128 223252
rect 342088 218074 342116 223246
rect 342456 220794 342484 231662
rect 343008 224534 343036 231662
rect 342996 224528 343048 224534
rect 342996 224470 343048 224476
rect 343364 224528 343416 224534
rect 343364 224470 343416 224476
rect 342444 220788 342496 220794
rect 342444 220730 342496 220736
rect 342720 220516 342772 220522
rect 342720 220458 342772 220464
rect 342732 219298 342760 220458
rect 342720 219292 342772 219298
rect 342720 219234 342772 219240
rect 342076 218068 342128 218074
rect 342076 218010 342128 218016
rect 343376 217002 343404 224470
rect 343640 220108 343692 220114
rect 343640 220050 343692 220056
rect 343652 218890 343680 220050
rect 343836 219978 343864 231662
rect 344664 222902 344692 231676
rect 345308 229770 345336 231676
rect 345860 231662 345966 231690
rect 345296 229764 345348 229770
rect 345296 229706 345348 229712
rect 345664 229764 345716 229770
rect 345664 229706 345716 229712
rect 344652 222896 344704 222902
rect 344652 222838 344704 222844
rect 345676 222154 345704 229706
rect 345860 227186 345888 231662
rect 345848 227180 345900 227186
rect 345848 227122 345900 227128
rect 346032 227180 346084 227186
rect 346032 227122 346084 227128
rect 345664 222148 345716 222154
rect 345664 222090 345716 222096
rect 344928 221876 344980 221882
rect 344928 221818 344980 221824
rect 343824 219972 343876 219978
rect 343824 219914 343876 219920
rect 343640 218884 343692 218890
rect 343640 218826 343692 218832
rect 344100 218340 344152 218346
rect 344100 218282 344152 218288
rect 344112 217002 344140 218282
rect 344940 217002 344968 221818
rect 345756 218068 345808 218074
rect 345756 218010 345808 218016
rect 345768 217002 345796 218010
rect 341904 216974 342148 217002
rect 342976 216974 343404 217002
rect 343804 216974 344140 217002
rect 344632 216974 344968 217002
rect 345460 216974 345796 217002
rect 346044 217002 346072 227122
rect 346596 224942 346624 231676
rect 347240 225894 347268 231676
rect 347228 225888 347280 225894
rect 347228 225830 347280 225836
rect 346584 224936 346636 224942
rect 346584 224878 346636 224884
rect 347044 224664 347096 224670
rect 347044 224606 347096 224612
rect 346216 222896 346268 222902
rect 346216 222838 346268 222844
rect 346228 218074 346256 222838
rect 347056 218346 347084 224606
rect 347884 220114 347912 231676
rect 348528 225622 348556 231676
rect 349172 227050 349200 231676
rect 349160 227044 349212 227050
rect 349160 226986 349212 226992
rect 348516 225616 348568 225622
rect 348516 225558 348568 225564
rect 349068 225616 349120 225622
rect 349068 225558 349120 225564
rect 347872 220108 347924 220114
rect 347872 220050 347924 220056
rect 347412 218884 347464 218890
rect 347412 218826 347464 218832
rect 347044 218340 347096 218346
rect 347044 218282 347096 218288
rect 346216 218068 346268 218074
rect 346216 218010 346268 218016
rect 347424 217002 347452 218826
rect 348884 218204 348936 218210
rect 348884 218146 348936 218152
rect 348240 218068 348292 218074
rect 348240 218010 348292 218016
rect 348252 217002 348280 218010
rect 348896 217002 348924 218146
rect 349080 218074 349108 225558
rect 349816 224262 349844 231676
rect 350460 229906 350488 231676
rect 350448 229900 350500 229906
rect 350448 229842 350500 229848
rect 349988 228948 350040 228954
rect 349988 228890 350040 228896
rect 349804 224256 349856 224262
rect 349804 224198 349856 224204
rect 349068 218068 349120 218074
rect 349068 218010 349120 218016
rect 350000 217002 350028 228890
rect 351104 228546 351132 231676
rect 351288 231662 351762 231690
rect 351932 231662 352406 231690
rect 352576 231662 353050 231690
rect 351288 229094 351316 231662
rect 351288 229066 351408 229094
rect 351092 228540 351144 228546
rect 351092 228482 351144 228488
rect 351184 227316 351236 227322
rect 351184 227258 351236 227264
rect 350356 225956 350408 225962
rect 350356 225898 350408 225904
rect 346044 216974 346288 217002
rect 347116 216974 347452 217002
rect 347944 216974 348280 217002
rect 348772 216974 348924 217002
rect 349600 216974 350028 217002
rect 350368 217002 350396 225898
rect 351196 219026 351224 227258
rect 351380 221610 351408 229066
rect 351932 226166 351960 231662
rect 352576 229094 352604 231662
rect 352392 229066 352604 229094
rect 351920 226160 351972 226166
rect 351920 226102 351972 226108
rect 351644 224256 351696 224262
rect 351644 224198 351696 224204
rect 351368 221604 351420 221610
rect 351368 221546 351420 221552
rect 351184 219020 351236 219026
rect 351184 218962 351236 218968
rect 351656 217002 351684 224198
rect 352392 220522 352420 229066
rect 352564 226160 352616 226166
rect 352564 226102 352616 226108
rect 352380 220516 352432 220522
rect 352380 220458 352432 220464
rect 352576 218754 352604 226102
rect 353680 223038 353708 231676
rect 353956 231662 354338 231690
rect 354692 231662 354982 231690
rect 353668 223032 353720 223038
rect 353668 222974 353720 222980
rect 353956 221746 353984 231662
rect 353944 221740 353996 221746
rect 353944 221682 353996 221688
rect 353392 221604 353444 221610
rect 353392 221546 353444 221552
rect 353208 220516 353260 220522
rect 353208 220458 353260 220464
rect 352564 218748 352616 218754
rect 352564 218690 352616 218696
rect 352380 218068 352432 218074
rect 352380 218010 352432 218016
rect 352392 217002 352420 218010
rect 353220 217002 353248 220458
rect 353404 218210 353432 221546
rect 354692 220250 354720 231662
rect 354864 230172 354916 230178
rect 354864 230114 354916 230120
rect 354876 225962 354904 230114
rect 355612 229770 355640 231676
rect 355600 229764 355652 229770
rect 355600 229706 355652 229712
rect 356256 227458 356284 231676
rect 356900 228818 356928 231676
rect 357072 229764 357124 229770
rect 357072 229706 357124 229712
rect 356888 228812 356940 228818
rect 356888 228754 356940 228760
rect 356244 227452 356296 227458
rect 356244 227394 356296 227400
rect 354864 225956 354916 225962
rect 354864 225898 354916 225904
rect 355324 225888 355376 225894
rect 355324 225830 355376 225836
rect 354680 220244 354732 220250
rect 354680 220186 354732 220192
rect 354312 220108 354364 220114
rect 354312 220050 354364 220056
rect 354036 218748 354088 218754
rect 354036 218690 354088 218696
rect 353392 218204 353444 218210
rect 353392 218146 353444 218152
rect 354048 217002 354076 218690
rect 354324 218074 354352 220050
rect 355336 219298 355364 225830
rect 355784 223032 355836 223038
rect 355784 222974 355836 222980
rect 354588 219292 354640 219298
rect 354588 219234 354640 219240
rect 355324 219292 355376 219298
rect 355324 219234 355376 219240
rect 354312 218068 354364 218074
rect 354312 218010 354364 218016
rect 354600 217002 354628 219234
rect 355796 217002 355824 222974
rect 356520 218068 356572 218074
rect 356520 218010 356572 218016
rect 356532 217002 356560 218010
rect 357084 217002 357112 229706
rect 357256 227044 357308 227050
rect 357256 226986 357308 226992
rect 357268 218074 357296 226986
rect 357544 221474 357572 231676
rect 358188 226166 358216 231676
rect 358832 228410 358860 231676
rect 359016 231662 359490 231690
rect 359752 231662 360134 231690
rect 358820 228404 358872 228410
rect 358820 228346 358872 228352
rect 358176 226160 358228 226166
rect 358176 226102 358228 226108
rect 357532 221468 357584 221474
rect 357532 221410 357584 221416
rect 358176 221468 358228 221474
rect 358176 221410 358228 221416
rect 357256 218068 357308 218074
rect 357256 218010 357308 218016
rect 358188 217002 358216 221410
rect 359016 220386 359044 231662
rect 359752 223174 359780 231662
rect 360764 230042 360792 231676
rect 360752 230036 360804 230042
rect 360752 229978 360804 229984
rect 361212 229900 361264 229906
rect 361212 229842 361264 229848
rect 361224 229094 361252 229842
rect 361408 229094 361436 231676
rect 361224 229066 361344 229094
rect 361408 229066 361528 229094
rect 359924 228404 359976 228410
rect 359924 228346 359976 228352
rect 359740 223168 359792 223174
rect 359740 223110 359792 223116
rect 359004 220380 359056 220386
rect 359004 220322 359056 220328
rect 358728 218204 358780 218210
rect 358728 218146 358780 218152
rect 358740 217002 358768 218146
rect 359936 217002 359964 228346
rect 361316 218074 361344 229066
rect 361500 225758 361528 229066
rect 361488 225752 361540 225758
rect 361488 225694 361540 225700
rect 362052 223310 362080 231676
rect 362696 228682 362724 231676
rect 362684 228676 362736 228682
rect 362684 228618 362736 228624
rect 362592 228540 362644 228546
rect 362592 228482 362644 228488
rect 362040 223304 362092 223310
rect 362040 223246 362092 223252
rect 362316 221740 362368 221746
rect 362316 221682 362368 221688
rect 361488 220244 361540 220250
rect 361488 220186 361540 220192
rect 360660 218068 360712 218074
rect 360660 218010 360712 218016
rect 361304 218068 361356 218074
rect 361304 218010 361356 218016
rect 360672 217002 360700 218010
rect 361500 217002 361528 220186
rect 362328 217002 362356 221682
rect 350368 216974 350428 217002
rect 351256 216974 351684 217002
rect 352084 216974 352420 217002
rect 352912 216974 353248 217002
rect 353740 216974 354076 217002
rect 354568 216974 354628 217002
rect 355396 216974 355824 217002
rect 356224 216974 356560 217002
rect 357052 216974 357112 217002
rect 357880 216974 358216 217002
rect 358708 216974 358768 217002
rect 359536 216974 359964 217002
rect 360364 216974 360700 217002
rect 361192 216974 361528 217002
rect 362020 216974 362356 217002
rect 362604 217002 362632 228482
rect 363340 227322 363368 231676
rect 363328 227316 363380 227322
rect 363328 227258 363380 227264
rect 363604 227316 363656 227322
rect 363604 227258 363656 227264
rect 363616 218890 363644 227258
rect 363984 224670 364012 231676
rect 364536 231662 364642 231690
rect 363972 224664 364024 224670
rect 363972 224606 364024 224612
rect 363788 224528 363840 224534
rect 363788 224470 363840 224476
rect 363604 218884 363656 218890
rect 363604 218826 363656 218832
rect 363800 218210 363828 224470
rect 364536 221882 364564 231662
rect 365272 224398 365300 231676
rect 365536 225752 365588 225758
rect 365536 225694 365588 225700
rect 365260 224392 365312 224398
rect 365260 224334 365312 224340
rect 364524 221876 364576 221882
rect 364524 221818 364576 221824
rect 363972 219156 364024 219162
rect 363972 219098 364024 219104
rect 363788 218204 363840 218210
rect 363788 218146 363840 218152
rect 363984 217002 364012 219098
rect 365352 218476 365404 218482
rect 365352 218418 365404 218424
rect 364800 218068 364852 218074
rect 364800 218010 364852 218016
rect 364812 217002 364840 218010
rect 365364 217002 365392 218418
rect 365548 218074 365576 225694
rect 365916 224806 365944 231676
rect 366560 227186 366588 231676
rect 366548 227180 366600 227186
rect 366548 227122 366600 227128
rect 367204 225622 367232 231676
rect 367480 231662 367862 231690
rect 367192 225616 367244 225622
rect 367192 225558 367244 225564
rect 365904 224800 365956 224806
rect 365904 224742 365956 224748
rect 366916 223304 366968 223310
rect 366916 223246 366968 223252
rect 366732 223168 366784 223174
rect 366732 223110 366784 223116
rect 365536 218068 365588 218074
rect 365536 218010 365588 218016
rect 366456 218068 366508 218074
rect 366456 218010 366508 218016
rect 366468 217002 366496 218010
rect 362604 216974 362848 217002
rect 363676 216974 364012 217002
rect 364504 216974 364840 217002
rect 365332 216974 365392 217002
rect 366160 216974 366496 217002
rect 366744 217002 366772 223110
rect 366928 218074 366956 223246
rect 367480 222902 367508 231662
rect 368492 227322 368520 231676
rect 369136 228954 369164 231676
rect 369780 229094 369808 231676
rect 369596 229066 369808 229094
rect 369964 231662 370438 231690
rect 369124 228948 369176 228954
rect 369124 228890 369176 228896
rect 368480 227316 368532 227322
rect 368480 227258 368532 227264
rect 367744 225004 367796 225010
rect 367744 224946 367796 224952
rect 367468 222896 367520 222902
rect 367468 222838 367520 222844
rect 367756 218754 367784 224946
rect 368204 224392 368256 224398
rect 368204 224334 368256 224340
rect 367744 218748 367796 218754
rect 367744 218690 367796 218696
rect 366916 218068 366968 218074
rect 366916 218010 366968 218016
rect 368216 217002 368244 224334
rect 369596 224262 369624 229066
rect 369768 227180 369820 227186
rect 369768 227122 369820 227128
rect 369584 224256 369636 224262
rect 369584 224198 369636 224204
rect 368940 218068 368992 218074
rect 368940 218010 368992 218016
rect 368952 217002 368980 218010
rect 369780 217002 369808 227122
rect 369964 221610 369992 231662
rect 371068 230178 371096 231676
rect 371436 231662 371726 231690
rect 371056 230172 371108 230178
rect 371056 230114 371108 230120
rect 371056 228676 371108 228682
rect 371056 228618 371108 228624
rect 369952 221604 370004 221610
rect 369952 221546 370004 221552
rect 370504 221604 370556 221610
rect 370504 221546 370556 221552
rect 370516 218482 370544 221546
rect 370504 218476 370556 218482
rect 370504 218418 370556 218424
rect 370596 218340 370648 218346
rect 370596 218282 370648 218288
rect 370608 217002 370636 218282
rect 366744 216974 366988 217002
rect 367816 216974 368244 217002
rect 368644 216974 368980 217002
rect 369472 216974 369808 217002
rect 370300 216974 370636 217002
rect 371068 217002 371096 228618
rect 371436 220522 371464 231662
rect 372356 225894 372384 231676
rect 372816 231662 373014 231690
rect 372344 225888 372396 225894
rect 372344 225830 372396 225836
rect 372344 224256 372396 224262
rect 372344 224198 372396 224204
rect 371424 220516 371476 220522
rect 371424 220458 371476 220464
rect 372356 217002 372384 224198
rect 372528 220380 372580 220386
rect 372528 220322 372580 220328
rect 372540 218074 372568 220322
rect 372816 220114 372844 231662
rect 373644 225010 373672 231676
rect 373816 228812 373868 228818
rect 373816 228754 373868 228760
rect 373632 225004 373684 225010
rect 373632 224946 373684 224952
rect 372804 220108 372856 220114
rect 372804 220050 372856 220056
rect 373632 219428 373684 219434
rect 373632 219370 373684 219376
rect 372528 218068 372580 218074
rect 372528 218010 372580 218016
rect 372988 218068 373040 218074
rect 372988 218010 373040 218016
rect 373000 217002 373028 218010
rect 373644 217002 373672 219370
rect 373828 218074 373856 228754
rect 374288 227050 374316 231676
rect 374564 231662 374946 231690
rect 374276 227044 374328 227050
rect 374276 226986 374328 226992
rect 374564 221474 374592 231662
rect 375288 225616 375340 225622
rect 375288 225558 375340 225564
rect 374552 221468 374604 221474
rect 374552 221410 374604 221416
rect 374000 221196 374052 221202
rect 374000 221138 374052 221144
rect 374012 219162 374040 221138
rect 374000 219156 374052 219162
rect 374000 219098 374052 219104
rect 375104 218204 375156 218210
rect 375104 218146 375156 218152
rect 373816 218068 373868 218074
rect 373816 218010 373868 218016
rect 374736 218068 374788 218074
rect 374736 218010 374788 218016
rect 374748 217002 374776 218010
rect 371068 216974 371128 217002
rect 371956 216974 372384 217002
rect 372784 216974 373028 217002
rect 373612 216974 373672 217002
rect 374440 216974 374776 217002
rect 375116 217002 375144 218146
rect 375300 218074 375328 225558
rect 375576 223038 375604 231676
rect 376024 230308 376076 230314
rect 376024 230250 376076 230256
rect 375564 223032 375616 223038
rect 375564 222974 375616 222980
rect 376036 221746 376064 230250
rect 376220 229770 376248 231676
rect 376208 229764 376260 229770
rect 376208 229706 376260 229712
rect 376864 228410 376892 231676
rect 377048 231662 377522 231690
rect 376852 228404 376904 228410
rect 376852 228346 376904 228352
rect 376484 227044 376536 227050
rect 376484 226986 376536 226992
rect 376024 221740 376076 221746
rect 376024 221682 376076 221688
rect 375472 221468 375524 221474
rect 375472 221410 375524 221416
rect 375484 218346 375512 221410
rect 375472 218340 375524 218346
rect 375472 218282 375524 218288
rect 375288 218068 375340 218074
rect 375288 218010 375340 218016
rect 376496 217002 376524 226986
rect 377048 223156 377076 231662
rect 377956 228948 378008 228954
rect 377956 228890 378008 228896
rect 376864 223128 377076 223156
rect 376864 220250 376892 223128
rect 376852 220244 376904 220250
rect 376852 220186 376904 220192
rect 377036 220244 377088 220250
rect 377036 220186 377088 220192
rect 377048 219434 377076 220186
rect 377968 219434 377996 228890
rect 378152 224534 378180 231676
rect 378796 229906 378824 231676
rect 378784 229900 378836 229906
rect 378784 229842 378836 229848
rect 379440 228546 379468 231676
rect 379428 228540 379480 228546
rect 379428 228482 379480 228488
rect 378968 228404 379020 228410
rect 378968 228346 379020 228352
rect 378140 224528 378192 224534
rect 378140 224470 378192 224476
rect 377036 219428 377088 219434
rect 377968 219406 378088 219434
rect 377036 219370 377088 219376
rect 377220 218340 377272 218346
rect 377220 218282 377272 218288
rect 377232 217002 377260 218282
rect 378060 217002 378088 219406
rect 378980 217002 379008 228346
rect 380084 225758 380112 231676
rect 380728 230314 380756 231676
rect 381096 231662 381386 231690
rect 380716 230308 380768 230314
rect 380716 230250 380768 230256
rect 380716 229764 380768 229770
rect 380716 229706 380768 229712
rect 380072 225752 380124 225758
rect 380072 225694 380124 225700
rect 380256 225752 380308 225758
rect 380256 225694 380308 225700
rect 379428 220108 379480 220114
rect 379428 220050 379480 220056
rect 379440 217002 379468 220050
rect 380268 219434 380296 225694
rect 380728 219434 380756 229706
rect 381096 221202 381124 231662
rect 382016 223310 382044 231676
rect 382660 229094 382688 231676
rect 382844 231662 383318 231690
rect 382844 229094 382872 231662
rect 382568 229066 382688 229094
rect 382752 229066 382872 229094
rect 382568 224398 382596 229066
rect 382556 224392 382608 224398
rect 382556 224334 382608 224340
rect 382004 223304 382056 223310
rect 382004 223246 382056 223252
rect 382096 223032 382148 223038
rect 382096 222974 382148 222980
rect 381084 221196 381136 221202
rect 381084 221138 381136 221144
rect 380176 219406 380296 219434
rect 380636 219406 380756 219434
rect 380176 218210 380204 219406
rect 380164 218204 380216 218210
rect 380164 218146 380216 218152
rect 380636 217002 380664 219406
rect 381912 218204 381964 218210
rect 381912 218146 381964 218152
rect 381360 218068 381412 218074
rect 381360 218010 381412 218016
rect 381372 217002 381400 218010
rect 381924 217002 381952 218146
rect 382108 218074 382136 222974
rect 382752 221746 382780 229066
rect 382924 224392 382976 224398
rect 382924 224334 382976 224340
rect 382740 221740 382792 221746
rect 382740 221682 382792 221688
rect 382740 221604 382792 221610
rect 382740 221546 382792 221552
rect 382096 218068 382148 218074
rect 382096 218010 382148 218016
rect 382752 217002 382780 221546
rect 382936 218210 382964 224334
rect 383948 223174 383976 231676
rect 384592 227186 384620 231676
rect 385236 228682 385264 231676
rect 385420 231662 385894 231690
rect 385224 228676 385276 228682
rect 385224 228618 385276 228624
rect 384580 227180 384632 227186
rect 384580 227122 384632 227128
rect 384764 226908 384816 226914
rect 384764 226850 384816 226856
rect 383936 223168 383988 223174
rect 383936 223110 383988 223116
rect 383568 219020 383620 219026
rect 383568 218962 383620 218968
rect 382924 218204 382976 218210
rect 382924 218146 382976 218152
rect 383580 217002 383608 218962
rect 384776 217002 384804 226850
rect 385420 220386 385448 231662
rect 385684 226364 385736 226370
rect 385684 226306 385736 226312
rect 385408 220380 385460 220386
rect 385408 220322 385460 220328
rect 385696 218346 385724 226306
rect 386328 222896 386380 222902
rect 386328 222838 386380 222844
rect 386144 218748 386196 218754
rect 386144 218690 386196 218696
rect 385684 218340 385736 218346
rect 385684 218282 385736 218288
rect 385500 218068 385552 218074
rect 385500 218010 385552 218016
rect 385512 217002 385540 218010
rect 386156 217002 386184 218690
rect 386340 218074 386368 222838
rect 386524 221474 386552 231676
rect 387168 228818 387196 231676
rect 387432 230376 387484 230382
rect 387432 230318 387484 230324
rect 387156 228812 387208 228818
rect 387156 228754 387208 228760
rect 387444 224262 387472 230318
rect 387812 225622 387840 231676
rect 388456 230382 388484 231676
rect 388640 231662 389114 231690
rect 388444 230376 388496 230382
rect 388444 230318 388496 230324
rect 388444 225888 388496 225894
rect 388444 225830 388496 225836
rect 387800 225616 387852 225622
rect 387800 225558 387852 225564
rect 387432 224256 387484 224262
rect 387432 224198 387484 224204
rect 387708 224256 387760 224262
rect 387708 224198 387760 224204
rect 386512 221468 386564 221474
rect 386512 221410 386564 221416
rect 387156 220992 387208 220998
rect 387156 220934 387208 220940
rect 386328 218068 386380 218074
rect 386328 218010 386380 218016
rect 387168 217002 387196 220934
rect 387720 217002 387748 224198
rect 388456 219026 388484 225830
rect 388640 220250 388668 231662
rect 389744 227050 389772 231676
rect 389916 229900 389968 229906
rect 389916 229842 389968 229848
rect 389732 227044 389784 227050
rect 389732 226986 389784 226992
rect 389928 220998 389956 229842
rect 390388 228954 390416 231676
rect 390376 228948 390428 228954
rect 390376 228890 390428 228896
rect 390192 228540 390244 228546
rect 390192 228482 390244 228488
rect 389916 220992 389968 220998
rect 389916 220934 389968 220940
rect 388628 220244 388680 220250
rect 388628 220186 388680 220192
rect 388812 219156 388864 219162
rect 388812 219098 388864 219104
rect 388444 219020 388496 219026
rect 388444 218962 388496 218968
rect 388824 217002 388852 219098
rect 390204 218074 390232 228482
rect 391032 225758 391060 231676
rect 391388 227180 391440 227186
rect 391388 227122 391440 227128
rect 391020 225752 391072 225758
rect 391020 225694 391072 225700
rect 390468 221468 390520 221474
rect 390468 221410 390520 221416
rect 389640 218068 389692 218074
rect 389640 218010 389692 218016
rect 390192 218068 390244 218074
rect 390192 218010 390244 218016
rect 389652 217002 389680 218010
rect 390480 217002 390508 221410
rect 391400 217002 391428 227122
rect 391676 226370 391704 231676
rect 392136 231662 392334 231690
rect 391664 226364 391716 226370
rect 391664 226306 391716 226312
rect 391756 225616 391808 225622
rect 391756 225558 391808 225564
rect 375116 216974 375268 217002
rect 376096 216974 376524 217002
rect 376924 216974 377260 217002
rect 377752 216974 378088 217002
rect 378580 216974 379008 217002
rect 379408 216974 379468 217002
rect 380236 216974 380664 217002
rect 381064 216974 381400 217002
rect 381892 216974 381952 217002
rect 382720 216974 382780 217002
rect 383548 216974 383608 217002
rect 384376 216974 384804 217002
rect 385204 216974 385540 217002
rect 386032 216974 386184 217002
rect 386860 216974 387196 217002
rect 387688 216974 387748 217002
rect 388516 216974 388852 217002
rect 389344 216974 389680 217002
rect 390172 216974 390508 217002
rect 391000 216974 391428 217002
rect 391768 217002 391796 225558
rect 392136 220114 392164 231662
rect 392964 223038 392992 231676
rect 393608 228410 393636 231676
rect 394252 229770 394280 231676
rect 394240 229764 394292 229770
rect 394240 229706 394292 229712
rect 393596 228404 393648 228410
rect 393596 228346 393648 228352
rect 393964 227928 394016 227934
rect 393964 227870 394016 227876
rect 392952 223032 393004 223038
rect 392952 222974 393004 222980
rect 392124 220108 392176 220114
rect 392124 220050 392176 220056
rect 393976 219162 394004 227870
rect 394516 224528 394568 224534
rect 394516 224470 394568 224476
rect 393964 219156 394016 219162
rect 393964 219098 394016 219104
rect 392952 218612 393004 218618
rect 392952 218554 393004 218560
rect 392964 217002 392992 218554
rect 394332 218204 394384 218210
rect 394332 218146 394384 218152
rect 393780 218068 393832 218074
rect 393780 218010 393832 218016
rect 393792 217002 393820 218010
rect 394344 217002 394372 218146
rect 394528 218074 394556 224470
rect 394896 221610 394924 231676
rect 395540 226914 395568 231676
rect 395712 227044 395764 227050
rect 395712 226986 395764 226992
rect 395528 226908 395580 226914
rect 395528 226850 395580 226856
rect 394884 221604 394936 221610
rect 394884 221546 394936 221552
rect 395724 219434 395752 226986
rect 396184 224398 396212 231676
rect 396552 231662 396842 231690
rect 396552 225894 396580 231662
rect 397472 227798 397500 231676
rect 396724 227792 396776 227798
rect 396724 227734 396776 227740
rect 397460 227792 397512 227798
rect 397460 227734 397512 227740
rect 396540 225888 396592 225894
rect 396540 225830 396592 225836
rect 396172 224392 396224 224398
rect 396172 224334 396224 224340
rect 395988 220108 396040 220114
rect 395988 220050 396040 220056
rect 395540 219406 395752 219434
rect 394516 218068 394568 218074
rect 394516 218010 394568 218016
rect 395540 217002 395568 219406
rect 396000 217002 396028 220050
rect 396736 218754 396764 227734
rect 398116 224262 398144 231676
rect 398392 231662 398774 231690
rect 398104 224256 398156 224262
rect 398104 224198 398156 224204
rect 398392 222902 398420 231662
rect 399404 229906 399432 231676
rect 399392 229900 399444 229906
rect 399392 229842 399444 229848
rect 399852 229764 399904 229770
rect 399852 229706 399904 229712
rect 398748 228268 398800 228274
rect 398748 228210 398800 228216
rect 398380 222896 398432 222902
rect 398380 222838 398432 222844
rect 398564 222896 398616 222902
rect 398564 222838 398616 222844
rect 397092 221604 397144 221610
rect 397092 221546 397144 221552
rect 396724 218748 396776 218754
rect 396724 218690 396776 218696
rect 397104 217002 397132 221546
rect 398576 218074 398604 222838
rect 397920 218068 397972 218074
rect 397920 218010 397972 218016
rect 398564 218068 398616 218074
rect 398564 218010 398616 218016
rect 397932 217002 397960 218010
rect 398760 217002 398788 228210
rect 399576 218068 399628 218074
rect 399576 218010 399628 218016
rect 399588 217002 399616 218010
rect 391768 216974 391828 217002
rect 392656 216974 392992 217002
rect 393484 216974 393820 217002
rect 394312 216974 394372 217002
rect 395140 216974 395568 217002
rect 395968 216974 396028 217002
rect 396796 216974 397132 217002
rect 397624 216974 397960 217002
rect 398452 216974 398788 217002
rect 399280 216974 399616 217002
rect 399864 217002 399892 229706
rect 400048 228546 400076 231676
rect 400036 228540 400088 228546
rect 400036 228482 400088 228488
rect 400036 228404 400088 228410
rect 400036 228346 400088 228352
rect 400048 218074 400076 228346
rect 400692 227186 400720 231676
rect 401336 227934 401364 231676
rect 401704 231662 401994 231690
rect 401324 227928 401376 227934
rect 401324 227870 401376 227876
rect 400864 227792 400916 227798
rect 400864 227734 400916 227740
rect 400680 227180 400732 227186
rect 400680 227122 400732 227128
rect 400876 218618 400904 227734
rect 401324 227180 401376 227186
rect 401324 227122 401376 227128
rect 400864 218612 400916 218618
rect 400864 218554 400916 218560
rect 400036 218068 400088 218074
rect 400036 218010 400088 218016
rect 401336 217002 401364 227122
rect 401704 221474 401732 231662
rect 402244 227928 402296 227934
rect 402244 227870 402296 227876
rect 401692 221468 401744 221474
rect 401692 221410 401744 221416
rect 402060 218884 402112 218890
rect 402060 218826 402112 218832
rect 402072 217002 402100 218826
rect 402256 218210 402284 227870
rect 402624 227798 402652 231676
rect 403268 227798 403296 231676
rect 403544 231662 403926 231690
rect 402612 227792 402664 227798
rect 402612 227734 402664 227740
rect 403256 227792 403308 227798
rect 403256 227734 403308 227740
rect 403544 225622 403572 231662
rect 403992 228676 404044 228682
rect 403992 228618 404044 228624
rect 403532 225616 403584 225622
rect 403532 225558 403584 225564
rect 402704 218748 402756 218754
rect 402704 218690 402756 218696
rect 402244 218204 402296 218210
rect 402244 218146 402296 218152
rect 402716 217002 402744 218690
rect 403716 218068 403768 218074
rect 403716 218010 403768 218016
rect 403728 217002 403756 218010
rect 399864 216974 400108 217002
rect 400936 216974 401364 217002
rect 401764 216974 402100 217002
rect 402592 216974 402744 217002
rect 403420 216974 403756 217002
rect 404004 217002 404032 228618
rect 404176 225004 404228 225010
rect 404176 224946 404228 224952
rect 404188 218074 404216 224946
rect 404556 224534 404584 231676
rect 404740 231662 405214 231690
rect 404544 224528 404596 224534
rect 404544 224470 404596 224476
rect 404740 220114 404768 231662
rect 405464 224256 405516 224262
rect 405464 224198 405516 224204
rect 404728 220108 404780 220114
rect 404728 220050 404780 220056
rect 404176 218068 404228 218074
rect 404176 218010 404228 218016
rect 405476 217002 405504 224198
rect 405844 222902 405872 231676
rect 406488 227050 406516 231676
rect 407146 231662 407344 231690
rect 406476 227044 406528 227050
rect 406476 226986 406528 226992
rect 407028 223304 407080 223310
rect 407028 223246 407080 223252
rect 405832 222896 405884 222902
rect 405832 222838 405884 222844
rect 406200 219564 406252 219570
rect 406200 219506 406252 219512
rect 406212 217002 406240 219506
rect 407040 217002 407068 223246
rect 407316 221610 407344 231662
rect 407776 228546 407804 231676
rect 407764 228540 407816 228546
rect 407764 228482 407816 228488
rect 408420 227186 408448 231676
rect 409064 228274 409092 231676
rect 409708 229770 409736 231676
rect 409696 229764 409748 229770
rect 409696 229706 409748 229712
rect 409604 228404 409656 228410
rect 409604 228346 409656 228352
rect 409052 228268 409104 228274
rect 409052 228210 409104 228216
rect 409144 227792 409196 227798
rect 409144 227734 409196 227740
rect 408408 227180 408460 227186
rect 408408 227122 408460 227128
rect 407764 226364 407816 226370
rect 407764 226306 407816 226312
rect 407304 221604 407356 221610
rect 407304 221546 407356 221552
rect 407580 219020 407632 219026
rect 407580 218962 407632 218968
rect 407592 217002 407620 218962
rect 407776 218890 407804 226306
rect 408408 221468 408460 221474
rect 408408 221410 408460 221416
rect 407764 218884 407816 218890
rect 407764 218826 407816 218832
rect 408420 217002 408448 221410
rect 409156 218754 409184 227734
rect 409144 218748 409196 218754
rect 409144 218690 409196 218696
rect 409616 217002 409644 228346
rect 410352 227798 410380 231676
rect 410800 229900 410852 229906
rect 410800 229842 410852 229848
rect 410812 229094 410840 229842
rect 410996 229094 411024 231676
rect 410812 229066 410932 229094
rect 410996 229066 411116 229094
rect 410340 227792 410392 227798
rect 410340 227734 410392 227740
rect 410904 218074 410932 229066
rect 411088 228682 411116 229066
rect 411076 228676 411128 228682
rect 411076 228618 411128 228624
rect 411076 228540 411128 228546
rect 411076 228482 411128 228488
rect 410340 218068 410392 218074
rect 410340 218010 410392 218016
rect 410892 218068 410944 218074
rect 410892 218010 410944 218016
rect 410352 217002 410380 218010
rect 411088 217002 411116 228482
rect 411640 226370 411668 231676
rect 411904 227792 411956 227798
rect 411904 227734 411956 227740
rect 411628 226364 411680 226370
rect 411628 226306 411680 226312
rect 411916 219026 411944 227734
rect 412284 225010 412312 231676
rect 412744 231662 412942 231690
rect 412548 227044 412600 227050
rect 412548 226986 412600 226992
rect 412272 225004 412324 225010
rect 412272 224946 412324 224952
rect 411904 219020 411956 219026
rect 411904 218962 411956 218968
rect 412560 218890 412588 226986
rect 412744 219570 412772 231662
rect 413572 227798 413600 231676
rect 413836 230240 413888 230246
rect 413836 230182 413888 230188
rect 413560 227792 413612 227798
rect 413560 227734 413612 227740
rect 412732 219564 412784 219570
rect 412732 219506 412784 219512
rect 413848 219434 413876 230182
rect 414216 224262 414244 231676
rect 414204 224256 414256 224262
rect 414204 224198 414256 224204
rect 414860 223310 414888 231676
rect 415504 228410 415532 231676
rect 416148 228546 416176 231676
rect 416792 229094 416820 231676
rect 417436 229906 417464 231676
rect 417712 231662 418094 231690
rect 418356 231662 418738 231690
rect 417424 229900 417476 229906
rect 417424 229842 417476 229848
rect 417712 229094 417740 231662
rect 416792 229066 416912 229094
rect 416136 228540 416188 228546
rect 416136 228482 416188 228488
rect 415492 228404 415544 228410
rect 415492 228346 415544 228352
rect 416688 227792 416740 227798
rect 416688 227734 416740 227740
rect 415308 223712 415360 223718
rect 415308 223654 415360 223660
rect 414848 223304 414900 223310
rect 414848 223246 414900 223252
rect 414480 220040 414532 220046
rect 414480 219982 414532 219988
rect 413756 219406 413876 219434
rect 411996 218884 412048 218890
rect 411996 218826 412048 218832
rect 412548 218884 412600 218890
rect 412548 218826 412600 218832
rect 412008 217002 412036 218826
rect 412548 218748 412600 218754
rect 412548 218690 412600 218696
rect 412560 217002 412588 218690
rect 413756 217002 413784 219406
rect 414492 217002 414520 219982
rect 415320 217002 415348 223654
rect 416504 222420 416556 222426
rect 416504 222362 416556 222368
rect 416136 218068 416188 218074
rect 416136 218010 416188 218016
rect 416148 217002 416176 218010
rect 404004 216974 404248 217002
rect 405076 216974 405504 217002
rect 405904 216974 406240 217002
rect 406732 216974 407068 217002
rect 407560 216974 407620 217002
rect 408388 216974 408448 217002
rect 409216 216974 409644 217002
rect 410044 216974 410380 217002
rect 410872 216974 411116 217002
rect 411700 216974 412036 217002
rect 412528 216974 412588 217002
rect 413356 216974 413784 217002
rect 414184 216974 414520 217002
rect 415012 216974 415348 217002
rect 415840 216974 416176 217002
rect 416516 217002 416544 222362
rect 416700 218074 416728 227734
rect 416884 221474 416912 229066
rect 417160 229066 417740 229094
rect 416872 221468 416924 221474
rect 416872 221410 416924 221416
rect 417160 218754 417188 229066
rect 418356 220046 418384 231662
rect 419368 227050 419396 231676
rect 420012 230246 420040 231676
rect 420000 230240 420052 230246
rect 420000 230182 420052 230188
rect 419632 229152 419684 229158
rect 419632 229094 419684 229100
rect 419356 227044 419408 227050
rect 419356 226986 419408 226992
rect 419448 226908 419500 226914
rect 419448 226850 419500 226856
rect 418344 220040 418396 220046
rect 418344 219982 418396 219988
rect 417792 219428 417844 219434
rect 417792 219370 417844 219376
rect 417148 218748 417200 218754
rect 417148 218690 417200 218696
rect 416688 218068 416740 218074
rect 416688 218010 416740 218016
rect 417804 217002 417832 219370
rect 419264 219156 419316 219162
rect 419264 219098 419316 219104
rect 418620 218068 418672 218074
rect 418620 218010 418672 218016
rect 418632 217002 418660 218010
rect 419276 217002 419304 219098
rect 419460 218074 419488 226850
rect 419644 223718 419672 229094
rect 420656 227798 420684 231676
rect 421024 231662 421314 231690
rect 420644 227792 420696 227798
rect 420644 227734 420696 227740
rect 420828 224256 420880 224262
rect 420828 224198 420880 224204
rect 419632 223712 419684 223718
rect 419632 223654 419684 223660
rect 420644 220856 420696 220862
rect 420644 220798 420696 220804
rect 419448 218068 419500 218074
rect 419448 218010 419500 218016
rect 420276 218068 420328 218074
rect 420276 218010 420328 218016
rect 420288 217002 420316 218010
rect 416516 216974 416668 217002
rect 417496 216974 417832 217002
rect 418324 216974 418660 217002
rect 419152 216974 419304 217002
rect 419980 216974 420316 217002
rect 420656 217002 420684 220798
rect 420840 218074 420868 224198
rect 421024 219502 421052 231662
rect 421944 229158 421972 231676
rect 422312 231662 422602 231690
rect 422864 231662 423246 231690
rect 421932 229152 421984 229158
rect 421932 229094 421984 229100
rect 422312 229094 422340 231662
rect 422220 229066 422340 229094
rect 422220 222426 422248 229066
rect 422208 222420 422260 222426
rect 422208 222362 422260 222368
rect 421932 220108 421984 220114
rect 421932 220050 421984 220056
rect 421012 219496 421064 219502
rect 421012 219438 421064 219444
rect 420828 218068 420880 218074
rect 420828 218010 420880 218016
rect 421944 217002 421972 220050
rect 422864 219434 422892 231662
rect 423496 229152 423548 229158
rect 423496 229094 423548 229100
rect 422680 219406 422892 219434
rect 422680 219162 422708 219406
rect 422668 219156 422720 219162
rect 422668 219098 422720 219104
rect 422760 218068 422812 218074
rect 422760 218010 422812 218016
rect 422772 217002 422800 218010
rect 423508 217002 423536 229094
rect 423876 220862 423904 231676
rect 424520 226914 424548 231676
rect 424508 226908 424560 226914
rect 424508 226850 424560 226856
rect 425164 224262 425192 231676
rect 425440 231662 425822 231690
rect 425152 224256 425204 224262
rect 425152 224198 425204 224204
rect 424968 222148 425020 222154
rect 424968 222090 425020 222096
rect 423864 220856 423916 220862
rect 423864 220798 423916 220804
rect 424416 218204 424468 218210
rect 424416 218146 424468 218152
rect 424428 217002 424456 218146
rect 424980 217002 425008 222090
rect 425440 218074 425468 231662
rect 426452 224942 426480 231676
rect 426820 231662 427110 231690
rect 426440 224936 426492 224942
rect 426440 224878 426492 224884
rect 426820 220114 426848 231662
rect 427740 229158 427768 231676
rect 427728 229152 427780 229158
rect 427728 229094 427780 229100
rect 428384 229094 428412 231676
rect 428752 231662 429042 231690
rect 429304 231662 429686 231690
rect 429948 231662 430330 231690
rect 430684 231662 430974 231690
rect 431236 231662 431618 231690
rect 432064 231662 432262 231690
rect 432708 231662 432906 231690
rect 433550 231662 433748 231690
rect 428384 229066 428504 229094
rect 426992 224936 427044 224942
rect 426992 224878 427044 224884
rect 426808 220108 426860 220114
rect 426808 220050 426860 220056
rect 426808 218340 426860 218346
rect 426808 218282 426860 218288
rect 425428 218068 425480 218074
rect 425428 218010 425480 218016
rect 426072 218068 426124 218074
rect 426072 218010 426124 218016
rect 426084 217002 426112 218010
rect 426820 217002 426848 218282
rect 427004 218210 427032 224878
rect 427820 224256 427872 224262
rect 427820 224198 427872 224204
rect 427832 219434 427860 224198
rect 427740 219406 427860 219434
rect 428280 219428 428332 219434
rect 426992 218204 427044 218210
rect 426992 218146 427044 218152
rect 427740 217002 427768 219406
rect 428280 219370 428332 219376
rect 428292 217002 428320 219370
rect 428476 218074 428504 229066
rect 428752 224262 428780 231662
rect 428740 224256 428792 224262
rect 428740 224198 428792 224204
rect 429304 222154 429332 231662
rect 429292 222148 429344 222154
rect 429292 222090 429344 222096
rect 429948 219434 429976 231662
rect 429580 219406 429976 219434
rect 430212 219428 430264 219434
rect 429580 218346 429608 219406
rect 430212 219370 430264 219376
rect 429568 218340 429620 218346
rect 429568 218282 429620 218288
rect 428464 218068 428516 218074
rect 428464 218010 428516 218016
rect 429108 218068 429160 218074
rect 429108 218010 429160 218016
rect 429120 217002 429148 218010
rect 430224 217002 430252 219370
rect 430684 218074 430712 231662
rect 431236 219434 431264 231662
rect 432064 219570 432092 231662
rect 432236 220516 432288 220522
rect 432236 220458 432288 220464
rect 432052 219564 432104 219570
rect 432052 219506 432104 219512
rect 432248 219434 432276 220458
rect 432708 219434 432736 231662
rect 433524 229832 433576 229838
rect 433524 229774 433576 229780
rect 433536 229094 433564 229774
rect 433720 229094 433748 231662
rect 434180 229838 434208 231676
rect 434168 229832 434220 229838
rect 434168 229774 434220 229780
rect 433536 229066 433656 229094
rect 433720 229066 433840 229094
rect 430960 219406 431264 219434
rect 431972 219406 432276 219434
rect 432696 219428 432748 219434
rect 430672 218068 430724 218074
rect 430672 218010 430724 218016
rect 430960 217002 430988 219406
rect 431972 218090 432000 219406
rect 432696 219370 432748 219376
rect 433248 218204 433300 218210
rect 433248 218146 433300 218152
rect 431880 218062 432000 218090
rect 432696 218068 432748 218074
rect 431880 217002 431908 218062
rect 432696 218010 432748 218016
rect 432708 217002 432736 218010
rect 433260 217002 433288 218146
rect 420656 216974 420808 217002
rect 421636 216974 421972 217002
rect 422464 216974 422800 217002
rect 423292 216974 423536 217002
rect 424120 216974 424456 217002
rect 424948 216974 425008 217002
rect 425776 216974 426112 217002
rect 426604 216974 426848 217002
rect 427432 216974 427768 217002
rect 428260 216974 428320 217002
rect 429088 216974 429148 217002
rect 429916 216974 430252 217002
rect 430744 216974 430988 217002
rect 431572 216974 431908 217002
rect 432400 216974 432736 217002
rect 433228 216974 433288 217002
rect 433628 217002 433656 229066
rect 433812 218074 433840 229066
rect 434824 220522 434852 231676
rect 435284 231662 435482 231690
rect 436126 231662 436416 231690
rect 434812 220516 434864 220522
rect 434812 220458 434864 220464
rect 435284 218210 435312 231662
rect 436388 224398 436416 231662
rect 436572 231662 436770 231690
rect 437032 231662 437414 231690
rect 437768 231662 438058 231690
rect 436572 229094 436600 231662
rect 436572 229066 436692 229094
rect 436376 224392 436428 224398
rect 436376 224334 436428 224340
rect 436284 224256 436336 224262
rect 436284 224198 436336 224204
rect 435272 218204 435324 218210
rect 435272 218146 435324 218152
rect 436008 218204 436060 218210
rect 436008 218146 436060 218152
rect 433800 218068 433852 218074
rect 433800 218010 433852 218016
rect 434996 218068 435048 218074
rect 434996 218010 435048 218016
rect 435008 217002 435036 218010
rect 436020 217002 436048 218146
rect 436296 218074 436324 224198
rect 436284 218068 436336 218074
rect 436284 218010 436336 218016
rect 436468 218068 436520 218074
rect 436468 218010 436520 218016
rect 433628 216974 434056 217002
rect 434884 216974 435036 217002
rect 435712 216974 436048 217002
rect 436480 217002 436508 218010
rect 436664 217138 436692 229066
rect 436836 224392 436888 224398
rect 436836 224334 436888 224340
rect 436848 218210 436876 224334
rect 437032 224262 437060 231662
rect 437020 224256 437072 224262
rect 437020 224198 437072 224204
rect 437768 219434 437796 231662
rect 438688 229838 438716 231676
rect 439332 230382 439360 231676
rect 439608 231662 439990 231690
rect 439320 230376 439372 230382
rect 439320 230318 439372 230324
rect 438676 229832 438728 229838
rect 438676 229774 438728 229780
rect 439320 229832 439372 229838
rect 439320 229774 439372 229780
rect 438952 224256 439004 224262
rect 438952 224198 439004 224204
rect 437492 219406 437796 219434
rect 436836 218204 436888 218210
rect 436836 218146 436888 218152
rect 437492 218074 437520 219406
rect 438964 218074 438992 224198
rect 437480 218068 437532 218074
rect 437480 218010 437532 218016
rect 438492 218068 438544 218074
rect 438492 218010 438544 218016
rect 438952 218068 439004 218074
rect 438952 218010 439004 218016
rect 436664 217110 436968 217138
rect 436940 217002 436968 217110
rect 438504 217002 438532 218010
rect 439332 217002 439360 229774
rect 439608 224262 439636 231662
rect 440332 230376 440384 230382
rect 440332 230318 440384 230324
rect 439596 224256 439648 224262
rect 439596 224198 439648 224204
rect 440148 218068 440200 218074
rect 440148 218010 440200 218016
rect 440160 217002 440188 218010
rect 436480 216974 436540 217002
rect 436940 216974 437368 217002
rect 438196 216974 438532 217002
rect 439024 216974 439360 217002
rect 439852 216974 440188 217002
rect 440344 217002 440372 230318
rect 440620 229094 440648 231676
rect 441264 229158 441292 231676
rect 441908 230450 441936 231676
rect 442092 231662 442566 231690
rect 443210 231662 443408 231690
rect 441896 230444 441948 230450
rect 441896 230386 441948 230392
rect 442092 230330 442120 231662
rect 441724 230302 442120 230330
rect 441252 229152 441304 229158
rect 441252 229094 441304 229100
rect 440620 229066 440740 229094
rect 440712 218074 440740 229066
rect 441724 219434 441752 230302
rect 442080 229152 442132 229158
rect 442080 229094 442132 229100
rect 441632 219406 441752 219434
rect 441632 218090 441660 219406
rect 440700 218068 440752 218074
rect 440700 218010 440752 218016
rect 441540 218062 441660 218090
rect 441540 217002 441568 218062
rect 440344 216974 440680 217002
rect 441508 216974 441568 217002
rect 442092 217002 442120 229094
rect 443380 217002 443408 231662
rect 443552 230444 443604 230450
rect 443552 230386 443604 230392
rect 442092 216974 442336 217002
rect 443164 216974 443408 217002
rect 443564 217002 443592 230386
rect 443840 230246 443868 231676
rect 444484 230450 444512 231676
rect 444668 231662 445142 231690
rect 444472 230444 444524 230450
rect 444472 230386 444524 230392
rect 444668 230330 444696 231662
rect 444484 230302 444696 230330
rect 443828 230240 443880 230246
rect 443828 230182 443880 230188
rect 444484 217002 444512 230302
rect 444656 230240 444708 230246
rect 444656 230182 444708 230188
rect 444668 229094 444696 230182
rect 445772 229094 445800 231676
rect 446416 229158 446444 231676
rect 446404 229152 446456 229158
rect 446404 229094 446456 229100
rect 444668 229066 445248 229094
rect 445772 229066 446076 229094
rect 445220 217002 445248 229066
rect 446048 217002 446076 229066
rect 447060 228818 447088 231676
rect 447244 231662 447718 231690
rect 447048 228812 447100 228818
rect 447048 228754 447100 228760
rect 447244 219434 447272 231662
rect 447600 230444 447652 230450
rect 447600 230386 447652 230392
rect 447152 219406 447272 219434
rect 447152 217870 447180 219406
rect 447140 217864 447192 217870
rect 447140 217806 447192 217812
rect 447612 217002 447640 230386
rect 448348 230330 448376 231676
rect 448348 230302 448744 230330
rect 448716 229094 448744 230302
rect 448992 229430 449020 231676
rect 449636 230382 449664 231676
rect 449624 230376 449676 230382
rect 449624 230318 449676 230324
rect 448980 229424 449032 229430
rect 448980 229366 449032 229372
rect 450280 229294 450308 231676
rect 450544 230376 450596 230382
rect 450544 230318 450596 230324
rect 450268 229288 450320 229294
rect 450268 229230 450320 229236
rect 448716 229066 449388 229094
rect 448520 229016 448572 229022
rect 448520 228958 448572 228964
rect 447784 217864 447836 217870
rect 447784 217806 447836 217812
rect 443564 216974 443992 217002
rect 444484 216974 444820 217002
rect 445220 216974 445648 217002
rect 446048 216974 446476 217002
rect 447304 216974 447640 217002
rect 447796 217002 447824 217806
rect 448532 217002 448560 228958
rect 449360 217002 449388 229066
rect 450176 228812 450228 228818
rect 450176 228754 450228 228760
rect 450188 217002 450216 228754
rect 450556 218414 450584 230318
rect 450924 229158 450952 231676
rect 451568 230382 451596 231676
rect 452226 231662 452608 231690
rect 451556 230376 451608 230382
rect 451556 230318 451608 230324
rect 451372 229424 451424 229430
rect 451372 229366 451424 229372
rect 450912 229152 450964 229158
rect 450912 229094 450964 229100
rect 451384 224262 451412 229366
rect 451832 229288 451884 229294
rect 451832 229230 451884 229236
rect 451372 224256 451424 224262
rect 451372 224198 451424 224204
rect 450544 218408 450596 218414
rect 450544 218350 450596 218356
rect 451844 217002 451872 229230
rect 452016 224256 452068 224262
rect 452016 224198 452068 224204
rect 452028 219434 452056 224198
rect 452580 221474 452608 231662
rect 452856 230246 452884 231676
rect 453304 230376 453356 230382
rect 453304 230318 453356 230324
rect 452844 230240 452896 230246
rect 452844 230182 452896 230188
rect 452752 229152 452804 229158
rect 452752 229094 452804 229100
rect 452568 221468 452620 221474
rect 452568 221410 452620 221416
rect 447796 216974 448132 217002
rect 448532 216974 448960 217002
rect 449360 216974 449788 217002
rect 450188 216974 450616 217002
rect 451444 216974 451872 217002
rect 451936 219406 452056 219434
rect 451936 217002 451964 219406
rect 452764 217002 452792 229094
rect 453316 218074 453344 230318
rect 453500 229974 453528 231676
rect 454144 230110 454172 231676
rect 454316 230240 454368 230246
rect 454316 230182 454368 230188
rect 454132 230104 454184 230110
rect 454132 230046 454184 230052
rect 453488 229968 453540 229974
rect 453488 229910 453540 229916
rect 453580 218408 453632 218414
rect 453580 218350 453632 218356
rect 453304 218068 453356 218074
rect 453304 218010 453356 218016
rect 453592 217002 453620 218350
rect 454328 217002 454356 230182
rect 454788 223582 454816 231676
rect 455432 230382 455460 231676
rect 455420 230376 455472 230382
rect 455420 230318 455472 230324
rect 455328 230104 455380 230110
rect 455328 230046 455380 230052
rect 454776 223576 454828 223582
rect 454776 223518 454828 223524
rect 455340 220794 455368 230046
rect 455788 229968 455840 229974
rect 455788 229910 455840 229916
rect 455800 229094 455828 229910
rect 456076 229094 456104 231676
rect 455800 229066 456012 229094
rect 456076 229066 456196 229094
rect 455328 220788 455380 220794
rect 455328 220730 455380 220736
rect 455420 218068 455472 218074
rect 455420 218010 455472 218016
rect 455432 217002 455460 218010
rect 455984 217002 456012 229066
rect 456168 224262 456196 229066
rect 456156 224256 456208 224262
rect 456156 224198 456208 224204
rect 456720 221610 456748 231676
rect 457168 230376 457220 230382
rect 457168 230318 457220 230324
rect 457180 229094 457208 230318
rect 457364 230042 457392 231676
rect 457352 230036 457404 230042
rect 457352 229978 457404 229984
rect 457180 229066 457668 229094
rect 456708 221604 456760 221610
rect 456708 221546 456760 221552
rect 456708 221468 456760 221474
rect 456708 221410 456760 221416
rect 456720 219434 456748 221410
rect 456720 219406 456840 219434
rect 456812 217002 456840 219406
rect 457640 217002 457668 229066
rect 458008 219298 458036 231676
rect 458652 225826 458680 231676
rect 459310 231662 459508 231690
rect 458640 225820 458692 225826
rect 458640 225762 458692 225768
rect 458548 220788 458600 220794
rect 458548 220730 458600 220736
rect 457996 219292 458048 219298
rect 457996 219234 458048 219240
rect 458560 217002 458588 220730
rect 459480 220250 459508 231662
rect 459744 224256 459796 224262
rect 459744 224198 459796 224204
rect 459468 220244 459520 220250
rect 459468 220186 459520 220192
rect 459756 217002 459784 224198
rect 459940 222902 459968 231676
rect 460584 223718 460612 231676
rect 461242 231662 461624 231690
rect 461886 231662 462176 231690
rect 461596 229094 461624 231662
rect 461596 229066 461992 229094
rect 460572 223712 460624 223718
rect 460572 223654 460624 223660
rect 460112 223576 460164 223582
rect 460112 223518 460164 223524
rect 459928 222896 459980 222902
rect 459928 222838 459980 222844
rect 451936 216974 452272 217002
rect 452764 216974 453100 217002
rect 453592 216974 453928 217002
rect 454328 216974 454756 217002
rect 455432 216974 455584 217002
rect 455984 216974 456412 217002
rect 456812 216974 457240 217002
rect 457640 216974 458068 217002
rect 458560 216974 458896 217002
rect 459724 216974 459784 217002
rect 460124 217002 460152 223518
rect 461768 221604 461820 221610
rect 461768 221546 461820 221552
rect 461124 219292 461176 219298
rect 461124 219234 461176 219240
rect 461136 217002 461164 219234
rect 461780 217002 461808 221546
rect 461964 218210 461992 229066
rect 462148 222154 462176 231662
rect 462516 229094 462544 231676
rect 462424 229066 462544 229094
rect 462424 224262 462452 229066
rect 462596 225820 462648 225826
rect 462596 225762 462648 225768
rect 462412 224256 462464 224262
rect 462412 224198 462464 224204
rect 462136 222148 462188 222154
rect 462136 222090 462188 222096
rect 461952 218204 462004 218210
rect 461952 218146 462004 218152
rect 462608 217002 462636 225762
rect 463160 225282 463188 231676
rect 463804 230382 463832 231676
rect 464462 231662 465028 231690
rect 465106 231662 465488 231690
rect 465750 231662 466040 231690
rect 463792 230376 463844 230382
rect 463792 230318 463844 230324
rect 464068 230036 464120 230042
rect 464068 229978 464120 229984
rect 463148 225276 463200 225282
rect 463148 225218 463200 225224
rect 462964 223712 463016 223718
rect 462964 223654 463016 223660
rect 462976 218074 463004 223654
rect 462964 218068 463016 218074
rect 462964 218010 463016 218016
rect 464080 217002 464108 229978
rect 465000 219638 465028 231662
rect 465460 230246 465488 231662
rect 465724 230376 465776 230382
rect 465724 230318 465776 230324
rect 465448 230240 465500 230246
rect 465448 230182 465500 230188
rect 465736 220794 465764 230318
rect 466012 228886 466040 231662
rect 466000 228880 466052 228886
rect 466000 228822 466052 228828
rect 466380 224874 466408 231676
rect 467038 231662 467328 231690
rect 467104 225276 467156 225282
rect 467104 225218 467156 225224
rect 466368 224868 466420 224874
rect 466368 224810 466420 224816
rect 466736 222896 466788 222902
rect 466736 222838 466788 222844
rect 465724 220788 465776 220794
rect 465724 220730 465776 220736
rect 465172 220244 465224 220250
rect 465172 220186 465224 220192
rect 464988 219632 465040 219638
rect 464988 219574 465040 219580
rect 464344 218068 464396 218074
rect 464344 218010 464396 218016
rect 460124 216974 460552 217002
rect 461136 216974 461380 217002
rect 461780 216974 462208 217002
rect 462608 216974 463036 217002
rect 463864 216974 464108 217002
rect 464356 217002 464384 218010
rect 465184 217002 465212 220186
rect 466000 218204 466052 218210
rect 466000 218146 466052 218152
rect 466012 217002 466040 218146
rect 466748 217002 466776 222838
rect 467116 218074 467144 225218
rect 467300 222902 467328 231662
rect 467668 227322 467696 231676
rect 468326 231662 468800 231690
rect 468970 231662 469168 231690
rect 467656 227316 467708 227322
rect 467656 227258 467708 227264
rect 467288 222896 467340 222902
rect 467288 222838 467340 222844
rect 468484 222148 468536 222154
rect 468484 222090 468536 222096
rect 467104 218068 467156 218074
rect 467104 218010 467156 218016
rect 467840 218068 467892 218074
rect 467840 218010 467892 218016
rect 467852 217002 467880 218010
rect 468496 217002 468524 222090
rect 468772 221610 468800 231662
rect 468760 221604 468812 221610
rect 468760 221546 468812 221552
rect 469140 220386 469168 231662
rect 469404 230240 469456 230246
rect 469404 230182 469456 230188
rect 469416 225622 469444 230182
rect 469600 229770 469628 231676
rect 469588 229764 469640 229770
rect 469588 229706 469640 229712
rect 469864 228880 469916 228886
rect 469864 228822 469916 228828
rect 469404 225616 469456 225622
rect 469404 225558 469456 225564
rect 469680 224256 469732 224262
rect 469680 224198 469732 224204
rect 469312 220788 469364 220794
rect 469312 220730 469364 220736
rect 469128 220380 469180 220386
rect 469128 220322 469180 220328
rect 469324 217002 469352 220730
rect 469692 217138 469720 224198
rect 469876 218550 469904 228822
rect 470244 228410 470272 231676
rect 470232 228404 470284 228410
rect 470232 228346 470284 228352
rect 470888 224262 470916 231676
rect 471546 231662 471928 231690
rect 471244 224868 471296 224874
rect 471244 224810 471296 224816
rect 470876 224256 470928 224262
rect 470876 224198 470928 224204
rect 469864 218544 469916 218550
rect 469864 218486 469916 218492
rect 470968 218544 471020 218550
rect 470968 218486 471020 218492
rect 469692 217110 470088 217138
rect 470060 217002 470088 217110
rect 470980 217002 471008 218486
rect 471256 218074 471284 224810
rect 471900 222154 471928 231662
rect 472176 225758 472204 231676
rect 472834 231662 473308 231690
rect 473478 231662 473768 231690
rect 472164 225752 472216 225758
rect 472164 225694 472216 225700
rect 471888 222148 471940 222154
rect 471888 222090 471940 222096
rect 473280 220250 473308 231662
rect 473544 225616 473596 225622
rect 473544 225558 473596 225564
rect 473268 220244 473320 220250
rect 473268 220186 473320 220192
rect 471980 219632 472032 219638
rect 471980 219574 472032 219580
rect 471244 218068 471296 218074
rect 471244 218010 471296 218016
rect 471992 217002 472020 219574
rect 472624 218068 472676 218074
rect 472624 218010 472676 218016
rect 472636 217002 472664 218010
rect 473556 217002 473584 225558
rect 473740 223582 473768 231662
rect 474108 227186 474136 231676
rect 474752 227798 474780 231676
rect 475410 231662 475976 231690
rect 474740 227792 474792 227798
rect 474740 227734 474792 227740
rect 474096 227180 474148 227186
rect 474096 227122 474148 227128
rect 473728 223576 473780 223582
rect 473728 223518 473780 223524
rect 475016 222896 475068 222902
rect 475016 222838 475068 222844
rect 474280 221604 474332 221610
rect 474280 221546 474332 221552
rect 474292 217002 474320 221546
rect 475028 217002 475056 222838
rect 475948 220114 475976 231662
rect 476040 230466 476068 231676
rect 476040 230450 476160 230466
rect 476040 230444 476172 230450
rect 476040 230438 476120 230444
rect 476120 230386 476172 230392
rect 476684 230042 476712 231676
rect 476672 230036 476724 230042
rect 476672 229978 476724 229984
rect 476764 229764 476816 229770
rect 476764 229706 476816 229712
rect 476580 227316 476632 227322
rect 476580 227258 476632 227264
rect 476120 220380 476172 220386
rect 476120 220322 476172 220328
rect 475936 220108 475988 220114
rect 475936 220050 475988 220056
rect 476132 217002 476160 220322
rect 476592 219434 476620 227258
rect 476776 220794 476804 229706
rect 477328 227050 477356 231676
rect 477972 230246 478000 231676
rect 478630 231662 478828 231690
rect 478604 230444 478656 230450
rect 478604 230386 478656 230392
rect 477960 230240 478012 230246
rect 477960 230182 478012 230188
rect 477316 227044 477368 227050
rect 477316 226986 477368 226992
rect 478616 225622 478644 230386
rect 478800 230330 478828 231662
rect 478800 230302 479012 230330
rect 478788 230240 478840 230246
rect 478788 230182 478840 230188
rect 478604 225616 478656 225622
rect 478604 225558 478656 225564
rect 477500 224256 477552 224262
rect 477500 224198 477552 224204
rect 476764 220788 476816 220794
rect 476764 220730 476816 220736
rect 476592 219406 476712 219434
rect 476684 217002 476712 219406
rect 477512 217002 477540 224198
rect 478800 221610 478828 230182
rect 478984 228546 479012 230302
rect 479260 229906 479288 231676
rect 479248 229900 479300 229906
rect 479248 229842 479300 229848
rect 478972 228540 479024 228546
rect 478972 228482 479024 228488
rect 479524 228404 479576 228410
rect 479524 228346 479576 228352
rect 479248 222148 479300 222154
rect 479248 222090 479300 222096
rect 478788 221604 478840 221610
rect 478788 221546 478840 221552
rect 478420 220788 478472 220794
rect 478420 220730 478472 220736
rect 478432 217002 478460 220730
rect 479260 217002 479288 222090
rect 479536 218346 479564 228346
rect 479904 223038 479932 231676
rect 480548 224398 480576 231676
rect 480720 230036 480772 230042
rect 480720 229978 480772 229984
rect 480732 226030 480760 229978
rect 481192 227322 481220 231676
rect 481836 230382 481864 231676
rect 482494 231662 482968 231690
rect 481824 230376 481876 230382
rect 481824 230318 481876 230324
rect 482744 227792 482796 227798
rect 482744 227734 482796 227740
rect 481180 227316 481232 227322
rect 481180 227258 481232 227264
rect 480720 226024 480772 226030
rect 480720 225966 480772 225972
rect 480812 225752 480864 225758
rect 480812 225694 480864 225700
rect 480536 224392 480588 224398
rect 480536 224334 480588 224340
rect 479892 223032 479944 223038
rect 479892 222974 479944 222980
rect 479524 218340 479576 218346
rect 479524 218282 479576 218288
rect 480352 218340 480404 218346
rect 480352 218282 480404 218288
rect 480364 217002 480392 218282
rect 480824 217002 480852 225694
rect 480996 223576 481048 223582
rect 480996 223518 481048 223524
rect 481008 218074 481036 223518
rect 482756 222329 482784 227734
rect 482742 222320 482798 222329
rect 482742 222255 482798 222264
rect 481732 220244 481784 220250
rect 481732 220186 481784 220192
rect 480996 218068 481048 218074
rect 480996 218010 481048 218016
rect 481744 217002 481772 220186
rect 482756 218074 482784 222255
rect 482940 220522 482968 231662
rect 483124 223174 483152 231676
rect 483782 231662 484348 231690
rect 484426 231662 484808 231690
rect 483112 223168 483164 223174
rect 483112 223110 483164 223116
rect 484320 221882 484348 231662
rect 484780 229770 484808 231662
rect 484768 229764 484820 229770
rect 484768 229706 484820 229712
rect 485056 228682 485084 231676
rect 485044 228676 485096 228682
rect 485044 228618 485096 228624
rect 484860 227180 484912 227186
rect 484860 227122 484912 227128
rect 484308 221876 484360 221882
rect 484308 221818 484360 221824
rect 484032 221468 484084 221474
rect 484032 221410 484084 221416
rect 482928 220516 482980 220522
rect 482928 220458 482980 220464
rect 482560 218068 482612 218074
rect 482560 218010 482612 218016
rect 482744 218068 482796 218074
rect 482744 218010 482796 218016
rect 482572 217002 482600 218010
rect 484044 217002 484072 221410
rect 484872 218754 484900 227122
rect 485700 220386 485728 231676
rect 485872 225616 485924 225622
rect 485872 225558 485924 225564
rect 485884 223689 485912 225558
rect 485870 223680 485926 223689
rect 485870 223615 485926 223624
rect 486344 222902 486372 231676
rect 486516 230376 486568 230382
rect 486516 230318 486568 230324
rect 486528 225894 486556 230318
rect 486988 228410 487016 231676
rect 487646 231662 488028 231690
rect 486976 228404 487028 228410
rect 486976 228346 487028 228352
rect 487804 226024 487856 226030
rect 487804 225966 487856 225972
rect 486516 225888 486568 225894
rect 486516 225830 486568 225836
rect 486606 223680 486662 223689
rect 486606 223615 486662 223624
rect 486332 222896 486384 222902
rect 486332 222838 486384 222844
rect 485688 220380 485740 220386
rect 485688 220322 485740 220328
rect 485872 220108 485924 220114
rect 485872 220050 485924 220056
rect 484860 218748 484912 218754
rect 484860 218690 484912 218696
rect 484872 217002 484900 218690
rect 485044 218068 485096 218074
rect 485044 218010 485096 218016
rect 464356 216974 464692 217002
rect 465184 216974 465520 217002
rect 466012 216974 466348 217002
rect 466748 216974 467176 217002
rect 467852 216974 468004 217002
rect 468496 216974 468832 217002
rect 469324 216974 469660 217002
rect 470060 216974 470488 217002
rect 470980 216974 471316 217002
rect 471992 216974 472144 217002
rect 472636 216974 472972 217002
rect 473556 216974 473800 217002
rect 474292 216974 474628 217002
rect 475028 216974 475456 217002
rect 476132 216974 476284 217002
rect 476684 216974 477112 217002
rect 477512 216974 477940 217002
rect 478432 216974 478768 217002
rect 479260 216974 479596 217002
rect 480364 216974 480424 217002
rect 480824 216974 481252 217002
rect 481744 216974 482080 217002
rect 482572 216974 482908 217002
rect 483736 216974 484072 217002
rect 484564 216974 484900 217002
rect 485056 217002 485084 218010
rect 485884 217002 485912 220050
rect 486620 217002 486648 223615
rect 487816 218113 487844 225966
rect 488000 225758 488028 231662
rect 488184 231662 488290 231690
rect 487988 225752 488040 225758
rect 487988 225694 488040 225700
rect 488184 220250 488212 231662
rect 488920 227186 488948 231676
rect 488908 227180 488960 227186
rect 488908 227122 488960 227128
rect 489000 227044 489052 227050
rect 489000 226986 489052 226992
rect 488172 220244 488224 220250
rect 488172 220186 488224 220192
rect 489012 219473 489040 226986
rect 489564 224262 489592 231676
rect 490208 229634 490236 231676
rect 490866 231662 491248 231690
rect 490564 229900 490616 229906
rect 490564 229842 490616 229848
rect 490196 229628 490248 229634
rect 490196 229570 490248 229576
rect 489552 224256 489604 224262
rect 489552 224198 489604 224204
rect 489184 221604 489236 221610
rect 489184 221546 489236 221552
rect 488998 219464 489054 219473
rect 488998 219399 489054 219408
rect 487802 218104 487858 218113
rect 487802 218039 487858 218048
rect 487816 217002 487844 218039
rect 489012 217002 489040 219399
rect 485056 216974 485392 217002
rect 485884 216974 486220 217002
rect 486620 216974 487048 217002
rect 487816 216974 487876 217002
rect 488704 216974 489040 217002
rect 489196 217002 489224 221546
rect 490576 218929 490604 229842
rect 491220 229094 491248 231662
rect 491220 229066 491340 229094
rect 490748 228540 490800 228546
rect 490748 228482 490800 228488
rect 490760 219201 490788 228482
rect 491312 225622 491340 229066
rect 491496 228546 491524 231676
rect 491680 231662 492154 231690
rect 492798 231662 493088 231690
rect 491484 228540 491536 228546
rect 491484 228482 491536 228488
rect 491300 225616 491352 225622
rect 491300 225558 491352 225564
rect 491680 220114 491708 231662
rect 492680 227316 492732 227322
rect 492680 227258 492732 227264
rect 491944 223032 491996 223038
rect 491944 222974 491996 222980
rect 491668 220108 491720 220114
rect 491668 220050 491720 220056
rect 490746 219192 490802 219201
rect 490746 219127 490802 219136
rect 490562 218920 490618 218929
rect 490562 218855 490618 218864
rect 490760 217002 490788 219127
rect 491206 218920 491262 218929
rect 491206 218855 491262 218864
rect 491220 217002 491248 218855
rect 491956 218657 491984 222974
rect 491942 218648 491998 218657
rect 491942 218583 491998 218592
rect 489196 216974 489532 217002
rect 490360 216974 490788 217002
rect 491188 216974 491248 217002
rect 491956 217002 491984 218583
rect 492692 218385 492720 227258
rect 493060 224670 493088 231662
rect 493428 229294 493456 231676
rect 494072 229906 494100 231676
rect 494348 231662 494730 231690
rect 494060 229900 494112 229906
rect 494060 229842 494112 229848
rect 493968 229628 494020 229634
rect 493968 229570 494020 229576
rect 493416 229288 493468 229294
rect 493416 229230 493468 229236
rect 493980 227458 494008 229570
rect 493968 227452 494020 227458
rect 493968 227394 494020 227400
rect 493048 224664 493100 224670
rect 493048 224606 493100 224612
rect 492864 224392 492916 224398
rect 492864 224334 492916 224340
rect 492678 218376 492734 218385
rect 492678 218311 492734 218320
rect 492876 217002 492904 224334
rect 494348 221746 494376 231662
rect 495360 227322 495388 231676
rect 495348 227316 495400 227322
rect 495348 227258 495400 227264
rect 496004 225894 496032 231676
rect 496188 231662 496662 231690
rect 494796 225888 494848 225894
rect 494796 225830 494848 225836
rect 495992 225888 496044 225894
rect 495992 225830 496044 225836
rect 494336 221740 494388 221746
rect 494336 221682 494388 221688
rect 494808 219201 494836 225830
rect 495808 223168 495860 223174
rect 495808 223110 495860 223116
rect 495348 220516 495400 220522
rect 495348 220458 495400 220464
rect 494794 219192 494850 219201
rect 494794 219127 494850 219136
rect 493874 217696 493930 217705
rect 493874 217631 493930 217640
rect 493888 217002 493916 217631
rect 494808 217002 494836 219127
rect 495360 218074 495388 220458
rect 495348 218068 495400 218074
rect 495348 218010 495400 218016
rect 495360 217002 495388 218010
rect 491956 216974 492016 217002
rect 492844 216974 492904 217002
rect 493672 216974 493916 217002
rect 494500 216974 494836 217002
rect 495328 216974 495388 217002
rect 495820 217002 495848 223110
rect 496188 221610 496216 231662
rect 496820 229764 496872 229770
rect 496820 229706 496872 229712
rect 496832 223961 496860 229706
rect 497292 224398 497320 231676
rect 497936 229158 497964 231676
rect 497924 229152 497976 229158
rect 497924 229094 497976 229100
rect 497280 224392 497332 224398
rect 497280 224334 497332 224340
rect 496818 223952 496874 223961
rect 496818 223887 496874 223896
rect 497830 223952 497886 223961
rect 497830 223887 497886 223896
rect 496912 221876 496964 221882
rect 496912 221818 496964 221824
rect 496176 221604 496228 221610
rect 496176 221546 496228 221552
rect 496924 219162 496952 221818
rect 496912 219156 496964 219162
rect 496912 219098 496964 219104
rect 496924 217002 496952 219098
rect 497844 217002 497872 223887
rect 498580 223446 498608 231676
rect 498844 228676 498896 228682
rect 498844 228618 498896 228624
rect 498568 223440 498620 223446
rect 498568 223382 498620 223388
rect 498856 217297 498884 228618
rect 499224 227050 499252 231676
rect 499868 230246 499896 231676
rect 499856 230240 499908 230246
rect 499856 230182 499908 230188
rect 500224 229288 500276 229294
rect 500224 229230 500276 229236
rect 499212 227044 499264 227050
rect 499212 226986 499264 226992
rect 499856 222896 499908 222902
rect 499856 222838 499908 222844
rect 499120 220380 499172 220386
rect 499120 220322 499172 220328
rect 498842 217288 498898 217297
rect 498842 217223 498898 217232
rect 498856 217002 498884 217223
rect 495820 216974 496156 217002
rect 496924 216974 496984 217002
rect 497812 216974 497872 217002
rect 498640 216974 498884 217002
rect 499132 217002 499160 220322
rect 499868 218958 499896 222838
rect 500236 220522 500264 229230
rect 500512 223038 500540 231676
rect 501156 226166 501184 231676
rect 501800 230042 501828 231676
rect 501788 230036 501840 230042
rect 501788 229978 501840 229984
rect 502444 228410 502472 231676
rect 503102 231662 503392 231690
rect 503364 229094 503392 231662
rect 503732 230382 503760 231676
rect 504390 231662 504680 231690
rect 503720 230376 503772 230382
rect 503720 230318 503772 230324
rect 504364 230240 504416 230246
rect 504364 230182 504416 230188
rect 503364 229066 503484 229094
rect 501328 228404 501380 228410
rect 501328 228346 501380 228352
rect 502432 228404 502484 228410
rect 502432 228346 502484 228352
rect 501144 226160 501196 226166
rect 501144 226102 501196 226108
rect 500500 223032 500552 223038
rect 500500 222974 500552 222980
rect 500224 220516 500276 220522
rect 500224 220458 500276 220464
rect 501340 219745 501368 228346
rect 503260 227180 503312 227186
rect 503260 227122 503312 227128
rect 501512 225752 501564 225758
rect 501512 225694 501564 225700
rect 501326 219736 501382 219745
rect 501326 219671 501382 219680
rect 500052 219286 500448 219314
rect 499856 218952 499908 218958
rect 499856 218894 499908 218900
rect 499868 217002 499896 218894
rect 500052 218657 500080 219286
rect 500420 219201 500448 219286
rect 500222 219192 500278 219201
rect 500222 219127 500278 219136
rect 500406 219192 500462 219201
rect 500406 219127 500462 219136
rect 500236 218657 500264 219127
rect 500038 218648 500094 218657
rect 500038 218583 500094 218592
rect 500222 218648 500278 218657
rect 500222 218583 500278 218592
rect 500224 218068 500276 218074
rect 500224 218010 500276 218016
rect 500236 217569 500264 218010
rect 500222 217560 500278 217569
rect 500222 217495 500278 217504
rect 501340 217002 501368 219671
rect 499132 216974 499468 217002
rect 499868 216974 500296 217002
rect 501124 216974 501368 217002
rect 501524 217002 501552 225694
rect 502432 220244 502484 220250
rect 502432 220186 502484 220192
rect 502444 218074 502472 220186
rect 502432 218068 502484 218074
rect 502432 218010 502484 218016
rect 502444 217002 502472 218010
rect 503272 217002 503300 227122
rect 503456 223310 503484 229066
rect 504088 224256 504140 224262
rect 504088 224198 504140 224204
rect 503444 223304 503496 223310
rect 503444 223246 503496 223252
rect 503718 217016 503774 217025
rect 501524 216974 501952 217002
rect 502444 216974 502780 217002
rect 503272 216974 503718 217002
rect 504100 217002 504128 224198
rect 504376 220386 504404 230182
rect 504652 224262 504680 231662
rect 505020 225758 505048 231676
rect 505664 230178 505692 231676
rect 505652 230172 505704 230178
rect 505652 230114 505704 230120
rect 506112 229900 506164 229906
rect 506112 229842 506164 229848
rect 505652 227452 505704 227458
rect 505652 227394 505704 227400
rect 505008 225752 505060 225758
rect 505008 225694 505060 225700
rect 504640 224256 504692 224262
rect 504640 224198 504692 224204
rect 504364 220380 504416 220386
rect 504364 220322 504416 220328
rect 504548 219360 504600 219366
rect 504548 219302 504600 219308
rect 504560 219201 504588 219302
rect 504546 219192 504602 219201
rect 504546 219127 504602 219136
rect 504730 219192 504786 219201
rect 504730 219127 504732 219136
rect 504784 219127 504786 219136
rect 504732 219098 504784 219104
rect 504730 218920 504786 218929
rect 504730 218855 504786 218864
rect 504744 218618 504772 218855
rect 504732 218612 504784 218618
rect 504732 218554 504784 218560
rect 505284 218612 505336 218618
rect 505284 218554 505336 218560
rect 505296 218385 505324 218554
rect 505282 218376 505338 218385
rect 505282 218311 505338 218320
rect 505664 218210 505692 227394
rect 505928 225616 505980 225622
rect 505928 225558 505980 225564
rect 505940 220017 505968 225558
rect 506124 225418 506152 229842
rect 506308 227186 506336 231676
rect 506480 228540 506532 228546
rect 506480 228482 506532 228488
rect 506296 227180 506348 227186
rect 506296 227122 506348 227128
rect 506112 225412 506164 225418
rect 506112 225354 506164 225360
rect 505926 220008 505982 220017
rect 505926 219943 505982 219952
rect 505652 218204 505704 218210
rect 505652 218146 505704 218152
rect 505664 217002 505692 218146
rect 504100 216974 504436 217002
rect 505264 216974 505692 217002
rect 505940 217002 505968 219943
rect 506294 219192 506350 219201
rect 506294 219127 506350 219136
rect 506308 218754 506336 219127
rect 506296 218748 506348 218754
rect 506296 218690 506348 218696
rect 506492 217002 506520 228482
rect 506952 224534 506980 231676
rect 507124 230376 507176 230382
rect 507124 230318 507176 230324
rect 506940 224528 506992 224534
rect 506940 224470 506992 224476
rect 507136 220250 507164 230318
rect 507596 229770 507624 231676
rect 507584 229764 507636 229770
rect 507584 229706 507636 229712
rect 508240 225622 508268 231676
rect 508228 225616 508280 225622
rect 508228 225558 508280 225564
rect 508596 224664 508648 224670
rect 508596 224606 508648 224612
rect 507766 220280 507822 220289
rect 507124 220244 507176 220250
rect 507766 220215 507822 220224
rect 507124 220186 507176 220192
rect 507780 220114 507808 220215
rect 507768 220108 507820 220114
rect 507768 220050 507820 220056
rect 507780 217002 507808 220050
rect 508608 217002 508636 224606
rect 508884 222902 508912 231676
rect 509528 229430 509556 231676
rect 509884 230036 509936 230042
rect 509884 229978 509936 229984
rect 509516 229424 509568 229430
rect 509516 229366 509568 229372
rect 508872 222896 508924 222902
rect 508872 222838 508924 222844
rect 509896 222154 509924 229978
rect 510172 228546 510200 231676
rect 510816 230382 510844 231676
rect 511474 231662 511856 231690
rect 511828 230518 511856 231662
rect 511816 230512 511868 230518
rect 511816 230454 511868 230460
rect 510804 230376 510856 230382
rect 510804 230318 510856 230324
rect 511816 230376 511868 230382
rect 511816 230318 511868 230324
rect 510160 228540 510212 228546
rect 510160 228482 510212 228488
rect 511448 227316 511500 227322
rect 511448 227258 511500 227264
rect 510344 225412 510396 225418
rect 510344 225354 510396 225360
rect 510356 224058 510384 225354
rect 510344 224052 510396 224058
rect 510344 223994 510396 224000
rect 509884 222148 509936 222154
rect 509884 222090 509936 222096
rect 509240 220516 509292 220522
rect 509240 220458 509292 220464
rect 508870 217832 508926 217841
rect 508870 217767 508926 217776
rect 508884 217025 508912 217767
rect 505940 216974 506092 217002
rect 506492 216974 506920 217002
rect 507748 216974 507808 217002
rect 508576 216974 508636 217002
rect 508870 217016 508926 217025
rect 503718 216951 503774 216960
rect 509252 217002 509280 220458
rect 510356 217002 510384 223994
rect 510712 221740 510764 221746
rect 510712 221682 510764 221688
rect 510724 220969 510752 221682
rect 510710 220960 510766 220969
rect 510710 220895 510766 220904
rect 509252 216974 509404 217002
rect 510232 216974 510384 217002
rect 510724 217002 510752 220895
rect 511460 217002 511488 227258
rect 511828 220114 511856 230318
rect 512104 227594 512132 231676
rect 512762 231662 513328 231690
rect 513406 231662 513696 231690
rect 512092 227588 512144 227594
rect 512092 227530 512144 227536
rect 512276 225888 512328 225894
rect 512276 225830 512328 225836
rect 512288 224233 512316 225830
rect 512274 224224 512330 224233
rect 512274 224159 512330 224168
rect 511816 220108 511868 220114
rect 511816 220050 511868 220056
rect 512288 217002 512316 224159
rect 513300 220522 513328 231662
rect 513668 229634 513696 231662
rect 513840 230172 513892 230178
rect 513840 230114 513892 230120
rect 513656 229628 513708 229634
rect 513656 229570 513708 229576
rect 513852 229094 513880 230114
rect 513760 229066 513880 229094
rect 513760 222018 513788 229066
rect 514036 228682 514064 231676
rect 514024 228676 514076 228682
rect 514024 228618 514076 228624
rect 514024 224392 514076 224398
rect 514024 224334 514076 224340
rect 513748 222012 513800 222018
rect 513748 221954 513800 221960
rect 513470 221776 513526 221785
rect 513470 221711 513526 221720
rect 513484 221610 513512 221711
rect 513472 221604 513524 221610
rect 513472 221546 513524 221552
rect 513288 220516 513340 220522
rect 513288 220458 513340 220464
rect 513484 217002 513512 221546
rect 514036 217002 514064 224334
rect 514680 223786 514708 231676
rect 515324 230178 515352 231676
rect 515312 230172 515364 230178
rect 515312 230114 515364 230120
rect 514852 229084 514904 229090
rect 514852 229026 514904 229032
rect 514864 223922 514892 229026
rect 514852 223916 514904 223922
rect 514852 223858 514904 223864
rect 515220 223916 515272 223922
rect 515220 223858 515272 223864
rect 514668 223780 514720 223786
rect 514668 223722 514720 223728
rect 514760 218952 514812 218958
rect 514760 218894 514812 218900
rect 514772 218657 514800 218894
rect 514758 218648 514814 218657
rect 514758 218583 514814 218592
rect 514942 218648 514998 218657
rect 514942 218583 514944 218592
rect 514996 218583 514998 218592
rect 514944 218554 514996 218560
rect 515232 217002 515260 223858
rect 515772 223440 515824 223446
rect 515772 223382 515824 223388
rect 515784 221241 515812 223382
rect 515968 223174 515996 231676
rect 516612 227730 516640 231676
rect 517256 229906 517284 231676
rect 517244 229900 517296 229906
rect 517244 229842 517296 229848
rect 516784 229764 516836 229770
rect 516784 229706 516836 229712
rect 516600 227724 516652 227730
rect 516600 227666 516652 227672
rect 516416 227044 516468 227050
rect 516416 226986 516468 226992
rect 515956 223168 516008 223174
rect 515956 223110 516008 223116
rect 515770 221232 515826 221241
rect 515770 221167 515826 221176
rect 510724 216974 511060 217002
rect 511460 216974 511888 217002
rect 512288 216974 512716 217002
rect 513484 216974 513544 217002
rect 514036 216974 514372 217002
rect 515200 216974 515260 217002
rect 515784 217002 515812 221167
rect 516428 217002 516456 226986
rect 516796 223446 516824 229706
rect 517900 226030 517928 231676
rect 518164 229424 518216 229430
rect 518164 229366 518216 229372
rect 517888 226024 517940 226030
rect 517888 225966 517940 225972
rect 516784 223440 516836 223446
rect 516784 223382 516836 223388
rect 518176 220726 518204 229366
rect 518544 228818 518572 231676
rect 518900 230308 518952 230314
rect 518900 230250 518952 230256
rect 518532 228812 518584 228818
rect 518532 228754 518584 228760
rect 518912 226302 518940 230250
rect 519188 230042 519216 231676
rect 519176 230036 519228 230042
rect 519176 229978 519228 229984
rect 518900 226296 518952 226302
rect 518900 226238 518952 226244
rect 519268 226160 519320 226166
rect 519268 226102 519320 226108
rect 518440 223032 518492 223038
rect 518440 222974 518492 222980
rect 518808 223032 518860 223038
rect 518808 222974 518860 222980
rect 518452 221513 518480 222974
rect 518820 222154 518848 222974
rect 518808 222148 518860 222154
rect 518808 222090 518860 222096
rect 518438 221504 518494 221513
rect 518438 221439 518494 221448
rect 518164 220720 518216 220726
rect 518164 220662 518216 220668
rect 517704 220380 517756 220386
rect 517704 220322 517756 220328
rect 517716 217002 517744 220322
rect 515784 216974 516028 217002
rect 516428 216974 516856 217002
rect 517684 216974 517744 217002
rect 518452 217002 518480 221439
rect 518806 220552 518862 220561
rect 518806 220487 518862 220496
rect 518820 220386 518848 220487
rect 518808 220380 518860 220386
rect 518808 220322 518860 220328
rect 519280 217002 519308 226102
rect 519542 224496 519598 224505
rect 519542 224431 519598 224440
rect 519556 223961 519584 224431
rect 519832 224398 519860 231676
rect 520476 230382 520504 231676
rect 520464 230376 520516 230382
rect 520464 230318 520516 230324
rect 521120 227458 521148 231676
rect 521568 230376 521620 230382
rect 521568 230318 521620 230324
rect 521292 228404 521344 228410
rect 521292 228346 521344 228352
rect 521108 227452 521160 227458
rect 521108 227394 521160 227400
rect 519820 224392 519872 224398
rect 519820 224334 519872 224340
rect 519542 223952 519598 223961
rect 519542 223887 519598 223896
rect 519820 222148 519872 222154
rect 519820 222090 519872 222096
rect 519832 217002 519860 222090
rect 521304 220862 521332 228346
rect 521292 220856 521344 220862
rect 521292 220798 521344 220804
rect 521304 217002 521332 220798
rect 521580 220386 521608 230318
rect 521764 228410 521792 231676
rect 522422 231662 522896 231690
rect 522488 229628 522540 229634
rect 522488 229570 522540 229576
rect 521752 228404 521804 228410
rect 521752 228346 521804 228352
rect 522500 223310 522528 229570
rect 521752 223304 521804 223310
rect 521752 223246 521804 223252
rect 522488 223304 522540 223310
rect 522488 223246 522540 223252
rect 521568 220380 521620 220386
rect 521568 220322 521620 220328
rect 518452 216974 518512 217002
rect 519280 216974 519340 217002
rect 519832 216974 520168 217002
rect 520996 216974 521332 217002
rect 521764 217002 521792 223246
rect 522868 221746 522896 231662
rect 523052 229770 523080 231676
rect 523040 229764 523092 229770
rect 523040 229706 523092 229712
rect 523696 227050 523724 231676
rect 523972 231662 524354 231690
rect 523684 227044 523736 227050
rect 523684 226986 523736 226992
rect 523040 224256 523092 224262
rect 523040 224198 523092 224204
rect 523052 222057 523080 224198
rect 523038 222048 523094 222057
rect 523038 221983 523094 221992
rect 523406 222048 523462 222057
rect 523406 221983 523462 221992
rect 522856 221740 522908 221746
rect 522856 221682 522908 221688
rect 521936 220244 521988 220250
rect 521936 220186 521988 220192
rect 521948 219502 521976 220186
rect 521936 219496 521988 219502
rect 521936 219438 521988 219444
rect 522580 219496 522632 219502
rect 522580 219438 522632 219444
rect 522592 217002 522620 219438
rect 523420 217002 523448 221983
rect 523972 221882 524000 231662
rect 524984 229158 525012 231676
rect 525156 230172 525208 230178
rect 525156 230114 525208 230120
rect 524972 229152 525024 229158
rect 524972 229094 525024 229100
rect 524144 225752 524196 225758
rect 524144 225694 524196 225700
rect 524156 224954 524184 225694
rect 524156 224926 524368 224954
rect 523960 221876 524012 221882
rect 523960 221818 524012 221824
rect 524340 219314 524368 224926
rect 525168 222766 525196 230114
rect 525628 225894 525656 231676
rect 525984 229900 526036 229906
rect 525984 229842 526036 229848
rect 525996 226166 526024 229842
rect 525984 226160 526036 226166
rect 525984 226102 526036 226108
rect 525616 225888 525668 225894
rect 525616 225830 525668 225836
rect 526272 224534 526300 231676
rect 526916 230450 526944 231676
rect 526904 230444 526956 230450
rect 526904 230386 526956 230392
rect 526444 227180 526496 227186
rect 526444 227122 526496 227128
rect 525800 224528 525852 224534
rect 525800 224470 525852 224476
rect 526260 224528 526312 224534
rect 526260 224470 526312 224476
rect 525156 222760 525208 222766
rect 525156 222702 525208 222708
rect 524788 222352 524840 222358
rect 524788 222294 524840 222300
rect 524800 222018 524828 222294
rect 524788 222012 524840 222018
rect 524788 221954 524840 221960
rect 524340 219286 524414 219314
rect 524052 219224 524104 219230
rect 524050 219192 524052 219201
rect 524104 219192 524106 219201
rect 524050 219127 524106 219136
rect 524234 219192 524290 219201
rect 524234 219127 524290 219136
rect 524248 219042 524276 219127
rect 524386 219042 524414 219286
rect 524064 219014 524276 219042
rect 524340 219014 524414 219042
rect 524064 218958 524092 219014
rect 524052 218952 524104 218958
rect 524052 218894 524104 218900
rect 524340 218770 524368 219014
rect 523972 218754 524276 218770
rect 523960 218748 524276 218754
rect 524012 218742 524276 218748
rect 524340 218742 524414 218770
rect 523960 218690 524012 218696
rect 524248 218657 524276 218742
rect 523774 218648 523830 218657
rect 523774 218583 523830 218592
rect 524234 218648 524290 218657
rect 524234 218583 524290 218592
rect 523788 218482 523816 218583
rect 524386 218498 524414 218742
rect 523776 218476 523828 218482
rect 523776 218418 523828 218424
rect 524340 218470 524414 218498
rect 524340 217002 524368 218470
rect 521764 216974 521824 217002
rect 522592 216974 522652 217002
rect 523420 216974 523480 217002
rect 524308 216974 524368 217002
rect 524800 217002 524828 221954
rect 525812 217870 525840 224470
rect 526456 220998 526484 227122
rect 527364 225616 527416 225622
rect 527364 225558 527416 225564
rect 527180 223440 527232 223446
rect 527180 223382 527232 223388
rect 527192 222494 527220 223382
rect 527180 222488 527232 222494
rect 527180 222430 527232 222436
rect 526444 220992 526496 220998
rect 526444 220934 526496 220940
rect 526456 219434 526484 220934
rect 526272 219406 526484 219434
rect 525800 217864 525852 217870
rect 525800 217806 525852 217812
rect 526272 217002 526300 219406
rect 526444 217864 526496 217870
rect 526444 217806 526496 217812
rect 524800 216974 525136 217002
rect 525964 216974 526300 217002
rect 526456 217002 526484 217806
rect 527192 217002 527220 222430
rect 527376 221134 527404 225558
rect 527560 224262 527588 231676
rect 528204 227322 528232 231676
rect 528560 230036 528612 230042
rect 528560 229978 528612 229984
rect 528192 227316 528244 227322
rect 528192 227258 528244 227264
rect 527548 224256 527600 224262
rect 527548 224198 527600 224204
rect 528572 223446 528600 229978
rect 528848 229906 528876 231676
rect 528836 229900 528888 229906
rect 528836 229842 528888 229848
rect 528560 223440 528612 223446
rect 528560 223382 528612 223388
rect 528928 222896 528980 222902
rect 528928 222838 528980 222844
rect 527364 221128 527416 221134
rect 527364 221070 527416 221076
rect 528008 221128 528060 221134
rect 528008 221070 528060 221076
rect 528020 217002 528048 221070
rect 528558 220280 528614 220289
rect 528558 220215 528614 220224
rect 528742 220280 528798 220289
rect 528742 220215 528798 220224
rect 528572 219978 528600 220215
rect 528560 219972 528612 219978
rect 528560 219914 528612 219920
rect 528756 219570 528784 220215
rect 528744 219564 528796 219570
rect 528744 219506 528796 219512
rect 528940 219434 528968 222838
rect 529492 222222 529520 231676
rect 530136 230382 530164 231676
rect 530794 231662 531176 231690
rect 531148 230518 531176 231662
rect 531136 230512 531188 230518
rect 531136 230454 531188 230460
rect 530124 230376 530176 230382
rect 530124 230318 530176 230324
rect 531228 230376 531280 230382
rect 531228 230318 531280 230324
rect 530952 228540 531004 228546
rect 530952 228482 531004 228488
rect 529848 225004 529900 225010
rect 529848 224946 529900 224952
rect 529480 222216 529532 222222
rect 529480 222158 529532 222164
rect 529860 220726 529888 224946
rect 530964 221270 530992 228482
rect 530952 221264 531004 221270
rect 530952 221206 531004 221212
rect 529848 220720 529900 220726
rect 529848 220662 529900 220668
rect 528848 219406 528968 219434
rect 529860 219434 529888 220662
rect 529860 219406 529980 219434
rect 528468 219224 528520 219230
rect 528282 219192 528338 219201
rect 528282 219127 528338 219136
rect 528466 219192 528468 219201
rect 528520 219192 528522 219201
rect 528466 219127 528522 219136
rect 528296 218890 528324 219127
rect 528284 218884 528336 218890
rect 528284 218826 528336 218832
rect 528284 218680 528336 218686
rect 528282 218648 528284 218657
rect 528336 218648 528338 218657
rect 528282 218583 528338 218592
rect 528466 218648 528522 218657
rect 528466 218583 528522 218592
rect 528650 218648 528706 218657
rect 528650 218583 528706 218592
rect 528480 218482 528508 218583
rect 528664 218482 528692 218583
rect 528468 218476 528520 218482
rect 528468 218418 528520 218424
rect 528652 218476 528704 218482
rect 528652 218418 528704 218424
rect 528848 217002 528876 219406
rect 529020 218884 529072 218890
rect 529020 218826 529072 218832
rect 529032 218657 529060 218826
rect 529018 218648 529074 218657
rect 529018 218583 529074 218592
rect 529952 217002 529980 219406
rect 530964 217002 530992 221206
rect 531240 220250 531268 230318
rect 531424 228546 531452 231676
rect 532082 231662 532556 231690
rect 531412 228540 531464 228546
rect 531412 228482 531464 228488
rect 531964 226296 532016 226302
rect 531964 226238 532016 226244
rect 531228 220244 531280 220250
rect 531228 220186 531280 220192
rect 531504 220108 531556 220114
rect 531504 220050 531556 220056
rect 526456 216974 526792 217002
rect 527192 216974 527620 217002
rect 528020 216974 528448 217002
rect 528848 216974 529276 217002
rect 529952 216974 530104 217002
rect 530932 216974 530992 217002
rect 531516 217002 531544 220050
rect 531976 218754 532004 226238
rect 532528 220114 532556 231662
rect 532712 229294 532740 231676
rect 532700 229288 532752 229294
rect 532700 229230 532752 229236
rect 533160 227588 533212 227594
rect 533160 227530 533212 227536
rect 533172 222986 533200 227530
rect 533356 227186 533384 231676
rect 533724 231662 534014 231690
rect 533344 227180 533396 227186
rect 533344 227122 533396 227128
rect 533172 222958 533384 222986
rect 533356 222086 533384 222958
rect 533344 222080 533396 222086
rect 532698 222048 532754 222057
rect 532698 221983 532754 221992
rect 532882 222048 532938 222057
rect 533344 222022 533396 222028
rect 532882 221983 532938 221992
rect 532712 221354 532740 221983
rect 532896 221513 532924 221983
rect 532882 221504 532938 221513
rect 532882 221439 532938 221448
rect 533066 221504 533122 221513
rect 533066 221439 533122 221448
rect 533080 221354 533108 221439
rect 532712 221326 533108 221354
rect 532516 220108 532568 220114
rect 532516 220050 532568 220056
rect 531964 218748 532016 218754
rect 531964 218690 532016 218696
rect 532608 218748 532660 218754
rect 532608 218690 532660 218696
rect 532620 217002 532648 218690
rect 531516 216974 531760 217002
rect 532588 216974 532648 217002
rect 533356 217002 533384 222022
rect 533724 221610 533752 231662
rect 534644 230042 534672 231676
rect 534816 230240 534868 230246
rect 534816 230182 534868 230188
rect 534632 230036 534684 230042
rect 534632 229978 534684 229984
rect 534632 229764 534684 229770
rect 534632 229706 534684 229712
rect 534644 224806 534672 229706
rect 534828 229094 534856 230182
rect 534828 229066 535132 229094
rect 534632 224800 534684 224806
rect 534632 224742 534684 224748
rect 534908 223304 534960 223310
rect 534908 223246 534960 223252
rect 533712 221604 533764 221610
rect 533712 221546 533764 221552
rect 534632 221468 534684 221474
rect 534632 221410 534684 221416
rect 534644 220726 534672 221410
rect 534632 220720 534684 220726
rect 534632 220662 534684 220668
rect 534632 220516 534684 220522
rect 534632 220458 534684 220464
rect 534078 220280 534134 220289
rect 534078 220215 534134 220224
rect 534262 220280 534318 220289
rect 534262 220215 534318 220224
rect 534092 219366 534120 220215
rect 534276 219978 534304 220215
rect 534264 219972 534316 219978
rect 534264 219914 534316 219920
rect 534080 219360 534132 219366
rect 534080 219302 534132 219308
rect 534262 219192 534318 219201
rect 534262 219127 534264 219136
rect 534316 219127 534318 219136
rect 534446 219192 534502 219201
rect 534446 219127 534502 219136
rect 534264 219098 534316 219104
rect 534080 218952 534132 218958
rect 534080 218894 534132 218900
rect 534092 218657 534120 218894
rect 534078 218648 534134 218657
rect 534078 218583 534134 218592
rect 534262 218648 534318 218657
rect 534262 218583 534264 218592
rect 534316 218583 534318 218592
rect 534264 218554 534316 218560
rect 534460 218482 534488 219127
rect 534448 218476 534500 218482
rect 534448 218418 534500 218424
rect 534644 217002 534672 220458
rect 534920 218346 534948 223246
rect 535104 220726 535132 229066
rect 535288 225622 535316 231676
rect 535460 230308 535512 230314
rect 535460 230250 535512 230256
rect 535472 229906 535500 230250
rect 535460 229900 535512 229906
rect 535460 229842 535512 229848
rect 535932 228682 535960 231676
rect 536576 229906 536604 231676
rect 536564 229900 536616 229906
rect 536564 229842 536616 229848
rect 536748 229288 536800 229294
rect 536748 229230 536800 229236
rect 535736 228676 535788 228682
rect 535736 228618 535788 228624
rect 535920 228676 535972 228682
rect 535920 228618 535972 228624
rect 535276 225616 535328 225622
rect 535276 225558 535328 225564
rect 535460 221604 535512 221610
rect 535460 221546 535512 221552
rect 535092 220720 535144 220726
rect 535092 220662 535144 220668
rect 535472 220590 535500 221546
rect 535748 220590 535776 228618
rect 536380 223780 536432 223786
rect 536380 223722 536432 223728
rect 535460 220584 535512 220590
rect 535460 220526 535512 220532
rect 535736 220584 535788 220590
rect 535736 220526 535788 220532
rect 534908 218340 534960 218346
rect 534908 218282 534960 218288
rect 533356 216974 533416 217002
rect 534244 216974 534672 217002
rect 534920 217002 534948 218282
rect 535748 217002 535776 220526
rect 536392 217002 536420 223722
rect 536760 223310 536788 229230
rect 536748 223304 536800 223310
rect 536748 223246 536800 223252
rect 537220 222902 537248 231676
rect 537864 225758 537892 231676
rect 538508 229770 538536 231676
rect 538692 231662 539166 231690
rect 538496 229764 538548 229770
rect 538496 229706 538548 229712
rect 537852 225752 537904 225758
rect 537852 225694 537904 225700
rect 538692 224954 538720 231662
rect 539600 230308 539652 230314
rect 539600 230250 539652 230256
rect 538864 227724 538916 227730
rect 538864 227666 538916 227672
rect 538508 224926 538720 224954
rect 538312 223168 538364 223174
rect 538312 223110 538364 223116
rect 537208 222896 537260 222902
rect 537208 222838 537260 222844
rect 537576 222760 537628 222766
rect 537576 222702 537628 222708
rect 537588 217002 537616 222702
rect 534920 216974 535072 217002
rect 535748 216974 535900 217002
rect 536392 216974 536728 217002
rect 537556 216974 537616 217002
rect 538324 217002 538352 223110
rect 538508 221610 538536 224926
rect 538680 222080 538732 222086
rect 538680 222022 538732 222028
rect 538692 221610 538720 222022
rect 538496 221604 538548 221610
rect 538496 221546 538548 221552
rect 538680 221604 538732 221610
rect 538680 221546 538732 221552
rect 538876 217002 538904 227666
rect 539612 226030 539640 230250
rect 543648 230172 543700 230178
rect 543648 230114 543700 230120
rect 541256 228812 541308 228818
rect 541256 228754 541308 228760
rect 539784 226296 539836 226302
rect 539784 226238 539836 226244
rect 539600 226024 539652 226030
rect 539600 225966 539652 225972
rect 539796 223786 539824 226238
rect 540612 226160 540664 226166
rect 540612 226102 540664 226108
rect 539784 223780 539836 223786
rect 539784 223722 539836 223728
rect 539048 223168 539100 223174
rect 539048 223110 539100 223116
rect 539060 222018 539088 223110
rect 539048 222012 539100 222018
rect 539048 221954 539100 221960
rect 539796 217002 539824 223722
rect 540624 219502 540652 226102
rect 540612 219496 540664 219502
rect 540612 219438 540664 219444
rect 540624 217002 540652 219438
rect 541268 217002 541296 228754
rect 542544 224392 542596 224398
rect 542544 224334 542596 224340
rect 542360 223440 542412 223446
rect 542360 223382 542412 223388
rect 542372 222766 542400 223382
rect 542360 222760 542412 222766
rect 542360 222702 542412 222708
rect 542372 217002 542400 222702
rect 542556 219910 542584 224334
rect 543660 223650 543688 230114
rect 552756 230036 552808 230042
rect 552756 229978 552808 229984
rect 549536 228948 549588 228954
rect 549536 228890 549588 228896
rect 545764 228404 545816 228410
rect 545764 228346 545816 228352
rect 544568 227452 544620 227458
rect 544568 227394 544620 227400
rect 544580 224954 544608 227394
rect 544580 224926 544700 224954
rect 543648 223644 543700 223650
rect 543648 223586 543700 223592
rect 543740 220720 543792 220726
rect 544476 220720 544528 220726
rect 543792 220668 544476 220674
rect 543740 220662 544528 220668
rect 543752 220646 544516 220662
rect 543752 220510 544516 220538
rect 543752 220454 543780 220510
rect 543740 220448 543792 220454
rect 543740 220390 543792 220396
rect 543738 220280 543794 220289
rect 543738 220215 543794 220224
rect 543922 220280 543978 220289
rect 543922 220215 543978 220224
rect 542544 219904 542596 219910
rect 542544 219846 542596 219852
rect 543096 219904 543148 219910
rect 543096 219846 543148 219852
rect 543108 217002 543136 219846
rect 543752 219774 543780 220215
rect 543740 219768 543792 219774
rect 543740 219710 543792 219716
rect 543936 219366 543964 220215
rect 543924 219360 543976 219366
rect 543924 219302 543976 219308
rect 543462 219192 543518 219201
rect 543462 219127 543518 219136
rect 543646 219192 543702 219201
rect 543646 219127 543702 219136
rect 543922 219192 543978 219201
rect 543922 219127 543978 219136
rect 544106 219192 544162 219201
rect 544106 219127 544162 219136
rect 544292 219156 544344 219162
rect 543476 218822 543504 219127
rect 543660 218958 543688 219127
rect 543936 218958 543964 219127
rect 543648 218952 543700 218958
rect 543648 218894 543700 218900
rect 543924 218952 543976 218958
rect 543924 218894 543976 218900
rect 543464 218816 543516 218822
rect 543464 218758 543516 218764
rect 543924 218816 543976 218822
rect 543924 218758 543976 218764
rect 543936 218657 543964 218758
rect 543462 218648 543518 218657
rect 543462 218583 543464 218592
rect 543516 218583 543518 218592
rect 543922 218648 543978 218657
rect 544120 218618 544148 219127
rect 544292 219098 544344 219104
rect 544304 218618 544332 219098
rect 543922 218583 543978 218592
rect 544108 218612 544160 218618
rect 543464 218554 543516 218560
rect 544108 218554 544160 218560
rect 544292 218612 544344 218618
rect 544292 218554 544344 218560
rect 544488 217002 544516 220510
rect 544672 219230 544700 224926
rect 545776 219638 545804 228346
rect 548524 227044 548576 227050
rect 548524 226986 548576 226992
rect 547420 224800 547472 224806
rect 547420 224742 547472 224748
rect 546500 221740 546552 221746
rect 546500 221682 546552 221688
rect 545764 219632 545816 219638
rect 545764 219574 545816 219580
rect 544660 219224 544712 219230
rect 544660 219166 544712 219172
rect 538324 216974 538384 217002
rect 538876 216974 539212 217002
rect 539796 216974 540040 217002
rect 540624 216974 540868 217002
rect 541268 216974 541696 217002
rect 542372 216974 542524 217002
rect 543108 216974 543352 217002
rect 544180 216974 544516 217002
rect 544672 217002 544700 219166
rect 545776 217002 545804 219574
rect 546512 217002 546540 221682
rect 547432 219094 547460 224742
rect 548536 221746 548564 226986
rect 549548 224398 549576 228890
rect 551008 225888 551060 225894
rect 551008 225830 551060 225836
rect 549536 224392 549588 224398
rect 549536 224334 549588 224340
rect 548984 221876 549036 221882
rect 548984 221818 549036 221824
rect 548524 221740 548576 221746
rect 548524 221682 548576 221688
rect 547420 219088 547472 219094
rect 547420 219030 547472 219036
rect 547432 217002 547460 219030
rect 548536 217002 548564 221682
rect 548708 220176 548760 220182
rect 548708 220118 548760 220124
rect 548720 219774 548748 220118
rect 548708 219768 548760 219774
rect 548708 219710 548760 219716
rect 544672 216974 545008 217002
rect 545776 216974 545836 217002
rect 546512 216974 546664 217002
rect 547432 216974 547492 217002
rect 548320 216974 548564 217002
rect 548996 217002 549024 221818
rect 549548 217002 549576 224334
rect 551020 219774 551048 225830
rect 551836 224800 551888 224806
rect 551836 224742 551888 224748
rect 551284 224528 551336 224534
rect 551284 224470 551336 224476
rect 551008 219768 551060 219774
rect 551008 219710 551060 219716
rect 551020 217002 551048 219710
rect 548996 216974 549148 217002
rect 549548 216974 549976 217002
rect 550804 216974 551048 217002
rect 551296 217002 551324 224470
rect 551848 220726 551876 224742
rect 552768 224534 552796 229978
rect 554056 228410 554084 240343
rect 554320 238740 554372 238746
rect 554320 238682 554372 238688
rect 554332 238241 554360 238682
rect 554318 238232 554374 238241
rect 554318 238167 554374 238176
rect 554504 236088 554556 236094
rect 554502 236056 554504 236065
rect 554556 236056 554558 236065
rect 554502 235991 554558 236000
rect 554412 234592 554464 234598
rect 554412 234534 554464 234540
rect 554424 233889 554452 234534
rect 554410 233880 554466 233889
rect 554410 233815 554466 233824
rect 554044 228404 554096 228410
rect 554044 228346 554096 228352
rect 553676 227316 553728 227322
rect 553676 227258 553728 227264
rect 552756 224528 552808 224534
rect 552756 224470 552808 224476
rect 552020 224256 552072 224262
rect 552020 224198 552072 224204
rect 551836 220720 551888 220726
rect 551836 220662 551888 220668
rect 551848 219450 551876 220662
rect 552032 220454 552060 224198
rect 553308 220584 553360 220590
rect 553308 220526 553360 220532
rect 553492 220584 553544 220590
rect 553492 220526 553544 220532
rect 552020 220448 552072 220454
rect 552020 220390 552072 220396
rect 552756 220448 552808 220454
rect 552756 220390 552808 220396
rect 551848 219422 552060 219450
rect 552032 217002 552060 219422
rect 552570 219192 552626 219201
rect 552570 219127 552626 219136
rect 552584 218958 552612 219127
rect 552572 218952 552624 218958
rect 552572 218894 552624 218900
rect 552768 217002 552796 220390
rect 553320 220289 553348 220526
rect 553122 220280 553178 220289
rect 553122 220215 553178 220224
rect 553306 220280 553362 220289
rect 553306 220215 553362 220224
rect 553136 219366 553164 220215
rect 553504 220046 553532 220526
rect 553492 220040 553544 220046
rect 553492 219982 553544 219988
rect 553124 219360 553176 219366
rect 553124 219302 553176 219308
rect 552938 219192 552994 219201
rect 552938 219127 552994 219136
rect 552952 218618 552980 219127
rect 553490 218920 553546 218929
rect 553490 218855 553546 218864
rect 553308 218816 553360 218822
rect 553308 218758 553360 218764
rect 553320 218657 553348 218758
rect 553504 218754 553532 218855
rect 553492 218748 553544 218754
rect 553492 218690 553544 218696
rect 553122 218648 553178 218657
rect 552940 218612 552992 218618
rect 553122 218583 553124 218592
rect 552940 218554 552992 218560
rect 553176 218583 553178 218592
rect 553306 218648 553362 218657
rect 553306 218583 553362 218592
rect 553124 218554 553176 218560
rect 553490 217832 553546 217841
rect 553490 217767 553546 217776
rect 553216 217592 553268 217598
rect 553214 217560 553216 217569
rect 553268 217560 553270 217569
rect 553214 217495 553270 217504
rect 553504 217025 553532 217767
rect 553490 217016 553546 217025
rect 551296 216974 551632 217002
rect 552032 216974 552460 217002
rect 552768 216974 553288 217002
rect 508870 216951 508926 216960
rect 553688 217002 553716 227258
rect 555436 227050 555464 244258
rect 555424 227044 555476 227050
rect 555424 226986 555476 226992
rect 555332 226024 555384 226030
rect 555332 225966 555384 225972
rect 555344 218958 555372 225966
rect 556816 224262 556844 251194
rect 558184 242208 558236 242214
rect 558184 242150 558236 242156
rect 558196 236094 558224 242150
rect 558184 236088 558236 236094
rect 558184 236030 558236 236036
rect 559576 230042 559604 256702
rect 559564 230036 559616 230042
rect 559564 229978 559616 229984
rect 559748 229900 559800 229906
rect 559748 229842 559800 229848
rect 558368 228540 558420 228546
rect 558368 228482 558420 228488
rect 558380 224954 558408 228482
rect 558380 224926 558592 224954
rect 558184 224800 558236 224806
rect 558184 224742 558236 224748
rect 558368 224800 558420 224806
rect 558368 224742 558420 224748
rect 558196 224534 558224 224742
rect 558000 224528 558052 224534
rect 558000 224470 558052 224476
rect 558184 224528 558236 224534
rect 558184 224470 558236 224476
rect 558012 224346 558040 224470
rect 558380 224346 558408 224742
rect 558012 224318 558408 224346
rect 556804 224256 556856 224262
rect 556804 224198 556856 224204
rect 557448 223644 557500 223650
rect 557448 223586 557500 223592
rect 555700 222216 555752 222222
rect 555700 222158 555752 222164
rect 553860 218952 553912 218958
rect 553858 218920 553860 218929
rect 555332 218952 555384 218958
rect 553912 218920 553914 218929
rect 555332 218894 555384 218900
rect 553858 218855 553914 218864
rect 553858 218648 553914 218657
rect 553858 218583 553860 218592
rect 553912 218583 553914 218592
rect 553860 218554 553912 218560
rect 554228 217592 554280 217598
rect 554226 217560 554228 217569
rect 554280 217560 554282 217569
rect 554226 217495 554282 217504
rect 555344 217002 555372 218894
rect 555712 217870 555740 222158
rect 556252 220312 556304 220318
rect 556252 220254 556304 220260
rect 555700 217864 555752 217870
rect 555700 217806 555752 217812
rect 553688 216974 554116 217002
rect 554944 216974 555372 217002
rect 555712 217002 555740 217806
rect 556264 217002 556292 220254
rect 557460 217002 557488 223586
rect 558564 220726 558592 224926
rect 559760 220726 559788 229842
rect 559932 223304 559984 223310
rect 559932 223246 559984 223252
rect 558000 220720 558052 220726
rect 558000 220662 558052 220668
rect 558552 220720 558604 220726
rect 558552 220662 558604 220668
rect 559748 220720 559800 220726
rect 559748 220662 559800 220668
rect 555712 216974 555772 217002
rect 556264 216974 556600 217002
rect 557428 216974 557488 217002
rect 558012 217002 558040 220662
rect 558564 220250 558592 220662
rect 558920 220584 558972 220590
rect 558920 220526 558972 220532
rect 558552 220244 558604 220250
rect 558552 220186 558604 220192
rect 558368 219224 558420 219230
rect 558368 219166 558420 219172
rect 558184 219088 558236 219094
rect 558184 219030 558236 219036
rect 558196 218618 558224 219030
rect 558184 218612 558236 218618
rect 558184 218554 558236 218560
rect 558380 218210 558408 219166
rect 558736 218884 558788 218890
rect 558736 218826 558788 218832
rect 558184 218204 558236 218210
rect 558184 218146 558236 218152
rect 558368 218204 558420 218210
rect 558368 218146 558420 218152
rect 558196 218090 558224 218146
rect 558748 218090 558776 218826
rect 558196 218062 558776 218090
rect 558932 217002 558960 220526
rect 559944 217002 559972 223246
rect 560760 221876 560812 221882
rect 560760 221818 560812 221824
rect 560772 221474 560800 221818
rect 560760 221468 560812 221474
rect 560760 221410 560812 221416
rect 560956 221406 560984 259422
rect 562324 252612 562376 252618
rect 562324 252554 562376 252560
rect 562336 229094 562364 252554
rect 567200 230036 567252 230042
rect 567200 229978 567252 229984
rect 565084 229764 565136 229770
rect 565084 229706 565136 229712
rect 562336 229066 562548 229094
rect 561312 227180 561364 227186
rect 561312 227122 561364 227128
rect 561324 224954 561352 227122
rect 561140 224926 561352 224954
rect 560944 221400 560996 221406
rect 560944 221342 560996 221348
rect 561140 217734 561168 224926
rect 562048 224800 562100 224806
rect 562048 224742 562100 224748
rect 561312 221876 561364 221882
rect 561312 221818 561364 221824
rect 561128 217728 561180 217734
rect 561128 217670 561180 217676
rect 561140 217274 561168 217670
rect 561048 217246 561168 217274
rect 561048 217002 561076 217246
rect 558012 216974 558256 217002
rect 558932 216974 559084 217002
rect 559912 216974 559972 217002
rect 560740 216974 561076 217002
rect 561324 217002 561352 221818
rect 562060 217002 562088 224742
rect 562520 220522 562548 229066
rect 563060 228676 563112 228682
rect 563060 228618 563112 228624
rect 563072 224954 563100 228618
rect 563520 225616 563572 225622
rect 563520 225558 563572 225564
rect 563532 224954 563560 225558
rect 563072 224926 563284 224954
rect 562508 220516 562560 220522
rect 562508 220458 562560 220464
rect 563256 219230 563284 224926
rect 563348 224926 563560 224954
rect 563348 220538 563376 224926
rect 565096 221882 565124 229706
rect 567212 229094 567240 229978
rect 568592 229094 568620 260850
rect 570616 234598 570644 261462
rect 571340 249076 571392 249082
rect 571340 249018 571392 249024
rect 570604 234592 570656 234598
rect 570604 234534 570656 234540
rect 571352 229094 571380 249018
rect 577516 238746 577544 261598
rect 645872 261526 645900 277766
rect 645860 261520 645912 261526
rect 645860 261462 645912 261468
rect 632704 246356 632756 246362
rect 632704 246298 632756 246304
rect 592684 245676 592736 245682
rect 592684 245618 592736 245624
rect 577504 238740 577556 238746
rect 577504 238682 577556 238688
rect 567212 229066 567976 229094
rect 568592 229066 569448 229094
rect 571352 229066 571932 229094
rect 566096 225752 566148 225758
rect 566096 225694 566148 225700
rect 565636 222896 565688 222902
rect 565636 222838 565688 222844
rect 565084 221876 565136 221882
rect 565084 221818 565136 221824
rect 563532 220918 563744 220946
rect 563532 220726 563560 220918
rect 563716 220810 563744 220918
rect 563716 220782 564480 220810
rect 563520 220720 563572 220726
rect 563520 220662 563572 220668
rect 563704 220652 563756 220658
rect 563704 220594 563756 220600
rect 563716 220538 563744 220594
rect 563348 220510 563744 220538
rect 563348 219722 563376 220510
rect 563348 219694 563468 219722
rect 563244 219224 563296 219230
rect 563244 219166 563296 219172
rect 562784 219156 562836 219162
rect 562784 219098 562836 219104
rect 563060 219156 563112 219162
rect 563060 219098 563112 219104
rect 562796 218929 562824 219098
rect 563072 219042 563100 219098
rect 563072 219014 563284 219042
rect 562782 218920 562838 218929
rect 562782 218855 562838 218864
rect 563058 218920 563114 218929
rect 563058 218855 563114 218864
rect 563072 218754 563100 218855
rect 563060 218748 563112 218754
rect 563060 218690 563112 218696
rect 563256 218385 563284 219014
rect 563058 218376 563114 218385
rect 563058 218311 563114 218320
rect 563242 218376 563298 218385
rect 563242 218311 563298 218320
rect 562876 217864 562928 217870
rect 562874 217832 562876 217841
rect 562928 217832 562930 217841
rect 562874 217767 562930 217776
rect 563072 217598 563100 218311
rect 563244 217728 563296 217734
rect 563244 217670 563296 217676
rect 563060 217592 563112 217598
rect 563060 217534 563112 217540
rect 563256 217297 563284 217670
rect 563058 217288 563114 217297
rect 563058 217223 563060 217232
rect 563112 217223 563114 217232
rect 563242 217288 563298 217297
rect 563242 217223 563298 217232
rect 563060 217194 563112 217200
rect 562692 217116 562744 217122
rect 562692 217058 562744 217064
rect 562704 217002 562732 217058
rect 563440 217002 563468 219694
rect 564452 219230 564480 220782
rect 563704 219224 563756 219230
rect 563704 219166 563756 219172
rect 564440 219224 564492 219230
rect 564440 219166 564492 219172
rect 565176 219224 565228 219230
rect 565176 219166 565228 219172
rect 561324 216974 561568 217002
rect 562060 216974 562732 217002
rect 563224 216974 563468 217002
rect 563716 217002 563744 219166
rect 565188 217938 565216 219166
rect 565176 217932 565228 217938
rect 565176 217874 565228 217880
rect 565188 217002 565216 217874
rect 563716 216974 564052 217002
rect 564880 216974 565216 217002
rect 565648 217002 565676 222838
rect 566108 217002 566136 225694
rect 567752 223304 567804 223310
rect 567752 223246 567804 223252
rect 567764 222222 567792 223246
rect 567752 222216 567804 222222
rect 567752 222158 567804 222164
rect 567292 221876 567344 221882
rect 567292 221818 567344 221824
rect 567016 219156 567068 219162
rect 567016 219098 567068 219104
rect 567304 219144 567332 221818
rect 567304 219116 567700 219144
rect 567028 218210 567056 219098
rect 567016 218204 567068 218210
rect 567016 218146 567068 218152
rect 567304 217002 567332 219116
rect 567672 219026 567700 219116
rect 567476 219020 567528 219026
rect 567476 218962 567528 218968
rect 567660 219020 567712 219026
rect 567660 218962 567712 218968
rect 567488 218210 567516 218962
rect 567752 218612 567804 218618
rect 567752 218554 567804 218560
rect 567764 218346 567792 218554
rect 567752 218340 567804 218346
rect 567752 218282 567804 218288
rect 567476 218204 567528 218210
rect 567476 218146 567528 218152
rect 567948 217002 567976 229066
rect 568672 221400 568724 221406
rect 568672 221342 568724 221348
rect 568120 218884 568172 218890
rect 568120 218826 568172 218832
rect 568304 218884 568356 218890
rect 568304 218826 568356 218832
rect 568132 218346 568160 218826
rect 568120 218340 568172 218346
rect 568120 218282 568172 218288
rect 568316 217938 568344 218826
rect 568304 217932 568356 217938
rect 568304 217874 568356 217880
rect 568684 217002 568712 221342
rect 569420 217002 569448 229066
rect 570328 224256 570380 224262
rect 570328 224198 570380 224204
rect 570340 217002 570368 224198
rect 571616 222896 571668 222902
rect 571616 222838 571668 222844
rect 571628 220658 571656 222838
rect 571616 220652 571668 220658
rect 571616 220594 571668 220600
rect 571340 220516 571392 220522
rect 571340 220458 571392 220464
rect 571352 217002 571380 220458
rect 571708 217388 571760 217394
rect 571708 217330 571760 217336
rect 571720 217025 571748 217330
rect 571706 217016 571762 217025
rect 565648 216974 565708 217002
rect 566108 216974 566536 217002
rect 567304 216974 567364 217002
rect 567948 216974 568192 217002
rect 568684 216974 569020 217002
rect 569420 216974 569848 217002
rect 570340 216974 570676 217002
rect 571352 216974 571504 217002
rect 553490 216951 553546 216960
rect 571904 217002 571932 229066
rect 581644 228404 581696 228410
rect 581644 228346 581696 228352
rect 579540 219406 579752 219434
rect 579540 219314 579568 219406
rect 579448 219298 579568 219314
rect 579724 219298 579752 219406
rect 579436 219292 579568 219298
rect 579488 219286 579568 219292
rect 579712 219292 579764 219298
rect 579436 219234 579488 219240
rect 579712 219234 579764 219240
rect 577504 219156 577556 219162
rect 577504 219098 577556 219104
rect 576044 219026 576624 219042
rect 572168 219020 572220 219026
rect 572168 218962 572220 218968
rect 576044 219020 576636 219026
rect 576044 219014 576584 219020
rect 572180 217938 572208 218962
rect 572444 218884 572496 218890
rect 572444 218826 572496 218832
rect 572456 218385 572484 218826
rect 572442 218376 572498 218385
rect 572442 218311 572498 218320
rect 576044 217938 576072 219014
rect 576584 218962 576636 218968
rect 576216 218884 576268 218890
rect 576584 218884 576636 218890
rect 576268 218844 576440 218872
rect 576216 218826 576268 218832
rect 576216 218748 576268 218754
rect 576216 218690 576268 218696
rect 576228 217938 576256 218690
rect 576412 218226 576440 218844
rect 576584 218826 576636 218832
rect 576596 218385 576624 218826
rect 576582 218376 576638 218385
rect 576582 218311 576638 218320
rect 576766 218376 576822 218385
rect 576766 218311 576822 218320
rect 576780 218226 576808 218311
rect 576412 218198 576808 218226
rect 572168 217932 572220 217938
rect 572168 217874 572220 217880
rect 576032 217932 576084 217938
rect 576032 217874 576084 217880
rect 576216 217932 576268 217938
rect 576216 217874 576268 217880
rect 572352 217796 572404 217802
rect 572352 217738 572404 217744
rect 576584 217796 576636 217802
rect 576584 217738 576636 217744
rect 572364 217297 572392 217738
rect 576596 217682 576624 217738
rect 576596 217654 576808 217682
rect 576780 217569 576808 217654
rect 577320 217660 577372 217666
rect 577320 217602 577372 217608
rect 576582 217560 576638 217569
rect 576582 217495 576584 217504
rect 576636 217495 576638 217504
rect 576766 217560 576822 217569
rect 576766 217495 576822 217504
rect 576952 217524 577004 217530
rect 576584 217466 576636 217472
rect 576952 217466 577004 217472
rect 572350 217288 572406 217297
rect 572350 217223 572406 217232
rect 572534 217288 572590 217297
rect 572534 217223 572590 217232
rect 575386 217288 575442 217297
rect 575386 217223 575442 217232
rect 572548 217122 572576 217223
rect 572536 217116 572588 217122
rect 572536 217058 572588 217064
rect 571904 216974 572332 217002
rect 571706 216951 571762 216960
rect 575400 216481 575428 217223
rect 576964 217025 576992 217466
rect 577136 217388 577188 217394
rect 577136 217330 577188 217336
rect 576950 217016 577006 217025
rect 576950 216951 577006 216960
rect 577148 216753 577176 217330
rect 577134 216744 577190 216753
rect 577134 216679 577190 216688
rect 575386 216472 575442 216481
rect 575386 216407 575442 216416
rect 577332 215150 577360 217602
rect 577320 215144 577372 215150
rect 577320 215086 577372 215092
rect 577516 214606 577544 219098
rect 577688 219020 577740 219026
rect 577688 218962 577740 218968
rect 577700 215966 577728 218962
rect 577872 218612 577924 218618
rect 577872 218554 577924 218560
rect 577688 215960 577740 215966
rect 577688 215902 577740 215908
rect 577884 215014 577912 218554
rect 578056 218476 578108 218482
rect 578056 218418 578108 218424
rect 577872 215008 577924 215014
rect 577872 214950 577924 214956
rect 578068 214878 578096 218418
rect 578240 217796 578292 217802
rect 578240 217738 578292 217744
rect 578056 214872 578108 214878
rect 578056 214814 578108 214820
rect 578252 214742 578280 217738
rect 578240 214736 578292 214742
rect 578240 214678 578292 214684
rect 577504 214600 577556 214606
rect 577504 214542 577556 214548
rect 578882 214024 578938 214033
rect 578882 213959 578938 213968
rect 578514 211712 578570 211721
rect 578514 211647 578570 211656
rect 578528 211206 578556 211647
rect 578516 211200 578568 211206
rect 578516 211142 578568 211148
rect 578424 209840 578476 209846
rect 578422 209808 578424 209817
rect 578476 209808 578478 209817
rect 578422 209743 578478 209752
rect 578896 208350 578924 213959
rect 580908 211200 580960 211206
rect 580908 211142 580960 211148
rect 580080 209840 580132 209846
rect 580080 209782 580132 209788
rect 578884 208344 578936 208350
rect 578884 208286 578936 208292
rect 580092 207670 580120 209782
rect 580264 208616 580316 208622
rect 580264 208558 580316 208564
rect 580080 207664 580132 207670
rect 580080 207606 580132 207612
rect 579526 207496 579582 207505
rect 579582 207454 579752 207482
rect 579526 207431 579582 207440
rect 579526 205864 579582 205873
rect 579526 205799 579528 205808
rect 579580 205799 579582 205808
rect 579528 205770 579580 205776
rect 579724 204270 579752 207454
rect 579712 204264 579764 204270
rect 579712 204206 579764 204212
rect 578514 203280 578570 203289
rect 578514 203215 578570 203224
rect 578528 202978 578556 203215
rect 578516 202972 578568 202978
rect 578516 202914 578568 202920
rect 578790 200832 578846 200841
rect 578790 200767 578846 200776
rect 578804 200190 578832 200767
rect 578792 200184 578844 200190
rect 578792 200126 578844 200132
rect 579526 198928 579582 198937
rect 579526 198863 579582 198872
rect 579540 198762 579568 198863
rect 579528 198756 579580 198762
rect 579528 198698 579580 198704
rect 578514 196480 578570 196489
rect 578514 196415 578570 196424
rect 578528 196042 578556 196415
rect 578516 196036 578568 196042
rect 578516 195978 578568 195984
rect 579526 194984 579582 194993
rect 579526 194919 579582 194928
rect 579540 194614 579568 194919
rect 579528 194608 579580 194614
rect 579528 194550 579580 194556
rect 579526 192264 579582 192273
rect 579526 192199 579582 192208
rect 579540 191894 579568 192199
rect 579528 191888 579580 191894
rect 579528 191830 579580 191836
rect 579526 190768 579582 190777
rect 579526 190703 579582 190712
rect 579540 190534 579568 190703
rect 579528 190528 579580 190534
rect 579528 190470 579580 190476
rect 579526 188048 579582 188057
rect 579526 187983 579582 187992
rect 579540 187746 579568 187983
rect 579528 187740 579580 187746
rect 579528 187682 579580 187688
rect 579528 186312 579580 186318
rect 579526 186280 579528 186289
rect 579580 186280 579582 186289
rect 579526 186215 579582 186224
rect 579528 184884 579580 184890
rect 579528 184826 579580 184832
rect 579540 184385 579568 184826
rect 579526 184376 579582 184385
rect 579526 184311 579582 184320
rect 579528 182164 579580 182170
rect 579528 182106 579580 182112
rect 579540 181937 579568 182106
rect 579526 181928 579582 181937
rect 579526 181863 579582 181872
rect 578792 180804 578844 180810
rect 578792 180746 578844 180752
rect 578804 180169 578832 180746
rect 578790 180160 578846 180169
rect 578790 180095 578846 180104
rect 578792 178084 578844 178090
rect 578792 178026 578844 178032
rect 578804 175137 578832 178026
rect 579528 177948 579580 177954
rect 579528 177890 579580 177896
rect 579540 177721 579568 177890
rect 579526 177712 579582 177721
rect 579526 177647 579582 177656
rect 578790 175128 578846 175137
rect 578790 175063 578846 175072
rect 578424 174548 578476 174554
rect 578424 174490 578476 174496
rect 578436 173505 578464 174490
rect 578422 173496 578478 173505
rect 578422 173431 578478 173440
rect 578240 173256 578292 173262
rect 578240 173198 578292 173204
rect 578252 171057 578280 173198
rect 578424 172508 578476 172514
rect 578424 172450 578476 172456
rect 578238 171048 578294 171057
rect 578238 170983 578294 170992
rect 578436 169289 578464 172450
rect 579804 171148 579856 171154
rect 579632 171106 579804 171134
rect 578422 169280 578478 169289
rect 578422 169215 578478 169224
rect 579632 168450 579660 171106
rect 579804 171090 579856 171096
rect 579540 168422 579660 168450
rect 579540 166977 579568 168422
rect 579526 166968 579582 166977
rect 579526 166903 579582 166912
rect 579528 166320 579580 166326
rect 579528 166262 579580 166268
rect 579344 164892 579396 164898
rect 579344 164834 579396 164840
rect 579356 162761 579384 164834
rect 579540 164529 579568 166262
rect 579526 164520 579582 164529
rect 579526 164455 579582 164464
rect 579342 162752 579398 162761
rect 579342 162687 579398 162696
rect 578240 162580 578292 162586
rect 578240 162522 578292 162528
rect 578252 159905 578280 162522
rect 578424 162172 578476 162178
rect 578424 162114 578476 162120
rect 578238 159896 578294 159905
rect 578238 159831 578294 159840
rect 578436 158409 578464 162114
rect 578422 158400 578478 158409
rect 578422 158335 578478 158344
rect 578516 157616 578568 157622
rect 578516 157558 578568 157564
rect 578528 155961 578556 157558
rect 578514 155952 578570 155961
rect 578514 155887 578570 155896
rect 578700 154216 578752 154222
rect 578700 154158 578752 154164
rect 578712 154057 578740 154158
rect 578698 154048 578754 154057
rect 578698 153983 578754 153992
rect 578240 152652 578292 152658
rect 578240 152594 578292 152600
rect 578252 151745 578280 152594
rect 578238 151736 578294 151745
rect 578238 151671 578294 151680
rect 578332 151088 578384 151094
rect 578332 151030 578384 151036
rect 578344 149705 578372 151030
rect 578330 149696 578386 149705
rect 578330 149631 578386 149640
rect 579528 148368 579580 148374
rect 579528 148310 579580 148316
rect 579540 147529 579568 148310
rect 579526 147520 579582 147529
rect 579526 147455 579582 147464
rect 578884 145580 578936 145586
rect 578884 145522 578936 145528
rect 578608 139324 578660 139330
rect 578608 139266 578660 139272
rect 578620 138825 578648 139266
rect 578606 138816 578662 138825
rect 578606 138751 578662 138760
rect 578896 136649 578924 145522
rect 579436 144696 579488 144702
rect 579434 144664 579436 144673
rect 579488 144664 579490 144673
rect 579434 144599 579490 144608
rect 579528 143472 579580 143478
rect 579528 143414 579580 143420
rect 579540 143041 579568 143414
rect 579526 143032 579582 143041
rect 579526 142967 579582 142976
rect 579528 140616 579580 140622
rect 579526 140584 579528 140593
rect 579580 140584 579582 140593
rect 579526 140519 579582 140528
rect 579528 138168 579580 138174
rect 579528 138110 579580 138116
rect 579068 137284 579120 137290
rect 579068 137226 579120 137232
rect 578882 136640 578938 136649
rect 578882 136575 578938 136584
rect 579080 132297 579108 137226
rect 579540 134473 579568 138110
rect 579526 134464 579582 134473
rect 579526 134399 579582 134408
rect 579066 132288 579122 132297
rect 579066 132223 579122 132232
rect 578700 131776 578752 131782
rect 578700 131718 578752 131724
rect 578712 129713 578740 131718
rect 578698 129704 578754 129713
rect 578698 129639 578754 129648
rect 578516 128036 578568 128042
rect 578516 127978 578568 127984
rect 578528 127809 578556 127978
rect 578514 127800 578570 127809
rect 578514 127735 578570 127744
rect 579068 127016 579120 127022
rect 579068 126958 579120 126964
rect 578884 122256 578936 122262
rect 578884 122198 578936 122204
rect 578516 121372 578568 121378
rect 578516 121314 578568 121320
rect 578528 121145 578556 121314
rect 578514 121136 578570 121145
rect 578514 121071 578570 121080
rect 578516 114504 578568 114510
rect 578514 114472 578516 114481
rect 578568 114472 578570 114481
rect 578514 114407 578570 114416
rect 578896 110401 578924 122198
rect 578882 110392 578938 110401
rect 578882 110327 578938 110336
rect 578332 108724 578384 108730
rect 578332 108666 578384 108672
rect 578344 108361 578372 108666
rect 578330 108352 578386 108361
rect 578330 108287 578386 108296
rect 579080 105913 579108 126958
rect 579528 125384 579580 125390
rect 579526 125352 579528 125361
rect 579580 125352 579582 125361
rect 579526 125287 579582 125296
rect 579252 124160 579304 124166
rect 579252 124102 579304 124108
rect 579264 123593 579292 124102
rect 579250 123584 579306 123593
rect 579250 123519 579306 123528
rect 579528 118448 579580 118454
rect 579526 118416 579528 118425
rect 579580 118416 579582 118425
rect 579526 118351 579582 118360
rect 579344 117224 579396 117230
rect 579344 117166 579396 117172
rect 579356 116929 579384 117166
rect 579342 116920 579398 116929
rect 579342 116855 579398 116864
rect 580276 114510 580304 208558
rect 580920 206922 580948 211142
rect 580908 206916 580960 206922
rect 580908 206858 580960 206864
rect 580448 202972 580500 202978
rect 580448 202914 580500 202920
rect 580460 200054 580488 202914
rect 580448 200048 580500 200054
rect 580448 199990 580500 199996
rect 580908 162920 580960 162926
rect 580908 162862 580960 162868
rect 580920 157622 580948 162862
rect 580908 157616 580960 157622
rect 580908 157558 580960 157564
rect 580448 137420 580500 137426
rect 580448 137362 580500 137368
rect 580460 128042 580488 137362
rect 580448 128036 580500 128042
rect 580448 127978 580500 127984
rect 580632 125656 580684 125662
rect 580632 125598 580684 125604
rect 580448 122120 580500 122126
rect 580448 122062 580500 122068
rect 580264 114504 580316 114510
rect 580264 114446 580316 114452
rect 579528 113144 579580 113150
rect 579528 113086 579580 113092
rect 579540 112713 579568 113086
rect 579526 112704 579582 112713
rect 579526 112639 579582 112648
rect 580264 106344 580316 106350
rect 580264 106286 580316 106292
rect 579066 105904 579122 105913
rect 579066 105839 579122 105848
rect 579436 105188 579488 105194
rect 579436 105130 579488 105136
rect 579252 103352 579304 103358
rect 579250 103320 579252 103329
rect 579304 103320 579306 103329
rect 579250 103255 579306 103264
rect 578332 101720 578384 101726
rect 578330 101688 578332 101697
rect 578384 101688 578386 101697
rect 578330 101623 578386 101632
rect 578606 99376 578662 99385
rect 578606 99311 578608 99320
rect 578660 99311 578662 99320
rect 578608 99282 578660 99288
rect 579252 98796 579304 98802
rect 579252 98738 579304 98744
rect 579264 97481 579292 98738
rect 579250 97472 579306 97481
rect 577688 97436 577740 97442
rect 579250 97407 579306 97416
rect 577688 97378 577740 97384
rect 577504 97300 577556 97306
rect 577504 97242 577556 97248
rect 312018 53108 314042 53122
rect 130384 52012 130436 52018
rect 130384 51954 130436 51960
rect 129372 51876 129424 51882
rect 129372 51818 129424 51824
rect 129186 51776 129242 51785
rect 129004 51740 129056 51746
rect 129186 51711 129242 51720
rect 129004 51682 129056 51688
rect 50528 50652 50580 50658
rect 50528 50594 50580 50600
rect 128452 50652 128504 50658
rect 128452 50594 128504 50600
rect 48964 49292 49016 49298
rect 48964 49234 49016 49240
rect 46388 49020 46440 49026
rect 46388 48962 46440 48968
rect 128464 48142 128492 50594
rect 128636 50380 128688 50386
rect 128636 50322 128688 50328
rect 128452 48136 128504 48142
rect 128452 48078 128504 48084
rect 128648 47870 128676 50322
rect 128820 49156 128872 49162
rect 128820 49098 128872 49104
rect 128636 47864 128688 47870
rect 128636 47806 128688 47812
rect 128832 44266 128860 49098
rect 129016 44946 129044 51682
rect 129004 44940 129056 44946
rect 129004 44882 129056 44888
rect 129200 44810 129228 51711
rect 129188 44804 129240 44810
rect 129188 44746 129240 44752
rect 129384 44674 129412 51818
rect 130396 51074 130424 51954
rect 306024 51746 306052 53108
rect 145380 51740 145432 51746
rect 145380 51682 145432 51688
rect 306012 51740 306064 51746
rect 306012 51682 306064 51688
rect 130396 51046 130700 51074
rect 129556 49292 129608 49298
rect 129556 49234 129608 49240
rect 129568 45082 129596 49234
rect 130476 49020 130528 49026
rect 130476 48962 130528 48968
rect 129556 45076 129608 45082
rect 129556 45018 129608 45024
rect 129372 44668 129424 44674
rect 129372 44610 129424 44616
rect 130488 44305 130516 48962
rect 130474 44296 130530 44305
rect 128820 44260 128872 44266
rect 130474 44231 130530 44240
rect 128820 44202 128872 44208
rect 130672 44130 130700 51046
rect 145392 50810 145420 51682
rect 145084 50782 145420 50810
rect 131028 50516 131080 50522
rect 131028 50458 131080 50464
rect 130660 44124 130712 44130
rect 130660 44066 130712 44072
rect 131040 43994 131068 50458
rect 308048 50289 308076 53108
rect 312018 53094 314056 53108
rect 316020 53094 318380 53122
rect 314028 50386 314056 53094
rect 318352 50522 318380 53094
rect 464988 52828 465040 52834
rect 464988 52770 465040 52776
rect 467012 52828 467064 52834
rect 467012 52770 467064 52776
rect 459020 52686 459324 52714
rect 457720 52284 457772 52290
rect 457720 52226 457772 52232
rect 318340 50516 318392 50522
rect 318340 50458 318392 50464
rect 314016 50380 314068 50386
rect 314016 50322 314068 50328
rect 308034 50280 308090 50289
rect 308034 50215 308090 50224
rect 131948 48136 132000 48142
rect 131948 48078 132000 48084
rect 131764 47864 131816 47870
rect 131764 47806 131816 47812
rect 131776 44742 131804 47806
rect 131764 44736 131816 44742
rect 131764 44678 131816 44684
rect 131960 44590 131988 48078
rect 457732 47705 457760 52226
rect 457904 52148 457956 52154
rect 457904 52090 457956 52096
rect 457916 47977 457944 52090
rect 458088 52012 458140 52018
rect 458088 51954 458140 51960
rect 458100 48249 458128 51954
rect 458272 50516 458324 50522
rect 458272 50458 458324 50464
rect 458086 48240 458142 48249
rect 458086 48175 458142 48184
rect 457902 47968 457958 47977
rect 457902 47903 457958 47912
rect 457718 47696 457774 47705
rect 457718 47631 457774 47640
rect 458284 46889 458312 50458
rect 458456 50380 458508 50386
rect 458456 50322 458508 50328
rect 458270 46880 458326 46889
rect 458270 46815 458326 46824
rect 142370 46702 142660 46730
rect 131948 44584 132000 44590
rect 131948 44526 132000 44532
rect 132592 44328 132644 44334
rect 132590 44296 132592 44305
rect 142632 44305 142660 46702
rect 458468 46617 458496 50322
rect 459020 47433 459048 52686
rect 459296 52578 459324 52686
rect 463608 52692 463660 52698
rect 463608 52634 463660 52640
rect 463620 52578 463648 52634
rect 459296 52550 459632 52578
rect 463312 52550 463648 52578
rect 463772 52562 464108 52578
rect 463772 52556 464120 52562
rect 463772 52550 464068 52556
rect 464068 52498 464120 52504
rect 459172 52426 459508 52442
rect 465000 52426 465028 52770
rect 466828 52692 466880 52698
rect 466828 52634 466880 52640
rect 466460 52556 466512 52562
rect 466460 52498 466512 52504
rect 465152 52426 465488 52442
rect 459172 52420 459520 52426
rect 459172 52414 459468 52420
rect 459468 52362 459520 52368
rect 464988 52420 465040 52426
rect 465152 52420 465500 52426
rect 465152 52414 465448 52420
rect 464988 52362 465040 52368
rect 465448 52362 465500 52368
rect 462594 52320 462650 52329
rect 459756 52290 460092 52306
rect 459744 52284 460092 52290
rect 459796 52278 460092 52284
rect 461932 52290 462268 52306
rect 461932 52284 462280 52290
rect 461932 52278 462228 52284
rect 459744 52226 459796 52232
rect 462392 52278 462594 52306
rect 465612 52290 465948 52306
rect 465612 52284 465960 52290
rect 465612 52278 465908 52284
rect 462594 52255 462650 52264
rect 462228 52226 462280 52232
rect 465908 52226 465960 52232
rect 462852 52154 463188 52170
rect 460848 52148 460900 52154
rect 462852 52148 463200 52154
rect 462852 52142 463148 52148
rect 460848 52090 460900 52096
rect 463148 52090 463200 52096
rect 460860 52034 460888 52090
rect 461766 52048 461822 52057
rect 460216 52018 460552 52034
rect 460204 52012 460552 52018
rect 460256 52006 460552 52012
rect 460860 52006 461012 52034
rect 461472 52006 461766 52034
rect 464232 52018 464568 52034
rect 464692 52018 465028 52034
rect 464232 52012 464580 52018
rect 464232 52006 464528 52012
rect 461766 51983 461822 51992
rect 460204 51954 460256 51960
rect 464692 52012 465040 52018
rect 464692 52006 464988 52012
rect 464528 51954 464580 51960
rect 464988 51954 465040 51960
rect 466472 51474 466500 52498
rect 466642 52320 466698 52329
rect 466642 52255 466698 52264
rect 466656 51649 466684 52255
rect 466642 51640 466698 51649
rect 466642 51575 466698 51584
rect 466460 51468 466512 51474
rect 466460 51410 466512 51416
rect 466840 50930 466868 52634
rect 467024 51066 467052 52770
rect 475384 52420 475436 52426
rect 475384 52362 475436 52368
rect 475568 52420 475620 52426
rect 475568 52362 475620 52368
rect 475396 51950 475424 52362
rect 475200 51944 475252 51950
rect 475200 51886 475252 51892
rect 475384 51944 475436 51950
rect 475384 51886 475436 51892
rect 475212 51474 475240 51886
rect 475200 51468 475252 51474
rect 475200 51410 475252 51416
rect 475580 51338 475608 52362
rect 475568 51332 475620 51338
rect 475568 51274 475620 51280
rect 467012 51060 467064 51066
rect 467012 51002 467064 51008
rect 466828 50924 466880 50930
rect 466828 50866 466880 50872
rect 544028 50386 544056 53108
rect 545684 53094 546020 53122
rect 547892 53094 548044 53122
rect 521108 50380 521160 50386
rect 521108 50322 521160 50328
rect 544016 50380 544068 50386
rect 544016 50322 544068 50328
rect 467012 49428 467064 49434
rect 467012 49370 467064 49376
rect 466644 49292 466696 49298
rect 466644 49234 466696 49240
rect 466460 49156 466512 49162
rect 466460 49098 466512 49104
rect 466472 48249 466500 49098
rect 466458 48240 466514 48249
rect 466458 48175 466514 48184
rect 466656 47977 466684 49234
rect 466828 49020 466880 49026
rect 466828 48962 466880 48968
rect 466642 47968 466698 47977
rect 466642 47903 466698 47912
rect 466840 47705 466868 48962
rect 466826 47696 466882 47705
rect 459172 47654 459232 47682
rect 459632 47654 459968 47682
rect 460092 47654 460152 47682
rect 460552 47654 460796 47682
rect 459006 47424 459062 47433
rect 459006 47359 459062 47368
rect 458454 46608 458510 46617
rect 458454 46543 458510 46552
rect 431222 44840 431278 44849
rect 431222 44775 431278 44784
rect 132644 44296 132646 44305
rect 132590 44231 132646 44240
rect 142618 44296 142674 44305
rect 142618 44231 142674 44240
rect 307298 44160 307354 44169
rect 307298 44095 307354 44104
rect 131028 43988 131080 43994
rect 131028 43930 131080 43936
rect 187332 43580 187384 43586
rect 187332 43522 187384 43528
rect 43628 42832 43680 42838
rect 43628 42774 43680 42780
rect 187344 42092 187372 43522
rect 194322 42120 194378 42129
rect 194074 42078 194322 42106
rect 307312 42106 307340 44095
rect 419722 43888 419778 43897
rect 419722 43823 419778 43832
rect 415398 43616 415454 43625
rect 415398 43551 415454 43560
rect 310428 42764 310480 42770
rect 310428 42706 310480 42712
rect 310440 42106 310468 42706
rect 415412 42364 415440 43551
rect 419736 42500 419764 43823
rect 431236 43654 431264 44775
rect 431224 43648 431276 43654
rect 439596 43648 439648 43654
rect 431224 43590 431276 43596
rect 439594 43616 439596 43625
rect 441620 43648 441672 43654
rect 439648 43616 439650 43625
rect 439594 43551 439650 43560
rect 441618 43616 441620 43625
rect 441672 43616 441674 43625
rect 441618 43551 441674 43560
rect 431224 42764 431276 42770
rect 431224 42706 431276 42712
rect 456064 42764 456116 42770
rect 456064 42706 456116 42712
rect 404452 42356 404504 42362
rect 404452 42298 404504 42304
rect 405556 42356 405608 42362
rect 405556 42298 405608 42304
rect 420736 42356 420788 42362
rect 420736 42298 420788 42304
rect 427084 42356 427136 42362
rect 427084 42298 427136 42304
rect 307004 42078 307340 42106
rect 310132 42078 310468 42106
rect 194322 42055 194378 42064
rect 361946 41848 362002 41857
rect 361790 41806 361946 41834
rect 365166 41848 365222 41857
rect 364918 41806 365166 41834
rect 361946 41783 362002 41792
rect 365166 41783 365222 41792
rect 404464 41478 404492 42298
rect 405568 42092 405596 42298
rect 416686 42256 416742 42265
rect 416686 42191 416742 42200
rect 416700 42106 416728 42191
rect 416622 42078 416728 42106
rect 420748 41478 420776 42298
rect 427096 41478 427124 42298
rect 431236 42090 431264 42706
rect 446402 42256 446458 42265
rect 446402 42191 446458 42200
rect 431224 42084 431276 42090
rect 431224 42026 431276 42032
rect 446416 41585 446444 42191
rect 456076 42090 456104 42706
rect 456064 42084 456116 42090
rect 456064 42026 456116 42032
rect 446402 41576 446458 41585
rect 446402 41511 446458 41520
rect 459204 41478 459232 47654
rect 459940 42106 459968 47654
rect 460124 44849 460152 47654
rect 460110 44840 460166 44849
rect 460110 44775 460166 44784
rect 460768 43353 460796 47654
rect 460998 47410 461026 47668
rect 461458 47410 461486 47668
rect 460952 47382 461026 47410
rect 461412 47382 461486 47410
rect 461596 47654 461932 47682
rect 462392 47654 462728 47682
rect 462852 47654 462912 47682
rect 460754 43344 460810 43353
rect 460754 43279 460810 43288
rect 460952 42401 460980 47382
rect 461412 42945 461440 47382
rect 461596 43625 461624 47654
rect 462700 43625 462728 47654
rect 462884 43897 462912 47654
rect 463068 47654 463312 47682
rect 462870 43888 462926 43897
rect 462870 43823 462926 43832
rect 461582 43616 461638 43625
rect 461582 43551 461638 43560
rect 462686 43616 462742 43625
rect 462686 43551 462742 43560
rect 461398 42936 461454 42945
rect 461398 42871 461454 42880
rect 463068 42770 463096 47654
rect 463758 47410 463786 47668
rect 463712 47382 463786 47410
rect 463896 47654 464232 47682
rect 464692 47654 464752 47682
rect 463712 44441 463740 47382
rect 463698 44432 463754 44441
rect 463698 44367 463754 44376
rect 463896 44169 463924 47654
rect 464724 44305 464752 47654
rect 465138 47410 465166 47668
rect 465092 47382 465166 47410
rect 465276 47654 465612 47682
rect 465092 46889 465120 47382
rect 465078 46880 465134 46889
rect 465078 46815 465134 46824
rect 465276 46617 465304 47654
rect 466826 47631 466882 47640
rect 467024 47433 467052 49370
rect 467010 47424 467066 47433
rect 467010 47359 467066 47368
rect 521120 47025 521148 50322
rect 545684 49473 545712 53094
rect 545670 49464 545726 49473
rect 545670 49399 545726 49408
rect 547892 47569 547920 53094
rect 550008 48929 550036 53108
rect 549994 48920 550050 48929
rect 549994 48855 550050 48864
rect 552032 47841 552060 53108
rect 553688 53094 554024 53122
rect 576124 53100 576176 53106
rect 553688 49201 553716 53094
rect 576124 53042 576176 53048
rect 572076 52284 572128 52290
rect 572076 52226 572128 52232
rect 571708 52080 571760 52086
rect 571708 52022 571760 52028
rect 571720 51474 571748 52022
rect 572088 51950 572116 52226
rect 576136 52154 576164 53042
rect 576124 52148 576176 52154
rect 576124 52090 576176 52096
rect 576308 52148 576360 52154
rect 576308 52090 576360 52096
rect 572076 51944 572128 51950
rect 572076 51886 572128 51892
rect 571708 51468 571760 51474
rect 571708 51410 571760 51416
rect 576320 51338 576348 52090
rect 576308 51332 576360 51338
rect 576308 51274 576360 51280
rect 577516 49434 577544 97242
rect 577700 52426 577728 97378
rect 579252 95192 579304 95198
rect 579252 95134 579304 95140
rect 579264 95033 579292 95134
rect 579250 95024 579306 95033
rect 579250 94959 579306 94968
rect 579448 93854 579476 105130
rect 579448 93826 579568 93854
rect 579344 93152 579396 93158
rect 579342 93120 579344 93129
rect 579396 93120 579398 93129
rect 579342 93055 579398 93064
rect 578240 91860 578292 91866
rect 578240 91802 578292 91808
rect 578252 90953 578280 91802
rect 578238 90944 578294 90953
rect 578238 90879 578294 90888
rect 579344 88324 579396 88330
rect 579344 88266 579396 88272
rect 579356 88097 579384 88266
rect 579342 88088 579398 88097
rect 579342 88023 579398 88032
rect 578792 86488 578844 86494
rect 578790 86456 578792 86465
rect 578844 86456 578846 86465
rect 578790 86391 578846 86400
rect 579344 84040 579396 84046
rect 579342 84008 579344 84017
rect 579396 84008 579398 84017
rect 579342 83943 579398 83952
rect 578700 82816 578752 82822
rect 578700 82758 578752 82764
rect 578712 82249 578740 82758
rect 578698 82240 578754 82249
rect 578698 82175 578754 82184
rect 578884 82136 578936 82142
rect 578884 82078 578936 82084
rect 578608 78260 578660 78266
rect 578608 78202 578660 78208
rect 578620 77897 578648 78202
rect 578606 77888 578662 77897
rect 578606 77823 578662 77832
rect 578700 77240 578752 77246
rect 578700 77182 578752 77188
rect 578712 74534 578740 77182
rect 578896 75721 578924 82078
rect 579540 80073 579568 93826
rect 579526 80064 579582 80073
rect 579526 79999 579582 80008
rect 580276 78266 580304 106286
rect 580460 99346 580488 122062
rect 580644 108730 580672 125598
rect 580632 108724 580684 108730
rect 580632 108666 580684 108672
rect 580448 99340 580500 99346
rect 580448 99282 580500 99288
rect 580632 98660 580684 98666
rect 580632 98602 580684 98608
rect 580644 86494 580672 98602
rect 581656 97986 581684 228346
rect 592696 220114 592724 245618
rect 621664 241528 621716 241534
rect 621664 241470 621716 241476
rect 619640 225004 619692 225010
rect 619640 224946 619692 224952
rect 598388 224664 598440 224670
rect 598388 224606 598440 224612
rect 593970 222320 594026 222329
rect 593970 222255 594026 222264
rect 592684 220108 592736 220114
rect 592684 220050 592736 220056
rect 582564 220040 582616 220046
rect 582378 220008 582434 220017
rect 582378 219943 582434 219952
rect 582562 220008 582564 220017
rect 582616 220008 582618 220017
rect 582562 219943 582618 219952
rect 582392 219858 582420 219943
rect 582392 219830 582788 219858
rect 582378 219736 582434 219745
rect 582760 219722 582788 219830
rect 582760 219694 582972 219722
rect 582378 219671 582434 219680
rect 582392 219586 582420 219671
rect 582392 219558 582512 219586
rect 582484 219366 582512 219558
rect 582472 219360 582524 219366
rect 582472 219302 582524 219308
rect 582380 218884 582432 218890
rect 582380 218826 582432 218832
rect 582392 218482 582420 218826
rect 582380 218476 582432 218482
rect 582380 218418 582432 218424
rect 582380 217252 582432 217258
rect 582380 217194 582432 217200
rect 582392 216753 582420 217194
rect 582564 216776 582616 216782
rect 582378 216744 582434 216753
rect 582378 216679 582434 216688
rect 582562 216744 582564 216753
rect 582616 216744 582618 216753
rect 582562 216679 582618 216688
rect 582944 216209 582972 219694
rect 583114 219464 583170 219473
rect 583114 219399 583170 219408
rect 583128 219230 583156 219399
rect 583116 219224 583168 219230
rect 583116 219166 583168 219172
rect 591580 217524 591632 217530
rect 591580 217466 591632 217472
rect 591592 217025 591620 217466
rect 591762 217288 591818 217297
rect 591762 217223 591818 217232
rect 591946 217288 592002 217297
rect 591946 217223 591948 217232
rect 591776 217122 591804 217223
rect 592000 217223 592002 217232
rect 591948 217194 592000 217200
rect 591764 217116 591816 217122
rect 591764 217058 591816 217064
rect 591578 217016 591634 217025
rect 591946 217016 592002 217025
rect 591578 216951 591634 216960
rect 591776 216974 591946 217002
rect 591776 216481 591804 216974
rect 591946 216951 592002 216960
rect 591762 216472 591818 216481
rect 591762 216407 591818 216416
rect 582930 216200 582986 216209
rect 582930 216135 582986 216144
rect 593984 210202 594012 222255
rect 594798 219736 594854 219745
rect 594798 219671 594854 219680
rect 594812 210202 594840 219671
rect 596824 219360 596876 219366
rect 596824 219302 596876 219308
rect 595902 218920 595958 218929
rect 595902 218855 595904 218864
rect 595956 218855 595958 218864
rect 596086 218920 596142 218929
rect 596086 218855 596142 218864
rect 595904 218826 595956 218832
rect 596100 218482 596128 218855
rect 596088 218476 596140 218482
rect 596088 218418 596140 218424
rect 594984 218204 595036 218210
rect 594984 218146 595036 218152
rect 594996 217326 595024 218146
rect 595720 217524 595772 217530
rect 595720 217466 595772 217472
rect 594984 217320 595036 217326
rect 594984 217262 595036 217268
rect 595168 217116 595220 217122
rect 595168 217058 595220 217064
rect 595180 210202 595208 217058
rect 595732 210202 595760 217466
rect 596270 216608 596326 216617
rect 596270 216543 596326 216552
rect 596284 210202 596312 216543
rect 596836 210202 596864 219302
rect 597560 218884 597612 218890
rect 597560 218826 597612 218832
rect 597572 217598 597600 218826
rect 597560 217592 597612 217598
rect 597560 217534 597612 217540
rect 597558 217152 597614 217161
rect 597558 217087 597614 217096
rect 597572 210202 597600 217087
rect 597926 216336 597982 216345
rect 597926 216271 597982 216280
rect 597940 210202 597968 216271
rect 598400 210202 598428 224606
rect 606758 224496 606814 224505
rect 606758 224431 606814 224440
rect 606772 223961 606800 224431
rect 617154 224224 617210 224233
rect 617154 224159 617210 224168
rect 615500 224052 615552 224058
rect 615500 223994 615552 224000
rect 606758 223952 606814 223961
rect 606758 223887 606814 223896
rect 611634 223680 611690 223689
rect 611634 223615 611690 223624
rect 600686 222048 600742 222057
rect 600686 221983 600742 221992
rect 604460 222012 604512 222018
rect 599030 221776 599086 221785
rect 599030 221711 599086 221720
rect 599044 214470 599072 221711
rect 599214 220960 599270 220969
rect 599214 220895 599270 220904
rect 599032 214464 599084 214470
rect 599032 214406 599084 214412
rect 599228 210202 599256 220895
rect 600412 220856 600464 220862
rect 600412 220798 600464 220804
rect 600424 214470 600452 220798
rect 599584 214464 599636 214470
rect 599584 214406 599636 214412
rect 600412 214464 600464 214470
rect 600412 214406 600464 214412
rect 599596 210202 599624 214406
rect 600504 214328 600556 214334
rect 600504 214270 600556 214276
rect 600516 210202 600544 214270
rect 593984 210174 594412 210202
rect 594812 210174 594964 210202
rect 595180 210174 595516 210202
rect 595732 210174 596068 210202
rect 596284 210174 596620 210202
rect 596836 210174 597172 210202
rect 597572 210174 597724 210202
rect 597940 210174 598276 210202
rect 598400 210174 598828 210202
rect 599228 210174 599380 210202
rect 599596 210174 599932 210202
rect 600484 210174 600544 210202
rect 600700 210066 600728 221983
rect 604460 221954 604512 221960
rect 603080 221604 603132 221610
rect 603080 221546 603132 221552
rect 601974 221504 602030 221513
rect 601974 221439 602030 221448
rect 600870 221232 600926 221241
rect 600870 221167 600926 221176
rect 600884 214334 600912 221167
rect 601792 220992 601844 220998
rect 601792 220934 601844 220940
rect 601240 214464 601292 214470
rect 601240 214406 601292 214412
rect 600872 214328 600924 214334
rect 600872 214270 600924 214276
rect 601252 210202 601280 214406
rect 601804 212430 601832 220934
rect 601792 212424 601844 212430
rect 601792 212366 601844 212372
rect 601988 210202 602016 221439
rect 603092 212430 603120 221546
rect 603356 221264 603408 221270
rect 603356 221206 603408 221212
rect 603368 212534 603396 221206
rect 603540 221128 603592 221134
rect 603540 221070 603592 221076
rect 603552 215294 603580 221070
rect 603276 212506 603396 212534
rect 603460 215266 603580 215294
rect 602344 212424 602396 212430
rect 602344 212366 602396 212372
rect 603080 212424 603132 212430
rect 603080 212366 603132 212372
rect 602356 210202 602384 212366
rect 603276 211070 603304 212506
rect 603264 211064 603316 211070
rect 603264 211006 603316 211012
rect 603460 210882 603488 215266
rect 604472 212430 604500 221954
rect 607220 221740 607272 221746
rect 607220 221682 607272 221688
rect 604642 220280 604698 220289
rect 604642 220215 604698 220224
rect 604000 212424 604052 212430
rect 604000 212366 604052 212372
rect 604460 212424 604512 212430
rect 604460 212366 604512 212372
rect 603632 211064 603684 211070
rect 603632 211006 603684 211012
rect 603276 210854 603488 210882
rect 603276 210202 603304 210854
rect 601252 210174 601588 210202
rect 601988 210174 602140 210202
rect 602356 210174 602692 210202
rect 603244 210174 603304 210202
rect 603644 210202 603672 211006
rect 604012 210202 604040 212366
rect 604656 210202 604684 220215
rect 605840 219904 605892 219910
rect 605840 219846 605892 219852
rect 605102 218648 605158 218657
rect 605102 218583 605158 218592
rect 605116 217734 605144 218583
rect 605104 217728 605156 217734
rect 605104 217670 605156 217676
rect 605104 212424 605156 212430
rect 605104 212366 605156 212372
rect 605116 210202 605144 212366
rect 603644 210174 603796 210202
rect 604012 210174 604348 210202
rect 604656 210174 604900 210202
rect 605116 210174 605452 210202
rect 605852 210118 605880 219846
rect 606668 219632 606720 219638
rect 606668 219574 606720 219580
rect 606024 219496 606076 219502
rect 606024 219438 606076 219444
rect 606036 215294 606064 219438
rect 605944 215266 606064 215294
rect 605944 210202 605972 215266
rect 606680 210202 606708 219574
rect 607232 210202 607260 221682
rect 611360 220652 611412 220658
rect 611360 220594 611412 220600
rect 610532 220516 610584 220522
rect 610532 220458 610584 220464
rect 608692 220380 608744 220386
rect 608692 220322 608744 220328
rect 607772 219768 607824 219774
rect 607772 219710 607824 219716
rect 607784 210202 607812 219710
rect 608704 210202 608732 220322
rect 609428 220244 609480 220250
rect 609428 220186 609480 220192
rect 608966 217832 609022 217841
rect 608966 217767 609022 217776
rect 608980 210202 609008 217767
rect 609440 210202 609468 220186
rect 610070 217560 610126 217569
rect 610070 217495 610126 217504
rect 610084 210202 610112 217495
rect 610544 210202 610572 220458
rect 611372 210202 611400 220594
rect 611648 210202 611676 223615
rect 611820 218748 611872 218754
rect 611820 218690 611872 218696
rect 611832 217462 611860 218690
rect 613016 218204 613068 218210
rect 613016 218146 613068 218152
rect 611820 217456 611872 217462
rect 611820 217398 611872 217404
rect 612280 215144 612332 215150
rect 612280 215086 612332 215092
rect 612292 210202 612320 215086
rect 612830 213208 612886 213217
rect 612830 213143 612886 213152
rect 612844 210202 612872 213143
rect 613028 212906 613056 218146
rect 614488 218000 614540 218006
rect 614488 217942 614540 217948
rect 614120 217728 614172 217734
rect 614120 217670 614172 217676
rect 613384 217592 613436 217598
rect 613384 217534 613436 217540
rect 613016 212900 613068 212906
rect 613016 212842 613068 212848
rect 613396 210202 613424 217534
rect 614132 210202 614160 217670
rect 614500 210202 614528 217942
rect 615512 214470 615540 223994
rect 616880 223916 616932 223922
rect 616880 223858 616932 223864
rect 615682 220280 615738 220289
rect 615682 220215 615738 220224
rect 615500 214464 615552 214470
rect 615500 214406 615552 214412
rect 615040 212900 615092 212906
rect 615040 212842 615092 212848
rect 615052 210202 615080 212842
rect 615696 210202 615724 220215
rect 616892 214606 616920 223858
rect 616880 214600 616932 214606
rect 616880 214542 616932 214548
rect 616144 214464 616196 214470
rect 616144 214406 616196 214412
rect 616156 210202 616184 214406
rect 617168 210202 617196 224159
rect 618260 223032 618312 223038
rect 618260 222974 618312 222980
rect 617706 220552 617762 220561
rect 617706 220487 617762 220496
rect 617340 214600 617392 214606
rect 617340 214542 617392 214548
rect 605944 210174 606004 210202
rect 606680 210174 607108 210202
rect 607232 210174 607660 210202
rect 607784 210174 608212 210202
rect 608704 210174 608764 210202
rect 608980 210174 609316 210202
rect 609440 210174 609868 210202
rect 610084 210174 610420 210202
rect 610544 210174 610972 210202
rect 611372 210174 611524 210202
rect 611648 210174 612076 210202
rect 612292 210174 612628 210202
rect 612844 210174 613180 210202
rect 613396 210174 613732 210202
rect 614132 210174 614284 210202
rect 614500 210174 614836 210202
rect 615052 210174 615388 210202
rect 615696 210174 615940 210202
rect 616156 210174 616492 210202
rect 617044 210174 617196 210202
rect 617352 210202 617380 214542
rect 617720 210202 617748 220487
rect 618272 210202 618300 222974
rect 618810 219464 618866 219473
rect 618810 219399 618866 219408
rect 618824 210202 618852 219399
rect 619652 214606 619680 224946
rect 620008 222488 620060 222494
rect 620008 222430 620060 222436
rect 619824 222352 619876 222358
rect 619824 222294 619876 222300
rect 619640 214600 619692 214606
rect 619640 214542 619692 214548
rect 619836 210202 619864 222294
rect 617352 210174 617596 210202
rect 617720 210174 618148 210202
rect 618272 210174 618700 210202
rect 618824 210174 619252 210202
rect 619804 210174 619864 210202
rect 620020 210202 620048 222430
rect 621676 214878 621704 241470
rect 625252 224528 625304 224534
rect 625252 224470 625304 224476
rect 622400 223780 622452 223786
rect 622400 223722 622452 223728
rect 621848 215008 621900 215014
rect 621848 214950 621900 214956
rect 621112 214872 621164 214878
rect 621112 214814 621164 214820
rect 621664 214872 621716 214878
rect 621664 214814 621716 214820
rect 620560 214600 620612 214606
rect 620560 214542 620612 214548
rect 620572 210202 620600 214542
rect 621124 210202 621152 214814
rect 621860 210202 621888 214950
rect 620020 210174 620356 210202
rect 620572 210174 620908 210202
rect 621124 210174 621460 210202
rect 621860 210174 622012 210202
rect 622412 210118 622440 223722
rect 622584 222760 622636 222766
rect 622584 222702 622636 222708
rect 622596 214606 622624 222702
rect 622768 222624 622820 222630
rect 622768 222566 622820 222572
rect 622584 214600 622636 214606
rect 622584 214542 622636 214548
rect 622780 210202 622808 222566
rect 623778 219192 623834 219201
rect 623778 219127 623834 219136
rect 622950 218648 623006 218657
rect 622950 218583 623006 218592
rect 622964 216102 622992 218583
rect 622952 216096 623004 216102
rect 622952 216038 623004 216044
rect 623792 214606 623820 219127
rect 624424 214736 624476 214742
rect 624424 214678 624476 214684
rect 623320 214600 623372 214606
rect 623320 214542 623372 214548
rect 623780 214600 623832 214606
rect 623780 214542 623832 214548
rect 622564 210174 622808 210202
rect 623332 210202 623360 214542
rect 623872 214464 623924 214470
rect 623872 214406 623924 214412
rect 623884 210202 623912 214406
rect 624436 210202 624464 214678
rect 625264 214606 625292 224470
rect 625436 224392 625488 224398
rect 625436 224334 625488 224340
rect 625252 214600 625304 214606
rect 625252 214542 625304 214548
rect 625448 210202 625476 224334
rect 630954 223952 631010 223961
rect 630954 223887 631010 223896
rect 626540 223644 626592 223650
rect 626540 223586 626592 223592
rect 626080 217320 626132 217326
rect 626080 217262 626132 217268
rect 625620 214600 625672 214606
rect 625620 214542 625672 214548
rect 623332 210174 623668 210202
rect 623884 210174 624220 210202
rect 624436 210174 624772 210202
rect 625324 210174 625476 210202
rect 625632 210202 625660 214542
rect 626092 210202 626120 217262
rect 626552 210202 626580 223586
rect 627092 222216 627144 222222
rect 627092 222158 627144 222164
rect 627104 210202 627132 222158
rect 630678 218920 630734 218929
rect 630678 218855 630734 218864
rect 629390 218104 629446 218113
rect 629390 218039 629446 218048
rect 628288 217456 628340 217462
rect 628288 217398 628340 217404
rect 627826 216880 627882 216889
rect 627826 216815 627882 216824
rect 627840 212650 627868 216815
rect 627840 212622 628052 212650
rect 628024 210202 628052 212622
rect 628300 210202 628328 217398
rect 628840 215960 628892 215966
rect 628840 215902 628892 215908
rect 628852 210202 628880 215902
rect 629404 210202 629432 218039
rect 629944 216096 629996 216102
rect 629944 216038 629996 216044
rect 629956 210202 629984 216038
rect 630692 210202 630720 218855
rect 630968 210202 630996 223887
rect 631600 214464 631652 214470
rect 631600 214406 631652 214412
rect 631612 210202 631640 214406
rect 632716 212770 632744 246298
rect 647252 242214 647280 277766
rect 648724 277394 648752 277780
rect 648632 277366 648752 277394
rect 648632 261662 648660 277366
rect 648620 261656 648672 261662
rect 648620 261598 648672 261604
rect 647240 242208 647292 242214
rect 647240 242150 647292 242156
rect 639602 230072 639658 230081
rect 639602 230007 639658 230016
rect 633716 227044 633768 227050
rect 633716 226986 633768 226992
rect 633440 220108 633492 220114
rect 633440 220050 633492 220056
rect 632888 214872 632940 214878
rect 632888 214814 632940 214820
rect 632704 212764 632756 212770
rect 632704 212706 632756 212712
rect 632900 210202 632928 214814
rect 633452 210202 633480 220050
rect 633728 210202 633756 226986
rect 636476 220108 636528 220114
rect 636476 220050 636528 220056
rect 636292 214600 636344 214606
rect 636292 214542 636344 214548
rect 635556 213512 635608 213518
rect 635556 213454 635608 213460
rect 634360 212764 634412 212770
rect 634360 212706 634412 212712
rect 634372 210202 634400 212706
rect 635568 210202 635596 213454
rect 625632 210174 625876 210202
rect 626092 210174 626428 210202
rect 626552 210174 626980 210202
rect 627104 210174 627532 210202
rect 628024 210174 628084 210202
rect 628300 210174 628636 210202
rect 628852 210174 629188 210202
rect 629404 210174 629740 210202
rect 629956 210174 630292 210202
rect 630692 210174 630844 210202
rect 630968 210174 631396 210202
rect 631612 210174 631948 210202
rect 632900 210174 633052 210202
rect 633452 210174 633604 210202
rect 633728 210174 634156 210202
rect 634372 210174 634708 210202
rect 635260 210174 635596 210202
rect 636304 210202 636332 214542
rect 636488 210202 636516 220050
rect 639616 214606 639644 230007
rect 650642 225584 650698 225593
rect 650642 225519 650698 225528
rect 649722 221504 649778 221513
rect 649722 221439 649778 221448
rect 644754 220416 644810 220425
rect 644754 220351 644810 220360
rect 643834 218920 643890 218929
rect 643834 218855 643890 218864
rect 640614 218648 640670 218657
rect 640614 218583 640670 218592
rect 639970 217832 640026 217841
rect 639970 217767 640026 217776
rect 639604 214600 639656 214606
rect 639604 214542 639656 214548
rect 638316 213920 638368 213926
rect 638316 213862 638368 213868
rect 638328 210202 638356 213862
rect 638868 213376 638920 213382
rect 638868 213318 638920 213324
rect 638880 210202 638908 213318
rect 639984 210202 640012 217767
rect 640628 213926 640656 218583
rect 643006 215928 643062 215937
rect 643006 215863 643062 215872
rect 640616 213920 640668 213926
rect 640616 213862 640668 213868
rect 641628 213784 641680 213790
rect 641628 213726 641680 213732
rect 640248 213648 640300 213654
rect 640248 213590 640300 213596
rect 640260 210202 640288 213590
rect 641640 210202 641668 213726
rect 642180 213240 642232 213246
rect 642180 213182 642232 213188
rect 642192 210202 642220 213182
rect 643020 210202 643048 215863
rect 643848 210202 643876 218855
rect 644570 217560 644626 217569
rect 644570 217495 644626 217504
rect 636304 210174 636364 210202
rect 636488 210174 636916 210202
rect 638020 210174 638356 210202
rect 638572 210174 638908 210202
rect 639676 210174 640012 210202
rect 640228 210174 640288 210202
rect 641332 210174 641668 210202
rect 641884 210174 642220 210202
rect 642988 210174 643048 210202
rect 643540 210174 643876 210202
rect 644584 210202 644612 217495
rect 644768 210202 644796 220351
rect 648618 219872 648674 219881
rect 648618 219807 648674 219816
rect 648252 218068 648304 218074
rect 648252 218010 648304 218016
rect 646594 216200 646650 216209
rect 646594 216135 646650 216144
rect 646608 210202 646636 216135
rect 647146 213208 647202 213217
rect 647146 213143 647202 213152
rect 647160 210202 647188 213143
rect 648264 210202 648292 218010
rect 648436 214736 648488 214742
rect 648436 214678 648488 214684
rect 644584 210174 644644 210202
rect 644768 210174 645196 210202
rect 646300 210174 646636 210202
rect 646852 210174 647188 210202
rect 647956 210174 648292 210202
rect 648448 210202 648476 214678
rect 648632 213926 648660 219807
rect 648620 213920 648672 213926
rect 648620 213862 648672 213868
rect 649264 213920 649316 213926
rect 649264 213862 649316 213868
rect 649276 210202 649304 213862
rect 649736 213654 649764 221439
rect 650460 213920 650512 213926
rect 650460 213862 650512 213868
rect 649724 213648 649776 213654
rect 649724 213590 649776 213596
rect 650472 210202 650500 213862
rect 650656 213790 650684 225519
rect 651286 219192 651342 219201
rect 651286 219127 651342 219136
rect 650644 213784 650696 213790
rect 650644 213726 650696 213732
rect 651300 210202 651328 219127
rect 651840 213648 651892 213654
rect 651840 213590 651892 213596
rect 651852 210202 651880 213590
rect 648448 210174 648508 210202
rect 649276 210174 649612 210202
rect 650164 210174 650500 210202
rect 651268 210174 651328 210202
rect 651820 210174 651880 210202
rect 605840 210112 605892 210118
rect 600700 210038 601036 210066
rect 605840 210054 605892 210060
rect 606208 210112 606260 210118
rect 622400 210112 622452 210118
rect 606260 210060 606556 210066
rect 606208 210054 606556 210060
rect 622400 210054 622452 210060
rect 622768 210112 622820 210118
rect 622820 210060 623116 210066
rect 622768 210054 623116 210060
rect 606220 210038 606556 210054
rect 622780 210038 623116 210054
rect 652036 209574 652064 338263
rect 652206 298480 652262 298489
rect 652206 298415 652262 298424
rect 652220 209710 652248 298415
rect 658936 233889 658964 390526
rect 659120 360097 659148 510614
rect 660316 411913 660344 550598
rect 661696 491609 661724 603094
rect 663076 535537 663104 656882
rect 664456 580145 664484 709310
rect 665836 626113 665864 749362
rect 666296 711657 666324 778359
rect 666480 755177 666508 879135
rect 668398 876344 668454 876353
rect 668398 876279 668454 876288
rect 667204 803208 667256 803214
rect 667204 803150 667256 803156
rect 666466 755168 666522 755177
rect 666466 755103 666522 755112
rect 666466 745512 666522 745521
rect 666466 745447 666522 745456
rect 666282 711648 666338 711657
rect 666282 711583 666338 711592
rect 666282 688664 666338 688673
rect 666282 688599 666338 688608
rect 665822 626104 665878 626113
rect 665822 626039 665878 626048
rect 666296 621217 666324 688599
rect 666480 665417 666508 745447
rect 667216 671129 667244 803150
rect 667846 780736 667902 780745
rect 667846 780671 667902 780680
rect 667662 742520 667718 742529
rect 667662 742455 667718 742464
rect 667202 671120 667258 671129
rect 667202 671055 667258 671064
rect 667676 665961 667704 742455
rect 667860 710297 667888 780671
rect 668412 754225 668440 876279
rect 669042 872536 669098 872545
rect 669042 872471 669098 872480
rect 668584 789404 668636 789410
rect 668584 789346 668636 789352
rect 668398 754216 668454 754225
rect 668398 754151 668454 754160
rect 668400 742756 668452 742762
rect 668400 742698 668452 742704
rect 668412 735321 668440 742698
rect 668398 735312 668454 735321
rect 668398 735247 668454 735256
rect 668214 731504 668270 731513
rect 668214 731439 668270 731448
rect 667846 710288 667902 710297
rect 667846 710223 667902 710232
rect 667846 705120 667902 705129
rect 667846 705055 667902 705064
rect 667662 665952 667718 665961
rect 667662 665887 667718 665896
rect 666466 665408 666522 665417
rect 666466 665343 666522 665352
rect 667204 628584 667256 628590
rect 667204 628526 667256 628532
rect 666282 621208 666338 621217
rect 666282 621143 666338 621152
rect 667018 593464 667074 593473
rect 667018 593399 667074 593408
rect 665824 590708 665876 590714
rect 665824 590650 665876 590656
rect 664442 580136 664498 580145
rect 664442 580071 664498 580080
rect 664444 576904 664496 576910
rect 664444 576846 664496 576852
rect 663062 535528 663118 535537
rect 663062 535463 663118 535472
rect 661868 523048 661920 523054
rect 661868 522990 661920 522996
rect 661682 491600 661738 491609
rect 661682 491535 661738 491544
rect 661684 456816 661736 456822
rect 661684 456758 661736 456764
rect 660302 411904 660358 411913
rect 660302 411839 660358 411848
rect 660304 378208 660356 378214
rect 660304 378150 660356 378156
rect 659106 360088 659162 360097
rect 659106 360023 659162 360032
rect 660316 234161 660344 378150
rect 661696 313585 661724 456758
rect 661880 406337 661908 522990
rect 663248 494760 663300 494766
rect 664456 494737 664484 576846
rect 663248 494702 663300 494708
rect 664442 494728 664498 494737
rect 663064 416832 663116 416838
rect 663064 416774 663116 416780
rect 661866 406328 661922 406337
rect 661866 406263 661922 406272
rect 661868 364404 661920 364410
rect 661868 364346 661920 364352
rect 661682 313576 661738 313585
rect 661682 313511 661738 313520
rect 660302 234152 660358 234161
rect 660302 234087 660358 234096
rect 658922 233880 658978 233889
rect 658922 233815 658978 233824
rect 661880 232558 661908 364346
rect 663076 268161 663104 416774
rect 663260 358601 663288 494702
rect 664442 494663 664498 494672
rect 665836 492153 665864 590650
rect 667032 528601 667060 593399
rect 667216 535265 667244 628526
rect 667662 603392 667718 603401
rect 667662 603327 667718 603336
rect 667386 564496 667442 564505
rect 667386 564431 667442 564440
rect 667202 535256 667258 535265
rect 667202 535191 667258 535200
rect 667018 528592 667074 528601
rect 667018 528527 667074 528536
rect 665822 492144 665878 492153
rect 665822 492079 665878 492088
rect 667400 485217 667428 564431
rect 667676 529961 667704 603327
rect 667662 529952 667718 529961
rect 667662 529887 667718 529896
rect 667386 485208 667442 485217
rect 667386 485143 667442 485152
rect 667204 484424 667256 484430
rect 667204 484366 667256 484372
rect 665824 470620 665876 470626
rect 665824 470562 665876 470568
rect 664444 404388 664496 404394
rect 664444 404330 664496 404336
rect 663246 358592 663302 358601
rect 663246 358527 663302 358536
rect 664456 271153 664484 404330
rect 665836 315489 665864 470562
rect 667216 360913 667244 484366
rect 667860 456249 667888 705055
rect 668030 693288 668086 693297
rect 668030 693223 668086 693232
rect 668044 619993 668072 693223
rect 668228 664193 668256 731439
rect 668400 669384 668452 669390
rect 668596 669361 668624 789346
rect 668768 775600 668820 775606
rect 668768 775542 668820 775548
rect 668780 742762 668808 775542
rect 669056 755449 669084 872471
rect 669042 755440 669098 755449
rect 669042 755375 669098 755384
rect 668768 742756 668820 742762
rect 668768 742698 668820 742704
rect 668858 738304 668914 738313
rect 668858 738239 668914 738248
rect 668872 731414 668900 738239
rect 669042 733816 669098 733825
rect 669042 733751 669098 733760
rect 668872 731386 668992 731414
rect 668766 730552 668822 730561
rect 668766 730487 668822 730496
rect 668400 669326 668452 669332
rect 668582 669352 668638 669361
rect 668214 664184 668270 664193
rect 668214 664119 668270 664128
rect 668412 643929 668440 669326
rect 668582 669287 668638 669296
rect 668780 666233 668808 730487
rect 668766 666224 668822 666233
rect 668766 666159 668822 666168
rect 668964 661745 668992 731386
rect 669056 673454 669084 733751
rect 669240 728249 669268 929455
rect 670606 928296 670662 928305
rect 670606 928231 670662 928240
rect 669778 864240 669834 864249
rect 669778 864175 669834 864184
rect 669792 750961 669820 864175
rect 669964 841832 670016 841838
rect 669964 841774 670016 841780
rect 669778 750952 669834 750961
rect 669778 750887 669834 750896
rect 669594 737080 669650 737089
rect 669594 737015 669650 737024
rect 669226 728240 669282 728249
rect 669226 728175 669282 728184
rect 669056 673426 669176 673454
rect 668950 661736 669006 661745
rect 668950 661671 669006 661680
rect 669148 661337 669176 673426
rect 669608 662017 669636 737015
rect 669778 730144 669834 730153
rect 669778 730079 669834 730088
rect 669594 662008 669650 662017
rect 669594 661943 669650 661952
rect 669134 661328 669190 661337
rect 669134 661263 669190 661272
rect 669792 659705 669820 730079
rect 669976 715737 670004 841774
rect 670422 780056 670478 780065
rect 670422 779991 670478 780000
rect 670436 779634 670464 779991
rect 670436 779606 670556 779634
rect 670330 779512 670386 779521
rect 670330 779447 670386 779456
rect 670146 775704 670202 775713
rect 670146 775639 670202 775648
rect 669962 715728 670018 715737
rect 669962 715663 670018 715672
rect 670160 710025 670188 775639
rect 670344 756254 670372 779447
rect 670528 756254 670556 779606
rect 670252 756226 670372 756254
rect 670436 756226 670556 756254
rect 670252 731414 670280 756226
rect 670436 731414 670464 756226
rect 670252 731386 670372 731414
rect 670436 731386 670556 731414
rect 670146 710016 670202 710025
rect 670146 709951 670202 709960
rect 670344 707985 670372 731386
rect 670330 707976 670386 707985
rect 670330 707911 670386 707920
rect 670528 707169 670556 731386
rect 670620 728906 670648 928231
rect 670790 865328 670846 865337
rect 670790 865263 670846 865272
rect 670804 754905 670832 865263
rect 670988 758713 671016 936391
rect 671986 935776 672042 935785
rect 671986 935711 672042 935720
rect 671344 895688 671396 895694
rect 671344 895630 671396 895636
rect 671158 775024 671214 775033
rect 671158 774959 671214 774968
rect 670974 758704 671030 758713
rect 670974 758639 671030 758648
rect 670974 758296 671030 758305
rect 670974 758231 671030 758240
rect 670790 754896 670846 754905
rect 670790 754831 670846 754840
rect 670620 728878 670832 728906
rect 670804 728657 670832 728878
rect 670790 728648 670846 728657
rect 670790 728583 670846 728592
rect 670790 714912 670846 714921
rect 670790 714847 670846 714856
rect 670514 707160 670570 707169
rect 670514 707095 670570 707104
rect 669964 696992 670016 696998
rect 669964 696934 670016 696940
rect 669778 659696 669834 659705
rect 669778 659631 669834 659640
rect 669226 654256 669282 654265
rect 669226 654191 669282 654200
rect 669042 645552 669098 645561
rect 669042 645487 669098 645496
rect 668398 643920 668454 643929
rect 668398 643855 668454 643864
rect 668584 643136 668636 643142
rect 668584 643078 668636 643084
rect 668030 619984 668086 619993
rect 668030 619919 668086 619928
rect 668398 601760 668454 601769
rect 668398 601695 668454 601704
rect 668412 527377 668440 601695
rect 668596 535945 668624 643078
rect 668858 638752 668914 638761
rect 668858 638687 668914 638696
rect 668872 574433 668900 638687
rect 669056 574841 669084 645487
rect 669042 574832 669098 574841
rect 669042 574767 669098 574776
rect 668858 574424 668914 574433
rect 668858 574359 668914 574368
rect 669240 574161 669268 654191
rect 669778 643512 669834 643521
rect 669778 643447 669834 643456
rect 669594 623928 669650 623937
rect 669594 623863 669650 623872
rect 669608 579057 669636 623863
rect 669594 579048 669650 579057
rect 669594 578983 669650 578992
rect 669594 577824 669650 577833
rect 669594 577759 669650 577768
rect 669226 574152 669282 574161
rect 669226 574087 669282 574096
rect 669042 557560 669098 557569
rect 669042 557495 669098 557504
rect 668582 535936 668638 535945
rect 668582 535871 668638 535880
rect 668398 527368 668454 527377
rect 668398 527303 668454 527312
rect 669056 485897 669084 557495
rect 669226 552664 669282 552673
rect 669226 552599 669282 552608
rect 669042 485888 669098 485897
rect 669042 485823 669098 485832
rect 669240 483993 669268 552599
rect 669412 536852 669464 536858
rect 669412 536794 669464 536800
rect 669226 483984 669282 483993
rect 669226 483919 669282 483928
rect 667846 456240 667902 456249
rect 667846 456175 667902 456184
rect 668584 444440 668636 444446
rect 668584 444382 668636 444388
rect 667202 360904 667258 360913
rect 667202 360839 667258 360848
rect 667204 350600 667256 350606
rect 667204 350542 667256 350548
rect 666652 324352 666704 324358
rect 666652 324294 666704 324300
rect 665822 315480 665878 315489
rect 665822 315415 665878 315424
rect 664442 271144 664498 271153
rect 664442 271079 664498 271088
rect 663062 268152 663118 268161
rect 663062 268087 663118 268096
rect 661868 232552 661920 232558
rect 661868 232494 661920 232500
rect 665088 232212 665140 232218
rect 665088 232154 665140 232160
rect 663798 231840 663854 231849
rect 663798 231775 663854 231784
rect 662050 231160 662106 231169
rect 662050 231095 662106 231104
rect 662236 231124 662288 231130
rect 660946 229800 661002 229809
rect 660946 229735 661002 229744
rect 653402 229120 653458 229129
rect 653402 229055 653458 229064
rect 652390 222864 652446 222873
rect 652390 222799 652446 222808
rect 652404 213518 652432 222799
rect 652942 221232 652998 221241
rect 652942 221167 652998 221176
rect 652760 214600 652812 214606
rect 652760 214542 652812 214548
rect 652392 213512 652444 213518
rect 652392 213454 652444 213460
rect 652772 210202 652800 214542
rect 652956 210338 652984 221167
rect 653126 220688 653182 220697
rect 653126 220623 653182 220632
rect 653140 213926 653168 220623
rect 653416 220114 653444 229055
rect 659568 227792 659620 227798
rect 659568 227734 659620 227740
rect 654782 226672 654838 226681
rect 654782 226607 654838 226616
rect 653404 220108 653456 220114
rect 653404 220050 653456 220056
rect 654796 218074 654824 226607
rect 658922 226400 658978 226409
rect 658922 226335 658978 226344
rect 656714 225040 656770 225049
rect 656714 224975 656770 224984
rect 656162 224496 656218 224505
rect 656162 224431 656218 224440
rect 654968 223644 655020 223650
rect 654968 223586 655020 223592
rect 654784 218068 654836 218074
rect 654784 218010 654836 218016
rect 653128 213920 653180 213926
rect 653128 213862 653180 213868
rect 652956 210310 653076 210338
rect 653048 210202 653076 210310
rect 654980 210202 655008 223586
rect 656176 215354 656204 224431
rect 656728 223650 656756 224975
rect 658186 223952 658242 223961
rect 658186 223887 658242 223896
rect 656898 223680 656954 223689
rect 656716 223644 656768 223650
rect 656898 223615 656954 223624
rect 656716 223586 656768 223592
rect 656912 222306 656940 223615
rect 657542 223136 657598 223145
rect 657542 223071 657598 223080
rect 656728 222278 656940 222306
rect 656530 217016 656586 217025
rect 656530 216951 656586 216960
rect 655428 215348 655480 215354
rect 655428 215290 655480 215296
rect 656164 215348 656216 215354
rect 656164 215290 656216 215296
rect 655440 210202 655468 215290
rect 656544 210202 656572 216951
rect 652772 210174 652924 210202
rect 653048 210174 653476 210202
rect 654580 210174 655008 210202
rect 655132 210174 655468 210202
rect 656236 210174 656572 210202
rect 656728 210202 656756 222278
rect 657556 213654 657584 223071
rect 657544 213648 657596 213654
rect 657544 213590 657596 213596
rect 658200 210202 658228 223887
rect 658936 214742 658964 226335
rect 658924 214736 658976 214742
rect 658924 214678 658976 214684
rect 659382 214568 659438 214577
rect 659382 214503 659438 214512
rect 658740 212764 658792 212770
rect 658740 212706 658792 212712
rect 658752 210202 658780 212706
rect 656728 210174 656788 210202
rect 657892 210174 658228 210202
rect 658444 210174 658780 210202
rect 659396 210202 659424 214503
rect 659580 212770 659608 227734
rect 660210 223408 660266 223417
rect 660210 223343 660266 223352
rect 660224 213382 660252 223343
rect 660960 213926 660988 229735
rect 660396 213920 660448 213926
rect 660396 213862 660448 213868
rect 660948 213920 661000 213926
rect 660948 213862 661000 213868
rect 660212 213376 660264 213382
rect 660212 213318 660264 213324
rect 659568 212764 659620 212770
rect 659568 212706 659620 212712
rect 660408 210202 660436 213862
rect 660948 213784 661000 213790
rect 660948 213726 661000 213732
rect 660960 210202 660988 213726
rect 661500 213172 661552 213178
rect 661500 213114 661552 213120
rect 661512 210202 661540 213114
rect 662064 210202 662092 231095
rect 662236 231066 662288 231072
rect 659396 210174 659548 210202
rect 660100 210174 660436 210202
rect 660652 210174 660988 210202
rect 661204 210174 661540 210202
rect 661756 210174 662092 210202
rect 662248 210202 662276 231066
rect 663062 230616 663118 230625
rect 663062 230551 663118 230560
rect 663076 215294 663104 230551
rect 663812 227746 663840 231775
rect 664442 230888 664498 230897
rect 664442 230823 664498 230832
rect 663628 227718 663840 227746
rect 663248 216164 663300 216170
rect 663248 216106 663300 216112
rect 663260 215294 663288 216106
rect 662984 215266 663104 215294
rect 663168 215266 663288 215294
rect 662984 213790 663012 215266
rect 662972 213784 663024 213790
rect 662972 213726 663024 213732
rect 663168 210202 663196 215266
rect 663628 210202 663656 227718
rect 664456 216170 664484 230823
rect 664444 216164 664496 216170
rect 664444 216106 664496 216112
rect 664810 213480 664866 213489
rect 664810 213415 664866 213424
rect 664260 213036 664312 213042
rect 664260 212978 664312 212984
rect 664272 210202 664300 212978
rect 664824 210202 664852 213415
rect 665100 213042 665128 232154
rect 665270 230344 665326 230353
rect 665270 230279 665326 230288
rect 665284 227798 665312 230279
rect 665272 227792 665324 227798
rect 665272 227734 665324 227740
rect 665822 225448 665878 225457
rect 665822 225383 665878 225392
rect 665454 220960 665510 220969
rect 665454 220895 665510 220904
rect 665088 213036 665140 213042
rect 665088 212978 665140 212984
rect 665468 212906 665496 220895
rect 665836 214606 665864 225383
rect 666282 215112 666338 215121
rect 666282 215047 666338 215056
rect 665824 214600 665876 214606
rect 665824 214542 665876 214548
rect 666296 213178 666324 215047
rect 666284 213172 666336 213178
rect 666284 213114 666336 213120
rect 665456 212900 665508 212906
rect 665456 212842 665508 212848
rect 662248 210174 662308 210202
rect 662860 210174 663196 210202
rect 663412 210174 663656 210202
rect 663964 210174 664300 210202
rect 664516 210174 664852 210202
rect 652208 209704 652260 209710
rect 652208 209646 652260 209652
rect 632152 209568 632204 209574
rect 652024 209568 652076 209574
rect 632204 209516 632500 209522
rect 632152 209510 632500 209516
rect 652024 209510 652076 209516
rect 632164 209494 632500 209510
rect 589464 208344 589516 208350
rect 589464 208286 589516 208292
rect 589476 208049 589504 208286
rect 589462 208040 589518 208049
rect 589462 207975 589518 207984
rect 589648 207664 589700 207670
rect 589648 207606 589700 207612
rect 589464 206916 589516 206922
rect 589464 206858 589516 206864
rect 589476 206417 589504 206858
rect 589462 206408 589518 206417
rect 589462 206343 589518 206352
rect 582380 205828 582432 205834
rect 582380 205770 582432 205776
rect 582392 202842 582420 205770
rect 589660 204785 589688 207606
rect 589646 204776 589702 204785
rect 589646 204711 589702 204720
rect 589464 204264 589516 204270
rect 589464 204206 589516 204212
rect 589476 203153 589504 204206
rect 589462 203144 589518 203153
rect 589462 203079 589518 203088
rect 582380 202836 582432 202842
rect 582380 202778 582432 202784
rect 589464 202836 589516 202842
rect 589464 202778 589516 202784
rect 589476 201521 589504 202778
rect 589462 201512 589518 201521
rect 589462 201447 589518 201456
rect 590384 200184 590436 200190
rect 590384 200126 590436 200132
rect 589464 200048 589516 200054
rect 589464 199990 589516 199996
rect 589476 199889 589504 199990
rect 589462 199880 589518 199889
rect 589462 199815 589518 199824
rect 589464 198756 589516 198762
rect 589464 198698 589516 198704
rect 589476 196625 589504 198698
rect 590396 198257 590424 200126
rect 590382 198248 590438 198257
rect 590382 198183 590438 198192
rect 589462 196616 589518 196625
rect 589462 196551 589518 196560
rect 589280 196036 589332 196042
rect 589280 195978 589332 195984
rect 589292 194993 589320 195978
rect 589278 194984 589334 194993
rect 589278 194919 589334 194928
rect 589464 194608 589516 194614
rect 589464 194550 589516 194556
rect 589476 193361 589504 194550
rect 589462 193352 589518 193361
rect 589462 193287 589518 193296
rect 589464 191888 589516 191894
rect 589464 191830 589516 191836
rect 589476 191729 589504 191830
rect 589462 191720 589518 191729
rect 589462 191655 589518 191664
rect 590568 190528 590620 190534
rect 590568 190470 590620 190476
rect 590580 190097 590608 190470
rect 590566 190088 590622 190097
rect 590566 190023 590622 190032
rect 589646 188456 589702 188465
rect 589646 188391 589702 188400
rect 589464 187740 589516 187746
rect 589464 187682 589516 187688
rect 589476 186833 589504 187682
rect 589462 186824 589518 186833
rect 589462 186759 589518 186768
rect 589660 186318 589688 188391
rect 589648 186312 589700 186318
rect 589648 186254 589700 186260
rect 589462 185192 589518 185201
rect 589462 185127 589518 185136
rect 589476 184890 589504 185127
rect 589464 184884 589516 184890
rect 589464 184826 589516 184832
rect 589462 183560 589518 183569
rect 589462 183495 589518 183504
rect 589476 182170 589504 183495
rect 589464 182164 589516 182170
rect 589464 182106 589516 182112
rect 590566 181928 590622 181937
rect 590566 181863 590622 181872
rect 590580 180810 590608 181863
rect 590568 180804 590620 180810
rect 590568 180746 590620 180752
rect 589646 180296 589702 180305
rect 589646 180231 589702 180240
rect 589462 178664 589518 178673
rect 589462 178599 589518 178608
rect 589476 178090 589504 178599
rect 589464 178084 589516 178090
rect 589464 178026 589516 178032
rect 589660 177954 589688 180231
rect 666664 178809 666692 324294
rect 667018 218104 667074 218113
rect 667018 218039 667074 218048
rect 667032 213217 667060 218039
rect 667018 213208 667074 213217
rect 667018 213143 667074 213152
rect 666836 209228 666888 209234
rect 666836 209170 666888 209176
rect 666650 178800 666706 178809
rect 666650 178735 666706 178744
rect 666848 178537 666876 209170
rect 667020 209092 667072 209098
rect 667020 209034 667072 209040
rect 666834 178528 666890 178537
rect 666834 178463 666890 178472
rect 589648 177948 589700 177954
rect 589648 177890 589700 177896
rect 589646 177032 589702 177041
rect 589646 176967 589702 176976
rect 589462 175400 589518 175409
rect 589462 175335 589464 175344
rect 589516 175335 589518 175344
rect 589464 175306 589516 175312
rect 582380 175296 582432 175302
rect 582380 175238 582432 175244
rect 582392 173262 582420 175238
rect 589660 174554 589688 176967
rect 589648 174548 589700 174554
rect 589648 174490 589700 174496
rect 589462 173768 589518 173777
rect 589462 173703 589518 173712
rect 582380 173256 582432 173262
rect 582380 173198 582432 173204
rect 589476 172582 589504 173703
rect 589464 172576 589516 172582
rect 589464 172518 589516 172524
rect 589462 172136 589518 172145
rect 589462 172071 589518 172080
rect 589476 171154 589504 172071
rect 589464 171148 589516 171154
rect 589464 171090 589516 171096
rect 589186 170504 589242 170513
rect 589186 170439 589242 170448
rect 582380 167068 582432 167074
rect 582380 167010 582432 167016
rect 582392 162586 582420 167010
rect 589200 166326 589228 170439
rect 589830 168872 589886 168881
rect 589830 168807 589886 168816
rect 589462 167240 589518 167249
rect 589462 167175 589518 167184
rect 589476 167074 589504 167175
rect 589464 167068 589516 167074
rect 589464 167010 589516 167016
rect 589188 166320 589240 166326
rect 589188 166262 589240 166268
rect 589646 165608 589702 165617
rect 589646 165543 589702 165552
rect 589462 163976 589518 163985
rect 589462 163911 589518 163920
rect 589476 162926 589504 163911
rect 589464 162920 589516 162926
rect 589464 162862 589516 162868
rect 582380 162580 582432 162586
rect 582380 162522 582432 162528
rect 589660 162178 589688 165543
rect 589844 164898 589872 168807
rect 589832 164892 589884 164898
rect 589832 164834 589884 164840
rect 590566 162344 590622 162353
rect 590566 162279 590622 162288
rect 589648 162172 589700 162178
rect 589648 162114 589700 162120
rect 589462 160712 589518 160721
rect 589462 160647 589518 160656
rect 589476 160138 589504 160647
rect 582380 160132 582432 160138
rect 582380 160074 582432 160080
rect 589464 160132 589516 160138
rect 589464 160074 589516 160080
rect 582392 152658 582420 160074
rect 590580 159390 590608 162279
rect 583760 159384 583812 159390
rect 583760 159326 583812 159332
rect 590568 159384 590620 159390
rect 590568 159326 590620 159332
rect 583772 154222 583800 159326
rect 588542 159080 588598 159089
rect 588542 159015 588598 159024
rect 587164 157412 587216 157418
rect 587164 157354 587216 157360
rect 585784 154624 585836 154630
rect 585784 154566 585836 154572
rect 583760 154216 583812 154222
rect 583760 154158 583812 154164
rect 584404 153264 584456 153270
rect 584404 153206 584456 153212
rect 582380 152652 582432 152658
rect 582380 152594 582432 152600
rect 583024 151836 583076 151842
rect 583024 151778 583076 151784
rect 583036 140622 583064 151778
rect 584416 143478 584444 153206
rect 585796 144702 585824 154566
rect 587176 148374 587204 157354
rect 588556 151094 588584 159015
rect 589278 157448 589334 157457
rect 589278 157383 589280 157392
rect 589332 157383 589334 157392
rect 589280 157354 589332 157360
rect 589462 155816 589518 155825
rect 589462 155751 589518 155760
rect 589476 154630 589504 155751
rect 589464 154624 589516 154630
rect 589464 154566 589516 154572
rect 589462 154184 589518 154193
rect 589462 154119 589518 154128
rect 589476 153270 589504 154119
rect 589464 153264 589516 153270
rect 589464 153206 589516 153212
rect 589462 152552 589518 152561
rect 589462 152487 589518 152496
rect 589476 151842 589504 152487
rect 589464 151836 589516 151842
rect 589464 151778 589516 151784
rect 588544 151088 588596 151094
rect 588544 151030 588596 151036
rect 589922 150920 589978 150929
rect 589922 150855 589978 150864
rect 589186 149288 589242 149297
rect 589186 149223 589242 149232
rect 587164 148368 587216 148374
rect 587164 148310 587216 148316
rect 585968 146328 586020 146334
rect 585968 146270 586020 146276
rect 585784 144696 585836 144702
rect 585784 144638 585836 144644
rect 584404 143472 584456 143478
rect 584404 143414 584456 143420
rect 583208 140820 583260 140826
rect 583208 140762 583260 140768
rect 583024 140616 583076 140622
rect 583024 140558 583076 140564
rect 581828 131912 581880 131918
rect 581828 131854 581880 131860
rect 581840 117230 581868 131854
rect 583220 125390 583248 140762
rect 584404 139460 584456 139466
rect 584404 139402 584456 139408
rect 583208 125384 583260 125390
rect 583208 125326 583260 125332
rect 583024 124908 583076 124914
rect 583024 124850 583076 124856
rect 581828 117224 581880 117230
rect 581828 117166 581880 117172
rect 581828 109744 581880 109750
rect 581828 109686 581880 109692
rect 581644 97980 581696 97986
rect 581644 97922 581696 97928
rect 580632 86488 580684 86494
rect 580632 86430 580684 86436
rect 581840 84046 581868 109686
rect 583036 103358 583064 124850
rect 584416 124166 584444 139402
rect 585980 138174 586008 146270
rect 588726 146024 588782 146033
rect 588726 145959 588782 145968
rect 587164 143608 587216 143614
rect 587164 143550 587216 143556
rect 585968 138168 586020 138174
rect 585968 138110 586020 138116
rect 585968 135312 586020 135318
rect 585968 135254 586020 135260
rect 584404 124160 584456 124166
rect 584404 124102 584456 124108
rect 584588 122868 584640 122874
rect 584588 122810 584640 122816
rect 583208 111104 583260 111110
rect 583208 111046 583260 111052
rect 583024 103352 583076 103358
rect 583024 103294 583076 103300
rect 583024 97572 583076 97578
rect 583024 97514 583076 97520
rect 581828 84040 581880 84046
rect 581828 83982 581880 83988
rect 581644 83496 581696 83502
rect 581644 83438 581696 83444
rect 580264 78260 580316 78266
rect 580264 78202 580316 78208
rect 579068 76560 579120 76566
rect 579068 76502 579120 76508
rect 578882 75712 578938 75721
rect 578882 75647 578938 75656
rect 578712 74506 578924 74534
rect 578516 62076 578568 62082
rect 578516 62018 578568 62024
rect 578528 61849 578556 62018
rect 578514 61840 578570 61849
rect 578514 61775 578570 61784
rect 577688 52420 577740 52426
rect 577688 52362 577740 52368
rect 578896 51474 578924 74506
rect 579080 64841 579108 76502
rect 579528 73160 579580 73166
rect 579526 73128 579528 73137
rect 579580 73128 579582 73137
rect 579526 73063 579582 73072
rect 581656 71534 581684 83438
rect 579252 71528 579304 71534
rect 579252 71470 579304 71476
rect 581644 71528 581696 71534
rect 581644 71470 581696 71476
rect 579264 71233 579292 71470
rect 579250 71224 579306 71233
rect 579250 71159 579306 71168
rect 579526 66328 579582 66337
rect 579526 66263 579528 66272
rect 579580 66263 579582 66272
rect 579528 66234 579580 66240
rect 579066 64832 579122 64841
rect 579066 64767 579122 64776
rect 579528 60716 579580 60722
rect 579528 60658 579580 60664
rect 579540 60353 579568 60658
rect 579526 60344 579582 60353
rect 579526 60279 579582 60288
rect 579528 57928 579580 57934
rect 579526 57896 579528 57905
rect 579580 57896 579582 57905
rect 579526 57831 579582 57840
rect 579528 56568 579580 56574
rect 579528 56510 579580 56516
rect 579540 56137 579568 56510
rect 579526 56128 579582 56137
rect 579526 56063 579582 56072
rect 583036 52154 583064 97514
rect 583220 82822 583248 111046
rect 583760 107704 583812 107710
rect 583760 107646 583812 107652
rect 583772 105194 583800 107646
rect 583760 105188 583812 105194
rect 583760 105130 583812 105136
rect 584600 101726 584628 122810
rect 585980 118454 586008 135254
rect 587176 131782 587204 143550
rect 588542 137864 588598 137873
rect 588542 137799 588598 137808
rect 587164 131776 587216 131782
rect 587164 131718 587216 131724
rect 587532 131164 587584 131170
rect 587532 131106 587584 131112
rect 587544 122262 587572 131106
rect 587532 122256 587584 122262
rect 587532 122198 587584 122204
rect 587348 121508 587400 121514
rect 587348 121450 587400 121456
rect 585968 118448 586020 118454
rect 585968 118390 586020 118396
rect 585784 117360 585836 117366
rect 585784 117302 585836 117308
rect 584588 101720 584640 101726
rect 584588 101662 584640 101668
rect 584404 101448 584456 101454
rect 584404 101390 584456 101396
rect 583208 82816 583260 82822
rect 583208 82758 583260 82764
rect 584416 73166 584444 101390
rect 585796 93158 585824 117302
rect 585968 116000 586020 116006
rect 585968 115942 586020 115948
rect 585784 93152 585836 93158
rect 585784 93094 585836 93100
rect 585980 91866 586008 115942
rect 587164 104916 587216 104922
rect 587164 104858 587216 104864
rect 585968 91860 586020 91866
rect 585968 91802 586020 91808
rect 584588 90364 584640 90370
rect 584588 90306 584640 90312
rect 584600 77246 584628 90306
rect 587176 82142 587204 104858
rect 587360 98802 587388 121450
rect 588556 121378 588584 137799
rect 588740 137290 588768 145959
rect 589200 145586 589228 149223
rect 589462 147656 589518 147665
rect 589462 147591 589518 147600
rect 589476 146334 589504 147591
rect 589464 146328 589516 146334
rect 589464 146270 589516 146276
rect 589188 145580 589240 145586
rect 589188 145522 589240 145528
rect 589462 144392 589518 144401
rect 589462 144327 589518 144336
rect 589476 143614 589504 144327
rect 589464 143608 589516 143614
rect 589464 143550 589516 143556
rect 589646 142760 589702 142769
rect 589646 142695 589702 142704
rect 589462 141128 589518 141137
rect 589462 141063 589518 141072
rect 589476 140826 589504 141063
rect 589464 140820 589516 140826
rect 589464 140762 589516 140768
rect 589462 139496 589518 139505
rect 589462 139431 589464 139440
rect 589516 139431 589518 139440
rect 589464 139402 589516 139408
rect 589660 137426 589688 142695
rect 589936 139330 589964 150855
rect 589924 139324 589976 139330
rect 589924 139266 589976 139272
rect 589648 137420 589700 137426
rect 589648 137362 589700 137368
rect 588728 137284 588780 137290
rect 588728 137226 588780 137232
rect 589462 136232 589518 136241
rect 589462 136167 589518 136176
rect 589476 135318 589504 136167
rect 589464 135312 589516 135318
rect 589464 135254 589516 135260
rect 590290 134600 590346 134609
rect 590290 134535 590346 134544
rect 589922 132968 589978 132977
rect 589922 132903 589978 132912
rect 589278 129704 589334 129713
rect 589278 129639 589334 129648
rect 589292 124914 589320 129639
rect 589462 128072 589518 128081
rect 589462 128007 589518 128016
rect 589476 127022 589504 128007
rect 589464 127016 589516 127022
rect 589464 126958 589516 126964
rect 589462 126440 589518 126449
rect 589462 126375 589518 126384
rect 589476 125662 589504 126375
rect 589464 125656 589516 125662
rect 589464 125598 589516 125604
rect 589280 124908 589332 124914
rect 589280 124850 589332 124856
rect 589738 124808 589794 124817
rect 589738 124743 589794 124752
rect 589462 123176 589518 123185
rect 589462 123111 589518 123120
rect 589476 122874 589504 123111
rect 589464 122868 589516 122874
rect 589464 122810 589516 122816
rect 589752 122126 589780 124743
rect 589740 122120 589792 122126
rect 589740 122062 589792 122068
rect 589278 121544 589334 121553
rect 589278 121479 589280 121488
rect 589332 121479 589334 121488
rect 589280 121450 589332 121456
rect 588544 121372 588596 121378
rect 588544 121314 588596 121320
rect 588726 119912 588782 119921
rect 588726 119847 588782 119856
rect 588544 113756 588596 113762
rect 588544 113698 588596 113704
rect 587348 98796 587400 98802
rect 587348 98738 587400 98744
rect 588556 88330 588584 113698
rect 588740 95198 588768 119847
rect 589462 118280 589518 118289
rect 589462 118215 589518 118224
rect 589476 117366 589504 118215
rect 589464 117360 589516 117366
rect 589464 117302 589516 117308
rect 589462 116648 589518 116657
rect 589462 116583 589518 116592
rect 589476 116006 589504 116583
rect 589464 116000 589516 116006
rect 589464 115942 589516 115948
rect 589554 115016 589610 115025
rect 589554 114951 589610 114960
rect 589568 113762 589596 114951
rect 589556 113756 589608 113762
rect 589556 113698 589608 113704
rect 589936 113150 589964 132903
rect 590304 131918 590332 134535
rect 667032 133113 667060 209034
rect 667216 181393 667244 350542
rect 668596 311953 668624 444382
rect 669424 403753 669452 536794
rect 669608 533089 669636 577759
rect 669792 570353 669820 643447
rect 669976 581097 670004 696934
rect 670422 684992 670478 685001
rect 670422 684927 670478 684936
rect 670238 668264 670294 668273
rect 670238 668199 670294 668208
rect 670252 630674 670280 668199
rect 670436 630674 670464 684927
rect 670804 669905 670832 714847
rect 670988 713697 671016 758231
rect 670974 713688 671030 713697
rect 670974 713623 671030 713632
rect 671172 705537 671200 774959
rect 671356 763745 671384 895630
rect 671802 869272 671858 869281
rect 671802 869207 671858 869216
rect 671342 763736 671398 763745
rect 671342 763671 671398 763680
rect 671434 759928 671490 759937
rect 671434 759863 671490 759872
rect 671448 757602 671476 759863
rect 671618 759112 671674 759121
rect 671618 759047 671674 759056
rect 671448 757574 671568 757602
rect 671342 757480 671398 757489
rect 671342 757415 671398 757424
rect 671356 721754 671384 757415
rect 671540 741074 671568 757574
rect 671264 721726 671384 721754
rect 671448 741046 671568 741074
rect 671264 715170 671292 721726
rect 671448 715329 671476 741046
rect 671434 715320 671490 715329
rect 671434 715255 671490 715264
rect 671264 715142 671384 715170
rect 671356 712881 671384 715142
rect 671632 714513 671660 759047
rect 671816 756254 671844 869207
rect 672000 757897 672028 935711
rect 672552 933201 672580 952167
rect 672736 947345 672764 975666
rect 675404 966521 675432 966723
rect 675390 966512 675446 966521
rect 675390 966447 675446 966456
rect 672998 966376 673054 966385
rect 672998 966311 673054 966320
rect 675114 966376 675170 966385
rect 675114 966311 675170 966320
rect 672722 947336 672778 947345
rect 672722 947271 672778 947280
rect 672722 938088 672778 938097
rect 672722 938023 672778 938032
rect 672538 933192 672594 933201
rect 672538 933127 672594 933136
rect 672354 787400 672410 787409
rect 672354 787335 672410 787344
rect 672368 785234 672396 787335
rect 672736 785234 672764 938023
rect 673012 932929 673040 966311
rect 675128 966090 675156 966311
rect 675128 966062 675418 966090
rect 674944 965421 675418 965449
rect 674378 962840 674434 962849
rect 674378 962775 674434 962784
rect 673182 960800 673238 960809
rect 673182 960735 673238 960744
rect 672998 932920 673054 932929
rect 672998 932855 673054 932864
rect 673196 930753 673224 960735
rect 674102 959304 674158 959313
rect 674102 959239 674158 959248
rect 673366 937408 673422 937417
rect 673366 937343 673422 937352
rect 673182 930744 673238 930753
rect 673182 930679 673238 930688
rect 673182 872264 673238 872273
rect 673182 872199 673238 872208
rect 672368 785206 672488 785234
rect 672736 785206 672856 785234
rect 672460 775574 672488 785206
rect 672630 783864 672686 783873
rect 672630 783799 672686 783808
rect 672460 775546 672580 775574
rect 671986 757888 672042 757897
rect 671986 757823 672042 757832
rect 671816 756226 672028 756254
rect 672000 751777 672028 756226
rect 671986 751768 672042 751777
rect 671986 751703 672042 751712
rect 672354 750136 672410 750145
rect 672354 750071 672410 750080
rect 671986 743472 672042 743481
rect 671986 743407 672042 743416
rect 671802 735584 671858 735593
rect 671802 735519 671858 735528
rect 671816 731414 671844 735519
rect 671816 731386 671936 731414
rect 671618 714504 671674 714513
rect 671618 714439 671674 714448
rect 671710 714096 671766 714105
rect 671710 714031 671766 714040
rect 671526 713280 671582 713289
rect 671526 713215 671582 713224
rect 671342 712872 671398 712881
rect 671342 712807 671398 712816
rect 671158 705528 671214 705537
rect 671158 705463 671214 705472
rect 671540 702434 671568 713215
rect 671724 702434 671752 714031
rect 671448 702406 671568 702434
rect 671632 702406 671752 702434
rect 671448 692774 671476 702406
rect 671632 692774 671660 702406
rect 671908 692774 671936 731386
rect 671356 692746 671476 692774
rect 671540 692746 671660 692774
rect 671816 692746 671936 692774
rect 670974 689072 671030 689081
rect 670974 689007 671030 689016
rect 670790 669896 670846 669905
rect 670790 669831 670846 669840
rect 670606 666632 670662 666641
rect 670606 666567 670662 666576
rect 670160 630646 670280 630674
rect 670344 630646 670464 630674
rect 670160 624345 670188 630646
rect 670146 624336 670202 624345
rect 670146 624271 670202 624280
rect 670344 622690 670372 630646
rect 670620 627914 670648 666567
rect 670790 647864 670846 647873
rect 670790 647799 670846 647808
rect 670252 622662 670372 622690
rect 670436 627886 670648 627914
rect 670252 621014 670280 622662
rect 670436 622577 670464 627886
rect 670606 624744 670662 624753
rect 670606 624679 670662 624688
rect 670422 622568 670478 622577
rect 670422 622503 670478 622512
rect 670620 621014 670648 624679
rect 670160 620986 670280 621014
rect 670436 620986 670648 621014
rect 670160 615777 670188 620986
rect 670146 615768 670202 615777
rect 670146 615703 670202 615712
rect 670436 605834 670464 620986
rect 670606 614952 670662 614961
rect 670606 614887 670662 614896
rect 670160 605806 670464 605834
rect 669962 581088 670018 581097
rect 669962 581023 670018 581032
rect 670160 580825 670188 605806
rect 670146 580816 670202 580825
rect 670146 580751 670202 580760
rect 670238 579456 670294 579465
rect 670238 579391 670294 579400
rect 669962 578640 670018 578649
rect 669962 578575 670018 578584
rect 669778 570344 669834 570353
rect 669778 570279 669834 570288
rect 669778 569528 669834 569537
rect 669778 569463 669834 569472
rect 669594 533080 669650 533089
rect 669594 533015 669650 533024
rect 669792 455161 669820 569463
rect 669976 534721 670004 578575
rect 670252 534993 670280 579391
rect 670422 553480 670478 553489
rect 670422 553415 670478 553424
rect 670238 534984 670294 534993
rect 670238 534919 670294 534928
rect 669962 534712 670018 534721
rect 669962 534647 670018 534656
rect 670436 482361 670464 553415
rect 670422 482352 670478 482361
rect 670422 482287 670478 482296
rect 670620 455433 670648 614887
rect 670804 571985 670832 647799
rect 670988 616593 671016 689007
rect 671356 688634 671384 692746
rect 671540 688634 671568 692746
rect 671816 688634 671844 692746
rect 671356 688606 671476 688634
rect 671540 688606 671660 688634
rect 671816 688606 671936 688634
rect 671250 670304 671306 670313
rect 671250 670239 671306 670248
rect 671264 625161 671292 670239
rect 671448 668545 671476 688606
rect 671632 669497 671660 688606
rect 671908 684298 671936 688606
rect 672000 684570 672028 743407
rect 672172 728476 672224 728482
rect 672172 728418 672224 728424
rect 672184 728249 672212 728418
rect 672368 728346 672396 750071
rect 672356 728340 672408 728346
rect 672356 728282 672408 728288
rect 672170 728240 672226 728249
rect 672170 728175 672226 728184
rect 672170 712464 672226 712473
rect 672170 712399 672226 712408
rect 672184 685874 672212 712399
rect 672552 710841 672580 775546
rect 672644 731414 672672 783799
rect 672828 759529 672856 785206
rect 672998 784272 673054 784281
rect 672998 784207 673054 784216
rect 672814 759520 672870 759529
rect 672814 759455 672870 759464
rect 672814 756256 672870 756265
rect 672814 756191 672870 756200
rect 672828 755177 672856 756191
rect 672814 755168 672870 755177
rect 672814 755103 672870 755112
rect 672814 734088 672870 734097
rect 672814 734023 672870 734032
rect 672644 731386 672764 731414
rect 672538 710832 672594 710841
rect 672538 710767 672594 710776
rect 672736 710682 672764 731386
rect 672552 710654 672764 710682
rect 672552 709481 672580 710654
rect 672538 709472 672594 709481
rect 672538 709407 672594 709416
rect 672538 698320 672594 698329
rect 672538 698255 672594 698264
rect 672354 696960 672410 696969
rect 672354 696895 672410 696904
rect 672184 685846 672304 685874
rect 672000 684542 672212 684570
rect 671908 684270 672028 684298
rect 671802 680096 671858 680105
rect 671802 680031 671858 680040
rect 671618 669488 671674 669497
rect 671618 669423 671674 669432
rect 671434 668536 671490 668545
rect 671434 668471 671490 668480
rect 671526 667992 671582 668001
rect 671526 667927 671582 667936
rect 671250 625152 671306 625161
rect 671250 625087 671306 625096
rect 671540 623529 671568 667927
rect 671526 623520 671582 623529
rect 671526 623455 671582 623464
rect 671158 622840 671214 622849
rect 671158 622775 671214 622784
rect 670974 616584 671030 616593
rect 670974 616519 671030 616528
rect 671172 578241 671200 622775
rect 671618 622296 671674 622305
rect 671618 622231 671674 622240
rect 671342 594824 671398 594833
rect 671342 594759 671398 594768
rect 671158 578232 671214 578241
rect 671158 578167 671214 578176
rect 670790 571976 670846 571985
rect 670790 571911 670846 571920
rect 670790 570752 670846 570761
rect 670790 570687 670846 570696
rect 670804 500993 670832 570687
rect 671158 548448 671214 548457
rect 671158 548383 671214 548392
rect 670974 532808 671030 532817
rect 670974 532743 671030 532752
rect 670790 500984 670846 500993
rect 670790 500919 670846 500928
rect 670988 489297 671016 532743
rect 670974 489288 671030 489297
rect 670974 489223 671030 489232
rect 671172 485625 671200 548383
rect 671356 524929 671384 594759
rect 671632 577425 671660 622231
rect 671816 620401 671844 680031
rect 672000 679946 672028 684270
rect 671908 679918 672028 679946
rect 671908 665802 671936 679918
rect 672184 676682 672212 684542
rect 672000 676654 672212 676682
rect 672000 665938 672028 676654
rect 672276 676214 672304 685846
rect 672184 676186 672304 676214
rect 672184 667457 672212 676186
rect 672170 667448 672226 667457
rect 672170 667383 672226 667392
rect 672000 665910 672212 665938
rect 671908 665774 672028 665802
rect 672000 665718 672028 665774
rect 671988 665712 672040 665718
rect 671988 665654 672040 665660
rect 672184 665530 672212 665910
rect 672000 665502 672212 665530
rect 672000 664465 672028 665502
rect 671986 664456 672042 664465
rect 671986 664391 672042 664400
rect 671986 661056 672042 661065
rect 671986 660991 672042 661000
rect 671802 620392 671858 620401
rect 671802 620327 671858 620336
rect 671618 577416 671674 577425
rect 671618 577351 671674 577360
rect 671802 577008 671858 577017
rect 671802 576943 671858 576952
rect 671816 567194 671844 576943
rect 671724 567166 671844 567194
rect 671724 538214 671752 567166
rect 671632 538186 671752 538214
rect 671632 531865 671660 538186
rect 671802 534304 671858 534313
rect 671802 534239 671858 534248
rect 671618 531856 671674 531865
rect 671618 531791 671674 531800
rect 671618 531448 671674 531457
rect 671618 531383 671674 531392
rect 671342 524920 671398 524929
rect 671342 524855 671398 524864
rect 671434 490512 671490 490521
rect 671434 490447 671490 490456
rect 671158 485616 671214 485625
rect 671158 485551 671214 485560
rect 670606 455424 670662 455433
rect 670606 455359 670662 455368
rect 669778 455152 669834 455161
rect 669778 455087 669834 455096
rect 669964 430636 670016 430642
rect 669964 430578 670016 430584
rect 669410 403744 669466 403753
rect 669410 403679 669466 403688
rect 668582 311944 668638 311953
rect 668582 311879 668638 311888
rect 667388 310548 667440 310554
rect 667388 310490 667440 310496
rect 667202 181384 667258 181393
rect 667202 181319 667258 181328
rect 667400 142769 667428 310490
rect 669226 302288 669282 302297
rect 669226 302223 669282 302232
rect 667572 284368 667624 284374
rect 667572 284310 667624 284316
rect 667386 142760 667442 142769
rect 667386 142695 667442 142704
rect 667584 135969 667612 284310
rect 668768 237448 668820 237454
rect 668768 237390 668820 237396
rect 668124 234592 668176 234598
rect 668124 234534 668176 234540
rect 668490 234560 668546 234569
rect 667940 231192 667992 231198
rect 667938 231160 667940 231169
rect 667992 231160 667994 231169
rect 667938 231095 667994 231104
rect 668136 230466 668164 234534
rect 668490 234495 668546 234504
rect 668306 231568 668362 231577
rect 668306 231503 668362 231512
rect 668320 230625 668348 231503
rect 668306 230616 668362 230625
rect 668306 230551 668362 230560
rect 668136 230438 668348 230466
rect 668124 230308 668176 230314
rect 668124 230250 668176 230256
rect 667940 225684 667992 225690
rect 667940 225626 667992 225632
rect 667952 223145 667980 225626
rect 667938 223136 667994 223145
rect 667938 223071 667994 223080
rect 667940 221264 667992 221270
rect 667938 221232 667940 221241
rect 667992 221232 667994 221241
rect 667938 221167 667994 221176
rect 667846 219464 667902 219473
rect 667846 219399 667902 219408
rect 667860 186314 667888 219399
rect 668136 192681 668164 230250
rect 668122 192672 668178 192681
rect 668122 192607 668178 192616
rect 668032 192500 668084 192506
rect 668032 192442 668084 192448
rect 668044 187649 668072 192442
rect 668030 187640 668086 187649
rect 668030 187575 668086 187584
rect 667768 186286 667888 186314
rect 667768 175001 667796 186286
rect 667940 184544 667992 184550
rect 667938 184512 667940 184521
rect 667992 184512 667994 184521
rect 667938 184447 667994 184456
rect 668320 182889 668348 230438
rect 668306 182880 668362 182889
rect 668306 182815 668362 182824
rect 667754 174992 667810 175001
rect 667754 174927 667810 174936
rect 667940 174888 667992 174894
rect 667940 174830 667992 174836
rect 667952 174729 667980 174830
rect 667938 174720 667994 174729
rect 667938 174655 667994 174664
rect 668032 169720 668084 169726
rect 668030 169688 668032 169697
rect 668084 169688 668086 169697
rect 668030 169623 668086 169632
rect 667940 165232 667992 165238
rect 667940 165174 667992 165180
rect 667952 164937 667980 165174
rect 667938 164928 667994 164937
rect 667938 164863 667994 164872
rect 667940 160064 667992 160070
rect 667938 160032 667940 160041
rect 667992 160032 667994 160041
rect 667938 159967 667994 159976
rect 668308 150272 668360 150278
rect 668306 150240 668308 150249
rect 668360 150240 668362 150249
rect 668306 150175 668362 150184
rect 668504 148617 668532 234495
rect 668780 153513 668808 237390
rect 669044 233028 669096 233034
rect 669044 232970 669096 232976
rect 669056 231962 669084 232970
rect 669056 231934 669176 231962
rect 668950 231840 669006 231849
rect 668950 231775 669006 231784
rect 668964 231305 668992 231775
rect 668950 231296 669006 231305
rect 668950 231231 669006 231240
rect 669148 229094 669176 231934
rect 668964 229066 669176 229094
rect 668964 224954 668992 229066
rect 668872 224926 668992 224954
rect 668872 215294 668900 224926
rect 669044 224868 669096 224874
rect 669044 224810 669096 224816
rect 669056 224369 669084 224810
rect 669042 224360 669098 224369
rect 669042 224295 669098 224304
rect 669042 221912 669098 221921
rect 669042 221847 669098 221856
rect 668872 215266 668992 215294
rect 668964 193214 668992 215266
rect 669056 212534 669084 221847
rect 669056 212506 669176 212534
rect 669148 209774 669176 212506
rect 669056 209746 669176 209774
rect 669056 200114 669084 209746
rect 669240 206553 669268 302223
rect 669976 275369 670004 430578
rect 671448 402529 671476 490447
rect 671632 488481 671660 531383
rect 671816 490929 671844 534239
rect 671802 490920 671858 490929
rect 671802 490855 671858 490864
rect 671802 489696 671858 489705
rect 671802 489631 671858 489640
rect 671618 488472 671674 488481
rect 671618 488407 671674 488416
rect 671434 402520 671490 402529
rect 671434 402455 671490 402464
rect 671816 401713 671844 489631
rect 672000 455705 672028 660991
rect 672170 648680 672226 648689
rect 672170 648615 672226 648624
rect 672184 579086 672212 648615
rect 672368 620673 672396 696895
rect 672552 621625 672580 698255
rect 672828 662561 672856 734023
rect 673012 709209 673040 784207
rect 673196 752593 673224 872199
rect 673380 760345 673408 937343
rect 674116 933881 674144 959239
rect 674392 949454 674420 962775
rect 674746 958352 674802 958361
rect 674746 958287 674802 958296
rect 674562 957128 674618 957137
rect 674562 957063 674618 957072
rect 674576 949454 674604 957063
rect 674760 954122 674788 958287
rect 674944 956354 674972 965421
rect 675298 964744 675354 964753
rect 675298 964679 675354 964688
rect 675312 963254 675340 964679
rect 675772 963393 675800 963595
rect 675758 963384 675814 963393
rect 675758 963319 675814 963328
rect 675220 963226 675340 963254
rect 675220 962418 675248 963226
rect 675496 962849 675524 963016
rect 675482 962840 675538 962849
rect 675482 962775 675538 962784
rect 675220 962390 675418 962418
rect 675128 961741 675418 961769
rect 675128 960809 675156 961741
rect 675114 960800 675170 960809
rect 675114 960735 675170 960744
rect 675114 959304 675170 959313
rect 675170 959262 675418 959290
rect 675114 959239 675170 959248
rect 675404 958361 675432 958732
rect 675390 958352 675446 958361
rect 675390 958287 675446 958296
rect 675772 957817 675800 958052
rect 675206 957808 675262 957817
rect 675206 957743 675262 957752
rect 675758 957808 675814 957817
rect 675758 957743 675814 957752
rect 674944 956326 675064 956354
rect 674300 949426 674420 949454
rect 674484 949426 674604 949454
rect 674668 954094 674788 954122
rect 674102 933872 674158 933881
rect 674102 933807 674158 933816
rect 674300 932657 674328 949426
rect 674286 932648 674342 932657
rect 674286 932583 674342 932592
rect 674484 930209 674512 949426
rect 674668 930481 674696 954094
rect 674838 953456 674894 953465
rect 674838 953391 674894 953400
rect 674654 930472 674710 930481
rect 674654 930407 674710 930416
rect 674470 930200 674526 930209
rect 674470 930135 674526 930144
rect 674852 928792 674880 953391
rect 675036 949454 675064 956326
rect 675220 955482 675248 957743
rect 675404 957137 675432 957440
rect 675390 957128 675446 957137
rect 675390 957063 675446 957072
rect 675758 956448 675814 956457
rect 675758 956383 675814 956392
rect 675772 956216 675800 956383
rect 675220 955454 675524 955482
rect 675496 955060 675524 955454
rect 675312 954366 675418 954394
rect 675312 953714 675340 954366
rect 675220 953686 675340 953714
rect 675220 951674 675248 953686
rect 675404 953465 675432 953768
rect 675390 953456 675446 953465
rect 675390 953391 675446 953400
rect 675404 952241 675432 952544
rect 675390 952232 675446 952241
rect 675390 952167 675446 952176
rect 675220 951646 675616 951674
rect 675390 951552 675446 951561
rect 675390 951487 675446 951496
rect 675404 949454 675432 951487
rect 675588 949454 675616 951646
rect 683302 950736 683358 950745
rect 683302 950671 683358 950680
rect 679622 949512 679678 949521
rect 675852 949476 675904 949482
rect 675036 949426 675156 949454
rect 675404 949426 675524 949454
rect 675588 949426 675852 949454
rect 675128 943934 675156 949426
rect 675496 943934 675524 949426
rect 679622 949447 679678 949456
rect 682384 949476 682436 949482
rect 675852 949418 675904 949424
rect 675128 943906 675432 943934
rect 675496 943906 675616 943934
rect 675206 937952 675262 937961
rect 675206 937887 675262 937896
rect 675220 937009 675248 937887
rect 675206 937000 675262 937009
rect 675206 936935 675262 936944
rect 675404 935513 675432 943906
rect 675390 935504 675446 935513
rect 675390 935439 675446 935448
rect 675588 934697 675616 943906
rect 676218 941760 676274 941769
rect 676218 941695 676274 941704
rect 676232 939321 676260 941695
rect 676218 939312 676274 939321
rect 676218 939247 676274 939256
rect 675574 934688 675630 934697
rect 675574 934623 675630 934632
rect 679636 934425 679664 949447
rect 682384 949418 682436 949424
rect 682396 935241 682424 949418
rect 683118 947336 683174 947345
rect 683118 947271 683174 947280
rect 683132 939729 683160 947271
rect 683118 939720 683174 939729
rect 683118 939655 683174 939664
rect 682382 935232 682438 935241
rect 682382 935167 682438 935176
rect 679622 934416 679678 934425
rect 679622 934351 679678 934360
rect 683316 932385 683344 950671
rect 703694 940508 703722 940644
rect 704154 940508 704182 940644
rect 704614 940508 704642 940644
rect 705074 940508 705102 940644
rect 705534 940508 705562 940644
rect 705994 940508 706022 940644
rect 706454 940508 706482 940644
rect 706914 940508 706942 940644
rect 707374 940508 707402 940644
rect 707834 940508 707862 940644
rect 708294 940508 708322 940644
rect 708754 940508 708782 940644
rect 709214 940508 709242 940644
rect 683302 932376 683358 932385
rect 683302 932311 683358 932320
rect 683118 929112 683174 929121
rect 683118 929047 683174 929056
rect 683132 928810 683160 929047
rect 675852 928804 675904 928810
rect 674852 928764 675852 928792
rect 675852 928746 675904 928752
rect 683120 928804 683172 928810
rect 683120 928746 683172 928752
rect 675298 879200 675354 879209
rect 675298 879135 675354 879144
rect 675312 877418 675340 879135
rect 675404 877418 675432 877540
rect 675312 877390 675432 877418
rect 675772 876625 675800 876860
rect 675758 876616 675814 876625
rect 675758 876551 675814 876560
rect 675114 876344 675170 876353
rect 675114 876279 675170 876288
rect 675128 873882 675156 876279
rect 675772 875945 675800 876248
rect 675758 875936 675814 875945
rect 675758 875871 675814 875880
rect 675404 874041 675432 874412
rect 675390 874032 675446 874041
rect 675390 873967 675446 873976
rect 675128 873854 675340 873882
rect 675312 873746 675340 873854
rect 675404 873746 675432 873868
rect 675312 873718 675432 873746
rect 675114 873216 675170 873225
rect 675170 873174 675418 873202
rect 675114 873151 675170 873160
rect 675114 872536 675170 872545
rect 675114 872471 675170 872480
rect 675128 870074 675156 872471
rect 675404 872273 675432 872576
rect 675390 872264 675446 872273
rect 675390 872199 675446 872208
rect 675128 870046 675418 870074
rect 674852 869502 675418 869530
rect 674852 868889 674880 869502
rect 674760 868861 674880 868889
rect 675312 868861 675418 868889
rect 674562 868456 674618 868465
rect 674562 868391 674618 868400
rect 674102 867232 674158 867241
rect 674102 867167 674158 867176
rect 673734 864920 673790 864929
rect 673734 864855 673790 864864
rect 673550 777472 673606 777481
rect 673550 777407 673606 777416
rect 673366 760336 673422 760345
rect 673366 760271 673422 760280
rect 673182 752584 673238 752593
rect 673182 752519 673238 752528
rect 673182 751360 673238 751369
rect 673182 751295 673238 751304
rect 673196 728142 673224 751295
rect 673366 739936 673422 739945
rect 673366 739871 673422 739880
rect 673184 728136 673236 728142
rect 673184 728078 673236 728084
rect 672998 709200 673054 709209
rect 672998 709135 673054 709144
rect 673182 697232 673238 697241
rect 673182 697167 673238 697176
rect 673000 665712 673052 665718
rect 672998 665680 673000 665689
rect 673052 665680 673054 665689
rect 672998 665615 673054 665624
rect 672814 662552 672870 662561
rect 672814 662487 672870 662496
rect 672722 648952 672778 648961
rect 672722 648887 672778 648896
rect 672736 640334 672764 648887
rect 672644 640306 672764 640334
rect 672644 630674 672672 640306
rect 672644 630646 672764 630674
rect 672538 621616 672594 621625
rect 672538 621551 672594 621560
rect 672736 621014 672764 630646
rect 672644 620986 672764 621014
rect 672354 620664 672410 620673
rect 672354 620599 672410 620608
rect 672446 608696 672502 608705
rect 672446 608631 672502 608640
rect 672460 607458 672488 608631
rect 672276 607430 672488 607458
rect 672276 579614 672304 607430
rect 672446 607336 672502 607345
rect 672446 607271 672502 607280
rect 672276 579586 672396 579614
rect 672172 579080 672224 579086
rect 672172 579022 672224 579028
rect 672368 574818 672396 579586
rect 672092 574790 672396 574818
rect 672092 567194 672120 574790
rect 672460 569954 672488 607271
rect 672644 575113 672672 620986
rect 673196 619721 673224 697167
rect 673380 663377 673408 739871
rect 673564 724305 673592 777407
rect 673748 772041 673776 864855
rect 673918 779240 673974 779249
rect 673918 779175 673974 779184
rect 673734 772032 673790 772041
rect 673734 771967 673790 771976
rect 673734 734360 673790 734369
rect 673734 734295 673790 734304
rect 673550 724296 673606 724305
rect 673550 724231 673606 724240
rect 673550 693560 673606 693569
rect 673550 693495 673606 693504
rect 673366 663368 673422 663377
rect 673366 663303 673422 663312
rect 673366 659968 673422 659977
rect 673366 659903 673422 659912
rect 673182 619712 673238 619721
rect 673182 619647 673238 619656
rect 672814 604888 672870 604897
rect 672814 604823 672870 604832
rect 672630 575104 672686 575113
rect 672630 575039 672686 575048
rect 672368 569926 672488 569954
rect 672368 567194 672396 569926
rect 672092 567166 672304 567194
rect 672368 567166 672488 567194
rect 672276 532545 672304 567166
rect 672262 532536 672318 532545
rect 672262 532471 672318 532480
rect 672460 529009 672488 567166
rect 672630 533488 672686 533497
rect 672630 533423 672686 533432
rect 672446 529000 672502 529009
rect 672446 528935 672502 528944
rect 672644 490113 672672 533423
rect 672828 530233 672856 604823
rect 672998 604344 673054 604353
rect 672998 604279 673054 604288
rect 673012 530641 673040 604279
rect 673380 601694 673408 659903
rect 673564 618633 673592 693495
rect 673748 682689 673776 734295
rect 673932 726889 673960 779175
rect 674116 753409 674144 867167
rect 674576 856994 674604 868391
rect 674760 856994 674788 868861
rect 674930 868728 674986 868737
rect 674930 868663 674986 868672
rect 675114 868728 675170 868737
rect 675114 868663 675170 868672
rect 674944 868034 674972 868663
rect 675128 868238 675156 868663
rect 675312 868465 675340 868861
rect 675298 868456 675354 868465
rect 675298 868391 675354 868400
rect 675128 868210 675418 868238
rect 674944 868006 675156 868034
rect 674930 866824 674986 866833
rect 674930 866759 674986 866768
rect 674484 856966 674604 856994
rect 674668 856966 674788 856994
rect 674944 856994 674972 866759
rect 675128 865858 675156 868006
rect 675298 867232 675354 867241
rect 675298 867167 675354 867176
rect 675312 867049 675340 867167
rect 675312 867021 675418 867049
rect 675128 865830 675418 865858
rect 675298 865328 675354 865337
rect 675298 865263 675354 865272
rect 675312 863818 675340 865263
rect 675496 864929 675524 865195
rect 675482 864920 675538 864929
rect 675482 864855 675538 864864
rect 675496 864249 675524 864552
rect 675482 864240 675538 864249
rect 675482 864175 675538 864184
rect 675312 863790 675432 863818
rect 675404 863328 675432 863790
rect 674944 856966 675340 856994
rect 674484 794894 674512 856966
rect 674668 794894 674696 856966
rect 675312 794894 675340 856966
rect 674484 794866 674604 794894
rect 674668 794866 674788 794894
rect 674286 788080 674342 788089
rect 674286 788015 674342 788024
rect 674300 765914 674328 788015
rect 674576 770681 674604 794866
rect 674562 770672 674618 770681
rect 674562 770607 674618 770616
rect 674300 765886 674696 765914
rect 674102 753400 674158 753409
rect 674102 753335 674158 753344
rect 674668 731414 674696 765886
rect 674760 757330 674788 794866
rect 675220 794866 675340 794894
rect 675220 786978 675248 794866
rect 675496 788089 675524 788324
rect 675482 788080 675538 788089
rect 675482 788015 675538 788024
rect 675496 787409 675524 787679
rect 675482 787400 675538 787409
rect 675482 787335 675538 787344
rect 675128 786950 675248 786978
rect 674930 786720 674986 786729
rect 674930 786655 674986 786664
rect 674944 782474 674972 786655
rect 675128 782474 675156 786950
rect 675404 786729 675432 787032
rect 675390 786720 675446 786729
rect 675390 786655 675446 786664
rect 674852 782446 674972 782474
rect 675036 782446 675156 782474
rect 675312 785182 675418 785210
rect 674852 776234 674880 782446
rect 675036 777209 675064 782446
rect 675312 780473 675340 785182
rect 675496 784281 675524 784652
rect 675482 784272 675538 784281
rect 675482 784207 675538 784216
rect 675496 783873 675524 783972
rect 675482 783864 675538 783873
rect 675482 783799 675538 783808
rect 675496 783057 675524 783360
rect 675482 783048 675538 783057
rect 675482 782983 675538 782992
rect 675496 780745 675524 780844
rect 675482 780736 675538 780745
rect 675482 780671 675538 780680
rect 675298 780464 675354 780473
rect 675298 780399 675354 780408
rect 675496 780065 675524 780300
rect 675482 780056 675538 780065
rect 675482 779991 675538 780000
rect 675496 779521 675524 779688
rect 675482 779512 675538 779521
rect 675482 779447 675538 779456
rect 675482 779240 675538 779249
rect 675482 779175 675538 779184
rect 675496 779008 675524 779175
rect 675298 778968 675354 778977
rect 675298 778903 675354 778912
rect 675022 777200 675078 777209
rect 675022 777135 675078 777144
rect 675312 777050 675340 778903
rect 675496 777481 675524 777852
rect 675482 777472 675538 777481
rect 675482 777407 675538 777416
rect 675312 777022 675432 777050
rect 675404 776628 675432 777022
rect 675482 776248 675538 776257
rect 674852 776206 675156 776234
rect 674930 775704 674986 775713
rect 674930 775639 674986 775648
rect 674944 774625 674972 775639
rect 674930 774616 674986 774625
rect 674930 774551 674986 774560
rect 675128 772814 675156 776206
rect 675482 776183 675538 776192
rect 675298 776112 675354 776121
rect 675298 776047 675354 776056
rect 675312 775588 675340 776047
rect 675496 776016 675524 776183
rect 675036 772786 675156 772814
rect 675220 775560 675340 775588
rect 675036 766601 675064 772786
rect 675022 766592 675078 766601
rect 675022 766527 675078 766536
rect 675220 765105 675248 775560
rect 675496 775033 675524 775336
rect 675482 775024 675538 775033
rect 675482 774959 675538 774968
rect 675482 774616 675538 774625
rect 675482 774551 675538 774560
rect 675496 774180 675524 774551
rect 675390 773392 675446 773401
rect 675390 773327 675446 773336
rect 675404 772814 675432 773327
rect 675404 772786 675892 772814
rect 675206 765096 675262 765105
rect 675206 765031 675262 765040
rect 674760 757302 674880 757330
rect 674852 757217 674880 757302
rect 674838 757208 674894 757217
rect 674838 757143 674894 757152
rect 675864 755857 675892 772786
rect 683210 772304 683266 772313
rect 683210 772239 683266 772248
rect 681002 768768 681058 768777
rect 681002 768703 681058 768712
rect 676770 761832 676826 761841
rect 676770 761767 676826 761776
rect 676034 757208 676090 757217
rect 676034 757143 676036 757152
rect 676088 757143 676090 757152
rect 676036 757114 676088 757120
rect 675850 755848 675906 755857
rect 675850 755783 675906 755792
rect 676784 754633 676812 761767
rect 681016 757081 681044 768703
rect 681002 757072 681058 757081
rect 681002 757007 681058 757016
rect 676770 754624 676826 754633
rect 676770 754559 676826 754568
rect 683224 753817 683252 772239
rect 683854 772032 683910 772041
rect 683854 771967 683910 771976
rect 683486 770672 683542 770681
rect 683486 770607 683542 770616
rect 683500 770054 683528 770607
rect 683500 770026 683620 770054
rect 683394 763736 683450 763745
rect 683394 763671 683450 763680
rect 683408 760753 683436 763671
rect 683394 760744 683450 760753
rect 683394 760679 683450 760688
rect 683396 757172 683448 757178
rect 683396 757114 683448 757120
rect 683210 753808 683266 753817
rect 683210 753743 683266 753752
rect 683408 752185 683436 757114
rect 683592 753001 683620 770026
rect 683868 756673 683896 771967
rect 703694 762076 703722 762212
rect 704154 762076 704182 762212
rect 704614 762076 704642 762212
rect 705074 762076 705102 762212
rect 705534 762076 705562 762212
rect 705994 762076 706022 762212
rect 706454 762076 706482 762212
rect 706914 762076 706942 762212
rect 707374 762076 707402 762212
rect 707834 762076 707862 762212
rect 708294 762076 708322 762212
rect 708754 762076 708782 762212
rect 709214 762076 709242 762212
rect 683854 756664 683910 756673
rect 683854 756599 683910 756608
rect 683578 752992 683634 753001
rect 683578 752927 683634 752936
rect 683394 752176 683450 752185
rect 683394 752111 683450 752120
rect 675298 745512 675354 745521
rect 675298 745447 675354 745456
rect 675114 743472 675170 743481
rect 675114 743407 675170 743416
rect 675128 742710 675156 743407
rect 675312 743322 675340 745447
rect 675312 743294 675418 743322
rect 675128 742682 675340 742710
rect 675312 742642 675340 742682
rect 675404 742642 675432 742696
rect 675312 742614 675432 742642
rect 674930 742520 674986 742529
rect 674930 742455 674986 742464
rect 674944 741074 674972 742455
rect 675312 742070 675432 742098
rect 675312 742030 675340 742070
rect 675128 742002 675340 742030
rect 675404 742016 675432 742070
rect 675128 741577 675156 742002
rect 675114 741568 675170 741577
rect 675114 741503 675170 741512
rect 674944 741046 675156 741074
rect 675128 740194 675156 741046
rect 675128 740166 675418 740194
rect 675298 739936 675354 739945
rect 675298 739871 675354 739880
rect 675312 738970 675340 739871
rect 675496 739401 675524 739636
rect 675482 739392 675538 739401
rect 675482 739327 675538 739336
rect 675404 738970 675432 739024
rect 675312 738942 675432 738970
rect 675206 738372 675262 738381
rect 675262 738330 675418 738358
rect 675206 738307 675262 738316
rect 675114 737080 675170 737089
rect 675114 737015 675170 737024
rect 675128 735333 675156 737015
rect 675404 735593 675432 735896
rect 675390 735584 675446 735593
rect 675390 735519 675446 735528
rect 674838 735312 674894 735321
rect 675128 735305 675418 735333
rect 674838 735247 674894 735256
rect 674852 734210 674880 735247
rect 675128 734658 675418 734686
rect 675128 734369 675156 734658
rect 675114 734360 675170 734369
rect 675114 734295 675170 734304
rect 674760 734182 674880 734210
rect 674760 733938 674788 734182
rect 674930 734088 674986 734097
rect 674930 734023 674986 734032
rect 674760 733910 674880 733938
rect 674852 731626 674880 733910
rect 674944 732850 674972 734023
rect 675128 734017 675418 734045
rect 675128 733825 675156 734017
rect 675114 733816 675170 733825
rect 675114 733751 675170 733760
rect 674944 732822 675418 732850
rect 675312 731734 675432 731762
rect 675312 731626 675340 731734
rect 674852 731598 675340 731626
rect 675404 731612 675432 731734
rect 675114 731504 675170 731513
rect 675114 731439 675170 731448
rect 674668 731386 674788 731414
rect 674378 728648 674434 728657
rect 674378 728583 674380 728592
rect 674432 728583 674434 728592
rect 674380 728554 674432 728560
rect 673918 726880 673974 726889
rect 673918 726815 673974 726824
rect 674760 726617 674788 731386
rect 675128 731218 675156 731439
rect 674944 731190 675156 731218
rect 674944 729178 674972 731190
rect 675128 730986 675418 731014
rect 675128 730561 675156 730986
rect 675114 730552 675170 730561
rect 675114 730487 675170 730496
rect 675128 730337 675418 730365
rect 675128 730153 675156 730337
rect 675114 730144 675170 730153
rect 675114 730079 675170 730088
rect 674944 729150 675418 729178
rect 683394 726880 683450 726889
rect 683394 726815 683450 726824
rect 674746 726608 674802 726617
rect 674746 726543 674802 726552
rect 681002 725792 681058 725801
rect 681002 725727 681058 725736
rect 677322 724296 677378 724305
rect 677322 724231 677324 724240
rect 677376 724231 677378 724240
rect 677324 724202 677376 724208
rect 681016 710841 681044 725727
rect 683212 724260 683264 724266
rect 683212 724202 683264 724208
rect 676034 710832 676090 710841
rect 676034 710767 676090 710776
rect 681002 710832 681058 710841
rect 681002 710767 681058 710776
rect 676048 709617 676076 710767
rect 676034 709608 676090 709617
rect 676034 709543 676090 709552
rect 675850 709472 675906 709481
rect 675850 709407 675906 709416
rect 675864 708801 675892 709407
rect 675850 708792 675906 708801
rect 675850 708727 675906 708736
rect 683224 708393 683252 724202
rect 683210 708384 683266 708393
rect 683210 708319 683266 708328
rect 683408 706761 683436 726815
rect 683762 726472 683818 726481
rect 683762 726407 683818 726416
rect 683776 711249 683804 726407
rect 703694 717196 703722 717264
rect 704154 717196 704182 717264
rect 704614 717196 704642 717264
rect 705074 717196 705102 717264
rect 705534 717196 705562 717264
rect 705994 717196 706022 717264
rect 706454 717196 706482 717264
rect 706914 717196 706942 717264
rect 707374 717196 707402 717264
rect 707834 717196 707862 717264
rect 708294 717196 708322 717264
rect 708754 717196 708782 717264
rect 709214 717196 709242 717264
rect 683762 711240 683818 711249
rect 683762 711175 683818 711184
rect 683394 706752 683450 706761
rect 683394 706687 683450 706696
rect 674470 706344 674526 706353
rect 674470 706279 674526 706288
rect 674102 690160 674158 690169
rect 674102 690095 674158 690104
rect 673734 682680 673790 682689
rect 673734 682615 673790 682624
rect 674116 678974 674144 690095
rect 674286 687304 674342 687313
rect 674286 687239 674342 687248
rect 674116 678946 674236 678974
rect 673826 645144 673882 645153
rect 673826 645079 673882 645088
rect 673550 618624 673606 618633
rect 673550 618559 673606 618568
rect 673642 604072 673698 604081
rect 673642 604007 673698 604016
rect 673196 601666 673408 601694
rect 673196 592034 673224 601666
rect 673460 598664 673512 598670
rect 673460 598606 673512 598612
rect 673472 592385 673500 598606
rect 673458 592376 673514 592385
rect 673656 592362 673684 604007
rect 673840 598670 673868 645079
rect 674208 642161 674236 678946
rect 674300 645854 674328 687239
rect 674484 645854 674512 706279
rect 675128 698329 675418 698337
rect 675114 698320 675418 698329
rect 675170 698309 675418 698320
rect 675114 698255 675170 698264
rect 675128 697666 675418 697694
rect 675128 697241 675156 697666
rect 675114 697232 675170 697241
rect 675114 697167 675170 697176
rect 675114 696960 675170 696969
rect 675114 696895 675170 696904
rect 675128 695209 675156 696895
rect 675404 696833 675432 697035
rect 675390 696824 675446 696833
rect 675390 696759 675446 696768
rect 675128 695181 675418 695209
rect 675680 694385 675708 694620
rect 675666 694376 675722 694385
rect 675666 694311 675722 694320
rect 675128 693994 675418 694022
rect 675128 693569 675156 693994
rect 675114 693560 675170 693569
rect 675114 693495 675170 693504
rect 675312 693382 675432 693410
rect 675312 693342 675340 693382
rect 675128 693314 675340 693342
rect 675404 693328 675432 693382
rect 674930 693288 674986 693297
rect 674930 693223 674986 693232
rect 674944 690894 674972 693223
rect 675128 693025 675156 693314
rect 675114 693016 675170 693025
rect 675114 692951 675170 692960
rect 674944 690866 675418 690894
rect 675404 690169 675432 690336
rect 675390 690160 675446 690169
rect 675390 690095 675446 690104
rect 675312 689710 675432 689738
rect 675312 689670 675340 689710
rect 674668 689642 675340 689670
rect 675404 689656 675432 689710
rect 674300 645826 674420 645854
rect 674484 645826 674604 645854
rect 674194 642152 674250 642161
rect 674392 642138 674420 645826
rect 674392 642110 674512 642138
rect 674194 642087 674250 642096
rect 674010 641744 674066 641753
rect 674010 641679 674066 641688
rect 673828 598664 673880 598670
rect 673828 598606 673880 598612
rect 673826 598360 673882 598369
rect 673826 598295 673882 598304
rect 673840 592482 673868 598295
rect 673828 592476 673880 592482
rect 673828 592418 673880 592424
rect 673656 592334 673868 592362
rect 673458 592311 673514 592320
rect 673552 592204 673604 592210
rect 673552 592146 673604 592152
rect 673196 592006 673408 592034
rect 673182 580816 673238 580825
rect 673182 580751 673238 580760
rect 673196 579873 673224 580751
rect 673182 579864 673238 579873
rect 673182 579799 673238 579808
rect 673184 579080 673236 579086
rect 673184 579022 673236 579028
rect 673196 573345 673224 579022
rect 673182 573336 673238 573345
rect 673182 573271 673238 573280
rect 673182 560144 673238 560153
rect 673182 560079 673238 560088
rect 672998 530632 673054 530641
rect 672998 530567 673054 530576
rect 672814 530224 672870 530233
rect 672814 530159 672870 530168
rect 672630 490104 672686 490113
rect 672630 490039 672686 490048
rect 673196 484809 673224 560079
rect 673182 484800 673238 484809
rect 673182 484735 673238 484744
rect 673380 456794 673408 592006
rect 673564 558906 673592 592146
rect 673840 592090 673868 592334
rect 673472 558878 673592 558906
rect 673656 592062 673868 592090
rect 673472 558090 673500 558878
rect 673656 558346 673684 592062
rect 674024 591297 674052 641679
rect 674484 641050 674512 642110
rect 674116 641022 674512 641050
rect 674116 636194 674144 641022
rect 674286 640792 674342 640801
rect 674576 640778 674604 645826
rect 674342 640750 674604 640778
rect 674286 640727 674342 640736
rect 674470 636304 674526 636313
rect 674470 636239 674526 636248
rect 674116 636166 674236 636194
rect 674208 635769 674236 636166
rect 674194 635760 674250 635769
rect 674194 635695 674250 635704
rect 674194 597408 674250 597417
rect 674194 597343 674250 597352
rect 674010 591288 674066 591297
rect 674010 591223 674066 591232
rect 673644 558340 673696 558346
rect 673644 558282 673696 558288
rect 674010 558104 674066 558113
rect 673472 558062 673684 558090
rect 673656 557870 673684 558062
rect 674010 558039 674066 558048
rect 673826 557968 673882 557977
rect 673826 557903 673882 557912
rect 673644 557864 673696 557870
rect 673644 557806 673696 557812
rect 673644 557728 673696 557734
rect 673696 557676 673776 557682
rect 673644 557670 673776 557676
rect 673656 557654 673776 557670
rect 673552 557456 673604 557462
rect 673472 557404 673552 557410
rect 673472 557398 673604 557404
rect 673472 557382 673592 557398
rect 673472 543734 673500 557382
rect 673748 549254 673776 557654
rect 673656 549226 673776 549254
rect 673656 545873 673684 549226
rect 673642 545864 673698 545873
rect 673642 545799 673698 545808
rect 673472 543706 673684 543734
rect 673656 528329 673684 543706
rect 673642 528320 673698 528329
rect 673642 528255 673698 528264
rect 673840 486169 673868 557903
rect 674024 487257 674052 558039
rect 674208 547097 674236 597343
rect 674484 589937 674512 636239
rect 674668 623257 674696 689642
rect 674930 689344 674986 689353
rect 674930 689279 674986 689288
rect 674944 688922 674972 689279
rect 675114 689072 675170 689081
rect 675170 689030 675418 689058
rect 675114 689007 675170 689016
rect 674944 688894 675156 688922
rect 674930 688664 674986 688673
rect 674930 688599 674986 688608
rect 674944 685998 674972 688599
rect 675128 686678 675156 688894
rect 675312 687806 675418 687834
rect 675312 687313 675340 687806
rect 675298 687304 675354 687313
rect 675298 687239 675354 687248
rect 675128 686650 675340 686678
rect 675312 686610 675340 686650
rect 675404 686610 675432 686664
rect 675312 686582 675432 686610
rect 674944 685970 675418 685998
rect 675114 685808 675170 685817
rect 675114 685743 675170 685752
rect 675128 676214 675156 685743
rect 675496 685001 675524 685372
rect 675482 684992 675538 685001
rect 675482 684927 675538 684936
rect 675312 684134 675418 684162
rect 675312 680105 675340 684134
rect 683118 682680 683174 682689
rect 683118 682615 683174 682624
rect 675298 680096 675354 680105
rect 675298 680031 675354 680040
rect 675128 676186 675248 676214
rect 674838 668808 674894 668817
rect 674838 668743 674894 668752
rect 674852 668273 674880 668743
rect 674838 668264 674894 668273
rect 674838 668199 674894 668208
rect 674838 664728 674894 664737
rect 674838 664663 674894 664672
rect 674852 664193 674880 664663
rect 674838 664184 674894 664193
rect 674838 664119 674894 664128
rect 674838 662280 674894 662289
rect 674838 662215 674894 662224
rect 674852 661745 674880 662215
rect 674838 661736 674894 661745
rect 674838 661671 674894 661680
rect 675220 650162 675248 676186
rect 676494 670304 676550 670313
rect 676494 670239 676550 670248
rect 676770 670304 676826 670313
rect 676770 670239 676826 670248
rect 676508 669905 676536 670239
rect 676494 669896 676550 669905
rect 676494 669831 676550 669840
rect 676784 669089 676812 670239
rect 676770 669080 676826 669089
rect 676770 669015 676826 669024
rect 676494 665816 676550 665825
rect 676494 665751 676550 665760
rect 676508 665009 676536 665751
rect 676494 665000 676550 665009
rect 676494 664935 676550 664944
rect 683132 662969 683160 682615
rect 683302 682408 683358 682417
rect 683302 682343 683358 682352
rect 683316 667049 683344 682343
rect 683486 681048 683542 681057
rect 683486 680983 683542 680992
rect 683302 667040 683358 667049
rect 683302 666975 683358 666984
rect 683500 664193 683528 680983
rect 703694 671908 703722 672044
rect 704154 671908 704182 672044
rect 704614 671908 704642 672044
rect 705074 671908 705102 672044
rect 705534 671908 705562 672044
rect 705994 671908 706022 672044
rect 706454 671908 706482 672044
rect 706914 671908 706942 672044
rect 707374 671908 707402 672044
rect 707834 671908 707862 672044
rect 708294 671908 708322 672044
rect 708754 671908 708782 672044
rect 709214 671908 709242 672044
rect 683486 664184 683542 664193
rect 683486 664119 683542 664128
rect 683118 662960 683174 662969
rect 683118 662895 683174 662904
rect 675390 660240 675446 660249
rect 675390 660175 675446 660184
rect 675404 659705 675432 660175
rect 675390 659696 675446 659705
rect 675390 659631 675446 659640
rect 675390 654256 675446 654265
rect 675390 654191 675446 654200
rect 675404 654134 675432 654191
rect 675312 654106 675432 654134
rect 675312 653018 675340 654106
rect 675312 652990 675432 653018
rect 675404 652460 675432 652990
rect 675588 652905 675616 653140
rect 675574 652896 675630 652905
rect 675574 652831 675630 652840
rect 675588 651545 675616 651848
rect 675574 651536 675630 651545
rect 675574 651471 675630 651480
rect 675220 650134 675340 650162
rect 675312 649994 675340 650134
rect 674852 649966 675340 649994
rect 674852 638217 674880 649966
rect 675404 649618 675432 650012
rect 674944 649590 675432 649618
rect 674944 647234 674972 649590
rect 675404 648961 675432 649468
rect 675390 648952 675446 648961
rect 675390 648887 675446 648896
rect 675128 648774 675418 648802
rect 675128 648689 675156 648774
rect 675114 648680 675170 648689
rect 675114 648615 675170 648624
rect 675404 647873 675432 648176
rect 675390 647864 675446 647873
rect 675390 647799 675446 647808
rect 674944 647206 675064 647234
rect 675036 645833 675064 647206
rect 675022 645824 675078 645833
rect 675022 645759 675078 645768
rect 675128 645646 675418 645674
rect 675128 645561 675156 645646
rect 675114 645552 675170 645561
rect 675114 645487 675170 645496
rect 675114 645144 675170 645153
rect 675170 645102 675418 645130
rect 675114 645079 675170 645088
rect 675772 644337 675800 644475
rect 675758 644328 675814 644337
rect 675758 644263 675814 644272
rect 675114 643920 675170 643929
rect 675114 643855 675170 643864
rect 675128 641458 675156 643855
rect 675312 643810 675418 643838
rect 675312 643521 675340 643810
rect 675298 643512 675354 643521
rect 675298 643447 675354 643456
rect 675312 642621 675418 642649
rect 675312 641753 675340 642621
rect 675298 641744 675354 641753
rect 675298 641679 675354 641688
rect 675128 641430 675418 641458
rect 675128 640781 675418 640809
rect 675128 640529 675156 640781
rect 675114 640520 675170 640529
rect 675114 640455 675170 640464
rect 675404 639849 675432 640152
rect 675390 639840 675446 639849
rect 675390 639775 675446 639784
rect 675496 638761 675524 638928
rect 675482 638752 675538 638761
rect 675482 638687 675538 638696
rect 674838 638208 674894 638217
rect 674838 638143 674894 638152
rect 675758 638208 675814 638217
rect 675758 638143 675814 638152
rect 674838 637936 674894 637945
rect 674838 637871 674894 637880
rect 674852 637786 674880 637871
rect 674852 637758 675156 637786
rect 674930 637664 674986 637673
rect 674930 637599 674986 637608
rect 674944 636217 674972 637599
rect 674930 636208 674986 636217
rect 674930 636143 674986 636152
rect 675128 626534 675156 637758
rect 675298 637664 675354 637673
rect 675298 637599 675354 637608
rect 675312 631417 675340 637599
rect 675772 637574 675800 638143
rect 676034 637936 676090 637945
rect 676034 637871 676090 637880
rect 675772 637546 675892 637574
rect 675482 636168 675538 636177
rect 675482 636103 675538 636112
rect 675298 631408 675354 631417
rect 675298 631343 675354 631352
rect 675496 626534 675524 636103
rect 675864 634234 675892 637546
rect 675852 634228 675904 634234
rect 675852 634170 675904 634176
rect 676048 631417 676076 637871
rect 683394 636848 683450 636857
rect 683394 636783 683450 636792
rect 683210 635488 683266 635497
rect 683210 635423 683266 635432
rect 683224 634814 683252 635423
rect 683408 634814 683436 636783
rect 683224 634786 683344 634814
rect 683408 634786 683528 634814
rect 682384 634228 682436 634234
rect 682384 634170 682436 634176
rect 676034 631408 676090 631417
rect 676034 631343 676090 631352
rect 674852 626506 675156 626534
rect 675220 626506 675524 626534
rect 674654 623248 674710 623257
rect 674654 623183 674710 623192
rect 674852 618338 674880 626506
rect 674852 618310 675064 618338
rect 674838 608696 674894 608705
rect 674838 608631 674894 608640
rect 674852 607073 674880 608631
rect 674838 607064 674894 607073
rect 674838 606999 674894 607008
rect 674838 601760 674894 601769
rect 674838 601695 674894 601704
rect 674852 600545 674880 601695
rect 674838 600536 674894 600545
rect 674838 600471 674894 600480
rect 674654 599856 674710 599865
rect 674654 599791 674710 599800
rect 674470 589928 674526 589937
rect 674470 589863 674526 589872
rect 674378 554432 674434 554441
rect 674378 554367 674434 554376
rect 674194 547088 674250 547097
rect 674194 547023 674250 547032
rect 674194 529408 674250 529417
rect 674194 529343 674250 529352
rect 674208 528601 674236 529343
rect 674194 528592 674250 528601
rect 674194 528527 674250 528536
rect 674010 487248 674066 487257
rect 674010 487183 674066 487192
rect 673826 486160 673882 486169
rect 673826 486095 673882 486104
rect 674392 483585 674420 554367
rect 674668 526969 674696 599791
rect 675036 599706 675064 618310
rect 675220 618254 675248 626506
rect 675574 623248 675630 623257
rect 675574 623183 675630 623192
rect 674944 599678 675064 599706
rect 675128 618226 675248 618254
rect 674944 599298 674972 599678
rect 675128 599570 675156 618226
rect 675588 617817 675616 623183
rect 675852 622872 675904 622878
rect 675850 622840 675852 622849
rect 676680 622872 676732 622878
rect 675904 622840 675906 622849
rect 675850 622775 675906 622784
rect 676402 622840 676458 622849
rect 676402 622775 676458 622784
rect 676678 622840 676680 622849
rect 676732 622840 676734 622849
rect 676678 622775 676734 622784
rect 676034 622568 676090 622577
rect 676416 622554 676444 622775
rect 676090 622526 676444 622554
rect 676034 622503 676090 622512
rect 682396 622033 682424 634170
rect 683118 628552 683174 628561
rect 683118 628487 683174 628496
rect 683132 625705 683160 628487
rect 683118 625696 683174 625705
rect 683118 625631 683174 625640
rect 682382 622024 682438 622033
rect 682382 621959 682438 621968
rect 676494 621616 676550 621625
rect 676494 621551 676550 621560
rect 676508 621217 676536 621551
rect 676494 621208 676550 621217
rect 676494 621143 676550 621152
rect 676494 620392 676550 620401
rect 676494 620327 676550 620336
rect 676508 619993 676536 620327
rect 676494 619984 676550 619993
rect 676494 619919 676550 619928
rect 683316 618361 683344 634786
rect 683302 618352 683358 618361
rect 683302 618287 683358 618296
rect 675574 617808 675630 617817
rect 675574 617743 675630 617752
rect 683500 617137 683528 634786
rect 703694 626892 703722 627028
rect 704154 626892 704182 627028
rect 704614 626892 704642 627028
rect 705074 626892 705102 627028
rect 705534 626892 705562 627028
rect 705994 626892 706022 627028
rect 706454 626892 706482 627028
rect 706914 626892 706942 627028
rect 707374 626892 707402 627028
rect 707834 626892 707862 627028
rect 708294 626892 708322 627028
rect 708754 626892 708782 627028
rect 709214 626892 709242 627028
rect 683486 617128 683542 617137
rect 683486 617063 683542 617072
rect 675496 607889 675524 608124
rect 675482 607880 675538 607889
rect 675482 607815 675538 607824
rect 675312 607465 675418 607493
rect 675312 607345 675340 607465
rect 675298 607336 675354 607345
rect 675298 607271 675354 607280
rect 675298 607064 675354 607073
rect 675298 606999 675354 607008
rect 675312 606846 675340 606999
rect 675312 606818 675418 606846
rect 675312 604982 675418 605010
rect 675312 604897 675340 604982
rect 675298 604888 675354 604897
rect 675298 604823 675354 604832
rect 675312 604438 675418 604466
rect 675312 604353 675340 604438
rect 675298 604344 675354 604353
rect 675298 604279 675354 604288
rect 675390 604072 675446 604081
rect 675390 604007 675446 604016
rect 675404 603772 675432 604007
rect 675298 603392 675354 603401
rect 675298 603327 675354 603336
rect 675312 601202 675340 603327
rect 675496 602993 675524 603160
rect 675482 602984 675538 602993
rect 675482 602919 675538 602928
rect 675312 601174 675432 601202
rect 675404 600644 675432 601174
rect 675298 600536 675354 600545
rect 675298 600471 675354 600480
rect 675128 599542 675248 599570
rect 675220 599434 675248 599542
rect 675312 599502 675340 600471
rect 675496 599865 675524 600100
rect 675482 599856 675538 599865
rect 675482 599791 675538 599800
rect 675312 599474 675418 599502
rect 674852 599270 674972 599298
rect 675128 599406 675248 599434
rect 674852 592657 674880 599270
rect 674838 592648 674894 592657
rect 674838 592583 674894 592592
rect 675128 592034 675156 599406
rect 675298 599312 675354 599321
rect 675298 599247 675354 599256
rect 675312 596442 675340 599247
rect 675496 598505 675524 598808
rect 675482 598496 675538 598505
rect 675482 598431 675538 598440
rect 675496 597417 675524 597652
rect 675482 597408 675538 597417
rect 675482 597343 675538 597352
rect 675312 596414 675418 596442
rect 675404 595377 675432 595816
rect 675390 595368 675446 595377
rect 675390 595303 675446 595312
rect 675496 594833 675524 595136
rect 675482 594824 675538 594833
rect 675482 594759 675538 594768
rect 675404 593473 675432 593980
rect 675390 593464 675446 593473
rect 675390 593399 675446 593408
rect 675574 593192 675630 593201
rect 675574 593127 675630 593136
rect 675298 592104 675354 592113
rect 675298 592039 675354 592048
rect 674944 592006 675156 592034
rect 674944 586514 674972 592006
rect 675312 586514 675340 592039
rect 674944 586486 675156 586514
rect 675312 586486 675432 586514
rect 675128 575521 675156 586486
rect 675114 575512 675170 575521
rect 675114 575447 675170 575456
rect 675404 572714 675432 586486
rect 675588 586265 675616 593127
rect 676034 592920 676090 592929
rect 676034 592855 676090 592864
rect 675850 592648 675906 592657
rect 675850 592583 675906 592592
rect 675864 591394 675892 592583
rect 675852 591388 675904 591394
rect 675852 591330 675904 591336
rect 675574 586256 675630 586265
rect 675574 586191 675630 586200
rect 676048 576609 676076 592855
rect 683394 592648 683450 592657
rect 683394 592583 683450 592592
rect 681002 591696 681058 591705
rect 681002 591631 681058 591640
rect 676034 576600 676090 576609
rect 676034 576535 676090 576544
rect 681016 576065 681044 591631
rect 682384 591388 682436 591394
rect 682384 591330 682436 591336
rect 681002 576056 681058 576065
rect 681002 575991 681058 576000
rect 676034 575104 676090 575113
rect 676034 575039 676090 575048
rect 676048 573753 676076 575039
rect 676034 573744 676090 573753
rect 676034 573679 676090 573688
rect 675220 572686 675432 572714
rect 674838 571160 674894 571169
rect 674838 571095 674894 571104
rect 674852 570353 674880 571095
rect 674838 570344 674894 570353
rect 674838 570279 674894 570288
rect 674838 559600 674894 559609
rect 674838 559535 674894 559544
rect 674852 553058 674880 559535
rect 675022 557560 675078 557569
rect 675022 557495 675078 557504
rect 675036 555801 675064 557495
rect 675022 555792 675078 555801
rect 675022 555727 675078 555736
rect 675220 554146 675248 572686
rect 682396 570761 682424 591330
rect 683408 571985 683436 592583
rect 683670 591288 683726 591297
rect 683670 591223 683726 591232
rect 683684 573209 683712 591223
rect 683854 589928 683910 589937
rect 683854 589863 683910 589872
rect 683868 576473 683896 589863
rect 703694 581740 703722 581876
rect 704154 581740 704182 581876
rect 704614 581740 704642 581876
rect 705074 581740 705102 581876
rect 705534 581740 705562 581876
rect 705994 581740 706022 581876
rect 706454 581740 706482 581876
rect 706914 581740 706942 581876
rect 707374 581740 707402 581876
rect 707834 581740 707862 581876
rect 708294 581740 708322 581876
rect 708754 581740 708782 581876
rect 709214 581740 709242 581876
rect 683854 576464 683910 576473
rect 683854 576399 683910 576408
rect 683670 573200 683726 573209
rect 683670 573135 683726 573144
rect 683394 571976 683450 571985
rect 683394 571911 683450 571920
rect 682382 570752 682438 570761
rect 682382 570687 682438 570696
rect 675390 564496 675446 564505
rect 675390 564431 675446 564440
rect 675404 564346 675432 564431
rect 675312 564318 675432 564346
rect 675312 562306 675340 564318
rect 675496 562737 675524 562904
rect 675482 562728 675538 562737
rect 675482 562663 675538 562672
rect 675312 562278 675418 562306
rect 675496 561241 675524 561612
rect 675482 561232 675538 561241
rect 675482 561167 675538 561176
rect 675390 560144 675446 560153
rect 675390 560079 675446 560088
rect 675404 559994 675432 560079
rect 675312 559966 675432 559994
rect 675312 559246 675340 559966
rect 675496 559609 675524 559776
rect 675482 559600 675538 559609
rect 675482 559535 675538 559544
rect 675312 559218 675418 559246
rect 675404 558113 675432 558620
rect 675390 558104 675446 558113
rect 675390 558039 675446 558048
rect 675404 557841 675432 557940
rect 675390 557832 675446 557841
rect 675390 557767 675446 557776
rect 675482 557560 675538 557569
rect 675312 557518 675482 557546
rect 675312 554933 675340 557518
rect 675482 557495 675538 557504
rect 675482 555792 675538 555801
rect 675482 555727 675538 555736
rect 675496 555492 675524 555727
rect 675312 554905 675418 554933
rect 675390 554432 675446 554441
rect 675390 554367 675446 554376
rect 675404 554268 675432 554367
rect 675036 554118 675248 554146
rect 675036 553394 675064 554118
rect 675206 554024 675262 554033
rect 675206 553959 675262 553968
rect 675036 553366 675156 553394
rect 674760 553030 674880 553058
rect 674760 552786 674788 553030
rect 674760 552758 674880 552786
rect 674852 546417 674880 552758
rect 675128 550225 675156 553366
rect 675220 552786 675248 553959
rect 675404 553489 675432 553656
rect 675390 553480 675446 553489
rect 675390 553415 675446 553424
rect 675220 552758 675340 552786
rect 675312 551253 675340 552758
rect 675482 552664 675538 552673
rect 675482 552599 675538 552608
rect 675496 552432 675524 552599
rect 675312 551225 675418 551253
rect 675772 550361 675800 550596
rect 675758 550352 675814 550361
rect 675758 550287 675814 550296
rect 675114 550216 675170 550225
rect 675114 550151 675170 550160
rect 675036 549937 675418 549965
rect 675036 547618 675064 549937
rect 675496 548457 675524 548760
rect 675482 548448 675538 548457
rect 675482 548383 675538 548392
rect 675850 547632 675906 547641
rect 675036 547590 675248 547618
rect 674838 546408 674894 546417
rect 674838 546343 674894 546352
rect 675220 546258 675248 547590
rect 675850 547567 675906 547576
rect 678242 547632 678298 547641
rect 678242 547567 678298 547576
rect 675864 546514 675892 547567
rect 675852 546508 675904 546514
rect 675852 546450 675904 546456
rect 675666 546408 675722 546417
rect 675666 546343 675722 546352
rect 675036 546230 675248 546258
rect 674838 545592 674894 545601
rect 674838 545527 674894 545536
rect 674852 540974 674880 545527
rect 674852 540946 674972 540974
rect 674654 526960 674710 526969
rect 674654 526895 674710 526904
rect 674944 509234 674972 540946
rect 674852 509206 674972 509234
rect 674852 502625 674880 509206
rect 674838 502616 674894 502625
rect 674838 502551 674894 502560
rect 675036 502466 675064 546230
rect 675298 546136 675354 546145
rect 675298 546071 675354 546080
rect 675312 545986 675340 546071
rect 674944 502438 675064 502466
rect 675128 545958 675340 545986
rect 674944 502217 674972 502438
rect 674930 502208 674986 502217
rect 674930 502143 674986 502152
rect 675128 487665 675156 545958
rect 675680 545578 675708 546343
rect 675312 545550 675708 545578
rect 675114 487656 675170 487665
rect 675114 487591 675170 487600
rect 675312 486441 675340 545550
rect 675758 534712 675814 534721
rect 675758 534647 675814 534656
rect 675772 534109 675800 534647
rect 675758 534100 675814 534109
rect 675758 534035 675814 534044
rect 675758 532536 675814 532545
rect 675758 532471 675814 532480
rect 675772 531661 675800 532471
rect 675758 531652 675814 531661
rect 675758 531587 675814 531596
rect 678256 531049 678284 547567
rect 683578 547360 683634 547369
rect 683578 547295 683634 547304
rect 681004 546508 681056 546514
rect 681004 546450 681056 546456
rect 681016 531457 681044 546450
rect 683302 545728 683358 545737
rect 683302 545663 683358 545672
rect 681002 531448 681058 531457
rect 681002 531383 681058 531392
rect 678242 531040 678298 531049
rect 678242 530975 678298 530984
rect 676034 530632 676090 530641
rect 676034 530567 676090 530576
rect 676048 528805 676076 530567
rect 676034 528796 676090 528805
rect 676034 528731 676090 528740
rect 683316 526561 683344 545663
rect 683592 527377 683620 547295
rect 683854 547088 683910 547097
rect 683854 547023 683910 547032
rect 683868 528193 683896 547023
rect 703694 536724 703722 536860
rect 704154 536724 704182 536860
rect 704614 536724 704642 536860
rect 705074 536724 705102 536860
rect 705534 536724 705562 536860
rect 705994 536724 706022 536860
rect 706454 536724 706482 536860
rect 706914 536724 706942 536860
rect 707374 536724 707402 536860
rect 707834 536724 707862 536860
rect 708294 536724 708322 536860
rect 708754 536724 708782 536860
rect 709214 536724 709242 536860
rect 683854 528184 683910 528193
rect 683854 528119 683910 528128
rect 683578 527368 683634 527377
rect 683578 527303 683634 527312
rect 683302 526552 683358 526561
rect 683302 526487 683358 526496
rect 683118 525736 683174 525745
rect 683118 525671 683174 525680
rect 677874 524512 677930 524521
rect 677874 524447 677930 524456
rect 676864 520328 676916 520334
rect 676864 520270 676916 520276
rect 675852 518832 675904 518838
rect 675852 518774 675904 518780
rect 675864 509234 675892 518774
rect 675496 509206 675892 509234
rect 675298 486432 675354 486441
rect 675298 486367 675354 486376
rect 674378 483576 674434 483585
rect 674378 483511 674434 483520
rect 673380 456766 673500 456794
rect 672906 456512 672962 456521
rect 672906 456447 672962 456456
rect 671986 455696 672042 455705
rect 671986 455631 672042 455640
rect 672078 455152 672134 455161
rect 672078 455087 672080 455096
rect 672132 455087 672134 455096
rect 672080 455058 672132 455064
rect 672920 454714 672948 456447
rect 673472 455870 673500 456766
rect 673946 456240 674002 456249
rect 673946 456175 673948 456184
rect 674000 456175 674002 456184
rect 673948 456146 674000 456152
rect 673828 456000 673880 456006
rect 673826 455968 673828 455977
rect 673880 455968 673882 455977
rect 673826 455903 673882 455912
rect 673460 455864 673512 455870
rect 673460 455806 673512 455812
rect 673596 455696 673652 455705
rect 673596 455631 673598 455640
rect 673650 455631 673652 455640
rect 673598 455602 673650 455608
rect 673274 455424 673330 455433
rect 673274 455359 673276 455368
rect 673328 455359 673330 455368
rect 673276 455330 673328 455336
rect 673386 455288 673442 455297
rect 673386 455223 673388 455232
rect 673440 455223 673442 455232
rect 673388 455194 673440 455200
rect 675496 454889 675524 509206
rect 676034 502616 676090 502625
rect 676034 502551 676090 502560
rect 676048 502382 676076 502551
rect 676036 502376 676088 502382
rect 676036 502318 676088 502324
rect 675850 502208 675906 502217
rect 675850 502143 675906 502152
rect 675864 500954 675892 502143
rect 676402 500984 676458 500993
rect 675852 500948 675904 500954
rect 676402 500919 676458 500928
rect 675852 500890 675904 500896
rect 676416 495434 676444 500919
rect 676876 495434 676904 520270
rect 677888 518838 677916 524447
rect 683132 520334 683160 525671
rect 683120 520328 683172 520334
rect 683120 520270 683172 520276
rect 677876 518832 677928 518838
rect 677876 518774 677928 518780
rect 683118 503704 683174 503713
rect 683118 503639 683174 503648
rect 678244 502376 678296 502382
rect 678244 502318 678296 502324
rect 676416 495406 676812 495434
rect 676876 495406 676996 495434
rect 676034 488064 676090 488073
rect 676034 487999 676090 488008
rect 675850 487248 675906 487257
rect 675850 487183 675906 487192
rect 675666 486160 675722 486169
rect 675666 486095 675722 486104
rect 675680 483177 675708 486095
rect 675864 484401 675892 487183
rect 675850 484392 675906 484401
rect 675850 484327 675906 484336
rect 675666 483168 675722 483177
rect 675666 483103 675722 483112
rect 675666 481944 675722 481953
rect 675666 481879 675722 481888
rect 673044 454880 673100 454889
rect 673044 454815 673046 454824
rect 673098 454815 673100 454824
rect 675482 454880 675538 454889
rect 675482 454815 675538 454824
rect 673046 454786 673098 454792
rect 672908 454708 672960 454714
rect 672908 454650 672960 454656
rect 673164 454640 673216 454646
rect 673162 454608 673164 454617
rect 673216 454608 673218 454617
rect 673162 454543 673218 454552
rect 672816 454232 672868 454238
rect 672814 454200 672816 454209
rect 672868 454200 672870 454209
rect 672814 454135 672870 454144
rect 672724 453960 672776 453966
rect 672722 453928 672724 453937
rect 672776 453928 672778 453937
rect 672722 453863 672778 453872
rect 675206 453928 675262 453937
rect 675680 453914 675708 481879
rect 675850 480720 675906 480729
rect 675850 480655 675906 480664
rect 675864 454209 675892 480655
rect 675850 454200 675906 454209
rect 675850 454135 675906 454144
rect 675262 453886 675708 453914
rect 675206 453863 675262 453872
rect 676048 453801 676076 487999
rect 676218 475416 676274 475425
rect 676218 475351 676274 475360
rect 676232 455977 676260 475351
rect 676218 455968 676274 455977
rect 676218 455903 676274 455912
rect 676784 454617 676812 495406
rect 676968 456521 676996 495406
rect 677506 492824 677562 492833
rect 677506 492759 677562 492768
rect 677520 491162 677548 492759
rect 677508 491156 677560 491162
rect 677508 491098 677560 491104
rect 678256 486849 678284 502318
rect 681004 500948 681056 500954
rect 681004 500890 681056 500896
rect 678242 486840 678298 486849
rect 678242 486775 678298 486784
rect 681016 481574 681044 500890
rect 683132 487257 683160 503639
rect 683302 494728 683358 494737
rect 683302 494663 683358 494672
rect 683316 491337 683344 494663
rect 703694 492796 703722 492864
rect 704154 492796 704182 492864
rect 704614 492796 704642 492864
rect 705074 492796 705102 492864
rect 705534 492796 705562 492864
rect 705994 492796 706022 492864
rect 706454 492796 706482 492864
rect 706914 492796 706942 492864
rect 707374 492796 707402 492864
rect 707834 492796 707862 492864
rect 708294 492796 708322 492864
rect 708754 492796 708782 492864
rect 709214 492796 709242 492864
rect 683302 491328 683358 491337
rect 683302 491263 683358 491272
rect 683304 491156 683356 491162
rect 683304 491098 683356 491104
rect 683118 487248 683174 487257
rect 683118 487183 683174 487192
rect 683316 482769 683344 491098
rect 683302 482760 683358 482769
rect 683302 482695 683358 482704
rect 681004 481568 681056 481574
rect 683120 481568 683172 481574
rect 681004 481510 681056 481516
rect 683118 481536 683120 481545
rect 683172 481536 683174 481545
rect 683118 481471 683174 481480
rect 676954 456512 677010 456521
rect 676954 456447 677010 456456
rect 676770 454608 676826 454617
rect 676770 454543 676826 454552
rect 676034 453792 676090 453801
rect 676034 453727 676090 453736
rect 683302 411904 683358 411913
rect 683302 411839 683358 411848
rect 676034 410544 676090 410553
rect 676034 410479 676090 410488
rect 674194 402248 674250 402257
rect 674194 402183 674250 402192
rect 671802 401704 671858 401713
rect 671802 401639 671858 401648
rect 672814 400480 672870 400489
rect 672814 400415 672870 400424
rect 672630 393952 672686 393961
rect 672630 393887 672686 393896
rect 671986 393544 672042 393553
rect 671986 393479 672042 393488
rect 671802 347712 671858 347721
rect 671802 347647 671858 347656
rect 670606 347304 670662 347313
rect 670606 347239 670662 347248
rect 669962 275360 670018 275369
rect 669962 275295 670018 275304
rect 670422 261624 670478 261633
rect 670422 261559 670478 261568
rect 670238 260400 670294 260409
rect 670238 260335 670294 260344
rect 670252 240281 670280 260335
rect 670436 247081 670464 261559
rect 670422 247072 670478 247081
rect 670422 247007 670478 247016
rect 670238 240272 670294 240281
rect 670238 240207 670294 240216
rect 669962 237144 670018 237153
rect 669962 237079 670018 237088
rect 669410 234968 669466 234977
rect 669410 234903 669466 234912
rect 669424 224954 669452 234903
rect 669596 234388 669648 234394
rect 669596 234330 669648 234336
rect 669424 224926 669544 224954
rect 669226 206544 669282 206553
rect 669226 206479 669282 206488
rect 669516 205634 669544 224926
rect 669424 205606 669544 205634
rect 669424 200114 669452 205606
rect 669056 200086 669176 200114
rect 668872 193186 668992 193214
rect 668872 183554 668900 193186
rect 669148 188494 669176 200086
rect 669240 200086 669452 200114
rect 669240 192522 669268 200086
rect 669240 192506 669360 192522
rect 669240 192500 669372 192506
rect 669240 192494 669320 192500
rect 669320 192442 669372 192448
rect 669136 188488 669188 188494
rect 669136 188430 669188 188436
rect 669318 188456 669374 188465
rect 669318 188391 669374 188400
rect 669332 188306 669360 188391
rect 669056 188278 669360 188306
rect 668872 183526 668992 183554
rect 668964 163305 668992 183526
rect 669056 176654 669084 188278
rect 669320 188216 669372 188222
rect 669148 188164 669320 188170
rect 669148 188158 669372 188164
rect 669148 188142 669360 188158
rect 669148 177290 669176 188142
rect 669608 184550 669636 234330
rect 669780 232892 669832 232898
rect 669780 232834 669832 232840
rect 669596 184544 669648 184550
rect 669596 184486 669648 184492
rect 669286 177398 669452 177426
rect 669286 177290 669314 177398
rect 669424 177313 669452 177398
rect 669148 177262 669314 177290
rect 669410 177304 669466 177313
rect 669410 177239 669466 177248
rect 669056 176626 669268 176654
rect 669240 168201 669268 176626
rect 669792 174894 669820 232834
rect 669780 174888 669832 174894
rect 669780 174830 669832 174836
rect 669778 168328 669834 168337
rect 669778 168263 669834 168272
rect 669226 168192 669282 168201
rect 669226 168127 669282 168136
rect 669134 164248 669190 164257
rect 669134 164183 669190 164192
rect 668950 163296 669006 163305
rect 668950 163231 669006 163240
rect 668766 153504 668822 153513
rect 668766 153439 668822 153448
rect 668766 153096 668822 153105
rect 668766 153031 668822 153040
rect 668490 148608 668546 148617
rect 668490 148543 668546 148552
rect 667938 137864 667994 137873
rect 667938 137799 667994 137808
rect 667570 135960 667626 135969
rect 667570 135895 667626 135904
rect 667952 135561 667980 137799
rect 667938 135552 667994 135561
rect 667938 135487 667994 135496
rect 667018 133104 667074 133113
rect 667018 133039 667074 133048
rect 590292 131912 590344 131918
rect 590292 131854 590344 131860
rect 590106 131336 590162 131345
rect 590106 131271 590162 131280
rect 590120 131170 590148 131271
rect 590108 131164 590160 131170
rect 590108 131106 590160 131112
rect 668780 125769 668808 153031
rect 669148 143721 669176 164183
rect 669134 143712 669190 143721
rect 669134 143647 669190 143656
rect 669226 141128 669282 141137
rect 669226 141063 669282 141072
rect 669240 138825 669268 141063
rect 669226 138816 669282 138825
rect 669226 138751 669282 138760
rect 668950 128344 669006 128353
rect 668950 128279 669006 128288
rect 668766 125760 668822 125769
rect 668766 125695 668822 125704
rect 668964 120873 668992 128279
rect 669226 122224 669282 122233
rect 669226 122159 669282 122168
rect 668950 120864 669006 120873
rect 668950 120799 669006 120808
rect 667940 120760 667992 120766
rect 667940 120702 667992 120708
rect 667952 119241 667980 120702
rect 667938 119232 667994 119241
rect 667938 119167 667994 119176
rect 667940 118108 667992 118114
rect 667940 118050 667992 118056
rect 667952 117609 667980 118050
rect 667938 117600 667994 117609
rect 667938 117535 667994 117544
rect 669240 114345 669268 122159
rect 669792 120766 669820 168263
rect 669976 160070 670004 237079
rect 670238 236872 670294 236881
rect 670238 236807 670294 236816
rect 670252 233034 670280 236807
rect 670620 234614 670648 347239
rect 671816 325689 671844 347647
rect 671802 325680 671858 325689
rect 671802 325615 671858 325624
rect 671710 261216 671766 261225
rect 671710 261151 671766 261160
rect 671526 260944 671582 260953
rect 671526 260879 671582 260888
rect 671342 256728 671398 256737
rect 671342 256663 671398 256672
rect 671068 237856 671120 237862
rect 671356 237833 671384 256663
rect 671540 246673 671568 260879
rect 671526 246664 671582 246673
rect 671526 246599 671582 246608
rect 671724 245313 671752 261151
rect 671710 245304 671766 245313
rect 671710 245239 671766 245248
rect 671068 237798 671120 237804
rect 671342 237824 671398 237833
rect 670436 234586 670648 234614
rect 670240 233028 670292 233034
rect 670240 232970 670292 232976
rect 670146 232792 670202 232801
rect 670146 232727 670202 232736
rect 670160 165238 670188 232727
rect 670436 229094 670464 234586
rect 671080 234569 671108 237798
rect 671342 237759 671398 237768
rect 671712 237584 671764 237590
rect 671712 237526 671764 237532
rect 671344 237176 671396 237182
rect 671344 237118 671396 237124
rect 671066 234560 671122 234569
rect 671066 234495 671122 234504
rect 670976 233912 671028 233918
rect 670976 233854 671028 233860
rect 670792 233368 670844 233374
rect 670792 233310 670844 233316
rect 670606 232520 670662 232529
rect 670606 232455 670662 232464
rect 670620 231854 670648 232455
rect 670344 229066 670464 229094
rect 670528 231826 670648 231854
rect 670344 223582 670372 229066
rect 670528 224890 670556 231826
rect 670804 229106 670832 233310
rect 670804 229078 670924 229106
rect 670700 226500 670752 226506
rect 670700 226442 670752 226448
rect 670712 226273 670740 226442
rect 670698 226264 670754 226273
rect 670698 226199 670754 226208
rect 670700 225480 670752 225486
rect 670698 225448 670700 225457
rect 670752 225448 670754 225457
rect 670698 225383 670754 225392
rect 670700 225072 670752 225078
rect 670698 225040 670700 225049
rect 670752 225040 670754 225049
rect 670698 224975 670754 224984
rect 670896 224954 670924 229078
rect 670988 225162 671016 233854
rect 671160 227996 671212 228002
rect 671160 227938 671212 227944
rect 671172 225729 671200 227938
rect 671158 225720 671214 225729
rect 671158 225655 671214 225664
rect 671158 225448 671214 225457
rect 671158 225383 671214 225392
rect 671172 225282 671200 225383
rect 671160 225276 671212 225282
rect 671160 225218 671212 225224
rect 670988 225134 671200 225162
rect 670896 224926 671108 224954
rect 670528 224862 670740 224890
rect 670516 223712 670568 223718
rect 670514 223680 670516 223689
rect 670568 223680 670570 223689
rect 670514 223615 670570 223624
rect 670332 223576 670384 223582
rect 670332 223518 670384 223524
rect 670712 223394 670740 224862
rect 670884 224664 670936 224670
rect 670882 224632 670884 224641
rect 670936 224632 670938 224641
rect 670882 224567 670938 224576
rect 670930 224120 670982 224126
rect 670930 224062 670982 224068
rect 670942 223961 670970 224062
rect 670928 223952 670984 223961
rect 670928 223887 670984 223896
rect 670712 223366 670832 223394
rect 670608 223304 670660 223310
rect 670608 223246 670660 223252
rect 670332 222216 670384 222222
rect 670332 222158 670384 222164
rect 670344 169726 670372 222158
rect 670620 220969 670648 223246
rect 670804 222222 670832 223366
rect 670792 222216 670844 222222
rect 670792 222158 670844 222164
rect 670790 222048 670846 222057
rect 670790 221983 670846 221992
rect 670804 221270 670832 221983
rect 670792 221264 670844 221270
rect 670792 221206 670844 221212
rect 670606 220960 670662 220969
rect 670606 220895 670662 220904
rect 670606 220688 670662 220697
rect 670606 220623 670662 220632
rect 670620 176497 670648 220623
rect 670790 220144 670846 220153
rect 670790 220079 670846 220088
rect 670606 176488 670662 176497
rect 670606 176423 670662 176432
rect 670804 175681 670832 220079
rect 671080 215294 671108 224926
rect 670988 215266 671108 215294
rect 670988 199209 671016 215266
rect 670974 199200 671030 199209
rect 670974 199135 671030 199144
rect 671172 194313 671200 225134
rect 671158 194304 671214 194313
rect 671158 194239 671214 194248
rect 670790 175672 670846 175681
rect 670790 175607 670846 175616
rect 670606 172000 670662 172009
rect 670606 171935 670662 171944
rect 670332 169720 670384 169726
rect 670332 169662 670384 169668
rect 670422 169552 670478 169561
rect 670422 169487 670478 169496
rect 670148 165232 670200 165238
rect 670148 165174 670200 165180
rect 670146 165064 670202 165073
rect 670146 164999 670202 165008
rect 669964 160064 670016 160070
rect 669964 160006 670016 160012
rect 669962 121408 670018 121417
rect 669962 121343 670018 121352
rect 669780 120760 669832 120766
rect 669780 120702 669832 120708
rect 669226 114336 669282 114345
rect 669226 114271 669282 114280
rect 590290 113384 590346 113393
rect 590290 113319 590346 113328
rect 589924 113144 589976 113150
rect 589924 113086 589976 113092
rect 589370 111752 589426 111761
rect 589370 111687 589426 111696
rect 589384 109750 589412 111687
rect 590304 111110 590332 113319
rect 669976 111450 670004 121343
rect 670160 118114 670188 164999
rect 670436 154873 670464 169487
rect 670422 154864 670478 154873
rect 670422 154799 670478 154808
rect 670620 149025 670648 171935
rect 671356 151814 671384 237118
rect 671528 237040 671580 237046
rect 671528 236982 671580 236988
rect 671540 231854 671568 236982
rect 671724 234569 671752 237526
rect 671710 234560 671766 234569
rect 671710 234495 671766 234504
rect 671712 234048 671764 234054
rect 671712 233990 671764 233996
rect 671448 231826 671568 231854
rect 671448 222194 671476 231826
rect 671724 229401 671752 233990
rect 671710 229392 671766 229401
rect 671710 229327 671766 229336
rect 671620 227656 671672 227662
rect 671620 227598 671672 227604
rect 671632 226953 671660 227598
rect 671804 227248 671856 227254
rect 671804 227190 671856 227196
rect 671816 227089 671844 227190
rect 671802 227080 671858 227089
rect 671802 227015 671858 227024
rect 671618 226944 671674 226953
rect 671618 226879 671674 226888
rect 671802 226672 671858 226681
rect 671802 226607 671804 226616
rect 671856 226607 671858 226616
rect 671804 226578 671856 226584
rect 671712 226296 671764 226302
rect 671632 226244 671712 226250
rect 671632 226238 671764 226244
rect 671632 226222 671752 226238
rect 671632 225162 671660 226222
rect 671802 226128 671858 226137
rect 671802 226063 671804 226072
rect 671856 226063 671858 226072
rect 671804 226034 671856 226040
rect 671820 225752 671872 225758
rect 671818 225720 671820 225729
rect 671872 225720 671874 225729
rect 671818 225655 671874 225664
rect 671802 225176 671858 225185
rect 671632 225134 671802 225162
rect 671802 225111 671858 225120
rect 671710 224904 671766 224913
rect 671710 224839 671766 224848
rect 671448 222166 671568 222194
rect 671540 158409 671568 222166
rect 671724 189417 671752 224839
rect 672000 211177 672028 393479
rect 672354 392320 672410 392329
rect 672354 392255 672410 392264
rect 672170 357096 672226 357105
rect 672170 357031 672226 357040
rect 672184 312497 672212 357031
rect 672170 312488 672226 312497
rect 672170 312423 672226 312432
rect 672368 235906 672396 392255
rect 672644 376281 672672 393887
rect 672630 376272 672686 376281
rect 672630 376207 672686 376216
rect 672630 356280 672686 356289
rect 672630 356215 672686 356224
rect 672644 311681 672672 356215
rect 672828 355881 672856 400415
rect 673182 399664 673238 399673
rect 673182 399599 673238 399608
rect 672998 397216 673054 397225
rect 672998 397151 673054 397160
rect 673012 378049 673040 397151
rect 672998 378040 673054 378049
rect 672998 377975 673054 377984
rect 673196 364334 673224 399599
rect 673366 396400 673422 396409
rect 673366 396335 673422 396344
rect 673380 382265 673408 396335
rect 673826 396128 673882 396137
rect 673826 396063 673882 396072
rect 673366 382256 673422 382265
rect 673366 382191 673422 382200
rect 673840 381449 673868 396063
rect 674010 395720 674066 395729
rect 674010 395655 674066 395664
rect 673826 381440 673882 381449
rect 673826 381375 673882 381384
rect 674024 375465 674052 395655
rect 674010 375456 674066 375465
rect 674010 375391 674066 375400
rect 673196 364306 673408 364334
rect 672814 355872 672870 355881
rect 672814 355807 672870 355816
rect 673182 355464 673238 355473
rect 673182 355399 673238 355408
rect 672814 351384 672870 351393
rect 672814 351319 672870 351328
rect 672828 337249 672856 351319
rect 672998 348936 673054 348945
rect 672998 348871 673054 348880
rect 672814 337240 672870 337249
rect 672814 337175 672870 337184
rect 673012 331537 673040 348871
rect 672998 331528 673054 331537
rect 672998 331463 673054 331472
rect 673196 325694 673224 355399
rect 673380 355065 673408 364306
rect 674208 357513 674236 402183
rect 674654 401432 674710 401441
rect 674654 401367 674710 401376
rect 674470 394496 674526 394505
rect 674470 394431 674526 394440
rect 674484 377777 674512 394431
rect 674470 377768 674526 377777
rect 674470 377703 674526 377712
rect 674194 357504 674250 357513
rect 674194 357439 674250 357448
rect 674668 356697 674696 401367
rect 676048 400217 676076 410479
rect 683118 406328 683174 406337
rect 683118 406263 683174 406272
rect 683132 403345 683160 406263
rect 683316 403753 683344 411839
rect 703694 404532 703722 404668
rect 704154 404532 704182 404668
rect 704614 404532 704642 404668
rect 705074 404532 705102 404668
rect 705534 404532 705562 404668
rect 705994 404532 706022 404668
rect 706454 404532 706482 404668
rect 706914 404532 706942 404668
rect 707374 404532 707402 404668
rect 707834 404532 707862 404668
rect 708294 404532 708322 404668
rect 708754 404532 708782 404668
rect 709214 404532 709242 404668
rect 683302 403744 683358 403753
rect 683302 403679 683358 403688
rect 683118 403336 683174 403345
rect 683118 403271 683174 403280
rect 676034 400208 676090 400217
rect 676034 400143 676090 400152
rect 676034 399392 676090 399401
rect 676034 399327 676090 399336
rect 675852 395752 675904 395758
rect 675036 395700 675852 395706
rect 675036 395694 675904 395700
rect 675036 395678 675892 395694
rect 675036 382582 675064 395678
rect 676048 395570 676076 399327
rect 676218 398440 676274 398449
rect 676218 398375 676274 398384
rect 675128 395542 676076 395570
rect 675128 384449 675156 395542
rect 676232 393314 676260 398375
rect 676402 398032 676458 398041
rect 676402 397967 676458 397976
rect 676416 395758 676444 397967
rect 681002 397624 681058 397633
rect 681002 397559 681058 397568
rect 676404 395752 676456 395758
rect 676404 395694 676456 395700
rect 675312 393286 676260 393314
rect 675312 386186 675340 393286
rect 681016 387705 681044 397559
rect 683026 392728 683082 392737
rect 683026 392663 683082 392672
rect 683040 389065 683068 392663
rect 683026 389056 683082 389065
rect 683026 388991 683082 389000
rect 681002 387696 681058 387705
rect 681002 387631 681058 387640
rect 675312 386158 675432 386186
rect 675404 385696 675432 386158
rect 675772 384985 675800 385084
rect 675758 384976 675814 384985
rect 675758 384911 675814 384920
rect 675128 384421 675418 384449
rect 675312 382622 675432 382650
rect 675312 382582 675340 382622
rect 675036 382554 675340 382582
rect 675404 382568 675432 382622
rect 675390 382256 675446 382265
rect 675390 382191 675446 382200
rect 675404 382024 675432 382191
rect 675114 381440 675170 381449
rect 675170 381398 675418 381426
rect 675114 381375 675170 381384
rect 675772 380633 675800 380732
rect 675758 380624 675814 380633
rect 675758 380559 675814 380568
rect 675758 378720 675814 378729
rect 675758 378655 675814 378664
rect 675772 378284 675800 378655
rect 675114 377768 675170 377777
rect 675170 377726 675340 377754
rect 675114 377703 675170 377712
rect 675312 377618 675340 377726
rect 675404 377618 675432 377740
rect 675312 377590 675432 377618
rect 675758 377360 675814 377369
rect 675758 377295 675814 377304
rect 675772 377060 675800 377295
rect 675206 376952 675262 376961
rect 675206 376887 675262 376896
rect 675220 373994 675248 376887
rect 675404 376281 675432 376448
rect 675390 376272 675446 376281
rect 675390 376207 675446 376216
rect 675390 375456 675446 375465
rect 675390 375391 675446 375400
rect 675404 375224 675432 375391
rect 675220 373966 675340 373994
rect 675312 373402 675340 373966
rect 675312 373374 675418 373402
rect 675666 373008 675722 373017
rect 675666 372943 675722 372952
rect 675680 372776 675708 372943
rect 675114 372600 675170 372609
rect 675114 372535 675170 372544
rect 675128 371566 675156 372535
rect 675128 371538 675418 371566
rect 675850 360904 675906 360913
rect 675850 360839 675906 360848
rect 675864 357921 675892 360839
rect 676034 360088 676090 360097
rect 676034 360023 676090 360032
rect 676048 358329 676076 360023
rect 703694 359380 703722 359516
rect 704154 359380 704182 359516
rect 704614 359380 704642 359516
rect 705074 359380 705102 359516
rect 705534 359380 705562 359516
rect 705994 359380 706022 359516
rect 706454 359380 706482 359516
rect 706914 359380 706942 359516
rect 707374 359380 707402 359516
rect 707834 359380 707862 359516
rect 708294 359380 708322 359516
rect 708754 359380 708782 359516
rect 709214 359380 709242 359516
rect 676034 358320 676090 358329
rect 676034 358255 676090 358264
rect 675850 357912 675906 357921
rect 675850 357847 675906 357856
rect 674654 356688 674710 356697
rect 674654 356623 674710 356632
rect 673366 355056 673422 355065
rect 673366 354991 673422 355000
rect 674654 354648 674710 354657
rect 674654 354583 674710 354592
rect 673366 353424 673422 353433
rect 673366 353359 673422 353368
rect 673380 340785 673408 353359
rect 674470 352608 674526 352617
rect 674470 352543 674526 352552
rect 674286 352200 674342 352209
rect 674286 352135 674342 352144
rect 673734 350568 673790 350577
rect 673734 350503 673790 350512
rect 673550 349480 673606 349489
rect 673550 349415 673606 349424
rect 673366 340776 673422 340785
rect 673366 340711 673422 340720
rect 673564 332761 673592 349415
rect 673550 332752 673606 332761
rect 673550 332687 673606 332696
rect 673748 331129 673776 350503
rect 674102 349752 674158 349761
rect 674102 349687 674158 349696
rect 673918 348528 673974 348537
rect 673918 348463 673974 348472
rect 673734 331120 673790 331129
rect 673734 331055 673790 331064
rect 673196 325666 673316 325694
rect 672814 312760 672870 312769
rect 672814 312695 672870 312704
rect 672630 311672 672686 311681
rect 672630 311607 672686 311616
rect 672630 304328 672686 304337
rect 672630 304263 672686 304272
rect 672644 287881 672672 304263
rect 672630 287872 672686 287881
rect 672630 287807 672686 287816
rect 672828 266937 672856 312695
rect 673090 311264 673146 311273
rect 673090 311199 673146 311208
rect 673104 267617 673132 311199
rect 673288 310865 673316 325666
rect 673274 310856 673330 310865
rect 673274 310791 673330 310800
rect 673734 305552 673790 305561
rect 673734 305487 673790 305496
rect 673550 304736 673606 304745
rect 673550 304671 673606 304680
rect 673274 303512 673330 303521
rect 673274 303447 673330 303456
rect 673090 267608 673146 267617
rect 673090 267543 673146 267552
rect 672814 266928 672870 266937
rect 672814 266863 672870 266872
rect 672814 266520 672870 266529
rect 672814 266455 672870 266464
rect 672630 257952 672686 257961
rect 672630 257887 672686 257896
rect 672644 257258 672672 257887
rect 672460 257230 672672 257258
rect 672460 253934 672488 257230
rect 672630 257136 672686 257145
rect 672630 257071 672686 257080
rect 672644 253934 672672 257071
rect 672460 253906 672580 253934
rect 672644 253906 672764 253934
rect 672552 242865 672580 253906
rect 672538 242856 672594 242865
rect 672538 242791 672594 242800
rect 672540 236496 672592 236502
rect 672540 236438 672592 236444
rect 672276 235878 672396 235906
rect 672156 230036 672208 230042
rect 672208 229984 672212 230024
rect 672156 229978 672212 229984
rect 672184 228698 672212 229978
rect 672092 228670 672212 228698
rect 672092 227712 672120 228670
rect 672276 228585 672304 235878
rect 672552 235226 672580 236438
rect 672368 235198 672580 235226
rect 672368 228834 672396 235198
rect 672540 235000 672592 235006
rect 672540 234942 672592 234948
rect 672552 230042 672580 234942
rect 672540 230036 672592 230042
rect 672540 229978 672592 229984
rect 672736 229786 672764 253906
rect 672828 231854 672856 266455
rect 673090 266112 673146 266121
rect 673090 266047 673146 266056
rect 673104 244274 673132 266047
rect 672920 244246 673132 244274
rect 672920 233730 672948 244246
rect 673092 236768 673144 236774
rect 673092 236710 673144 236716
rect 672920 233714 672994 233730
rect 672920 233708 673006 233714
rect 672920 233702 672954 233708
rect 672954 233650 673006 233656
rect 673104 233322 673132 236710
rect 673288 236586 673316 303447
rect 673564 290601 673592 304671
rect 673550 290592 673606 290601
rect 673550 290527 673606 290536
rect 673748 285569 673776 305487
rect 673734 285560 673790 285569
rect 673734 285495 673790 285504
rect 673642 259720 673698 259729
rect 673472 259678 673642 259706
rect 673472 245857 673500 259678
rect 673642 259655 673698 259664
rect 673642 258496 673698 258505
rect 673642 258431 673698 258440
rect 673458 245848 673514 245857
rect 673458 245783 673514 245792
rect 673526 237144 673582 237153
rect 673526 237079 673582 237088
rect 673540 236910 673568 237079
rect 673414 236904 673466 236910
rect 673412 236872 673414 236881
rect 673528 236904 673580 236910
rect 673466 236872 673468 236881
rect 673528 236846 673580 236852
rect 673412 236807 673468 236816
rect 673012 233294 673132 233322
rect 673196 236558 673316 236586
rect 673012 233238 673040 233294
rect 673000 233232 673052 233238
rect 673000 233174 673052 233180
rect 673196 231854 673224 236558
rect 673458 236328 673514 236337
rect 673458 236263 673514 236272
rect 673472 236162 673500 236263
rect 673460 236156 673512 236162
rect 673460 236098 673512 236104
rect 673460 235952 673512 235958
rect 673460 235894 673512 235900
rect 673472 235634 673500 235894
rect 673472 235606 673592 235634
rect 673368 235544 673420 235550
rect 673368 235486 673420 235492
rect 673380 232898 673408 235486
rect 673368 232892 673420 232898
rect 673368 232834 673420 232840
rect 673564 232642 673592 235606
rect 673380 232614 673592 232642
rect 673380 232529 673408 232614
rect 673366 232520 673422 232529
rect 673366 232455 673422 232464
rect 673460 232008 673512 232014
rect 673460 231950 673512 231956
rect 672828 231849 672948 231854
rect 672828 231840 672962 231849
rect 672828 231826 672906 231840
rect 672906 231775 672962 231784
rect 673104 231826 673224 231854
rect 672644 229758 672764 229786
rect 672368 228806 672580 228834
rect 672262 228576 672318 228585
rect 672262 228511 672318 228520
rect 672092 227684 672488 227712
rect 672172 227452 672224 227458
rect 672172 227394 672224 227400
rect 672184 227338 672212 227394
rect 672092 227310 672212 227338
rect 672092 226114 672120 227310
rect 672262 227080 672318 227089
rect 672262 227015 672264 227024
rect 672316 227015 672318 227024
rect 672264 226986 672316 226992
rect 672264 226908 672316 226914
rect 672264 226850 672316 226856
rect 672276 226545 672304 226850
rect 672262 226536 672318 226545
rect 672262 226471 672318 226480
rect 672092 226086 672212 226114
rect 672184 226001 672212 226086
rect 672170 225992 672226 226001
rect 672170 225927 672226 225936
rect 672170 224632 672226 224641
rect 672170 224567 672226 224576
rect 672184 217025 672212 224567
rect 672170 217016 672226 217025
rect 672170 216951 672226 216960
rect 672170 211440 672226 211449
rect 672170 211375 672226 211384
rect 671986 211168 672042 211177
rect 671986 211103 672042 211112
rect 672184 211018 672212 211375
rect 671908 210990 672212 211018
rect 671908 205634 671936 210990
rect 672262 210216 672318 210225
rect 672262 210151 672318 210160
rect 672078 209400 672134 209409
rect 672078 209335 672134 209344
rect 671908 205606 672028 205634
rect 672000 192409 672028 205606
rect 672092 197690 672120 209335
rect 672276 200841 672304 210151
rect 672262 200832 672318 200841
rect 672262 200767 672318 200776
rect 672092 197662 672212 197690
rect 672184 197577 672212 197662
rect 672170 197568 672226 197577
rect 672170 197503 672226 197512
rect 671986 192400 672042 192409
rect 671986 192335 672042 192344
rect 672460 191570 672488 227684
rect 672184 191542 672488 191570
rect 671710 189408 671766 189417
rect 671710 189343 671766 189352
rect 672184 188306 672212 191542
rect 672552 188465 672580 228806
rect 672644 215294 672672 229758
rect 673104 228528 673132 231826
rect 673472 231334 673500 231950
rect 673656 231849 673684 258431
rect 673752 236292 673804 236298
rect 673752 236234 673804 236240
rect 673764 236065 673792 236234
rect 673750 236056 673806 236065
rect 673750 235991 673806 236000
rect 673932 234614 673960 348463
rect 674116 335889 674144 349687
rect 674300 336705 674328 352135
rect 674286 336696 674342 336705
rect 674286 336631 674342 336640
rect 674102 335880 674158 335889
rect 674102 335815 674158 335824
rect 674484 333985 674512 352543
rect 674470 333976 674526 333985
rect 674470 333911 674526 333920
rect 674668 316034 674696 354583
rect 676034 353016 676090 353025
rect 676090 352974 676260 353002
rect 676034 352951 676090 352960
rect 675942 349208 675998 349217
rect 676232 349194 676260 352974
rect 675998 349166 676260 349194
rect 675942 349143 675998 349152
rect 675114 340776 675170 340785
rect 675114 340711 675170 340720
rect 675128 340558 675156 340711
rect 675128 340530 675340 340558
rect 675312 340490 675340 340530
rect 675404 340490 675432 340544
rect 675312 340462 675432 340490
rect 675758 340232 675814 340241
rect 675758 340167 675814 340176
rect 675772 339864 675800 340167
rect 675666 339416 675722 339425
rect 675666 339351 675722 339360
rect 675680 339252 675708 339351
rect 675574 337784 675630 337793
rect 675574 337719 675630 337728
rect 675588 337416 675616 337719
rect 675114 337240 675170 337249
rect 675114 337175 675170 337184
rect 675128 336857 675156 337175
rect 675128 336829 675418 336857
rect 675312 336178 675418 336206
rect 675312 335345 675340 336178
rect 675482 335880 675538 335889
rect 675482 335815 675538 335824
rect 675496 335580 675524 335815
rect 675298 335336 675354 335345
rect 675298 335271 675354 335280
rect 675114 333976 675170 333985
rect 675114 333911 675170 333920
rect 675128 333078 675156 333911
rect 675128 333050 675418 333078
rect 675114 332752 675170 332761
rect 675114 332687 675170 332696
rect 675128 332534 675156 332687
rect 675128 332506 675418 332534
rect 675758 332344 675814 332353
rect 675758 332279 675814 332288
rect 675772 331875 675800 332279
rect 675114 331528 675170 331537
rect 675114 331463 675170 331472
rect 675128 331242 675156 331463
rect 675128 331214 675418 331242
rect 675114 331120 675170 331129
rect 675114 331055 675170 331064
rect 675128 330049 675156 331055
rect 675128 330021 675418 330049
rect 675758 328400 675814 328409
rect 675758 328335 675814 328344
rect 675772 328168 675800 328335
rect 675128 327542 675418 327570
rect 675128 325689 675156 327542
rect 675390 326904 675446 326913
rect 675390 326839 675446 326848
rect 675404 326332 675432 326839
rect 675114 325680 675170 325689
rect 675114 325615 675170 325624
rect 674484 316006 674696 316034
rect 674484 310049 674512 316006
rect 676034 315480 676090 315489
rect 676034 315415 676090 315424
rect 676048 313313 676076 315415
rect 703694 314364 703722 314500
rect 704154 314364 704182 314500
rect 704614 314364 704642 314500
rect 705074 314364 705102 314500
rect 705534 314364 705562 314500
rect 705994 314364 706022 314500
rect 706454 314364 706482 314500
rect 706914 314364 706942 314500
rect 707374 314364 707402 314500
rect 707834 314364 707862 314500
rect 708294 314364 708322 314500
rect 708754 314364 708782 314500
rect 709214 314364 709242 314500
rect 676034 313304 676090 313313
rect 676034 313239 676090 313248
rect 674654 313032 674710 313041
rect 674654 312967 674710 312976
rect 674668 311953 674696 312967
rect 674838 312760 674894 312769
rect 674838 312695 674894 312704
rect 674852 312089 674880 312695
rect 674838 312080 674894 312089
rect 674838 312015 674894 312024
rect 674654 311944 674710 311953
rect 674654 311879 674710 311888
rect 674654 310448 674710 310457
rect 674654 310383 674710 310392
rect 674470 310040 674526 310049
rect 674470 309975 674526 309984
rect 674194 309632 674250 309641
rect 674194 309567 674250 309576
rect 674208 265033 674236 309567
rect 674378 303920 674434 303929
rect 674378 303855 674434 303864
rect 674392 286657 674420 303855
rect 674668 292574 674696 310383
rect 675114 309224 675170 309233
rect 675114 309159 675170 309168
rect 675128 302410 675156 309159
rect 676034 308408 676090 308417
rect 676090 308366 676260 308394
rect 676034 308343 676090 308352
rect 675390 308000 675446 308009
rect 675390 307935 675446 307944
rect 675036 302382 675156 302410
rect 675036 299474 675064 302382
rect 675036 299446 675156 299474
rect 674838 297120 674894 297129
rect 674838 297055 674894 297064
rect 674576 292546 674696 292574
rect 674378 286648 674434 286657
rect 674378 286583 674434 286592
rect 674576 265849 674604 292546
rect 674852 288130 674880 297055
rect 675128 294250 675156 299446
rect 675404 296721 675432 307935
rect 676232 305266 676260 308366
rect 681002 307592 681058 307601
rect 681002 307527 681058 307536
rect 678242 307184 678298 307193
rect 678242 307119 678298 307128
rect 675864 305238 676260 305266
rect 675864 302234 675892 305238
rect 675772 302206 675892 302234
rect 675390 296712 675446 296721
rect 675390 296647 675446 296656
rect 675772 296313 675800 302206
rect 675944 298104 675996 298110
rect 675944 298046 675996 298052
rect 675956 297673 675984 298046
rect 675942 297664 675998 297673
rect 675942 297599 675998 297608
rect 678256 297401 678284 307119
rect 678978 306368 679034 306377
rect 678978 306303 679034 306312
rect 678992 298110 679020 306303
rect 678980 298104 679032 298110
rect 678980 298046 679032 298052
rect 678242 297392 678298 297401
rect 678242 297327 678298 297336
rect 676218 297120 676274 297129
rect 681016 297090 681044 307527
rect 683026 302696 683082 302705
rect 683026 302631 683082 302640
rect 683040 299441 683068 302631
rect 683026 299432 683082 299441
rect 683026 299367 683082 299376
rect 676218 297055 676220 297064
rect 676272 297055 676274 297064
rect 681004 297084 681056 297090
rect 676220 297026 676272 297032
rect 681004 297026 681056 297032
rect 675758 296304 675814 296313
rect 675758 296239 675814 296248
rect 675758 295896 675814 295905
rect 675758 295831 675814 295840
rect 675772 295528 675800 295831
rect 675758 295216 675814 295225
rect 675758 295151 675814 295160
rect 675772 294879 675800 295151
rect 675128 294222 675418 294250
rect 675390 292904 675446 292913
rect 675390 292839 675446 292848
rect 675404 292400 675432 292839
rect 675574 292088 675630 292097
rect 675574 292023 675630 292032
rect 675588 291856 675616 292023
rect 675758 291544 675814 291553
rect 675758 291479 675814 291488
rect 675772 291176 675800 291479
rect 675114 290592 675170 290601
rect 675170 290550 675418 290578
rect 675114 290527 675170 290536
rect 674852 288102 675064 288130
rect 675036 288062 675064 288102
rect 675312 288102 675432 288130
rect 675312 288062 675340 288102
rect 675036 288034 675340 288062
rect 675404 288048 675432 288102
rect 675114 287872 675170 287881
rect 675114 287807 675170 287816
rect 675128 287518 675156 287807
rect 675128 287490 675418 287518
rect 675758 287056 675814 287065
rect 675758 286991 675814 287000
rect 675772 286892 675800 286991
rect 675390 286648 675446 286657
rect 675390 286583 675446 286592
rect 675404 286212 675432 286583
rect 675114 285560 675170 285569
rect 675114 285495 675170 285504
rect 675128 285070 675156 285495
rect 675128 285042 675340 285070
rect 675312 285002 675340 285042
rect 675404 285002 675432 285056
rect 675312 284974 675432 285002
rect 675758 283656 675814 283665
rect 675758 283591 675814 283600
rect 675772 283220 675800 283591
rect 675666 282840 675722 282849
rect 675666 282775 675722 282784
rect 675680 282540 675708 282775
rect 675680 281217 675708 281355
rect 675666 281208 675722 281217
rect 675666 281143 675722 281152
rect 683302 275360 683358 275369
rect 683302 275295 683358 275304
rect 683118 271144 683174 271153
rect 683118 271079 683174 271088
rect 683132 268161 683160 271079
rect 683316 268569 683344 275295
rect 703694 269348 703722 269484
rect 704154 269348 704182 269484
rect 704614 269348 704642 269484
rect 705074 269348 705102 269484
rect 705534 269348 705562 269484
rect 705994 269348 706022 269484
rect 706454 269348 706482 269484
rect 706914 269348 706942 269484
rect 707374 269348 707402 269484
rect 707834 269348 707862 269484
rect 708294 269348 708322 269484
rect 708754 269348 708782 269484
rect 709214 269348 709242 269484
rect 683302 268560 683358 268569
rect 683302 268495 683358 268504
rect 683118 268152 683174 268161
rect 683118 268087 683174 268096
rect 675022 267608 675078 267617
rect 675022 267543 675078 267552
rect 675036 266665 675064 267543
rect 675022 266656 675078 266665
rect 675022 266591 675078 266600
rect 674562 265840 674618 265849
rect 674562 265775 674618 265784
rect 674562 265432 674618 265441
rect 674562 265367 674618 265376
rect 674194 265024 674250 265033
rect 674194 264959 674250 264968
rect 674378 264616 674434 264625
rect 674378 264551 674434 264560
rect 674102 258904 674158 258913
rect 674102 258839 674158 258848
rect 674116 241505 674144 258839
rect 674102 241496 674158 241505
rect 674102 241431 674158 241440
rect 674088 235680 674140 235686
rect 674140 235628 674144 235668
rect 674088 235622 674144 235628
rect 674116 235142 674144 235622
rect 674104 235136 674156 235142
rect 674104 235078 674156 235084
rect 674196 234864 674248 234870
rect 674196 234806 674248 234812
rect 673932 234586 674144 234614
rect 673828 234252 673880 234258
rect 673828 234194 673880 234200
rect 673642 231840 673698 231849
rect 673642 231775 673698 231784
rect 673460 231328 673512 231334
rect 673460 231270 673512 231276
rect 673840 230314 673868 234194
rect 673948 233232 674000 233238
rect 674000 233180 674052 233186
rect 673948 233174 674052 233180
rect 673960 233158 674052 233174
rect 673828 230308 673880 230314
rect 673828 230250 673880 230256
rect 673458 230072 673514 230081
rect 673276 230036 673328 230042
rect 673458 230007 673514 230016
rect 673826 230072 673882 230081
rect 673826 230007 673882 230016
rect 673276 229978 673328 229984
rect 673288 229537 673316 229978
rect 673274 229528 673330 229537
rect 673472 229498 673500 230007
rect 673840 229838 673868 230007
rect 673828 229832 673880 229838
rect 673828 229774 673880 229780
rect 674024 229650 674052 233158
rect 674116 231690 674144 234586
rect 674208 231854 674236 234806
rect 674392 234614 674420 264551
rect 674576 244274 674604 265367
rect 675022 264208 675078 264217
rect 675022 264143 675078 264152
rect 674838 262032 674894 262041
rect 674838 261967 674894 261976
rect 674852 261225 674880 261967
rect 674838 261216 674894 261225
rect 674838 261151 674894 261160
rect 675036 258074 675064 264143
rect 678242 263256 678298 263265
rect 678242 263191 678298 263200
rect 676402 262848 676458 262857
rect 676402 262783 676458 262792
rect 676218 262440 676274 262449
rect 676218 262375 676274 262384
rect 676232 261225 676260 262375
rect 676218 261216 676274 261225
rect 676218 261151 676274 261160
rect 676416 260234 676444 262783
rect 675852 260228 675904 260234
rect 675852 260170 675904 260176
rect 676404 260228 676456 260234
rect 676404 260170 676456 260176
rect 675666 259176 675722 259185
rect 675666 259111 675722 259120
rect 675680 258233 675708 259111
rect 675666 258224 675722 258233
rect 675666 258159 675722 258168
rect 675864 258074 675892 260170
rect 674944 258046 675064 258074
rect 675496 258046 675892 258074
rect 674944 251174 674972 258046
rect 675298 257544 675354 257553
rect 675298 257479 675354 257488
rect 675312 256737 675340 257479
rect 675298 256728 675354 256737
rect 675298 256663 675354 256672
rect 675496 253934 675524 258046
rect 675312 253906 675524 253934
rect 675312 251174 675340 253906
rect 678256 252278 678284 263191
rect 675852 252272 675904 252278
rect 675496 252220 675852 252226
rect 675496 252214 675904 252220
rect 678244 252272 678296 252278
rect 678244 252214 678296 252220
rect 675496 252198 675892 252214
rect 675496 251258 675524 252198
rect 675484 251252 675536 251258
rect 675484 251194 675536 251200
rect 674944 251146 675064 251174
rect 675036 249393 675064 251146
rect 675220 251146 675340 251174
rect 674838 249384 674894 249393
rect 674838 249319 674894 249328
rect 675022 249384 675078 249393
rect 675022 249319 675078 249328
rect 674852 245426 674880 249319
rect 675022 248432 675078 248441
rect 675022 248367 675078 248376
rect 675036 245585 675064 248367
rect 675220 247398 675248 251146
rect 675484 250980 675536 250986
rect 675484 250922 675536 250928
rect 675496 250512 675524 250922
rect 675758 250336 675814 250345
rect 675758 250271 675814 250280
rect 675772 249900 675800 250271
rect 675390 249384 675446 249393
rect 675390 249319 675446 249328
rect 675404 249220 675432 249319
rect 675220 247370 675418 247398
rect 675298 247072 675354 247081
rect 675298 247007 675354 247016
rect 675312 246854 675340 247007
rect 675312 246826 675418 246854
rect 675298 246664 675354 246673
rect 675298 246599 675354 246608
rect 675312 246213 675340 246599
rect 675312 246185 675418 246213
rect 675298 245848 675354 245857
rect 675298 245783 675354 245792
rect 675022 245576 675078 245585
rect 675312 245562 675340 245783
rect 675312 245534 675418 245562
rect 675022 245511 675078 245520
rect 674852 245398 675156 245426
rect 674746 245304 674802 245313
rect 674746 245239 674802 245248
rect 674930 245304 674986 245313
rect 674930 245239 674986 245248
rect 674760 245154 674788 245239
rect 674760 245126 674880 245154
rect 674576 244246 674788 244274
rect 674536 235000 674588 235006
rect 674534 234968 674536 234977
rect 674588 234968 674590 234977
rect 674534 234903 674590 234912
rect 674392 234586 674604 234614
rect 674576 233481 674604 234586
rect 674760 234433 674788 244246
rect 674852 236382 674880 245126
rect 674944 241890 674972 245239
rect 675128 243085 675156 245398
rect 675128 243057 675418 243085
rect 675114 242856 675170 242865
rect 675114 242791 675170 242800
rect 675128 242533 675156 242791
rect 675128 242505 675418 242533
rect 674944 241862 675418 241890
rect 675114 241496 675170 241505
rect 675114 241431 675170 241440
rect 675128 241245 675156 241431
rect 675128 241217 675418 241245
rect 675114 240272 675170 240281
rect 675114 240207 675170 240216
rect 675128 240054 675156 240207
rect 675128 240026 675418 240054
rect 675390 238640 675446 238649
rect 675390 238575 675446 238584
rect 675404 238204 675432 238575
rect 675390 237824 675446 237833
rect 675390 237759 675446 237768
rect 675404 237524 675432 237759
rect 674852 236354 675418 236382
rect 674746 234424 674802 234433
rect 674746 234359 674802 234368
rect 675850 234424 675906 234433
rect 675850 234359 675852 234368
rect 675904 234359 675906 234368
rect 681004 234388 681056 234394
rect 675852 234330 675904 234336
rect 681004 234330 681056 234336
rect 674748 233912 674800 233918
rect 675096 233912 675148 233918
rect 674800 233872 675096 233900
rect 674748 233854 674800 233860
rect 675096 233854 675148 233860
rect 675236 233912 675288 233918
rect 675288 233872 676076 233900
rect 675236 233854 675288 233860
rect 675852 233776 675904 233782
rect 674852 233724 675852 233730
rect 674852 233718 675904 233724
rect 674852 233714 675892 233718
rect 674840 233708 675892 233714
rect 674892 233702 675892 233708
rect 674840 233650 674892 233656
rect 675116 233640 675168 233646
rect 675852 233640 675904 233646
rect 675168 233600 675852 233628
rect 675116 233582 675168 233588
rect 675852 233582 675904 233588
rect 675852 233504 675904 233510
rect 674562 233472 674618 233481
rect 674562 233407 674618 233416
rect 675850 233472 675852 233481
rect 675904 233472 675906 233481
rect 675850 233407 675906 233416
rect 676048 233374 676076 233872
rect 677692 233640 677744 233646
rect 677692 233582 677744 233588
rect 676036 233368 676088 233374
rect 676036 233310 676088 233316
rect 675852 232552 675904 232558
rect 675496 232500 675852 232506
rect 675496 232494 675904 232500
rect 675496 232490 675892 232494
rect 675484 232484 675892 232490
rect 675536 232478 675892 232484
rect 675484 232426 675536 232432
rect 674208 231826 674328 231854
rect 674116 231674 674212 231690
rect 674116 231668 674224 231674
rect 674116 231662 674172 231668
rect 674172 231610 674224 231616
rect 674300 230466 674328 231826
rect 674470 231840 674526 231849
rect 674470 231775 674526 231784
rect 674484 231674 674512 231775
rect 675180 231736 675232 231742
rect 675180 231678 675232 231684
rect 674472 231668 674524 231674
rect 674472 231610 674524 231616
rect 675192 231577 675220 231678
rect 675178 231568 675234 231577
rect 675070 231532 675122 231538
rect 675178 231503 675234 231512
rect 675070 231474 675122 231480
rect 674956 231328 675008 231334
rect 675082 231305 675110 231474
rect 674956 231270 675008 231276
rect 675068 231296 675124 231305
rect 674968 231146 674996 231270
rect 675068 231231 675124 231240
rect 674968 231130 675892 231146
rect 674968 231124 675904 231130
rect 674968 231118 675852 231124
rect 675852 231066 675904 231072
rect 675022 231024 675078 231033
rect 674484 230982 675022 231010
rect 674484 230858 674512 230982
rect 675022 230959 675078 230968
rect 676034 231024 676090 231033
rect 676034 230959 676090 230968
rect 674732 230920 674784 230926
rect 674730 230888 674732 230897
rect 674784 230888 674786 230897
rect 674472 230852 674524 230858
rect 674730 230823 674786 230832
rect 674472 230794 674524 230800
rect 674610 230716 674662 230722
rect 674610 230658 674662 230664
rect 674396 230648 674448 230654
rect 674448 230596 674558 230602
rect 674396 230590 674558 230596
rect 674408 230574 674558 230590
rect 674116 230438 674328 230466
rect 674116 229922 674144 230438
rect 674394 230344 674450 230353
rect 674530 230330 674558 230574
rect 674622 230466 674650 230658
rect 674622 230438 674880 230466
rect 674654 230344 674710 230353
rect 674530 230302 674654 230330
rect 674394 230279 674396 230288
rect 674448 230279 674450 230288
rect 674654 230279 674710 230288
rect 674396 230250 674448 230256
rect 674116 229894 674236 229922
rect 674024 229622 674144 229650
rect 673948 229560 674000 229566
rect 673932 229508 673948 229514
rect 673932 229502 674000 229508
rect 673274 229463 673330 229472
rect 673460 229492 673512 229498
rect 673460 229434 673512 229440
rect 673932 229486 673988 229502
rect 673460 229288 673512 229294
rect 673460 229230 673512 229236
rect 673472 229129 673500 229230
rect 673458 229120 673514 229129
rect 673458 229055 673514 229064
rect 673598 228948 673650 228954
rect 673650 228908 673776 228936
rect 673598 228890 673650 228896
rect 673368 228880 673420 228886
rect 673366 228848 673368 228857
rect 673420 228848 673422 228857
rect 673366 228783 673422 228792
rect 672736 228500 673132 228528
rect 673386 228576 673442 228585
rect 673386 228511 673388 228520
rect 672736 220130 672764 228500
rect 673440 228511 673442 228520
rect 673388 228482 673440 228488
rect 673058 228398 673592 228426
rect 673058 228138 673086 228398
rect 673276 228336 673328 228342
rect 673328 228296 673500 228324
rect 673276 228278 673328 228284
rect 673046 228132 673098 228138
rect 673046 228074 673098 228080
rect 672954 227724 673006 227730
rect 672954 227666 673006 227672
rect 672966 227474 672994 227666
rect 672966 227446 673224 227474
rect 672998 227080 673054 227089
rect 672998 227015 673054 227024
rect 673012 222578 673040 227015
rect 673196 226817 673224 227446
rect 673162 226808 673224 226817
rect 673218 226766 673224 226808
rect 673162 226743 673218 226752
rect 673472 225434 673500 228296
rect 673196 225406 673500 225434
rect 673196 224856 673224 225406
rect 673196 224828 673408 224856
rect 673182 223952 673238 223961
rect 673182 223887 673238 223896
rect 673012 222550 673132 222578
rect 672736 220102 672856 220130
rect 672828 215294 672856 220102
rect 673104 219314 673132 222550
rect 673012 219286 673132 219314
rect 673012 216209 673040 219286
rect 673196 219201 673224 223887
rect 673380 221513 673408 224828
rect 673366 221504 673422 221513
rect 673366 221439 673422 221448
rect 673564 221241 673592 228398
rect 673748 227089 673776 228908
rect 673734 227080 673790 227089
rect 673932 227066 673960 229486
rect 673932 227038 674052 227066
rect 673734 227015 673790 227024
rect 673734 226264 673790 226273
rect 673734 226199 673790 226208
rect 673748 225729 673776 226199
rect 673734 225720 673790 225729
rect 673734 225655 673790 225664
rect 673734 225448 673790 225457
rect 673734 225383 673790 225392
rect 673748 222057 673776 225383
rect 674024 224954 674052 227038
rect 673932 224926 674052 224954
rect 673932 222873 673960 224926
rect 673918 222864 673974 222873
rect 673918 222799 673974 222808
rect 673734 222048 673790 222057
rect 673734 221983 673790 221992
rect 673550 221232 673606 221241
rect 673550 221167 673606 221176
rect 673458 220416 673514 220425
rect 673458 220351 673514 220360
rect 673472 219881 673500 220351
rect 673458 219872 673514 219881
rect 673458 219807 673514 219816
rect 673182 219192 673238 219201
rect 673182 219127 673238 219136
rect 672998 216200 673054 216209
rect 672998 216135 673054 216144
rect 673366 215792 673422 215801
rect 673366 215727 673422 215736
rect 672644 215266 672764 215294
rect 672828 215266 672948 215294
rect 672538 188456 672594 188465
rect 672538 188391 672594 188400
rect 672184 188278 672488 188306
rect 672078 183560 672134 183569
rect 672078 183495 672134 183504
rect 671894 169960 671950 169969
rect 671894 169895 671950 169904
rect 671710 166968 671766 166977
rect 671710 166903 671766 166912
rect 671526 158400 671582 158409
rect 671526 158335 671582 158344
rect 670804 151786 671384 151814
rect 670804 150278 670832 151786
rect 670792 150272 670844 150278
rect 670792 150214 670844 150220
rect 670606 149016 670662 149025
rect 670606 148951 670662 148960
rect 671342 131744 671398 131753
rect 671342 131679 671398 131688
rect 670148 118108 670200 118114
rect 670148 118050 670200 118056
rect 671356 113174 671384 131679
rect 671526 130928 671582 130937
rect 671526 130863 671582 130872
rect 670804 113146 671384 113174
rect 667940 111444 667992 111450
rect 667940 111386 667992 111392
rect 669964 111444 670016 111450
rect 669964 111386 670016 111392
rect 590292 111104 590344 111110
rect 667952 111081 667980 111386
rect 590292 111046 590344 111052
rect 667938 111072 667994 111081
rect 667938 111007 667994 111016
rect 668582 111072 668638 111081
rect 668582 111007 668638 111016
rect 590106 110120 590162 110129
rect 590106 110055 590162 110064
rect 589372 109744 589424 109750
rect 589372 109686 589424 109692
rect 589462 108488 589518 108497
rect 589462 108423 589518 108432
rect 589476 107710 589504 108423
rect 589464 107704 589516 107710
rect 589464 107646 589516 107652
rect 589462 106856 589518 106865
rect 589462 106791 589518 106800
rect 589476 106350 589504 106791
rect 589464 106344 589516 106350
rect 589464 106286 589516 106292
rect 589830 105224 589886 105233
rect 589830 105159 589886 105168
rect 589844 104922 589872 105159
rect 589832 104916 589884 104922
rect 589832 104858 589884 104864
rect 589922 101960 589978 101969
rect 589922 101895 589978 101904
rect 588728 95192 588780 95198
rect 588728 95134 588780 95140
rect 588544 88324 588596 88330
rect 588544 88266 588596 88272
rect 589936 83502 589964 101895
rect 590120 98666 590148 110055
rect 667938 109304 667994 109313
rect 667938 109239 667994 109248
rect 590290 103592 590346 103601
rect 590290 103527 590346 103536
rect 590304 101454 590332 103527
rect 666650 102844 666706 102853
rect 666650 102779 666706 102788
rect 666664 102377 666692 102779
rect 666650 102368 666706 102377
rect 666650 102303 666706 102312
rect 590292 101448 590344 101454
rect 590292 101390 590344 101396
rect 624792 100156 624844 100162
rect 624792 100098 624844 100104
rect 595272 100014 595608 100042
rect 596192 100014 596344 100042
rect 596744 100014 597080 100042
rect 597572 100014 597816 100042
rect 598216 100014 598552 100042
rect 598952 100014 599288 100042
rect 599504 100014 600024 100042
rect 600424 100014 600760 100042
rect 600884 100014 601496 100042
rect 601896 100014 602232 100042
rect 602356 100014 602968 100042
rect 603092 100014 603704 100042
rect 590108 98660 590160 98666
rect 590108 98602 590160 98608
rect 595272 98122 595300 100014
rect 595260 98116 595312 98122
rect 595260 98058 595312 98064
rect 592684 97980 592736 97986
rect 592684 97922 592736 97928
rect 590108 97708 590160 97714
rect 590108 97650 590160 97656
rect 590120 90370 590148 97650
rect 590108 90364 590160 90370
rect 590108 90306 590160 90312
rect 589924 83496 589976 83502
rect 589924 83438 589976 83444
rect 587164 82136 587216 82142
rect 587164 82078 587216 82084
rect 588544 79348 588596 79354
rect 588544 79290 588596 79296
rect 584588 77240 584640 77246
rect 584588 77182 584640 77188
rect 584404 73160 584456 73166
rect 584404 73102 584456 73108
rect 583024 52148 583076 52154
rect 583024 52090 583076 52096
rect 578884 51468 578936 51474
rect 578884 51410 578936 51416
rect 588556 50930 588584 79290
rect 592696 51610 592724 97922
rect 592868 97844 592920 97850
rect 592868 97786 592920 97792
rect 592880 79354 592908 97786
rect 595272 93854 595300 98058
rect 596192 97578 596220 100014
rect 596180 97572 596232 97578
rect 596180 97514 596232 97520
rect 596744 97442 596772 100014
rect 597572 97986 597600 100014
rect 597560 97980 597612 97986
rect 597560 97922 597612 97928
rect 598216 97850 598244 100014
rect 598204 97844 598256 97850
rect 598204 97786 598256 97792
rect 596732 97436 596784 97442
rect 596732 97378 596784 97384
rect 598952 94586 598980 100014
rect 596824 94580 596876 94586
rect 596824 94522 596876 94528
rect 598940 94580 598992 94586
rect 598940 94522 598992 94528
rect 595272 93826 595484 93854
rect 595456 80714 595484 93826
rect 595444 80708 595496 80714
rect 595444 80650 595496 80656
rect 592868 79348 592920 79354
rect 592868 79290 592920 79296
rect 592684 51604 592736 51610
rect 592684 51546 592736 51552
rect 596836 51066 596864 94522
rect 599504 84194 599532 100014
rect 600424 97714 600452 100014
rect 600412 97708 600464 97714
rect 600412 97650 600464 97656
rect 600884 84194 600912 100014
rect 601896 97306 601924 100014
rect 601884 97300 601936 97306
rect 601884 97242 601936 97248
rect 602356 84194 602384 100014
rect 599136 84166 599532 84194
rect 600332 84166 600912 84194
rect 601712 84166 602384 84194
rect 596824 51060 596876 51066
rect 596824 51002 596876 51008
rect 588544 50924 588596 50930
rect 588544 50866 588596 50872
rect 577504 49428 577556 49434
rect 577504 49370 577556 49376
rect 599136 49298 599164 84166
rect 600332 51814 600360 84166
rect 600320 51808 600372 51814
rect 600320 51750 600372 51756
rect 599124 49292 599176 49298
rect 599124 49234 599176 49240
rect 553674 49192 553730 49201
rect 601712 49162 601740 84166
rect 603092 51921 603120 100014
rect 604426 99770 604454 100028
rect 605176 100014 605512 100042
rect 605912 100014 606248 100042
rect 606648 100014 606984 100042
rect 607384 100014 607720 100042
rect 608120 100014 608548 100042
rect 608856 100014 609192 100042
rect 609592 100014 609928 100042
rect 610328 100014 610664 100042
rect 604426 99742 604500 99770
rect 603078 51912 603134 51921
rect 603078 51847 603134 51856
rect 604472 51649 604500 99742
rect 605484 97442 605512 100014
rect 605472 97436 605524 97442
rect 605472 97378 605524 97384
rect 606220 96762 606248 100014
rect 606208 96756 606260 96762
rect 606208 96698 606260 96704
rect 606956 91798 606984 100014
rect 607128 96756 607180 96762
rect 607128 96698 607180 96704
rect 606944 91792 606996 91798
rect 606944 91734 606996 91740
rect 607140 75342 607168 96698
rect 607692 94518 607720 100014
rect 607680 94512 607732 94518
rect 607680 94454 607732 94460
rect 608520 84182 608548 100014
rect 609164 95946 609192 100014
rect 609152 95940 609204 95946
rect 609152 95882 609204 95888
rect 609900 85542 609928 100014
rect 610636 96762 610664 100014
rect 611050 99770 611078 100028
rect 611800 100014 612136 100042
rect 612536 100014 612688 100042
rect 613272 100014 613608 100042
rect 611004 99742 611078 99770
rect 610624 96756 610676 96762
rect 610624 96698 610676 96704
rect 611004 91050 611032 99742
rect 612108 96966 612136 100014
rect 612660 97306 612688 100014
rect 613384 97436 613436 97442
rect 613384 97378 613436 97384
rect 612648 97300 612700 97306
rect 612648 97242 612700 97248
rect 612096 96960 612148 96966
rect 612096 96902 612148 96908
rect 612648 96960 612700 96966
rect 612648 96902 612700 96908
rect 611176 96756 611228 96762
rect 611176 96698 611228 96704
rect 611188 93158 611216 96698
rect 612002 95840 612058 95849
rect 612002 95775 612058 95784
rect 611176 93152 611228 93158
rect 611176 93094 611228 93100
rect 610992 91044 611044 91050
rect 610992 90986 611044 90992
rect 609888 85536 609940 85542
rect 609888 85478 609940 85484
rect 608508 84176 608560 84182
rect 608508 84118 608560 84124
rect 607128 75336 607180 75342
rect 607128 75278 607180 75284
rect 612016 62082 612044 95775
rect 612660 79354 612688 96902
rect 612648 79348 612700 79354
rect 612648 79290 612700 79296
rect 613396 75206 613424 97378
rect 613580 96898 613608 100014
rect 613994 99770 614022 100028
rect 614744 100014 615080 100042
rect 615480 100014 615816 100042
rect 616216 100014 616552 100042
rect 616952 100014 617288 100042
rect 617688 100014 618024 100042
rect 618424 100014 618760 100042
rect 619160 100014 619588 100042
rect 619896 100014 620232 100042
rect 620632 100014 620968 100042
rect 621368 100014 621704 100042
rect 622104 100014 622348 100042
rect 622840 100014 623176 100042
rect 623576 100014 623728 100042
rect 624312 100014 624648 100042
rect 614856 99952 614908 99958
rect 614856 99894 614908 99900
rect 613994 99742 614068 99770
rect 613568 96892 613620 96898
rect 613568 96834 613620 96840
rect 614040 79490 614068 99742
rect 614028 79484 614080 79490
rect 614028 79426 614080 79432
rect 613384 75200 613436 75206
rect 613384 75142 613436 75148
rect 612004 62076 612056 62082
rect 612004 62018 612056 62024
rect 614868 57934 614896 99894
rect 615052 97034 615080 100014
rect 615040 97028 615092 97034
rect 615040 96970 615092 96976
rect 615040 96892 615092 96898
rect 615040 96834 615092 96840
rect 615052 77994 615080 96834
rect 615788 96830 615816 100014
rect 616144 97028 616196 97034
rect 616144 96970 616196 96976
rect 615776 96824 615828 96830
rect 615776 96766 615828 96772
rect 615040 77988 615092 77994
rect 615040 77930 615092 77936
rect 616156 76702 616184 96970
rect 616524 95062 616552 100014
rect 617260 96966 617288 100014
rect 617248 96960 617300 96966
rect 617248 96902 617300 96908
rect 616512 95056 616564 95062
rect 616512 94998 616564 95004
rect 617996 92478 618024 100014
rect 618732 97986 618760 100014
rect 618720 97980 618772 97986
rect 618720 97922 618772 97928
rect 618168 96960 618220 96966
rect 618168 96902 618220 96908
rect 617984 92472 618036 92478
rect 617984 92414 618036 92420
rect 618180 91050 618208 96902
rect 618904 96824 618956 96830
rect 618904 96766 618956 96772
rect 617524 91044 617576 91050
rect 617524 90986 617576 90992
rect 618168 91044 618220 91050
rect 618168 90986 618220 90992
rect 617536 88330 617564 90986
rect 617524 88324 617576 88330
rect 617524 88266 617576 88272
rect 618916 80850 618944 96766
rect 619560 93838 619588 100014
rect 620204 97442 620232 100014
rect 620192 97436 620244 97442
rect 620192 97378 620244 97384
rect 620284 97300 620336 97306
rect 620284 97242 620336 97248
rect 619548 93832 619600 93838
rect 619548 93774 619600 93780
rect 618904 80844 618956 80850
rect 618904 80786 618956 80792
rect 617522 77344 617578 77353
rect 617522 77279 617578 77288
rect 616144 76696 616196 76702
rect 616144 76638 616196 76644
rect 614856 57928 614908 57934
rect 614856 57870 614908 57876
rect 617536 53106 617564 77279
rect 618904 75676 618956 75682
rect 618904 75618 618956 75624
rect 617524 53100 617576 53106
rect 617524 53042 617576 53048
rect 604458 51640 604514 51649
rect 604458 51575 604514 51584
rect 553674 49127 553730 49136
rect 601700 49156 601752 49162
rect 601700 49098 601752 49104
rect 618916 49026 618944 75618
rect 620296 75478 620324 97242
rect 620940 95198 620968 100014
rect 621676 97306 621704 100014
rect 622320 99346 622348 100014
rect 622308 99340 622360 99346
rect 622308 99282 622360 99288
rect 623148 97578 623176 100014
rect 623700 99210 623728 100014
rect 623688 99204 623740 99210
rect 623688 99146 623740 99152
rect 623136 97572 623188 97578
rect 623136 97514 623188 97520
rect 621664 97300 621716 97306
rect 621664 97242 621716 97248
rect 624620 96898 624648 100014
rect 624608 96892 624660 96898
rect 624608 96834 624660 96840
rect 621664 95940 621716 95946
rect 621664 95882 621716 95888
rect 620928 95192 620980 95198
rect 620928 95134 620980 95140
rect 620928 94512 620980 94518
rect 620928 94454 620980 94460
rect 620940 89690 620968 94454
rect 620928 89684 620980 89690
rect 620928 89626 620980 89632
rect 621676 85406 621704 95882
rect 623228 95056 623280 95062
rect 623228 94998 623280 95004
rect 622400 93152 622452 93158
rect 622400 93094 622452 93100
rect 622412 86358 622440 93094
rect 623240 89554 623268 94998
rect 623228 89548 623280 89554
rect 623228 89490 623280 89496
rect 622400 86352 622452 86358
rect 622400 86294 622452 86300
rect 621664 85400 621716 85406
rect 621664 85342 621716 85348
rect 624804 84194 624832 100098
rect 625034 99770 625062 100028
rect 625784 100014 626120 100042
rect 626520 100014 626856 100042
rect 627256 100014 627592 100042
rect 627992 100014 628328 100042
rect 628728 100014 629064 100042
rect 629464 100014 629800 100042
rect 630200 100014 630536 100042
rect 630936 100014 631272 100042
rect 631672 100014 631916 100042
rect 632408 100014 632744 100042
rect 633144 100014 633388 100042
rect 633880 100014 634216 100042
rect 634616 100014 634768 100042
rect 635352 100014 635596 100042
rect 625034 99742 625108 99770
rect 625080 99074 625108 99742
rect 625068 99068 625120 99074
rect 625068 99010 625120 99016
rect 625804 97980 625856 97986
rect 625804 97922 625856 97928
rect 625816 92041 625844 97922
rect 626092 97714 626120 100014
rect 626080 97708 626132 97714
rect 626080 97650 626132 97656
rect 625988 97436 626040 97442
rect 625988 97378 626040 97384
rect 626000 93673 626028 97378
rect 626828 97034 626856 100014
rect 627564 98938 627592 100014
rect 627552 98932 627604 98938
rect 627552 98874 627604 98880
rect 628300 97850 628328 100014
rect 629036 98802 629064 100014
rect 629024 98796 629076 98802
rect 629024 98738 629076 98744
rect 629772 97986 629800 100014
rect 630508 98530 630536 100014
rect 630772 99340 630824 99346
rect 630772 99282 630824 99288
rect 630496 98524 630548 98530
rect 630496 98466 630548 98472
rect 629760 97980 629812 97986
rect 629760 97922 629812 97928
rect 628288 97844 628340 97850
rect 628288 97786 628340 97792
rect 629300 97300 629352 97306
rect 629300 97242 629352 97248
rect 626816 97028 626868 97034
rect 626816 96970 626868 96976
rect 629312 95826 629340 97242
rect 630784 95826 630812 99282
rect 629280 95798 629340 95826
rect 630752 95798 630812 95826
rect 631244 95470 631272 100014
rect 631416 98252 631468 98258
rect 631416 98194 631468 98200
rect 631428 97850 631456 98194
rect 631416 97844 631468 97850
rect 631416 97786 631468 97792
rect 631888 97306 631916 100014
rect 632060 97572 632112 97578
rect 632060 97514 632112 97520
rect 631876 97300 631928 97306
rect 631876 97242 631928 97248
rect 632072 95826 632100 97514
rect 632716 97442 632744 100014
rect 633360 97850 633388 100014
rect 633532 99204 633584 99210
rect 633532 99146 633584 99152
rect 633348 97844 633400 97850
rect 633348 97786 633400 97792
rect 632704 97436 632756 97442
rect 632704 97378 632756 97384
rect 633544 95826 633572 99146
rect 634188 97170 634216 100014
rect 634740 97578 634768 100014
rect 634728 97572 634780 97578
rect 634728 97514 634780 97520
rect 634176 97164 634228 97170
rect 634176 97106 634228 97112
rect 635004 96892 635056 96898
rect 635004 96834 635056 96840
rect 635016 95826 635044 96834
rect 635568 96393 635596 100014
rect 635752 100014 636088 100042
rect 636824 100014 637068 100042
rect 635554 96384 635610 96393
rect 635554 96319 635610 96328
rect 635752 96121 635780 100014
rect 636292 99068 636344 99074
rect 636292 99010 636344 99016
rect 635738 96112 635794 96121
rect 635738 96047 635794 96056
rect 636304 95826 636332 99010
rect 637040 96937 637068 100014
rect 637546 99770 637574 100028
rect 638296 100014 638632 100042
rect 637546 99742 637620 99770
rect 637026 96928 637082 96937
rect 637026 96863 637082 96872
rect 637592 96218 637620 99742
rect 637764 97708 637816 97714
rect 637764 97650 637816 97656
rect 637580 96212 637632 96218
rect 637580 96154 637632 96160
rect 637776 95826 637804 97650
rect 638604 96762 638632 100014
rect 639018 99770 639046 100028
rect 639768 100014 640104 100042
rect 639018 99742 639092 99770
rect 638592 96756 638644 96762
rect 638592 96698 638644 96704
rect 639064 96626 639092 99742
rect 639236 97028 639288 97034
rect 639236 96970 639288 96976
rect 639052 96620 639104 96626
rect 639052 96562 639104 96568
rect 639248 95826 639276 96970
rect 640076 96490 640104 100014
rect 640490 99770 640518 100028
rect 641240 100014 641576 100042
rect 640490 99742 640564 99770
rect 640064 96484 640116 96490
rect 640064 96426 640116 96432
rect 640536 96354 640564 99742
rect 640708 98932 640760 98938
rect 640708 98874 640760 98880
rect 640524 96348 640576 96354
rect 640524 96290 640576 96296
rect 640720 95826 640748 98874
rect 641548 96082 641576 100014
rect 641962 99770 641990 100028
rect 642712 100014 643048 100042
rect 641962 99742 642036 99770
rect 642008 96121 642036 99742
rect 642180 98252 642232 98258
rect 642180 98194 642232 98200
rect 641994 96112 642050 96121
rect 641536 96076 641588 96082
rect 641994 96047 642050 96056
rect 641536 96018 641588 96024
rect 642192 95826 642220 98194
rect 643020 97714 643048 100014
rect 643434 99770 643462 100028
rect 644184 100014 644336 100042
rect 643434 99742 643508 99770
rect 643008 97708 643060 97714
rect 643008 97650 643060 97656
rect 632072 95798 632224 95826
rect 633544 95798 633696 95826
rect 635016 95798 635168 95826
rect 636304 95798 636640 95826
rect 637776 95798 638112 95826
rect 639248 95798 639584 95826
rect 640720 95798 641056 95826
rect 642192 95798 642528 95826
rect 643480 95470 643508 99742
rect 643652 98796 643704 98802
rect 643652 98738 643704 98744
rect 643664 95826 643692 98738
rect 644308 97034 644336 100014
rect 644906 99770 644934 100028
rect 645656 100014 645808 100042
rect 644906 99742 644980 99770
rect 644296 97028 644348 97034
rect 644296 96970 644348 96976
rect 644952 95946 644980 99742
rect 645308 98048 645360 98054
rect 645308 97990 645360 97996
rect 645124 96484 645176 96490
rect 645124 96426 645176 96432
rect 644940 95940 644992 95946
rect 644940 95882 644992 95888
rect 643664 95798 644000 95826
rect 645136 95810 645164 96426
rect 645320 95826 645348 97990
rect 645780 96490 645808 100014
rect 646378 99770 646406 100028
rect 647114 99770 647142 100028
rect 647864 100014 648292 100042
rect 648600 100014 648936 100042
rect 649336 100014 649764 100042
rect 650072 100014 650408 100042
rect 650808 100014 651328 100042
rect 651544 100014 651880 100042
rect 652280 100014 652616 100042
rect 653016 100014 653352 100042
rect 653752 100014 653996 100042
rect 654488 100014 654824 100042
rect 646378 99742 646452 99770
rect 647114 99742 647188 99770
rect 645768 96484 645820 96490
rect 645768 96426 645820 96432
rect 645124 95804 645176 95810
rect 645320 95798 645472 95826
rect 645124 95746 645176 95752
rect 646424 95674 646452 99742
rect 647160 98666 647188 99742
rect 647148 98660 647200 98666
rect 647148 98602 647200 98608
rect 646596 98524 646648 98530
rect 646596 98466 646648 98472
rect 646608 95826 646636 98466
rect 647608 97164 647660 97170
rect 647608 97106 647660 97112
rect 647240 96756 647292 96762
rect 647240 96698 647292 96704
rect 647252 96234 647280 96698
rect 647422 96384 647478 96393
rect 647422 96319 647478 96328
rect 647252 96206 647372 96234
rect 646608 95798 646944 95826
rect 646412 95668 646464 95674
rect 646412 95610 646464 95616
rect 631232 95464 631284 95470
rect 631232 95406 631284 95412
rect 643468 95464 643520 95470
rect 643468 95406 643520 95412
rect 647148 95260 647200 95266
rect 647148 95202 647200 95208
rect 626448 95192 626500 95198
rect 626448 95134 626500 95140
rect 626460 94489 626488 95134
rect 647160 95033 647188 95202
rect 647146 95024 647202 95033
rect 647146 94959 647202 94968
rect 647344 94874 647372 96206
rect 647252 94846 647372 94874
rect 626446 94480 626502 94489
rect 626446 94415 626502 94424
rect 626448 93832 626500 93838
rect 626448 93774 626500 93780
rect 625986 93664 626042 93673
rect 625986 93599 626042 93608
rect 626460 92857 626488 93774
rect 626446 92848 626502 92857
rect 626446 92783 626502 92792
rect 626448 92472 626500 92478
rect 626448 92414 626500 92420
rect 625802 92032 625858 92041
rect 625802 91967 625858 91976
rect 626264 91792 626316 91798
rect 626264 91734 626316 91740
rect 625436 89684 625488 89690
rect 625436 89626 625488 89632
rect 625448 88777 625476 89626
rect 625434 88768 625490 88777
rect 625434 88703 625490 88712
rect 626276 87961 626304 91734
rect 626460 91225 626488 92414
rect 647252 91730 647280 94846
rect 647240 91724 647292 91730
rect 647240 91666 647292 91672
rect 626446 91216 626502 91225
rect 626446 91151 626502 91160
rect 626448 91044 626500 91050
rect 626448 90986 626500 90992
rect 626460 90409 626488 90986
rect 626446 90400 626502 90409
rect 626446 90335 626502 90344
rect 626446 89584 626502 89593
rect 626446 89519 626448 89528
rect 626500 89519 626502 89528
rect 626448 89490 626500 89496
rect 626448 88324 626500 88330
rect 626448 88266 626500 88272
rect 626262 87952 626318 87961
rect 626262 87887 626318 87896
rect 626460 87145 626488 88266
rect 626446 87136 626502 87145
rect 626446 87071 626502 87080
rect 626448 86352 626500 86358
rect 626446 86320 626448 86329
rect 626500 86320 626502 86329
rect 626446 86255 626502 86264
rect 626448 85536 626500 85542
rect 626446 85504 626448 85513
rect 626500 85504 626502 85513
rect 626446 85439 626502 85448
rect 625252 85400 625304 85406
rect 625252 85342 625304 85348
rect 625264 84697 625292 85342
rect 625250 84688 625306 84697
rect 625250 84623 625306 84632
rect 647436 84194 647464 96319
rect 647620 95198 647648 97106
rect 648068 95940 648120 95946
rect 648068 95882 648120 95888
rect 648080 95538 648108 95882
rect 648068 95532 648120 95538
rect 648068 95474 648120 95480
rect 647884 95464 647936 95470
rect 647884 95406 647936 95412
rect 647608 95192 647660 95198
rect 647608 95134 647660 95140
rect 647896 86766 647924 95406
rect 648264 94790 648292 100014
rect 648620 97300 648672 97306
rect 648620 97242 648672 97248
rect 648436 96348 648488 96354
rect 648436 96290 648488 96296
rect 648448 95946 648476 96290
rect 648436 95940 648488 95946
rect 648436 95882 648488 95888
rect 648252 94784 648304 94790
rect 648252 94726 648304 94732
rect 648632 92041 648660 97242
rect 648908 96354 648936 100014
rect 649080 97572 649132 97578
rect 649080 97514 649132 97520
rect 648896 96348 648948 96354
rect 648896 96290 648948 96296
rect 648618 92032 648674 92041
rect 648618 91967 648674 91976
rect 649092 89714 649120 97514
rect 649264 96620 649316 96626
rect 649264 96562 649316 96568
rect 649276 90710 649304 96562
rect 649264 90704 649316 90710
rect 649264 90646 649316 90652
rect 648908 89686 649120 89714
rect 647884 86760 647936 86766
rect 647884 86702 647936 86708
rect 624436 84166 624832 84194
rect 625804 84176 625856 84182
rect 622032 77308 622084 77314
rect 622032 77250 622084 77256
rect 621664 75948 621716 75954
rect 621664 75890 621716 75896
rect 620284 75472 620336 75478
rect 620284 75414 620336 75420
rect 621676 56574 621704 75890
rect 622044 75682 622072 77250
rect 622032 75676 622084 75682
rect 622032 75618 622084 75624
rect 623044 66292 623096 66298
rect 623044 66234 623096 66240
rect 621664 56568 621716 56574
rect 621664 56510 621716 56516
rect 618904 49020 618956 49026
rect 618904 48962 618956 48968
rect 552018 47832 552074 47841
rect 552018 47767 552074 47776
rect 547878 47560 547934 47569
rect 547878 47495 547934 47504
rect 521106 47016 521162 47025
rect 521106 46951 521162 46960
rect 465262 46608 465318 46617
rect 465262 46543 465318 46552
rect 623056 46510 623084 66234
rect 624436 60722 624464 84166
rect 625804 84118 625856 84124
rect 647252 84166 647464 84194
rect 625816 83881 625844 84118
rect 625802 83872 625858 83881
rect 625802 83807 625858 83816
rect 628746 83328 628802 83337
rect 628746 83263 628802 83272
rect 628760 80986 628788 83263
rect 629206 81696 629262 81705
rect 629206 81631 629262 81640
rect 628748 80980 628800 80986
rect 628748 80922 628800 80928
rect 629220 80034 629248 81631
rect 632808 80974 633144 81002
rect 642456 80980 642508 80986
rect 629208 80028 629260 80034
rect 629208 79970 629260 79976
rect 631048 78124 631100 78130
rect 631048 78066 631100 78072
rect 625802 77752 625858 77761
rect 625802 77687 625858 77696
rect 624424 60716 624476 60722
rect 624424 60658 624476 60664
rect 625816 52290 625844 77687
rect 631060 77450 631088 78066
rect 631048 77444 631100 77450
rect 631048 77386 631100 77392
rect 628472 77308 628524 77314
rect 628472 77250 628524 77256
rect 628484 75954 628512 77250
rect 628472 75948 628524 75954
rect 628472 75890 628524 75896
rect 628484 75290 628512 75890
rect 631060 75290 631088 77386
rect 632808 77314 632836 80974
rect 643080 80974 643140 81002
rect 642456 80922 642508 80928
rect 636752 80708 636804 80714
rect 636752 80650 636804 80656
rect 633440 80028 633492 80034
rect 633440 79970 633492 79976
rect 633452 78266 633480 79970
rect 633898 78568 633954 78577
rect 633898 78503 633954 78512
rect 633440 78260 633492 78266
rect 633440 78202 633492 78208
rect 633912 77353 633940 78503
rect 633898 77344 633954 77353
rect 632796 77308 632848 77314
rect 633898 77279 633954 77288
rect 632796 77250 632848 77256
rect 633912 75290 633940 77279
rect 636764 75290 636792 80650
rect 639602 77752 639658 77761
rect 639602 77687 639658 77696
rect 639616 75290 639644 77687
rect 642468 75290 642496 80922
rect 643112 78130 643140 80974
rect 646044 79484 646096 79490
rect 646044 79426 646096 79432
rect 645308 78260 645360 78266
rect 645308 78202 645360 78208
rect 643100 78124 643152 78130
rect 643100 78066 643152 78072
rect 645320 75290 645348 78202
rect 628176 75262 628512 75290
rect 631028 75262 631088 75290
rect 633880 75262 633940 75290
rect 636732 75262 636792 75290
rect 639584 75262 639644 75290
rect 642436 75262 642496 75290
rect 645288 75262 645348 75290
rect 646056 74534 646084 79426
rect 646320 79348 646372 79354
rect 646320 79290 646372 79296
rect 646056 74506 646176 74534
rect 646148 67153 646176 74506
rect 646134 67144 646190 67153
rect 646134 67079 646190 67088
rect 646332 59401 646360 79290
rect 646872 76696 646924 76702
rect 646872 76638 646924 76644
rect 646504 75336 646556 75342
rect 646504 75278 646556 75284
rect 646516 74225 646544 75278
rect 646502 74216 646558 74225
rect 646502 74151 646558 74160
rect 646884 68989 646912 76638
rect 646870 68980 646926 68989
rect 646870 68915 646926 68924
rect 646318 59392 646374 59401
rect 646318 59327 646374 59336
rect 647252 57361 647280 84166
rect 648908 82249 648936 89686
rect 649736 88806 649764 100014
rect 650184 97436 650236 97442
rect 650184 97378 650236 97384
rect 650000 95192 650052 95198
rect 650000 95134 650052 95140
rect 649724 88800 649776 88806
rect 649724 88742 649776 88748
rect 650012 84697 650040 95134
rect 650196 89593 650224 97378
rect 650380 97306 650408 100014
rect 650552 97844 650604 97850
rect 650552 97786 650604 97792
rect 650368 97300 650420 97306
rect 650368 97242 650420 97248
rect 650182 89584 650238 89593
rect 650182 89519 650238 89528
rect 650564 87145 650592 97786
rect 651300 93566 651328 100014
rect 651852 97578 651880 100014
rect 651840 97572 651892 97578
rect 651840 97514 651892 97520
rect 652588 96490 652616 100014
rect 653324 96626 653352 100014
rect 653968 97850 653996 100014
rect 653956 97844 654008 97850
rect 653956 97786 654008 97792
rect 654796 96898 654824 100014
rect 655210 99770 655238 100028
rect 655808 100014 655960 100042
rect 656696 100014 656848 100042
rect 657432 100014 657768 100042
rect 655210 99742 655284 99770
rect 655060 97844 655112 97850
rect 655060 97786 655112 97792
rect 654784 96892 654836 96898
rect 654784 96834 654836 96840
rect 653312 96620 653364 96626
rect 653312 96562 653364 96568
rect 652024 96484 652076 96490
rect 652024 96426 652076 96432
rect 652576 96484 652628 96490
rect 652576 96426 652628 96432
rect 651288 93560 651340 93566
rect 651288 93502 651340 93508
rect 650550 87136 650606 87145
rect 650550 87071 650606 87080
rect 652036 86222 652064 96426
rect 652208 95804 652260 95810
rect 652208 95746 652260 95752
rect 652220 86494 652248 95746
rect 653404 95668 653456 95674
rect 653404 95610 653456 95616
rect 653416 86902 653444 95610
rect 654784 94784 654836 94790
rect 654784 94726 654836 94732
rect 654796 93854 654824 94726
rect 655072 94217 655100 97786
rect 655256 96762 655284 99742
rect 655428 96892 655480 96898
rect 655428 96834 655480 96840
rect 655244 96756 655296 96762
rect 655244 96698 655296 96704
rect 655058 94208 655114 94217
rect 655058 94143 655114 94152
rect 655440 93854 655468 96834
rect 654796 93826 654916 93854
rect 654692 91724 654744 91730
rect 654692 91666 654744 91672
rect 654704 91497 654732 91666
rect 654690 91488 654746 91497
rect 654690 91423 654746 91432
rect 653404 86896 653456 86902
rect 653404 86838 653456 86844
rect 652208 86488 652260 86494
rect 652208 86430 652260 86436
rect 654888 86358 654916 93826
rect 655256 93826 655468 93854
rect 655256 88330 655284 93826
rect 655428 93560 655480 93566
rect 655428 93502 655480 93508
rect 655440 93401 655468 93502
rect 655426 93392 655482 93401
rect 655426 93327 655482 93336
rect 655428 90704 655480 90710
rect 655426 90672 655428 90681
rect 655480 90672 655482 90681
rect 655426 90607 655482 90616
rect 655808 89865 655836 100014
rect 656820 97170 656848 100014
rect 656808 97164 656860 97170
rect 656808 97106 656860 97112
rect 656164 95804 656216 95810
rect 656164 95746 656216 95752
rect 655794 89856 655850 89865
rect 655794 89791 655850 89800
rect 655244 88324 655296 88330
rect 655244 88266 655296 88272
rect 656176 86630 656204 95746
rect 657740 95132 657768 100014
rect 658154 99770 658182 100028
rect 658904 100014 659240 100042
rect 659640 100014 659976 100042
rect 660376 100014 660712 100042
rect 658154 99742 658228 99770
rect 658200 97442 658228 99742
rect 659212 97850 659240 100014
rect 659200 97844 659252 97850
rect 659200 97786 659252 97792
rect 659948 97714 659976 100014
rect 659752 97708 659804 97714
rect 659752 97650 659804 97656
rect 659936 97708 659988 97714
rect 659936 97650 659988 97656
rect 659568 97572 659620 97578
rect 659568 97514 659620 97520
rect 658188 97436 658240 97442
rect 658188 97378 658240 97384
rect 658280 97300 658332 97306
rect 658280 97242 658332 97248
rect 658292 95132 658320 97242
rect 658832 97028 658884 97034
rect 658832 96970 658884 96976
rect 658844 95132 658872 96970
rect 659580 95132 659608 97514
rect 659764 95146 659792 97650
rect 660684 96898 660712 100014
rect 661960 98660 662012 98666
rect 661960 98602 662012 98608
rect 661408 97164 661460 97170
rect 661408 97106 661460 97112
rect 660672 96892 660724 96898
rect 660672 96834 660724 96840
rect 660672 96212 660724 96218
rect 660672 96154 660724 96160
rect 659764 95118 660146 95146
rect 660684 95132 660712 96154
rect 661420 95132 661448 97106
rect 661972 95132 662000 98602
rect 663892 97844 663944 97850
rect 663892 97786 663944 97792
rect 663064 97436 663116 97442
rect 663064 97378 663116 97384
rect 662512 96756 662564 96762
rect 662512 96698 662564 96704
rect 662524 95132 662552 96698
rect 663076 95132 663104 97378
rect 663248 96892 663300 96898
rect 663248 96834 663300 96840
rect 658556 88800 658608 88806
rect 662328 88800 662380 88806
rect 658608 88748 658858 88754
rect 658556 88742 658858 88748
rect 658568 88726 658858 88742
rect 661986 88748 662328 88754
rect 661986 88742 662380 88748
rect 661986 88726 662368 88742
rect 658306 88330 658504 88346
rect 658306 88324 658516 88330
rect 658306 88318 658464 88324
rect 658464 88266 658516 88272
rect 657188 86902 657216 88196
rect 657176 86896 657228 86902
rect 657176 86838 657228 86844
rect 656164 86624 656216 86630
rect 656164 86566 656216 86572
rect 654876 86352 654928 86358
rect 654876 86294 654928 86300
rect 657740 86222 657768 88196
rect 659580 86970 659608 88196
rect 659568 86964 659620 86970
rect 659568 86906 659620 86912
rect 660132 86494 660160 88196
rect 660684 86630 660712 88196
rect 661420 86766 661448 88196
rect 661408 86760 661460 86766
rect 661408 86702 661460 86708
rect 660672 86624 660724 86630
rect 660672 86566 660724 86572
rect 660120 86488 660172 86494
rect 660120 86430 660172 86436
rect 662524 86358 662552 88196
rect 663260 86970 663288 96834
rect 663708 96076 663760 96082
rect 663708 96018 663760 96024
rect 663720 95962 663748 96018
rect 663720 95934 663840 95962
rect 663812 92970 663840 95934
rect 663720 92942 663840 92970
rect 663720 92857 663748 92942
rect 663706 92848 663762 92857
rect 663706 92783 663762 92792
rect 663904 88806 663932 97786
rect 665364 97708 665416 97714
rect 665364 97650 665416 97656
rect 665180 96620 665232 96626
rect 665180 96562 665232 96568
rect 664168 96484 664220 96490
rect 664168 96426 664220 96432
rect 664180 90681 664208 96426
rect 664352 96348 664404 96354
rect 664352 96290 664404 96296
rect 664166 90672 664222 90681
rect 664166 90607 664222 90616
rect 664364 89865 664392 96290
rect 664536 95940 664588 95946
rect 664536 95882 664588 95888
rect 664548 91769 664576 95882
rect 664534 91760 664590 91769
rect 664534 91695 664590 91704
rect 664350 89856 664406 89865
rect 664350 89791 664406 89800
rect 665192 89049 665220 96562
rect 665376 93401 665404 97650
rect 665362 93392 665418 93401
rect 665362 93327 665418 93336
rect 665178 89040 665234 89049
rect 665178 88975 665234 88984
rect 663892 88800 663944 88806
rect 663892 88742 663944 88748
rect 663248 86964 663300 86970
rect 663248 86906 663300 86912
rect 662512 86352 662564 86358
rect 662512 86294 662564 86300
rect 652024 86216 652076 86222
rect 652024 86158 652076 86164
rect 657728 86216 657780 86222
rect 657728 86158 657780 86164
rect 649998 84688 650054 84697
rect 649998 84623 650054 84632
rect 666664 84194 666692 102303
rect 667952 100162 667980 109239
rect 668400 106208 668452 106214
rect 668122 106176 668178 106185
rect 668122 106111 668178 106120
rect 668398 106176 668400 106185
rect 668452 106176 668454 106185
rect 668398 106111 668454 106120
rect 667940 100156 667992 100162
rect 667940 100098 667992 100104
rect 668136 100026 668164 106111
rect 668596 104417 668624 111007
rect 670804 106214 670832 113146
rect 671540 107817 671568 130863
rect 671724 115841 671752 166903
rect 671908 151881 671936 169895
rect 671894 151872 671950 151881
rect 671894 151807 671950 151816
rect 672092 140457 672120 183495
rect 672460 177993 672488 188278
rect 672446 177984 672502 177993
rect 672446 177919 672502 177928
rect 672538 175264 672594 175273
rect 672538 175199 672594 175208
rect 672078 140448 672134 140457
rect 672078 140383 672134 140392
rect 672552 130529 672580 175199
rect 672736 153105 672764 215266
rect 672920 209681 672948 215266
rect 673182 214160 673238 214169
rect 673182 214095 673238 214104
rect 672906 209672 672962 209681
rect 672906 209607 672962 209616
rect 672906 200832 672962 200841
rect 672906 200767 672962 200776
rect 672722 153096 672778 153105
rect 672722 153031 672778 153040
rect 672538 130520 672594 130529
rect 672538 130455 672594 130464
rect 672354 126032 672410 126041
rect 672354 125967 672410 125976
rect 671710 115832 671766 115841
rect 671710 115767 671766 115776
rect 672368 111489 672396 125967
rect 672920 124137 672948 200767
rect 673196 197713 673224 214095
rect 673380 201385 673408 215727
rect 673642 215384 673698 215393
rect 673642 215319 673698 215328
rect 673366 201376 673422 201385
rect 673366 201311 673422 201320
rect 673656 200841 673684 215319
rect 674116 213466 674144 229622
rect 673748 213438 674144 213466
rect 673748 213058 673776 213438
rect 674208 213194 674236 229894
rect 674852 229809 674880 230438
rect 675114 230072 675170 230081
rect 675170 230042 675892 230058
rect 675170 230036 675904 230042
rect 675170 230030 675852 230036
rect 675114 230007 675170 230016
rect 675852 229978 675904 229984
rect 674838 229800 674894 229809
rect 674838 229735 674894 229744
rect 676048 229634 676076 230959
rect 676862 230344 676918 230353
rect 676862 230279 676918 230288
rect 676496 230036 676548 230042
rect 676496 229978 676548 229984
rect 676036 229628 676088 229634
rect 676036 229570 676088 229576
rect 675114 229528 675170 229537
rect 675170 229498 675892 229514
rect 675170 229492 675904 229498
rect 675170 229486 675852 229492
rect 675114 229463 675170 229472
rect 675852 229434 675904 229440
rect 675114 228848 675170 228857
rect 675114 228783 675170 228792
rect 674746 226536 674802 226545
rect 674746 226471 674802 226480
rect 674378 225720 674434 225729
rect 674378 225655 674434 225664
rect 674392 220697 674420 225655
rect 674562 225176 674618 225185
rect 674562 225111 674618 225120
rect 674378 220688 674434 220697
rect 674378 220623 674434 220632
rect 674378 220416 674434 220425
rect 674576 220402 674604 225111
rect 674760 222194 674788 226471
rect 674954 225992 675010 226001
rect 674434 220374 674604 220402
rect 674668 222166 674788 222194
rect 674944 225936 674954 225978
rect 674944 225927 675010 225936
rect 674378 220351 674434 220360
rect 674668 218113 674696 222166
rect 674654 218104 674710 218113
rect 674654 218039 674710 218048
rect 674944 217682 674972 225927
rect 675128 223417 675156 228783
rect 676218 227080 676274 227089
rect 676218 227015 676274 227024
rect 675298 226808 675354 226817
rect 675298 226743 675354 226752
rect 675114 223408 675170 223417
rect 675114 223343 675170 223352
rect 675312 218906 675340 226743
rect 675574 224360 675630 224369
rect 675574 224295 675630 224304
rect 675588 218929 675616 224295
rect 675852 220108 675904 220114
rect 675852 220050 675904 220056
rect 674852 217654 674972 217682
rect 675128 218878 675340 218906
rect 675574 218920 675630 218929
rect 674852 217569 674880 217654
rect 674838 217560 674894 217569
rect 674838 217495 674894 217504
rect 674562 216608 674618 216617
rect 674562 216543 674618 216552
rect 674576 215294 674604 216543
rect 675128 216073 675156 218878
rect 675574 218855 675630 218864
rect 675864 216322 675892 220050
rect 676232 219586 676260 227015
rect 676508 220114 676536 229978
rect 676680 229492 676732 229498
rect 676680 229434 676732 229440
rect 676496 220108 676548 220114
rect 676496 220050 676548 220056
rect 676048 219558 676260 219586
rect 676048 218385 676076 219558
rect 676220 219428 676272 219434
rect 676220 219370 676272 219376
rect 676034 218376 676090 218385
rect 676034 218311 676090 218320
rect 676034 217832 676090 217841
rect 676034 217767 676090 217776
rect 675404 216294 675892 216322
rect 675114 216064 675170 216073
rect 675114 215999 675170 216008
rect 675404 215294 675432 216294
rect 675574 216200 675630 216209
rect 675574 216135 675630 216144
rect 674484 215266 674604 215294
rect 675036 215266 675432 215294
rect 674208 213166 674420 213194
rect 673748 213030 674052 213058
rect 673826 211168 673882 211177
rect 673826 211103 673882 211112
rect 673840 203969 673868 211103
rect 674024 210338 674052 213030
rect 674024 210310 674328 210338
rect 674010 208312 674066 208321
rect 674010 208247 674066 208256
rect 673826 203960 673882 203969
rect 673826 203895 673882 203904
rect 673642 200832 673698 200841
rect 673642 200767 673698 200776
rect 673182 197704 673238 197713
rect 673182 197639 673238 197648
rect 674024 195974 674052 208247
rect 674300 205634 674328 210310
rect 673932 195946 674052 195974
rect 674116 205606 674328 205634
rect 673366 174448 673422 174457
rect 673366 174383 673422 174392
rect 673182 169144 673238 169153
rect 673182 169079 673238 169088
rect 673196 152561 673224 169079
rect 673182 152552 673238 152561
rect 673182 152487 673238 152496
rect 673380 129713 673408 174383
rect 673932 172961 673960 195946
rect 673918 172952 673974 172961
rect 673918 172887 673974 172896
rect 674116 154601 674144 205606
rect 674392 195974 674420 213166
rect 674484 212534 674512 215266
rect 674838 214704 674894 214713
rect 674838 214639 674894 214648
rect 674654 213752 674710 213761
rect 674654 213687 674710 213696
rect 674668 212534 674696 213687
rect 674484 212506 674604 212534
rect 674668 212506 674788 212534
rect 674576 209681 674604 212506
rect 674562 209672 674618 209681
rect 674562 209607 674618 209616
rect 674760 202874 674788 212506
rect 674852 207210 674880 214639
rect 675036 207369 675064 215266
rect 675588 212534 675616 216135
rect 675852 215144 675904 215150
rect 675850 215112 675852 215121
rect 675904 215112 675906 215121
rect 675850 215047 675906 215056
rect 675758 214704 675814 214713
rect 676048 214690 676076 217767
rect 675814 214662 676076 214690
rect 675758 214639 675814 214648
rect 676034 214568 676090 214577
rect 676034 214503 676090 214512
rect 675852 214464 675904 214470
rect 675850 214432 675852 214441
rect 675904 214432 675906 214441
rect 675850 214367 675906 214376
rect 676048 213586 676076 214503
rect 676036 213580 676088 213586
rect 676036 213522 676088 213528
rect 675850 213480 675906 213489
rect 676232 213466 676260 219370
rect 676692 215294 676720 229434
rect 675906 213438 676260 213466
rect 676324 215266 676720 215294
rect 675850 213415 675906 213424
rect 675220 212506 675616 212534
rect 675022 207360 675078 207369
rect 675022 207295 675078 207304
rect 674852 207182 675064 207210
rect 675036 205034 675064 207182
rect 674668 202846 674788 202874
rect 674852 205006 675064 205034
rect 674852 202874 674880 205006
rect 675220 204762 675248 212506
rect 676324 211177 676352 215266
rect 676876 215150 676904 230279
rect 677416 229628 677468 229634
rect 677416 229570 677468 229576
rect 676864 215144 676916 215150
rect 676864 215086 676916 215092
rect 677428 214470 677456 229570
rect 677416 214464 677468 214470
rect 677416 214406 677468 214412
rect 677048 213580 677100 213586
rect 677048 213522 677100 213528
rect 677060 211449 677088 213522
rect 676770 211440 676826 211449
rect 676770 211375 676826 211384
rect 677046 211440 677102 211449
rect 677046 211375 677102 211384
rect 676310 211168 676366 211177
rect 676310 211103 676366 211112
rect 675482 209672 675538 209681
rect 675312 209630 675482 209658
rect 675312 205170 675340 209630
rect 675482 209607 675538 209616
rect 676784 208321 676812 211375
rect 677704 209409 677732 233582
rect 677876 233368 677928 233374
rect 677876 233310 677928 233316
rect 677690 209400 677746 209409
rect 677690 209335 677746 209344
rect 676770 208312 676826 208321
rect 676770 208247 676826 208256
rect 677888 206417 677916 233310
rect 678612 231124 678664 231130
rect 678612 231066 678664 231072
rect 678624 219434 678652 231066
rect 681016 220697 681044 234330
rect 683302 234152 683358 234161
rect 683302 234087 683358 234096
rect 683120 233436 683172 233442
rect 683120 233378 683172 233384
rect 683132 221513 683160 233378
rect 683316 223553 683344 234087
rect 683670 233880 683726 233889
rect 683670 233815 683726 233824
rect 683488 232552 683540 232558
rect 683488 232494 683540 232500
rect 683302 223544 683358 223553
rect 683302 223479 683358 223488
rect 683500 222737 683528 232494
rect 683684 223145 683712 233815
rect 684500 233300 684552 233306
rect 684500 233242 684552 233248
rect 683670 223136 683726 223145
rect 683670 223071 683726 223080
rect 683486 222728 683542 222737
rect 683486 222663 683542 222672
rect 683118 221504 683174 221513
rect 683118 221439 683174 221448
rect 681002 220688 681058 220697
rect 681002 220623 681058 220632
rect 684512 219881 684540 233242
rect 703694 224196 703722 224264
rect 704154 224196 704182 224264
rect 704614 224196 704642 224264
rect 705074 224196 705102 224264
rect 705534 224196 705562 224264
rect 705994 224196 706022 224264
rect 706454 224196 706482 224264
rect 706914 224196 706942 224264
rect 707374 224196 707402 224264
rect 707834 224196 707862 224264
rect 708294 224196 708322 224264
rect 708754 224196 708782 224264
rect 709214 224196 709242 224264
rect 684498 219872 684554 219881
rect 684498 219807 684554 219816
rect 678612 219428 678664 219434
rect 678612 219370 678664 219376
rect 679622 219056 679678 219065
rect 679622 218991 679678 219000
rect 679636 207097 679664 218991
rect 683302 213344 683358 213353
rect 683302 213279 683358 213288
rect 683118 212528 683174 212537
rect 683118 212463 683174 212472
rect 683132 211177 683160 212463
rect 683118 211168 683174 211177
rect 683118 211103 683174 211112
rect 683316 210361 683344 213279
rect 683302 210352 683358 210361
rect 683302 210287 683358 210296
rect 679622 207088 679678 207097
rect 679622 207023 679678 207032
rect 677874 206408 677930 206417
rect 677874 206343 677930 206352
rect 675758 205592 675814 205601
rect 675758 205527 675814 205536
rect 675772 205323 675800 205527
rect 675312 205142 675432 205170
rect 675220 204734 675340 204762
rect 675312 202874 675340 204734
rect 675404 204680 675432 205142
rect 675666 204232 675722 204241
rect 675666 204167 675722 204176
rect 675680 204035 675708 204167
rect 674852 202846 674972 202874
rect 674668 196081 674696 202846
rect 674944 202609 674972 202846
rect 675220 202846 675340 202874
rect 674930 202600 674986 202609
rect 674930 202535 674986 202544
rect 675220 202450 675248 202846
rect 675390 202600 675446 202609
rect 675390 202535 675446 202544
rect 675128 202422 675248 202450
rect 675128 201634 675156 202422
rect 675404 202195 675432 202535
rect 675312 201742 675432 201770
rect 675312 201634 675340 201742
rect 675128 201606 675340 201634
rect 675404 201620 675432 201742
rect 675114 201376 675170 201385
rect 675114 201311 675170 201320
rect 675128 201022 675156 201311
rect 675128 200994 675418 201022
rect 674838 200832 674894 200841
rect 674838 200767 674894 200776
rect 675758 200832 675814 200841
rect 675758 200767 675814 200776
rect 674852 199866 674880 200767
rect 675772 200328 675800 200767
rect 674852 199838 674972 199866
rect 674654 196072 674710 196081
rect 674654 196007 674710 196016
rect 674944 195974 674972 199838
rect 675390 198384 675446 198393
rect 675390 198319 675446 198328
rect 675404 197880 675432 198319
rect 675482 197704 675538 197713
rect 675482 197639 675538 197648
rect 675496 197336 675524 197639
rect 675758 197160 675814 197169
rect 675758 197095 675814 197104
rect 675772 196656 675800 197095
rect 675206 196072 675262 196081
rect 675262 196030 675418 196058
rect 675206 196007 675262 196016
rect 674300 195946 674420 195974
rect 674852 195946 674972 195974
rect 674300 179489 674328 195946
rect 674852 194834 674880 195946
rect 674852 194806 675418 194834
rect 675666 193216 675722 193225
rect 675666 193151 675722 193160
rect 675680 192984 675708 193151
rect 675114 192400 675170 192409
rect 675170 192358 675340 192386
rect 675114 192335 675170 192344
rect 675312 192250 675340 192358
rect 675404 192250 675432 192372
rect 675312 192222 675432 192250
rect 675758 191584 675814 191593
rect 675758 191519 675814 191528
rect 675772 191148 675800 191519
rect 675850 181384 675906 181393
rect 675850 181319 675906 181328
rect 674286 179480 674342 179489
rect 674286 179415 674342 179424
rect 675864 178129 675892 181319
rect 703694 179180 703722 179316
rect 704154 179180 704182 179316
rect 704614 179180 704642 179316
rect 705074 179180 705102 179316
rect 705534 179180 705562 179316
rect 705994 179180 706022 179316
rect 706454 179180 706482 179316
rect 706914 179180 706942 179316
rect 707374 179180 707402 179316
rect 707834 179180 707862 179316
rect 708294 179180 708322 179316
rect 708754 179180 708782 179316
rect 709214 179180 709242 179316
rect 676034 178800 676090 178809
rect 676034 178735 676090 178744
rect 675850 178120 675906 178129
rect 675850 178055 675906 178064
rect 676048 177721 676076 178735
rect 676034 177712 676090 177721
rect 676034 177647 676090 177656
rect 674286 176896 674342 176905
rect 674286 176831 674342 176840
rect 674102 154592 674158 154601
rect 674102 154527 674158 154536
rect 674300 132161 674328 176831
rect 674654 176080 674710 176089
rect 674654 176015 674710 176024
rect 674470 168736 674526 168745
rect 674470 168671 674526 168680
rect 674484 151065 674512 168671
rect 674470 151056 674526 151065
rect 674470 150991 674526 151000
rect 674286 132152 674342 132161
rect 674286 132087 674342 132096
rect 674668 131345 674696 176015
rect 676034 173224 676090 173233
rect 676090 173182 676260 173210
rect 676034 173159 676090 173168
rect 674838 172816 674894 172825
rect 674838 172751 674894 172760
rect 674852 157593 674880 172751
rect 675022 171184 675078 171193
rect 675022 171119 675078 171128
rect 675036 166994 675064 171119
rect 676232 169674 676260 173182
rect 681002 171592 681058 171601
rect 681002 171527 681058 171536
rect 676586 170776 676642 170785
rect 676586 170711 676642 170720
rect 675864 169646 676260 169674
rect 675864 166994 675892 169646
rect 676034 167920 676090 167929
rect 676034 167855 676090 167864
rect 674944 166966 675064 166994
rect 675496 166966 675892 166994
rect 674944 164234 674972 166966
rect 674944 164206 675064 164234
rect 674838 157584 674894 157593
rect 674838 157519 674894 157528
rect 675036 156657 675064 164206
rect 675206 161392 675262 161401
rect 675206 161327 675262 161336
rect 675220 159678 675248 161327
rect 675496 161106 675524 166966
rect 676048 165073 676076 167855
rect 676600 166433 676628 170711
rect 676586 166424 676642 166433
rect 676586 166359 676642 166368
rect 676034 165064 676090 165073
rect 676034 164999 676090 165008
rect 681016 162586 681044 171527
rect 675852 162580 675904 162586
rect 675852 162522 675904 162528
rect 681004 162580 681056 162586
rect 681004 162522 681056 162528
rect 675864 161401 675892 162522
rect 675850 161392 675906 161401
rect 675850 161327 675906 161336
rect 675312 161078 675524 161106
rect 675312 160290 675340 161078
rect 675404 160290 675432 160344
rect 675312 160262 675432 160290
rect 675220 159650 675418 159678
rect 675758 159352 675814 159361
rect 675758 159287 675814 159296
rect 675772 159052 675800 159287
rect 675482 157584 675538 157593
rect 675482 157519 675538 157528
rect 675496 157216 675524 157519
rect 675036 156629 675418 156657
rect 675758 156360 675814 156369
rect 675758 156295 675814 156304
rect 675772 155992 675800 156295
rect 675128 155366 675340 155394
rect 675128 154873 675156 155366
rect 675312 155258 675340 155366
rect 675404 155258 675432 155380
rect 675312 155230 675432 155258
rect 675114 154864 675170 154873
rect 675114 154799 675170 154808
rect 675312 152850 675418 152878
rect 675312 151609 675340 152850
rect 675482 152552 675538 152561
rect 675482 152487 675538 152496
rect 675496 152320 675524 152487
rect 675482 151872 675538 151881
rect 675482 151807 675538 151816
rect 675496 151675 675524 151807
rect 675298 151600 675354 151609
rect 675298 151535 675354 151544
rect 675114 151056 675170 151065
rect 675170 151014 675418 151042
rect 675114 150991 675170 151000
rect 675666 150376 675722 150385
rect 675666 150311 675722 150320
rect 675680 149835 675708 150311
rect 675298 149016 675354 149025
rect 675298 148951 675354 148960
rect 675312 146690 675340 148951
rect 675758 148472 675814 148481
rect 675758 148407 675814 148416
rect 675772 147968 675800 148407
rect 675666 147656 675722 147665
rect 675666 147591 675722 147600
rect 675680 147356 675708 147591
rect 675312 146662 675432 146690
rect 675404 146132 675432 146662
rect 683302 142760 683358 142769
rect 683302 142695 683358 142704
rect 683118 135960 683174 135969
rect 683118 135895 683174 135904
rect 683132 132705 683160 135895
rect 683316 133113 683344 142695
rect 703694 133892 703722 134028
rect 704154 133892 704182 134028
rect 704614 133892 704642 134028
rect 705074 133892 705102 134028
rect 705534 133892 705562 134028
rect 705994 133892 706022 134028
rect 706454 133892 706482 134028
rect 706914 133892 706942 134028
rect 707374 133892 707402 134028
rect 707834 133892 707862 134028
rect 708294 133892 708322 134028
rect 708754 133892 708782 134028
rect 709214 133892 709242 134028
rect 683302 133104 683358 133113
rect 683302 133039 683358 133048
rect 683118 132696 683174 132705
rect 683118 132631 683174 132640
rect 674654 131336 674710 131345
rect 674654 131271 674710 131280
rect 676218 130248 676274 130257
rect 676218 130183 676274 130192
rect 673366 129704 673422 129713
rect 673366 129639 673422 129648
rect 674102 129296 674158 129305
rect 674102 129231 674158 129240
rect 673182 124400 673238 124409
rect 673182 124335 673238 124344
rect 672906 124128 672962 124137
rect 672906 124063 672962 124072
rect 672906 123856 672962 123865
rect 672906 123791 672962 123800
rect 672722 123176 672778 123185
rect 672722 123111 672778 123120
rect 672538 122768 672594 122777
rect 672538 122703 672594 122712
rect 672552 112713 672580 122703
rect 672736 122233 672764 123111
rect 672722 122224 672778 122233
rect 672722 122159 672778 122168
rect 672920 118694 672948 123791
rect 672736 118666 672948 118694
rect 672736 117994 672764 118666
rect 672736 117966 672856 117994
rect 672538 112704 672594 112713
rect 672538 112639 672594 112648
rect 672354 111480 672410 111489
rect 672354 111415 672410 111424
rect 671526 107808 671582 107817
rect 671526 107743 671582 107752
rect 672828 106321 672856 117966
rect 673196 110401 673224 124335
rect 673366 123584 673422 123593
rect 673366 123519 673422 123528
rect 673182 110392 673238 110401
rect 673182 110327 673238 110336
rect 672814 106312 672870 106321
rect 672814 106247 672870 106256
rect 670792 106208 670844 106214
rect 670792 106150 670844 106156
rect 673380 105641 673408 123519
rect 674116 111081 674144 129231
rect 676232 128217 676260 130183
rect 674286 128208 674342 128217
rect 674286 128143 674342 128152
rect 676218 128208 676274 128217
rect 676218 128143 676274 128152
rect 676862 128208 676918 128217
rect 676862 128143 676918 128152
rect 674102 111072 674158 111081
rect 674102 111007 674158 111016
rect 673366 105632 673422 105641
rect 673366 105567 673422 105576
rect 668582 104408 668638 104417
rect 668582 104343 668638 104352
rect 668596 103514 668624 104343
rect 668320 103486 668624 103514
rect 668124 100020 668176 100026
rect 668124 99962 668176 99968
rect 668320 95849 668348 103486
rect 674300 102377 674328 128143
rect 674838 127664 674894 127673
rect 674838 127599 674894 127608
rect 674654 125624 674710 125633
rect 674654 125559 674710 125568
rect 674470 125216 674526 125225
rect 674470 125151 674526 125160
rect 674484 104666 674512 125151
rect 674668 110786 674696 125559
rect 674852 112010 674880 127599
rect 675022 126440 675078 126449
rect 675022 126375 675078 126384
rect 675036 114493 675064 126375
rect 676876 117337 676904 128143
rect 679622 127800 679678 127809
rect 679622 127735 679678 127744
rect 676862 117328 676918 117337
rect 675852 117292 675904 117298
rect 679636 117298 679664 127735
rect 676862 117263 676918 117272
rect 679624 117292 679676 117298
rect 675852 117234 675904 117240
rect 679624 117234 679676 117240
rect 675864 117178 675892 117234
rect 675312 117150 675892 117178
rect 675312 115138 675340 117150
rect 675312 115110 675418 115138
rect 675036 114465 675418 114493
rect 675312 113818 675418 113846
rect 675312 113121 675340 113818
rect 675298 113112 675354 113121
rect 675298 113047 675354 113056
rect 674852 111982 675418 112010
rect 675114 111480 675170 111489
rect 675170 111438 675418 111466
rect 675114 111415 675170 111424
rect 675312 110894 675432 110922
rect 675312 110786 675340 110894
rect 674668 110758 675340 110786
rect 675404 110772 675432 110894
rect 675114 110392 675170 110401
rect 675114 110327 675170 110336
rect 675128 110174 675156 110327
rect 675128 110146 675418 110174
rect 675758 108216 675814 108225
rect 675758 108151 675814 108160
rect 675772 107644 675800 108151
rect 675312 107222 675432 107250
rect 675312 107114 675340 107222
rect 675128 107086 675340 107114
rect 675404 107100 675432 107222
rect 675128 106321 675156 107086
rect 675114 106312 675170 106321
rect 675114 106247 675170 106256
rect 675772 106185 675800 106488
rect 675758 106176 675814 106185
rect 675758 106111 675814 106120
rect 675312 105862 675432 105890
rect 675312 105822 675340 105862
rect 675128 105794 675340 105822
rect 675404 105808 675432 105862
rect 675128 105641 675156 105794
rect 675114 105632 675170 105641
rect 675114 105567 675170 105576
rect 674484 104638 675340 104666
rect 675312 104530 675340 104638
rect 675404 104530 675432 104652
rect 675312 104502 675432 104530
rect 675666 103184 675722 103193
rect 675666 103119 675722 103128
rect 675680 102816 675708 103119
rect 675666 102504 675722 102513
rect 675666 102439 675722 102448
rect 674286 102368 674342 102377
rect 674286 102303 674342 102312
rect 675680 102136 675708 102439
rect 675758 101416 675814 101425
rect 675758 101351 675814 101360
rect 675772 100980 675800 101351
rect 668306 95840 668362 95849
rect 668306 95775 668362 95784
rect 666572 84166 666692 84194
rect 648894 82240 648950 82249
rect 648894 82175 648950 82184
rect 648988 80844 649040 80850
rect 648988 80786 649040 80792
rect 648804 75472 648856 75478
rect 648804 75414 648856 75420
rect 648816 64874 648844 75414
rect 649000 71777 649028 80786
rect 649172 77988 649224 77994
rect 649172 77930 649224 77936
rect 648986 71768 649042 71777
rect 648986 71703 649042 71712
rect 648632 64846 648844 64874
rect 648632 62121 648660 64846
rect 649184 64433 649212 77930
rect 666572 76566 666600 84166
rect 666560 76560 666612 76566
rect 666560 76502 666612 76508
rect 662604 75200 662656 75206
rect 662604 75142 662656 75148
rect 649170 64424 649226 64433
rect 649170 64359 649226 64368
rect 648618 62112 648674 62121
rect 648618 62047 648674 62056
rect 647238 57352 647294 57361
rect 647238 57287 647294 57296
rect 625804 52284 625856 52290
rect 625804 52226 625856 52232
rect 662418 48512 662474 48521
rect 662418 48447 662474 48456
rect 661590 47789 661646 47798
rect 661590 47724 661646 47733
rect 661604 46510 661632 47724
rect 623044 46504 623096 46510
rect 623044 46446 623096 46452
rect 661592 46504 661644 46510
rect 661592 46446 661644 46452
rect 464710 44296 464766 44305
rect 464710 44231 464766 44240
rect 463882 44160 463938 44169
rect 463882 44095 463938 44104
rect 465814 43616 465870 43625
rect 465814 43551 465870 43560
rect 463698 42936 463754 42945
rect 463698 42871 463754 42880
rect 463056 42764 463108 42770
rect 463056 42706 463108 42712
rect 460938 42392 460994 42401
rect 463712 42378 463740 42871
rect 465828 42500 465856 43551
rect 471058 43344 471114 43353
rect 471058 43279 471114 43288
rect 463712 42350 464036 42378
rect 460938 42327 460994 42336
rect 471072 42106 471100 43279
rect 518806 42800 518862 42809
rect 518806 42735 518862 42744
rect 518820 42364 518848 42735
rect 662432 42231 662460 48447
rect 662616 47433 662644 75142
rect 662602 47424 662658 47433
rect 662602 47359 662658 47368
rect 662420 42225 662472 42231
rect 662420 42167 662472 42173
rect 515402 42120 515458 42129
rect 459940 42078 460368 42106
rect 471072 42078 471408 42106
rect 515154 42078 515402 42106
rect 520922 42120 520978 42129
rect 520674 42078 520922 42106
rect 515402 42055 515458 42064
rect 522118 42120 522174 42129
rect 521870 42078 522118 42106
rect 520922 42055 520978 42064
rect 526442 42120 526498 42129
rect 526194 42078 526442 42106
rect 522118 42055 522174 42064
rect 529570 42120 529626 42129
rect 529322 42078 529570 42106
rect 526442 42055 526498 42064
rect 529570 42055 529626 42064
rect 404452 41472 404504 41478
rect 404452 41414 404504 41420
rect 420736 41472 420788 41478
rect 420736 41414 420788 41420
rect 427084 41472 427136 41478
rect 427084 41414 427136 41420
rect 459192 41472 459244 41478
rect 459192 41414 459244 41420
rect 141698 40488 141754 40497
rect 141698 40423 141754 40432
rect 141712 39984 141740 40423
<< via2 >>
rect 202694 1007412 202750 1007448
rect 202694 1007392 202696 1007412
rect 202696 1007392 202748 1007412
rect 202748 1007392 202750 1007412
rect 153750 1006596 153806 1006632
rect 153750 1006576 153752 1006596
rect 153752 1006576 153804 1006596
rect 153804 1006576 153806 1006596
rect 102322 1006460 102378 1006496
rect 102322 1006440 102324 1006460
rect 102324 1006440 102376 1006460
rect 102376 1006440 102378 1006460
rect 81254 995696 81310 995752
rect 86498 995560 86554 995616
rect 87786 995560 87842 995616
rect 90178 995560 90234 995616
rect 77206 995288 77262 995344
rect 84474 995016 84530 995072
rect 81990 994744 82046 994800
rect 85026 994472 85082 994528
rect 92478 997192 92534 997248
rect 92662 996920 92718 996976
rect 92478 996376 92534 996432
rect 89350 995016 89406 995072
rect 101954 1006324 102010 1006360
rect 101954 1006304 101956 1006324
rect 101956 1006304 102008 1006324
rect 102008 1006304 102010 1006324
rect 103978 1006188 104034 1006224
rect 103978 1006168 103980 1006188
rect 103980 1006168 104032 1006188
rect 104032 1006168 104034 1006188
rect 107658 1006188 107714 1006224
rect 107658 1006168 107660 1006188
rect 107660 1006168 107712 1006188
rect 107712 1006168 107714 1006188
rect 98274 1006052 98330 1006088
rect 98274 1006032 98276 1006052
rect 98276 1006032 98328 1006052
rect 98328 1006032 98330 1006052
rect 100298 1002652 100354 1002688
rect 100298 1002632 100300 1002652
rect 100300 1002632 100352 1002652
rect 100352 1002632 100354 1002652
rect 94502 996648 94558 996704
rect 85670 994200 85726 994256
rect 95146 994200 95202 994256
rect 42154 968768 42210 968824
rect 42154 967544 42210 967600
rect 42798 967544 42854 967600
rect 41970 967136 42026 967192
rect 42430 966728 42486 966784
rect 44546 968768 44602 968824
rect 43442 966728 43498 966784
rect 42430 964688 42486 964744
rect 42430 963872 42486 963928
rect 44362 964688 44418 964744
rect 44178 963872 44234 963928
rect 42430 963328 42486 963384
rect 43166 963328 43222 963384
rect 42430 963056 42486 963112
rect 41786 962104 41842 962160
rect 41786 959792 41842 959848
rect 41786 959112 41842 959168
rect 42982 963056 43038 963112
rect 42430 958704 42486 958760
rect 42062 957888 42118 957944
rect 41786 955440 41842 955496
rect 28538 952856 28594 952912
rect 28538 942656 28594 942712
rect 39302 952176 39358 952232
rect 37922 938984 37978 939040
rect 36542 938406 36598 938462
rect 42062 951904 42118 951960
rect 40038 951768 40094 951824
rect 39302 937352 39358 937408
rect 41418 951632 41474 951688
rect 41234 943064 41290 943120
rect 41234 941840 41290 941896
rect 41142 939392 41198 939448
rect 40958 938406 41014 938462
rect 40038 934496 40094 934552
rect 42062 937760 42118 937816
rect 42062 935720 42118 935776
rect 43718 958704 43774 958760
rect 43442 952856 43498 952912
rect 43534 940208 43590 940264
rect 43166 934904 43222 934960
rect 42982 934088 43038 934144
rect 42246 932864 42302 932920
rect 43350 932048 43406 932104
rect 41694 911920 41750 911976
rect 41510 911648 41566 911704
rect 42936 892472 42992 892528
rect 43074 891948 43130 891984
rect 43074 891928 43076 891948
rect 43076 891928 43128 891948
rect 43128 891928 43130 891948
rect 41602 885400 41658 885456
rect 41418 885128 41474 885184
rect 41234 817264 41290 817320
rect 41234 816448 41290 816504
rect 42062 884584 42118 884640
rect 41786 814000 41842 814056
rect 40958 813184 41014 813240
rect 40774 812776 40830 812832
rect 39302 811552 39358 811608
rect 33046 811144 33102 811200
rect 41142 812368 41198 812424
rect 42982 810328 43038 810384
rect 41970 808288 42026 808344
rect 41786 807200 41842 807256
rect 40958 805568 41014 805624
rect 42246 806656 42302 806712
rect 41970 805024 42026 805080
rect 41602 801660 41604 801680
rect 41604 801660 41656 801680
rect 41656 801660 41658 801680
rect 41602 801624 41658 801660
rect 41786 800264 41842 800320
rect 41786 799856 41842 799912
rect 42798 807880 42854 807936
rect 42614 801624 42670 801680
rect 42154 797272 42210 797328
rect 42154 796184 42210 796240
rect 42062 794960 42118 795016
rect 41786 794416 41842 794472
rect 41786 793736 41842 793792
rect 42706 794960 42762 795016
rect 43166 809512 43222 809568
rect 43166 796184 43222 796240
rect 42246 792512 42302 792568
rect 42430 792240 42486 792296
rect 42154 789384 42210 789440
rect 42798 789384 42854 789440
rect 42338 789112 42394 789168
rect 42614 788704 42670 788760
rect 42246 788160 42302 788216
rect 42430 788160 42486 788216
rect 42798 788568 42854 788624
rect 35806 773880 35862 773936
rect 35346 769392 35402 769448
rect 35530 768984 35586 769040
rect 35806 769004 35862 769040
rect 35806 768984 35808 769004
rect 35808 768984 35860 769004
rect 35860 768984 35862 769004
rect 35622 768168 35678 768224
rect 31022 767760 31078 767816
rect 35806 767760 35862 767816
rect 35162 766944 35218 767000
rect 35806 763292 35862 763328
rect 35806 763272 35808 763292
rect 35808 763272 35860 763292
rect 35860 763272 35862 763292
rect 36542 759056 36598 759112
rect 43074 766672 43130 766728
rect 41326 765312 41382 765368
rect 42522 765312 42578 765368
rect 42798 764632 42854 764688
rect 40314 757968 40370 758024
rect 39302 757696 39358 757752
rect 42154 757832 42210 757888
rect 40314 757424 40370 757480
rect 41786 755384 41842 755440
rect 42062 754024 42118 754080
rect 42246 753616 42302 753672
rect 41970 752936 42026 752992
rect 42614 753344 42670 753400
rect 42246 751984 42302 752040
rect 42062 751712 42118 751768
rect 41786 751032 41842 751088
rect 41786 750352 41842 750408
rect 42246 749400 42302 749456
rect 42430 749264 42486 749320
rect 42246 746544 42302 746600
rect 41970 746000 42026 746056
rect 42062 745456 42118 745512
rect 42430 746272 42486 746328
rect 42798 751712 42854 751768
rect 43074 749264 43130 749320
rect 42614 745456 42670 745512
rect 42706 745048 42762 745104
rect 42706 743008 42762 743064
rect 35806 730904 35862 730960
rect 41326 726416 41382 726472
rect 41142 726008 41198 726064
rect 39302 725192 39358 725248
rect 36542 724784 36598 724840
rect 31666 724376 31722 724432
rect 34518 723968 34574 724024
rect 34150 720316 34206 720352
rect 34150 720296 34152 720316
rect 34152 720296 34204 720316
rect 34204 720296 34206 720316
rect 31666 715400 31722 715456
rect 40682 723152 40738 723208
rect 40314 715128 40370 715184
rect 38658 714448 38714 714504
rect 41326 725600 41382 725656
rect 41142 721712 41198 721768
rect 43074 719752 43130 719808
rect 41878 719480 41934 719536
rect 42522 719480 42578 719536
rect 41694 719072 41750 719128
rect 42338 715128 42394 715184
rect 40682 714176 40738 714232
rect 41510 714176 41566 714232
rect 42062 714448 42118 714504
rect 41786 713904 41842 713960
rect 41786 713496 41842 713552
rect 42154 711320 42210 711376
rect 42154 711048 42210 711104
rect 42706 719072 42762 719128
rect 42614 711320 42670 711376
rect 41786 709824 41842 709880
rect 42246 709144 42302 709200
rect 42062 708464 42118 708520
rect 42062 707784 42118 707840
rect 42062 706696 42118 706752
rect 42246 705472 42302 705528
rect 41786 704248 41842 704304
rect 42890 710776 42946 710832
rect 42890 708464 42946 708520
rect 42430 702344 42486 702400
rect 42246 702072 42302 702128
rect 42062 701800 42118 701856
rect 42706 701800 42762 701856
rect 42614 701528 42670 701584
rect 35622 691328 35678 691384
rect 41418 689288 41474 689344
rect 35806 687656 35862 687712
rect 35622 687248 35678 687304
rect 35806 683188 35862 683224
rect 35806 683168 35808 683188
rect 35808 683168 35860 683188
rect 35860 683168 35862 683188
rect 35438 682760 35494 682816
rect 35622 682352 35678 682408
rect 35806 681980 35808 682000
rect 35808 681980 35860 682000
rect 35860 681980 35862 682000
rect 35806 681944 35862 681980
rect 32402 681536 32458 681592
rect 31022 681128 31078 681184
rect 35162 680720 35218 680776
rect 31022 672696 31078 672752
rect 41694 681844 41696 681864
rect 41696 681844 41748 681864
rect 41748 681844 41750 681864
rect 41694 681808 41750 681844
rect 41786 678544 41842 678600
rect 41326 677048 41382 677104
rect 42522 681808 42578 681864
rect 42798 679904 42854 679960
rect 41326 672424 41382 672480
rect 41326 671064 41382 671120
rect 39670 670928 39726 670984
rect 42154 672152 42210 672208
rect 41786 670656 41842 670712
rect 41786 670248 41842 670304
rect 42614 671064 42670 671120
rect 41786 669024 41842 669080
rect 42246 668888 42302 668944
rect 42246 667800 42302 667856
rect 41970 667664 42026 667720
rect 42246 667528 42302 667584
rect 42062 666984 42118 667040
rect 42062 666576 42118 666632
rect 42062 665624 42118 665680
rect 41786 665352 41842 665408
rect 42154 665080 42210 665136
rect 42154 664808 42210 664864
rect 41970 663992 42026 664048
rect 43074 676640 43130 676696
rect 42890 666576 42946 666632
rect 42522 662904 42578 662960
rect 42706 662768 42762 662824
rect 42338 662496 42394 662552
rect 42154 661000 42210 661056
rect 42154 660456 42210 660512
rect 42706 659776 42762 659832
rect 42154 658960 42210 659016
rect 42338 658552 42394 658608
rect 42154 657328 42210 657384
rect 42522 658280 42578 658336
rect 42706 657328 42762 657384
rect 35806 646720 35862 646776
rect 35806 644680 35862 644736
rect 41786 641620 41842 641676
rect 41786 641144 41842 641200
rect 35622 639784 35678 639840
rect 35806 639376 35862 639432
rect 35806 638560 35862 638616
rect 32402 638152 32458 638208
rect 42338 633800 42394 633856
rect 36542 630672 36598 630728
rect 42154 624416 42210 624472
rect 42430 624416 42486 624472
rect 42246 623736 42302 623792
rect 42062 623328 42118 623384
rect 42062 620880 42118 620936
rect 42706 620336 42762 620392
rect 42246 619656 42302 619712
rect 42522 618568 42578 618624
rect 42062 618296 42118 618352
rect 42246 617616 42302 617672
rect 42062 617072 42118 617128
rect 42062 616528 42118 616584
rect 42522 616528 42578 616584
rect 42154 615848 42210 615904
rect 42890 616120 42946 616176
rect 42614 615440 42670 615496
rect 42246 615168 42302 615224
rect 41786 614080 41842 614136
rect 43718 936128 43774 936184
rect 45558 943472 45614 943528
rect 44822 941432 44878 941488
rect 44546 936944 44602 937000
rect 44362 935312 44418 935368
rect 44178 933680 44234 933736
rect 46938 933272 46994 933328
rect 44086 892764 44142 892800
rect 44086 892744 44088 892764
rect 44088 892744 44140 892764
rect 44140 892744 44142 892764
rect 44086 892200 44142 892256
rect 44178 816040 44234 816096
rect 43534 814816 43590 814872
rect 43534 807608 43590 807664
rect 43718 806248 43774 806304
rect 45006 815224 45062 815280
rect 44362 814408 44418 814464
rect 44178 773200 44234 773256
rect 44638 813592 44694 813648
rect 44454 771976 44510 772032
rect 44270 771568 44326 771624
rect 44270 770344 44326 770400
rect 43902 763000 43958 763056
rect 44822 809920 44878 809976
rect 44822 792240 44878 792296
rect 44822 772792 44878 772848
rect 44638 770752 44694 770808
rect 44638 766264 44694 766320
rect 44638 754840 44694 754896
rect 45190 810736 45246 810792
rect 45374 799040 45430 799096
rect 45374 797272 45430 797328
rect 45190 788160 45246 788216
rect 45006 772384 45062 772440
rect 45006 771160 45062 771216
rect 44822 730088 44878 730144
rect 44638 729680 44694 729736
rect 44454 729272 44510 729328
rect 44270 727640 44326 727696
rect 44454 723560 44510 723616
rect 44178 722744 44234 722800
rect 44178 707784 44234 707840
rect 44454 705472 44510 705528
rect 45558 764224 45614 764280
rect 45190 728864 45246 728920
rect 45006 728456 45062 728512
rect 44914 721112 44970 721168
rect 44638 686840 44694 686896
rect 44362 686432 44418 686488
rect 44178 679496 44234 679552
rect 44178 667528 44234 667584
rect 44546 679088 44602 679144
rect 44730 677864 44786 677920
rect 44546 661000 44602 661056
rect 44362 643592 44418 643648
rect 44178 636520 44234 636576
rect 44362 636248 44418 636304
rect 44178 635296 44234 635352
rect 44086 625232 44142 625288
rect 44546 635704 44602 635760
rect 44362 624416 44418 624472
rect 44178 620880 44234 620936
rect 44546 619656 44602 619712
rect 44086 616120 44142 616176
rect 43074 611904 43130 611960
rect 43929 611904 43985 611960
rect 45374 721520 45430 721576
rect 45374 710776 45430 710832
rect 45190 686024 45246 686080
rect 45282 685616 45338 685672
rect 45098 643320 45154 643376
rect 42522 610952 42578 611008
rect 44500 610952 44556 611008
rect 45282 643048 45338 643104
rect 45374 642504 45430 642560
rect 46202 754024 46258 754080
rect 45742 728048 45798 728104
rect 46110 727368 46166 727424
rect 45742 685208 45798 685264
rect 45926 684800 45982 684856
rect 45742 683984 45798 684040
rect 46110 684392 46166 684448
rect 46110 680312 46166 680368
rect 46110 660456 46166 660512
rect 45926 642232 45982 642288
rect 45742 641416 45798 641472
rect 45926 641144 45982 641200
rect 45742 633392 45798 633448
rect 45098 600480 45154 600536
rect 44638 600072 44694 600128
rect 42982 596944 43038 597000
rect 42154 596808 42210 596864
rect 41234 595992 41290 596048
rect 33046 595584 33102 595640
rect 31022 594360 31078 594416
rect 35162 595176 35218 595232
rect 40682 594768 40738 594824
rect 40498 593136 40554 593192
rect 39946 590688 40002 590744
rect 40498 589600 40554 589656
rect 40314 589328 40370 589384
rect 40406 586472 40462 586528
rect 41694 594496 41750 594552
rect 41786 593544 41842 593600
rect 40682 584568 40738 584624
rect 41786 592728 41842 592784
rect 41786 592320 41842 592376
rect 41786 589464 41842 589520
rect 42614 594496 42670 594552
rect 42798 593952 42854 594008
rect 42062 586744 42118 586800
rect 42522 586472 42578 586528
rect 41694 584840 41750 584896
rect 41786 584296 41842 584352
rect 42338 581712 42394 581768
rect 41970 581440 42026 581496
rect 42246 580760 42302 580816
rect 42430 580760 42486 580816
rect 41970 580216 42026 580272
rect 41786 578176 41842 578232
rect 41786 577496 41842 577552
rect 42154 577088 42210 577144
rect 41970 576544 42026 576600
rect 42154 574096 42210 574152
rect 44454 591912 44510 591968
rect 43442 591504 43498 591560
rect 43166 584840 43222 584896
rect 43166 580760 43222 580816
rect 42890 577904 42946 577960
rect 42706 577496 42762 577552
rect 42614 573280 42670 573336
rect 42522 572056 42578 572112
rect 41786 570152 41842 570208
rect 42338 569200 42394 569256
rect 35806 558048 35862 558104
rect 42062 558456 42118 558512
rect 42062 557504 42118 557560
rect 35806 554804 35862 554840
rect 35806 554784 35808 554804
rect 35808 554784 35860 554804
rect 35860 554784 35862 554804
rect 35806 553560 35862 553616
rect 33782 551928 33838 551984
rect 31758 548086 31814 548142
rect 41326 552744 41382 552800
rect 41694 551792 41750 551848
rect 43074 551520 43130 551576
rect 41786 550704 41842 550760
rect 40498 549888 40554 549944
rect 41234 548140 41290 548142
rect 41234 548088 41236 548140
rect 41236 548088 41288 548140
rect 41288 548088 41290 548140
rect 41234 548086 41290 548088
rect 41970 550296 42026 550352
rect 41786 548392 41842 548448
rect 41694 548140 41750 548176
rect 41694 548120 41696 548140
rect 41696 548120 41748 548140
rect 41748 548120 41750 548140
rect 40498 545400 40554 545456
rect 42890 548392 42946 548448
rect 41970 545672 42026 545728
rect 41786 541048 41842 541104
rect 41786 540640 41842 540696
rect 42614 540232 42670 540288
rect 42246 538192 42302 538248
rect 42062 537920 42118 537976
rect 42614 537920 42670 537976
rect 42614 537376 42670 537432
rect 42246 536288 42302 536344
rect 41786 535200 41842 535256
rect 42522 534248 42578 534304
rect 42430 533296 42486 533352
rect 42706 532616 42762 532672
rect 42430 530168 42486 530224
rect 42062 529896 42118 529952
rect 41878 529352 41934 529408
rect 42706 529896 42762 529952
rect 42706 529624 42762 529680
rect 41326 425992 41382 426048
rect 40958 425584 41014 425640
rect 33782 424360 33838 424416
rect 41786 422728 41842 422784
rect 41142 418784 41198 418840
rect 41786 418512 41842 418568
rect 42798 423952 42854 424008
rect 42522 419872 42578 419928
rect 42062 411848 42118 411904
rect 42614 411848 42670 411904
rect 41786 409400 41842 409456
rect 42430 408448 42486 408504
rect 42430 407768 42486 407824
rect 42062 406680 42118 406736
rect 41786 406272 41842 406328
rect 42430 405592 42486 405648
rect 41786 403824 41842 403880
rect 42338 402872 42394 402928
rect 42430 402464 42486 402520
rect 41786 401920 41842 401976
rect 42430 399744 42486 399800
rect 43258 420688 43314 420744
rect 43074 419192 43130 419248
rect 41786 398792 41842 398848
rect 42062 387640 42118 387696
rect 41878 387232 41934 387288
rect 41142 387096 41198 387152
rect 42062 386688 42118 386744
rect 41878 386416 41934 386472
rect 42062 386416 42118 386472
rect 35438 383016 35494 383072
rect 35622 382608 35678 382664
rect 35806 382200 35862 382256
rect 35530 381384 35586 381440
rect 35806 381384 35862 381440
rect 35806 376488 35862 376544
rect 41510 382236 41512 382256
rect 41512 382236 41564 382256
rect 41564 382236 41566 382256
rect 41510 382200 41566 382236
rect 42798 382200 42854 382256
rect 41326 378528 41382 378584
rect 42338 378528 42394 378584
rect 40038 376896 40094 376952
rect 39578 375672 39634 375728
rect 37922 371320 37978 371376
rect 41786 368600 41842 368656
rect 42430 366968 42486 367024
rect 42430 365744 42486 365800
rect 41786 364248 41842 364304
rect 42430 364248 42486 364304
rect 41786 363704 41842 363760
rect 41786 362888 41842 362944
rect 41786 360032 41842 360088
rect 42154 359896 42210 359952
rect 41786 358672 41842 358728
rect 42430 357312 42486 357368
rect 42338 355952 42394 356008
rect 41878 355680 41934 355736
rect 43074 355544 43130 355600
rect 43626 590280 43682 590336
rect 44454 581032 44510 581088
rect 45374 599664 45430 599720
rect 44822 599256 44878 599312
rect 44638 557232 44694 557288
rect 46110 640872 46166 640928
rect 45926 598848 45982 598904
rect 45006 598440 45062 598496
rect 44822 556416 44878 556472
rect 48962 942248 49018 942304
rect 50342 940616 50398 940672
rect 51722 939800 51778 939856
rect 47582 891928 47638 891984
rect 47766 817672 47822 817728
rect 50342 816856 50398 816912
rect 47582 711048 47638 711104
rect 99470 1002516 99526 1002552
rect 99470 1002496 99472 1002516
rect 99472 1002496 99524 1002516
rect 99524 1002496 99526 1002516
rect 98274 1001972 98330 1002008
rect 98274 1001952 98276 1001972
rect 98276 1001952 98328 1001972
rect 98328 1001952 98330 1001972
rect 99102 1002108 99158 1002144
rect 99102 1002088 99104 1002108
rect 99104 1002088 99156 1002108
rect 99156 1002088 99158 1002108
rect 100298 1002380 100354 1002416
rect 100298 1002360 100300 1002380
rect 100300 1002360 100352 1002380
rect 100352 1002360 100354 1002380
rect 101126 1002244 101182 1002280
rect 101126 1002224 101128 1002244
rect 101128 1002224 101180 1002244
rect 101180 1002224 101182 1002244
rect 101126 1001952 101182 1002008
rect 98642 995832 98698 995888
rect 104806 1006052 104862 1006088
rect 104806 1006032 104808 1006052
rect 104808 1006032 104860 1006052
rect 104860 1006032 104862 1006052
rect 108486 1006052 108542 1006088
rect 108486 1006032 108488 1006052
rect 108488 1006032 108540 1006052
rect 108540 1006032 108542 1006052
rect 101954 1002108 102010 1002144
rect 101954 1002088 101956 1002108
rect 101956 1002088 102008 1002108
rect 102008 1002088 102010 1002108
rect 101402 995288 101458 995344
rect 97446 994744 97502 994800
rect 106830 1002652 106886 1002688
rect 106830 1002632 106832 1002652
rect 106832 1002632 106884 1002652
rect 106884 1002632 106886 1002652
rect 103150 1002516 103206 1002552
rect 103150 1002496 103152 1002516
rect 103152 1002496 103204 1002516
rect 103204 1002496 103206 1002516
rect 108026 1002516 108082 1002552
rect 108026 1002496 108028 1002516
rect 108028 1002496 108080 1002516
rect 108080 1002496 108082 1002516
rect 106002 1002380 106058 1002416
rect 106002 1002360 106004 1002380
rect 106004 1002360 106056 1002380
rect 106056 1002360 106058 1002380
rect 105634 1002244 105690 1002280
rect 105634 1002224 105636 1002244
rect 105636 1002224 105688 1002244
rect 105688 1002224 105690 1002244
rect 106830 1002108 106886 1002144
rect 106830 1002088 106832 1002108
rect 106832 1002088 106884 1002108
rect 106884 1002088 106886 1002108
rect 103150 1001972 103206 1002008
rect 103150 1001952 103152 1001972
rect 103152 1001952 103204 1001972
rect 103204 1001952 103206 1001972
rect 103978 1001952 104034 1002008
rect 106002 1001972 106058 1002008
rect 106002 1001952 106004 1001972
rect 106004 1001952 106056 1001972
rect 106056 1001952 106058 1001972
rect 97262 994472 97318 994528
rect 108854 1002244 108910 1002280
rect 108854 1002224 108856 1002244
rect 108856 1002224 108908 1002244
rect 108908 1002224 108910 1002244
rect 108854 1001972 108910 1002008
rect 108854 1001952 108856 1001972
rect 108856 1001952 108908 1001972
rect 108908 1001952 108910 1001972
rect 109682 1002108 109738 1002144
rect 109682 1002088 109684 1002108
rect 109684 1002088 109736 1002108
rect 109736 1002088 109738 1002108
rect 117226 997192 117282 997248
rect 116306 996920 116362 996976
rect 143814 997192 143870 997248
rect 143998 996648 144054 996704
rect 143998 996124 144054 996160
rect 143998 996104 144000 996124
rect 144000 996104 144052 996124
rect 144052 996104 144054 996124
rect 140410 995696 140466 995752
rect 141054 995696 141110 995752
rect 143630 995696 143686 995752
rect 136270 995560 136326 995616
rect 126242 995288 126298 995344
rect 124862 995016 124918 995072
rect 129094 994744 129150 994800
rect 132774 994200 132830 994256
rect 141698 995424 141754 995480
rect 141514 995288 141570 995344
rect 142066 995288 142122 995344
rect 137098 994472 137154 994528
rect 142066 994472 142122 994528
rect 139398 993928 139454 993984
rect 142342 993948 142398 993984
rect 142342 993928 142344 993948
rect 142344 993928 142396 993948
rect 142396 993928 142398 993948
rect 133878 993656 133934 993712
rect 144826 996920 144882 996976
rect 152094 1006460 152150 1006496
rect 152094 1006440 152096 1006460
rect 152096 1006440 152148 1006460
rect 152148 1006440 152150 1006460
rect 157430 1006460 157486 1006496
rect 157430 1006440 157432 1006460
rect 157432 1006440 157484 1006460
rect 157484 1006440 157486 1006460
rect 151726 1006324 151782 1006360
rect 151726 1006304 151728 1006324
rect 151728 1006304 151780 1006324
rect 151780 1006304 151782 1006324
rect 158258 1006324 158314 1006360
rect 158258 1006304 158260 1006324
rect 158260 1006304 158312 1006324
rect 158312 1006304 158314 1006324
rect 150898 1006188 150954 1006224
rect 150898 1006168 150900 1006188
rect 150900 1006168 150952 1006188
rect 150952 1006168 150954 1006188
rect 160282 1006188 160338 1006224
rect 160282 1006168 160284 1006188
rect 160284 1006168 160336 1006188
rect 160336 1006168 160338 1006188
rect 150070 1006052 150126 1006088
rect 150070 1006032 150072 1006052
rect 150072 1006032 150124 1006052
rect 150124 1006032 150126 1006052
rect 159454 1006052 159510 1006088
rect 159454 1006032 159456 1006052
rect 159456 1006032 159508 1006052
rect 159508 1006032 159510 1006052
rect 152922 1005372 152978 1005408
rect 152922 1005352 152924 1005372
rect 152924 1005352 152976 1005372
rect 152976 1005352 152978 1005372
rect 145562 993928 145618 993984
rect 142066 993692 142068 993712
rect 142068 993692 142120 993712
rect 142120 993692 142122 993712
rect 142066 993656 142122 993692
rect 142250 993676 142306 993712
rect 142250 993656 142252 993676
rect 142252 993656 142304 993676
rect 142304 993656 142306 993676
rect 144366 993656 144422 993712
rect 147678 996376 147734 996432
rect 149242 1001972 149298 1002008
rect 149242 1001952 149244 1001972
rect 149244 1001952 149296 1001972
rect 149296 1001952 149298 1001972
rect 152922 1005100 152978 1005136
rect 152922 1005080 152924 1005100
rect 152924 1005080 152976 1005100
rect 152976 1005080 152978 1005100
rect 149702 994472 149758 994528
rect 153750 1004964 153806 1005000
rect 153750 1004944 153752 1004964
rect 153752 1004944 153804 1004964
rect 153804 1004944 153806 1004964
rect 158626 1004964 158682 1005000
rect 158626 1004944 158628 1004964
rect 158628 1004944 158680 1004964
rect 158680 1004944 158682 1004964
rect 150898 1002108 150954 1002144
rect 150898 1002088 150900 1002108
rect 150900 1002088 150952 1002108
rect 150952 1002088 150954 1002108
rect 160650 1004828 160706 1004864
rect 160650 1004808 160652 1004828
rect 160652 1004808 160704 1004828
rect 160704 1004808 160706 1004828
rect 154118 1004692 154174 1004728
rect 154118 1004672 154120 1004692
rect 154120 1004672 154172 1004692
rect 154172 1004672 154174 1004692
rect 161110 1004692 161166 1004728
rect 161110 1004672 161112 1004692
rect 161112 1004672 161164 1004692
rect 161164 1004672 161166 1004692
rect 155774 1002516 155830 1002552
rect 155774 1002496 155776 1002516
rect 155776 1002496 155828 1002516
rect 155828 1002496 155830 1002516
rect 151726 1002244 151782 1002280
rect 151726 1002224 151728 1002244
rect 151728 1002224 151780 1002244
rect 151780 1002224 151782 1002244
rect 156602 1002380 156658 1002416
rect 156602 1002360 156604 1002380
rect 156604 1002360 156656 1002380
rect 156656 1002360 156658 1002380
rect 155774 1002244 155830 1002280
rect 155774 1002224 155776 1002244
rect 155776 1002224 155828 1002244
rect 155828 1002224 155830 1002244
rect 156602 1002108 156658 1002144
rect 156602 1002088 156604 1002108
rect 156604 1002088 156656 1002108
rect 156656 1002088 156658 1002108
rect 154578 1001972 154634 1002008
rect 154578 1001952 154580 1001972
rect 154580 1001952 154632 1001972
rect 154632 1001952 154634 1001972
rect 154946 1001972 155002 1002008
rect 154946 1001952 154948 1001972
rect 154948 1001952 155000 1001972
rect 155000 1001952 155002 1001972
rect 155130 995560 155186 995616
rect 155130 995016 155186 995072
rect 151082 994744 151138 994800
rect 157798 1001972 157854 1002008
rect 157798 1001952 157800 1001972
rect 157800 1001952 157852 1001972
rect 157852 1001952 157854 1001972
rect 149886 994200 149942 994256
rect 170310 997192 170366 997248
rect 195058 996376 195114 996432
rect 189446 995696 189502 995752
rect 190458 995696 190514 995752
rect 172426 995288 172482 995344
rect 184478 995016 184534 995072
rect 187606 995288 187662 995344
rect 184846 994744 184902 994800
rect 188158 994472 188214 994528
rect 190366 995016 190422 995072
rect 190550 995016 190606 995072
rect 195426 996648 195482 996704
rect 189078 994200 189134 994256
rect 183834 993520 183890 993576
rect 196806 996376 196862 996432
rect 505374 1007140 505430 1007176
rect 505374 1007120 505376 1007140
rect 505376 1007120 505428 1007140
rect 505428 1007120 505430 1007140
rect 357714 1006868 357770 1006904
rect 428002 1006884 428004 1006904
rect 428004 1006884 428056 1006904
rect 428056 1006884 428058 1006904
rect 357714 1006848 357716 1006868
rect 357716 1006848 357768 1006868
rect 357768 1006848 357770 1006868
rect 428002 1006848 428058 1006884
rect 505374 1006884 505376 1006904
rect 505376 1006884 505428 1006904
rect 505428 1006884 505430 1006904
rect 505374 1006848 505430 1006884
rect 360198 1006732 360254 1006768
rect 360198 1006712 360200 1006732
rect 360200 1006712 360252 1006732
rect 360252 1006712 360254 1006732
rect 210054 1006460 210110 1006496
rect 210054 1006440 210056 1006460
rect 210056 1006440 210108 1006460
rect 210108 1006440 210110 1006460
rect 306930 1006460 306986 1006496
rect 306930 1006440 306932 1006460
rect 306932 1006440 306984 1006460
rect 306984 1006440 306986 1006460
rect 201038 1006052 201094 1006088
rect 201038 1006032 201040 1006052
rect 201040 1006032 201092 1006052
rect 201092 1006032 201094 1006052
rect 202694 998708 202750 998744
rect 202694 998688 202696 998708
rect 202696 998688 202748 998708
rect 202748 998688 202750 998708
rect 200670 998028 200726 998064
rect 200670 998008 200672 998028
rect 200672 998008 200724 998028
rect 200724 998008 200726 998028
rect 201866 998164 201922 998200
rect 201866 998144 201868 998164
rect 201868 998144 201920 998164
rect 201920 998144 201922 998164
rect 200210 997228 200212 997248
rect 200212 997228 200264 997248
rect 200264 997228 200266 997248
rect 200210 997192 200266 997228
rect 200946 995696 201002 995752
rect 200762 994744 200818 994800
rect 198002 994472 198058 994528
rect 196622 994200 196678 994256
rect 202510 995832 202566 995888
rect 205546 1001972 205602 1002008
rect 205546 1001952 205548 1001972
rect 205548 1001952 205600 1001972
rect 205600 1001952 205602 1001972
rect 203890 998844 203946 998880
rect 203890 998824 203892 998844
rect 203892 998824 203944 998844
rect 203944 998824 203946 998844
rect 203890 998572 203946 998608
rect 203890 998552 203892 998572
rect 203892 998552 203944 998572
rect 203944 998552 203946 998572
rect 205546 998028 205602 998064
rect 205546 998008 205548 998028
rect 205548 998008 205600 998028
rect 205600 998008 205602 998028
rect 204718 997892 204774 997928
rect 204718 997872 204720 997892
rect 204720 997872 204772 997892
rect 204772 997872 204774 997892
rect 210422 1006324 210478 1006360
rect 210422 1006304 210424 1006324
rect 210424 1006304 210476 1006324
rect 210476 1006304 210478 1006324
rect 256146 1006324 256202 1006360
rect 256146 1006304 256148 1006324
rect 256148 1006304 256200 1006324
rect 256200 1006304 256202 1006324
rect 208398 1006188 208454 1006224
rect 208398 1006168 208400 1006188
rect 208400 1006168 208452 1006188
rect 208452 1006168 208454 1006188
rect 209226 1006052 209282 1006088
rect 209226 1006032 209228 1006052
rect 209228 1006032 209280 1006052
rect 209280 1006032 209282 1006052
rect 208398 1005116 208400 1005136
rect 208400 1005116 208452 1005136
rect 208452 1005116 208454 1005136
rect 208398 1005080 208454 1005116
rect 207570 1004980 207572 1005000
rect 207572 1004980 207624 1005000
rect 207624 1004980 207626 1005000
rect 207570 1004944 207626 1004980
rect 209226 1004828 209282 1004864
rect 209226 1004808 209228 1004828
rect 209228 1004808 209280 1004828
rect 209280 1004808 209282 1004828
rect 207202 1002496 207258 1002552
rect 206374 1002108 206430 1002144
rect 206374 1002088 206376 1002108
rect 206376 1002088 206428 1002108
rect 206428 1002088 206430 1002108
rect 206742 1001972 206798 1002008
rect 206742 1001952 206744 1001972
rect 206744 1001952 206796 1001972
rect 206796 1001952 206798 1001972
rect 207202 1002224 207258 1002280
rect 203522 995288 203578 995344
rect 210882 1002108 210938 1002144
rect 210882 1002088 210884 1002108
rect 210884 1002088 210936 1002108
rect 210936 1002088 210938 1002108
rect 211250 1002516 211306 1002552
rect 211250 1002496 211252 1002516
rect 211252 1002496 211304 1002516
rect 211304 1002496 211306 1002516
rect 211250 1002244 211306 1002280
rect 211250 1002224 211252 1002244
rect 211252 1002224 211304 1002244
rect 211304 1002224 211306 1002244
rect 212538 1004692 212594 1004728
rect 212538 1004672 212540 1004692
rect 212540 1004672 212592 1004692
rect 212592 1004672 212594 1004692
rect 212078 1001972 212134 1002008
rect 212078 1001952 212080 1001972
rect 212080 1001952 212132 1001972
rect 212132 1001952 212134 1001972
rect 202142 993520 202198 993576
rect 191838 992840 191894 992896
rect 240874 995696 240930 995752
rect 244094 995696 244150 995752
rect 246578 995696 246634 995752
rect 228362 995016 228418 995072
rect 236550 994744 236606 994800
rect 239586 994472 239642 994528
rect 238666 994200 238722 994256
rect 241978 995424 242034 995480
rect 243818 995424 243874 995480
rect 244002 995288 244058 995344
rect 240046 993928 240102 993984
rect 246946 996376 247002 996432
rect 247130 995288 247186 995344
rect 246946 994472 247002 994528
rect 255318 1006188 255374 1006224
rect 255318 1006168 255320 1006188
rect 255320 1006168 255372 1006188
rect 255372 1006168 255374 1006188
rect 261850 1006188 261906 1006224
rect 261850 1006168 261852 1006188
rect 261852 1006168 261904 1006188
rect 261904 1006168 261906 1006188
rect 252466 1006052 252522 1006088
rect 252466 1006032 252468 1006052
rect 252468 1006032 252520 1006052
rect 252520 1006032 252522 1006052
rect 260194 1006052 260250 1006088
rect 260194 1006032 260196 1006052
rect 260196 1006032 260248 1006052
rect 260248 1006032 260250 1006052
rect 263046 1004964 263102 1005000
rect 263046 1004944 263048 1004964
rect 263048 1004944 263100 1004964
rect 263100 1004944 263102 1004964
rect 256146 1002652 256202 1002688
rect 256146 1002632 256148 1002652
rect 256148 1002632 256200 1002652
rect 256200 1002632 256202 1002652
rect 250626 997192 250682 997248
rect 251638 996684 251640 996704
rect 251640 996684 251692 996704
rect 251692 996684 251694 996704
rect 251638 996648 251694 996684
rect 250442 995968 250498 996024
rect 252466 997772 252468 997792
rect 252468 997772 252520 997792
rect 252520 997772 252522 997792
rect 252466 997736 252522 997772
rect 254490 1002516 254546 1002552
rect 254490 1002496 254492 1002516
rect 254492 1002496 254544 1002516
rect 254544 1002496 254546 1002516
rect 261022 1002380 261078 1002416
rect 261022 1002360 261024 1002380
rect 261024 1002360 261076 1002380
rect 261076 1002360 261078 1002380
rect 262678 1002244 262734 1002280
rect 262678 1002224 262680 1002244
rect 262680 1002224 262732 1002244
rect 262732 1002224 262734 1002244
rect 254122 1002108 254178 1002144
rect 254122 1002088 254124 1002108
rect 254124 1002088 254176 1002108
rect 254176 1002088 254178 1002108
rect 263874 1002108 263930 1002144
rect 263874 1002088 263876 1002108
rect 263876 1002088 263928 1002108
rect 263928 1002088 263930 1002108
rect 255318 1001972 255374 1002008
rect 255318 1001952 255320 1001972
rect 255320 1001952 255372 1001972
rect 255372 1001952 255374 1001972
rect 263506 1001972 263562 1002008
rect 263506 1001952 263508 1001972
rect 263508 1001952 263560 1001972
rect 263560 1001952 263562 1001972
rect 259366 998300 259422 998336
rect 259366 998280 259368 998300
rect 259368 998280 259420 998300
rect 259420 998280 259422 998300
rect 253662 998164 253718 998200
rect 253662 998144 253664 998164
rect 253664 998144 253716 998164
rect 253716 998144 253718 998164
rect 258170 998164 258226 998200
rect 258170 998144 258172 998164
rect 258172 998144 258224 998164
rect 258224 998144 258226 998164
rect 257342 998044 257344 998064
rect 257344 998044 257396 998064
rect 257396 998044 257398 998064
rect 253662 997908 253664 997928
rect 253664 997908 253716 997928
rect 253716 997908 253718 997928
rect 253662 997872 253718 997908
rect 251822 994744 251878 994800
rect 257342 998008 257398 998044
rect 256514 997908 256516 997928
rect 256516 997908 256568 997928
rect 256568 997908 256570 997928
rect 256514 997872 256570 997908
rect 256974 997736 257030 997792
rect 258170 997872 258226 997928
rect 258998 997736 259054 997792
rect 259826 998044 259828 998064
rect 259828 998044 259880 998064
rect 259880 998044 259882 998064
rect 259826 998008 259882 998044
rect 260194 997908 260196 997928
rect 260196 997908 260248 997928
rect 260248 997908 260250 997928
rect 260194 997872 260250 997908
rect 261850 997736 261906 997792
rect 254766 994200 254822 994256
rect 249062 993928 249118 993984
rect 251454 992840 251510 992896
rect 298098 997872 298154 997928
rect 282734 995696 282790 995752
rect 287978 995696 288034 995752
rect 291750 995696 291806 995752
rect 293498 995696 293554 995752
rect 295062 995696 295118 995752
rect 296166 995560 296222 995616
rect 279422 995016 279478 995072
rect 286230 995288 286286 995344
rect 290278 994744 290334 994800
rect 290830 994200 290886 994256
rect 298742 996920 298798 996976
rect 299386 996512 299442 996568
rect 299386 996240 299442 996296
rect 299386 995696 299442 995752
rect 299202 995560 299258 995616
rect 299846 995968 299902 996024
rect 361394 1006324 361450 1006360
rect 361394 1006304 361396 1006324
rect 361396 1006304 361448 1006324
rect 361448 1006304 361450 1006324
rect 306102 1006188 306158 1006224
rect 306102 1006168 306104 1006188
rect 306104 1006168 306156 1006188
rect 306156 1006168 306158 1006188
rect 357346 1006188 357402 1006224
rect 357346 1006168 357348 1006188
rect 357348 1006168 357400 1006188
rect 357400 1006168 357402 1006188
rect 301686 1006032 301742 1006088
rect 303250 1006052 303306 1006088
rect 303250 1006032 303252 1006052
rect 303252 1006032 303304 1006052
rect 303304 1006032 303306 1006052
rect 300306 996376 300362 996432
rect 300122 994200 300178 994256
rect 304078 1006052 304134 1006088
rect 304078 1006032 304080 1006052
rect 304080 1006032 304132 1006052
rect 304132 1006032 304134 1006052
rect 311806 1006032 311862 1006088
rect 314658 1006052 314714 1006088
rect 314658 1006032 314660 1006052
rect 314660 1006032 314712 1006052
rect 314712 1006032 314714 1006052
rect 354862 1006032 354918 1006088
rect 356886 1006052 356942 1006088
rect 356886 1006032 356888 1006052
rect 356888 1006032 356940 1006052
rect 356940 1006032 356942 1006052
rect 304078 1005796 304080 1005816
rect 304080 1005796 304132 1005816
rect 304132 1005796 304134 1005816
rect 304078 1005760 304134 1005796
rect 313830 1004964 313886 1005000
rect 313830 1004944 313832 1004964
rect 313832 1004944 313884 1004964
rect 313884 1004944 313886 1004964
rect 314658 1004828 314714 1004864
rect 314658 1004808 314660 1004828
rect 314660 1004808 314712 1004828
rect 314712 1004808 314714 1004828
rect 315486 1004692 315542 1004728
rect 315486 1004672 315488 1004692
rect 315488 1004672 315540 1004692
rect 315540 1004672 315542 1004692
rect 304906 1002108 304962 1002144
rect 304906 1002088 304908 1002108
rect 304908 1002088 304960 1002108
rect 304960 1002088 304962 1002108
rect 310150 1002108 310206 1002144
rect 310150 1002088 310152 1002108
rect 310152 1002088 310204 1002108
rect 310204 1002088 310206 1002108
rect 310978 1001972 311034 1002008
rect 310978 1001952 310980 1001972
rect 310980 1001952 311032 1001972
rect 311032 1001952 311034 1001972
rect 308954 998572 309010 998608
rect 308954 998552 308956 998572
rect 308956 998552 309008 998572
rect 309008 998552 309010 998572
rect 301686 995968 301742 996024
rect 307298 998436 307354 998472
rect 307298 998416 307300 998436
rect 307300 998416 307352 998436
rect 307352 998416 307354 998436
rect 303250 997872 303306 997928
rect 302882 995696 302938 995752
rect 303250 997228 303252 997248
rect 303252 997228 303304 997248
rect 303304 997228 303306 997248
rect 303250 997192 303306 997228
rect 306102 998300 306158 998336
rect 306102 998280 306104 998300
rect 306104 998280 306156 998300
rect 306156 998280 306158 998300
rect 308126 998164 308182 998200
rect 308126 998144 308128 998164
rect 308128 998144 308180 998164
rect 308180 998144 308182 998164
rect 305274 997892 305330 997928
rect 305274 997872 305276 997892
rect 305276 997872 305328 997892
rect 305328 997872 305330 997892
rect 306930 998028 306986 998064
rect 306930 998008 306932 998028
rect 306932 998008 306984 998028
rect 306984 998008 306986 998028
rect 310610 998028 310666 998064
rect 310610 998008 310612 998028
rect 310612 998008 310664 998028
rect 310664 998008 310666 998028
rect 307758 997736 307814 997792
rect 308954 997892 309010 997928
rect 308954 997872 308956 997892
rect 308956 997872 309008 997892
rect 309008 997872 309010 997892
rect 310610 997736 310666 997792
rect 307022 994744 307078 994800
rect 354034 1001972 354090 1002008
rect 354034 1001952 354036 1001972
rect 354036 1001952 354088 1001972
rect 354088 1001952 354090 1001972
rect 360566 1005524 360568 1005544
rect 360568 1005524 360620 1005544
rect 360620 1005524 360622 1005544
rect 360566 1005488 360622 1005524
rect 358542 1005388 358544 1005408
rect 358544 1005388 358596 1005408
rect 358596 1005388 358598 1005408
rect 358542 1005352 358598 1005388
rect 357714 1005252 357716 1005272
rect 357716 1005252 357768 1005272
rect 357768 1005252 357770 1005272
rect 357714 1005216 357770 1005252
rect 355690 1004828 355746 1004864
rect 355690 1004808 355692 1004828
rect 355692 1004808 355744 1004828
rect 355744 1004808 355746 1004828
rect 356518 1004692 356574 1004728
rect 356518 1004672 356520 1004692
rect 356520 1004672 356572 1004692
rect 356572 1004672 356574 1004692
rect 360566 1003892 360568 1003912
rect 360568 1003892 360620 1003912
rect 360620 1003892 360622 1003912
rect 360566 1003856 360622 1003892
rect 355690 1003332 355746 1003368
rect 355690 1003312 355692 1003332
rect 355692 1003312 355744 1003332
rect 355744 1003312 355746 1003332
rect 358542 1002532 358544 1002552
rect 358544 1002532 358596 1002552
rect 358596 1002532 358598 1002552
rect 358542 1002496 358598 1002532
rect 359370 1002244 359426 1002280
rect 359370 1002224 359372 1002244
rect 359372 1002224 359424 1002244
rect 359424 1002224 359426 1002244
rect 359370 1001972 359426 1002008
rect 359370 1001952 359372 1001972
rect 359372 1001952 359424 1001972
rect 359424 1001952 359426 1001972
rect 361394 1004964 361450 1005000
rect 361394 1004944 361396 1004964
rect 361396 1004944 361448 1004964
rect 361448 1004944 361450 1004964
rect 363418 1006052 363474 1006088
rect 363418 1006032 363420 1006052
rect 363420 1006032 363472 1006052
rect 363472 1006032 363474 1006052
rect 362590 1004828 362646 1004864
rect 362590 1004808 362592 1004828
rect 362592 1004808 362644 1004828
rect 362644 1004808 362646 1004828
rect 364246 1004692 364302 1004728
rect 364246 1004672 364248 1004692
rect 364248 1004672 364300 1004692
rect 364300 1004672 364302 1004692
rect 365074 1002260 365076 1002280
rect 365076 1002260 365128 1002280
rect 365128 1002260 365130 1002280
rect 365074 1002224 365130 1002260
rect 365074 1001988 365076 1002008
rect 365076 1001988 365128 1002008
rect 365128 1001988 365130 1002008
rect 365074 1001952 365130 1001988
rect 365902 1002124 365904 1002144
rect 365904 1002124 365956 1002144
rect 365956 1002124 365958 1002144
rect 365902 1002088 365958 1002124
rect 430854 1006748 430856 1006768
rect 430856 1006748 430908 1006768
rect 430908 1006748 430910 1006768
rect 430854 1006712 430910 1006748
rect 506202 1006748 506204 1006768
rect 506204 1006748 506256 1006768
rect 506256 1006748 506258 1006768
rect 430026 1006476 430028 1006496
rect 430028 1006476 430080 1006496
rect 430080 1006476 430082 1006496
rect 430026 1006440 430082 1006476
rect 429198 1006324 429254 1006360
rect 429198 1006304 429200 1006324
rect 429200 1006304 429252 1006324
rect 429252 1006304 429254 1006324
rect 373262 998280 373318 998336
rect 372342 997192 372398 997248
rect 372526 996376 372582 996432
rect 372342 995968 372398 996024
rect 374642 994880 374698 994936
rect 380898 995424 380954 995480
rect 383382 996648 383438 996704
rect 383198 995696 383254 995752
rect 399942 996920 399998 996976
rect 400126 996376 400182 996432
rect 431682 1006440 431738 1006496
rect 431682 1006204 431684 1006224
rect 431684 1006204 431736 1006224
rect 431736 1006204 431738 1006224
rect 431682 1006168 431738 1006204
rect 421838 1006032 421894 1006088
rect 428370 1006052 428426 1006088
rect 428370 1006032 428372 1006052
rect 428372 1006032 428424 1006052
rect 428424 1006032 428426 1006052
rect 385682 995696 385738 995752
rect 386694 995696 386750 995752
rect 387890 995696 387946 995752
rect 388166 995696 388222 995752
rect 391938 995696 391994 995752
rect 396538 995696 396594 995752
rect 416134 995696 416190 995752
rect 382278 995152 382334 995208
rect 395158 994880 395214 994936
rect 415398 995444 415454 995480
rect 415398 995424 415400 995444
rect 415400 995424 415452 995444
rect 415452 995424 415454 995444
rect 425518 1005660 425520 1005680
rect 425520 1005660 425572 1005680
rect 425572 1005660 425574 1005680
rect 425518 1005624 425574 1005660
rect 427174 1005524 427176 1005544
rect 427176 1005524 427228 1005544
rect 427228 1005524 427230 1005544
rect 427174 1005488 427230 1005524
rect 428370 1005388 428372 1005408
rect 428372 1005388 428424 1005408
rect 428424 1005388 428426 1005408
rect 428370 1005352 428426 1005388
rect 423494 1005252 423496 1005272
rect 423496 1005252 423548 1005272
rect 423548 1005252 423550 1005272
rect 423494 1005216 423550 1005252
rect 431222 1004964 431278 1005000
rect 431222 1004944 431224 1004964
rect 431224 1004944 431276 1004964
rect 431276 1004944 431278 1004964
rect 422666 1004828 422722 1004864
rect 422666 1004808 422668 1004828
rect 422668 1004808 422720 1004828
rect 422720 1004808 422722 1004828
rect 432050 1004828 432106 1004864
rect 432050 1004808 432052 1004828
rect 432052 1004808 432104 1004828
rect 432104 1004808 432106 1004828
rect 430026 1004692 430082 1004728
rect 430026 1004672 430028 1004692
rect 430028 1004672 430080 1004692
rect 430080 1004672 430082 1004692
rect 424690 1004028 424692 1004048
rect 424692 1004028 424744 1004048
rect 424744 1004028 424746 1004048
rect 424690 1003992 424746 1004028
rect 426346 1003892 426348 1003912
rect 426348 1003892 426400 1003912
rect 426400 1003892 426402 1003912
rect 426346 1003856 426402 1003892
rect 423494 1002532 423496 1002552
rect 423496 1002532 423548 1002552
rect 423548 1002532 423550 1002552
rect 423494 1002496 423550 1002532
rect 425518 1002108 425574 1002144
rect 425518 1002088 425520 1002108
rect 425520 1002088 425572 1002108
rect 425572 1002088 425574 1002108
rect 427542 1002108 427598 1002144
rect 427542 1002088 427544 1002108
rect 427544 1002088 427596 1002108
rect 427596 1002088 427598 1002108
rect 421470 1001972 421526 1002008
rect 424322 1001988 424324 1002008
rect 424324 1001988 424376 1002008
rect 424376 1001988 424378 1002008
rect 421470 1001952 421472 1001972
rect 421472 1001952 421524 1001972
rect 421524 1001952 421526 1001972
rect 424322 1001952 424378 1001988
rect 425150 1001952 425206 1002008
rect 426346 1001952 426402 1002008
rect 429198 1001972 429254 1002008
rect 429198 1001952 429200 1001972
rect 429200 1001952 429252 1001972
rect 429252 1001952 429254 1001972
rect 433338 1002108 433394 1002144
rect 433338 1002088 433340 1002108
rect 433340 1002088 433392 1002108
rect 433392 1002088 433394 1002108
rect 432878 1001972 432934 1002008
rect 432878 1001952 432880 1001972
rect 432880 1001952 432932 1001972
rect 432932 1001952 432934 1001972
rect 506202 1006712 506258 1006748
rect 508226 1006460 508282 1006496
rect 508226 1006440 508228 1006460
rect 508228 1006440 508280 1006460
rect 508280 1006440 508282 1006460
rect 439686 996920 439742 996976
rect 439870 996376 439926 996432
rect 460938 995560 460994 995616
rect 458822 994472 458878 994528
rect 467102 998144 467158 998200
rect 507030 1006188 507086 1006224
rect 507030 1006168 507032 1006188
rect 507032 1006168 507084 1006188
rect 507084 1006168 507086 1006188
rect 498842 1006052 498898 1006088
rect 498842 1006032 498844 1006052
rect 498844 1006032 498896 1006052
rect 498896 1006032 498898 1006052
rect 502522 1006052 502578 1006088
rect 502522 1006032 502524 1006052
rect 502524 1006032 502576 1006052
rect 502576 1006032 502578 1006052
rect 509054 1006052 509110 1006088
rect 509054 1006032 509056 1006052
rect 509056 1006032 509108 1006052
rect 509108 1006032 509110 1006052
rect 505006 1005660 505008 1005680
rect 505008 1005660 505060 1005680
rect 505060 1005660 505062 1005680
rect 505006 1005624 505062 1005660
rect 502154 1005388 502156 1005408
rect 502156 1005388 502208 1005408
rect 502208 1005388 502210 1005408
rect 502154 1005352 502210 1005388
rect 499670 1005252 499672 1005272
rect 499672 1005252 499724 1005272
rect 499724 1005252 499726 1005272
rect 499670 1005216 499726 1005252
rect 500498 1005100 500554 1005136
rect 500498 1005080 500500 1005100
rect 500500 1005080 500552 1005100
rect 500552 1005080 500554 1005100
rect 500498 1004828 500554 1004864
rect 500498 1004808 500500 1004828
rect 500500 1004808 500552 1004828
rect 500552 1004808 500554 1004828
rect 471242 995968 471298 996024
rect 469862 995016 469918 995072
rect 469218 994744 469274 994800
rect 472254 996648 472310 996704
rect 472438 995696 472494 995752
rect 488998 996920 489054 996976
rect 494058 996376 494114 996432
rect 474002 995696 474058 995752
rect 474738 995696 474794 995752
rect 477038 995696 477094 995752
rect 481454 995696 481510 995752
rect 482742 995696 482798 995752
rect 485594 995696 485650 995752
rect 487986 995696 488042 995752
rect 488906 995696 488962 995752
rect 471886 994200 471942 994256
rect 477682 995424 477738 995480
rect 476762 994200 476818 994256
rect 482282 994744 482338 994800
rect 501326 1004692 501382 1004728
rect 501326 1004672 501328 1004692
rect 501328 1004672 501380 1004692
rect 501380 1004672 501382 1004692
rect 498474 1001972 498530 1002008
rect 498474 1001952 498476 1001972
rect 498476 1001952 498528 1001972
rect 498528 1001952 498530 1001972
rect 504546 1003892 504548 1003912
rect 504548 1003892 504600 1003912
rect 504600 1003892 504602 1003912
rect 504546 1003856 504602 1003892
rect 503350 1002380 503406 1002416
rect 503350 1002360 503352 1002380
rect 503352 1002360 503404 1002380
rect 503404 1002360 503406 1002380
rect 504178 1002244 504234 1002280
rect 504178 1002224 504180 1002244
rect 504180 1002224 504232 1002244
rect 504232 1002224 504234 1002244
rect 501694 1001972 501750 1002008
rect 501694 1001952 501696 1001972
rect 501696 1001952 501748 1001972
rect 501748 1001952 501750 1001972
rect 502522 1002108 502578 1002144
rect 502522 1002088 502524 1002108
rect 502524 1002088 502576 1002108
rect 502576 1002088 502578 1002108
rect 503350 1001972 503406 1002008
rect 503350 1001952 503352 1001972
rect 503352 1001952 503404 1001972
rect 503404 1001952 503406 1001972
rect 502062 995560 502118 995616
rect 502062 995016 502118 995072
rect 507858 1004828 507914 1004864
rect 507858 1004808 507860 1004828
rect 507860 1004808 507912 1004828
rect 507912 1004808 507914 1004828
rect 507398 1004692 507454 1004728
rect 507398 1004672 507400 1004692
rect 507400 1004672 507452 1004692
rect 507452 1004672 507454 1004692
rect 506202 1001952 506258 1002008
rect 554778 1006884 554780 1006904
rect 554780 1006884 554832 1006904
rect 554832 1006884 554834 1006904
rect 509882 1002108 509938 1002144
rect 509882 1002088 509884 1002108
rect 509884 1002088 509936 1002108
rect 509936 1002088 509938 1002108
rect 510342 1001972 510398 1002008
rect 510342 1001952 510344 1001972
rect 510344 1001952 510396 1001972
rect 510396 1001952 510398 1001972
rect 468482 993928 468538 993984
rect 481086 993928 481142 993984
rect 516690 996648 516746 996704
rect 516874 996376 516930 996432
rect 517334 996920 517390 996976
rect 517150 995832 517206 995888
rect 516966 995560 517022 995616
rect 516690 995288 516746 995344
rect 554778 1006848 554834 1006884
rect 555974 1006748 555976 1006768
rect 555976 1006748 556028 1006768
rect 556028 1006748 556030 1006768
rect 555974 1006712 556030 1006748
rect 518898 996104 518954 996160
rect 559654 1006460 559710 1006496
rect 559654 1006440 559656 1006460
rect 559656 1006440 559708 1006460
rect 559708 1006440 559710 1006460
rect 556802 1006188 556858 1006224
rect 556802 1006168 556804 1006188
rect 556804 1006168 556856 1006188
rect 556856 1006168 556858 1006188
rect 551098 1006032 551154 1006088
rect 555146 1006052 555202 1006088
rect 555146 1006032 555148 1006052
rect 555148 1006032 555200 1006052
rect 555200 1006032 555202 1006052
rect 520922 995016 520978 995072
rect 520186 994744 520242 994800
rect 553122 1005388 553124 1005408
rect 553124 1005388 553176 1005408
rect 553176 1005388 553178 1005408
rect 553122 1005352 553178 1005388
rect 551466 1005252 551468 1005272
rect 551468 1005252 551520 1005272
rect 551520 1005252 551522 1005272
rect 551466 1005216 551522 1005252
rect 555974 1004828 556030 1004864
rect 555974 1004808 555976 1004828
rect 555976 1004808 556028 1004828
rect 556028 1004808 556030 1004828
rect 552294 1003892 552296 1003912
rect 552296 1003892 552348 1003912
rect 552348 1003892 552350 1003912
rect 552294 1003856 552350 1003892
rect 553950 1002244 554006 1002280
rect 553950 1002224 553952 1002244
rect 553952 1002224 554004 1002244
rect 554004 1002224 554006 1002244
rect 550270 1001172 550272 1001192
rect 550272 1001172 550324 1001192
rect 550324 1001172 550326 1001192
rect 550270 1001136 550326 1001172
rect 552294 998436 552350 998472
rect 552294 998416 552296 998436
rect 552296 998416 552348 998436
rect 552348 998416 552350 998436
rect 551466 998028 551522 998064
rect 551466 998008 551468 998028
rect 551468 998008 551520 998028
rect 551520 998008 551522 998028
rect 524050 997192 524106 997248
rect 540886 996920 540942 996976
rect 524050 996648 524106 996704
rect 524786 995696 524842 995752
rect 532146 995696 532202 995752
rect 532790 995696 532846 995752
rect 535918 995696 535974 995752
rect 538218 995696 538274 995752
rect 529846 995424 529902 995480
rect 530214 995460 530216 995480
rect 530216 995460 530268 995480
rect 530268 995460 530270 995480
rect 530214 995424 530270 995460
rect 526350 994744 526406 994800
rect 536746 994744 536802 994800
rect 538034 994472 538090 994528
rect 553122 997892 553178 997928
rect 553122 997872 553124 997892
rect 553124 997872 553176 997892
rect 553176 997872 553178 997892
rect 553950 1001952 554006 1002008
rect 554778 1001952 554834 1002008
rect 557170 1006052 557226 1006088
rect 557170 1006032 557172 1006052
rect 557172 1006032 557224 1006052
rect 557224 1006032 557226 1006052
rect 557630 1004692 557686 1004728
rect 557630 1004672 557632 1004692
rect 557632 1004672 557684 1004692
rect 557684 1004672 557686 1004692
rect 557998 1002380 558054 1002416
rect 557998 1002360 558000 1002380
rect 558000 1002360 558052 1002380
rect 558052 1002360 558054 1002380
rect 560850 1004692 560906 1004728
rect 560850 1004672 560852 1004692
rect 560852 1004672 560904 1004692
rect 560904 1004672 560906 1004692
rect 558826 1002652 558882 1002688
rect 558826 1002632 558828 1002652
rect 558828 1002632 558880 1002652
rect 558880 1002632 558882 1002652
rect 558826 1001972 558882 1002008
rect 558826 1001952 558828 1001972
rect 558828 1001952 558880 1001972
rect 558880 1001952 558882 1001972
rect 560850 1002516 560906 1002552
rect 560850 1002496 560852 1002516
rect 560852 1002496 560904 1002516
rect 560904 1002496 560906 1002516
rect 560482 1002244 560538 1002280
rect 560482 1002224 560484 1002244
rect 560484 1002224 560536 1002244
rect 560536 1002224 560538 1002244
rect 560022 1002108 560078 1002144
rect 560022 1002088 560024 1002108
rect 560024 1002088 560076 1002108
rect 560076 1002088 560078 1002108
rect 561678 1001972 561734 1002008
rect 561678 1001952 561680 1001972
rect 561680 1001952 561732 1001972
rect 561732 1001952 561734 1001972
rect 570786 994744 570842 994800
rect 590566 996940 590622 996976
rect 590566 996920 590568 996940
rect 590568 996920 590620 996940
rect 590620 996920 590622 996940
rect 590566 996648 590622 996704
rect 590750 996376 590806 996432
rect 590566 995016 590622 995072
rect 622398 995968 622454 996024
rect 620282 995424 620338 995480
rect 626630 995696 626686 995752
rect 627182 995696 627238 995752
rect 627918 995696 627974 995752
rect 633990 995696 634046 995752
rect 635830 995696 635886 995752
rect 642086 995696 642142 995752
rect 631506 995424 631562 995480
rect 634542 994744 634598 994800
rect 576306 990936 576362 990992
rect 660578 995035 660634 995072
rect 660578 995016 660580 995035
rect 660580 995016 660632 995035
rect 660632 995016 660634 995035
rect 62118 975976 62174 976032
rect 651654 975840 651710 975896
rect 62118 962920 62174 962976
rect 651470 962512 651526 962568
rect 62118 949864 62174 949920
rect 652206 949320 652262 949376
rect 651470 936128 651526 936184
rect 661682 957752 661738 957808
rect 660302 941704 660358 941760
rect 665822 939800 665878 939856
rect 672538 952176 672594 952232
rect 669962 938440 670018 938496
rect 668582 937624 668638 937680
rect 667202 937080 667258 937136
rect 670974 936400 671030 936456
rect 658922 935992 658978 936048
rect 669226 929464 669282 929520
rect 62118 923752 62174 923808
rect 651470 922664 651526 922720
rect 62118 910696 62174 910752
rect 652390 909492 652446 909528
rect 652390 909472 652392 909492
rect 652392 909472 652444 909492
rect 652444 909472 652446 909492
rect 62118 897776 62174 897832
rect 651470 896144 651526 896200
rect 55862 892744 55918 892800
rect 54482 892472 54538 892528
rect 53286 892200 53342 892256
rect 651654 882816 651710 882872
rect 62118 871664 62174 871720
rect 651470 869624 651526 869680
rect 62118 858608 62174 858664
rect 651470 856296 651526 856352
rect 62118 845552 62174 845608
rect 53102 799040 53158 799096
rect 651838 842968 651894 843024
rect 62762 832496 62818 832552
rect 62118 819440 62174 819496
rect 62118 806520 62174 806576
rect 62118 793620 62174 793656
rect 62118 793600 62120 793620
rect 62120 793600 62172 793620
rect 62172 793600 62174 793620
rect 54482 774288 54538 774344
rect 51722 773472 51778 773528
rect 50342 730496 50398 730552
rect 48962 669296 49018 669352
rect 47306 637880 47362 637936
rect 47122 637608 47178 637664
rect 47122 618568 47178 618624
rect 47306 615576 47362 615632
rect 46110 598032 46166 598088
rect 47766 636928 47822 636984
rect 51722 691328 51778 691384
rect 51722 646584 51778 646640
rect 651470 829776 651526 829832
rect 651470 816448 651526 816504
rect 651470 803276 651526 803312
rect 651470 803256 651472 803276
rect 651472 803256 651524 803276
rect 651524 803256 651526 803276
rect 651470 789928 651526 789984
rect 62762 788568 62818 788624
rect 62762 780408 62818 780464
rect 62118 767372 62174 767408
rect 62118 767352 62120 767372
rect 62120 767352 62172 767372
rect 62172 767352 62174 767372
rect 62118 754296 62174 754352
rect 652390 776600 652446 776656
rect 651470 763292 651526 763328
rect 651470 763272 651472 763292
rect 651472 763272 651524 763292
rect 651524 763272 651526 763292
rect 651470 750080 651526 750136
rect 62762 743008 62818 743064
rect 62118 741240 62174 741296
rect 651838 736752 651894 736808
rect 55862 730088 55918 730144
rect 62762 728184 62818 728240
rect 62118 715264 62174 715320
rect 62118 702208 62174 702264
rect 54482 688064 54538 688120
rect 53102 644680 53158 644736
rect 50342 626592 50398 626648
rect 47766 618296 47822 618352
rect 51722 601704 51778 601760
rect 48962 601296 49018 601352
rect 651470 723424 651526 723480
rect 660302 778912 660358 778968
rect 658922 715944 658978 716000
rect 652574 710232 652630 710288
rect 652390 696940 652392 696960
rect 652392 696940 652444 696960
rect 652444 696940 652446 696960
rect 652390 696904 652446 696940
rect 62762 689424 62818 689480
rect 62118 689152 62174 689208
rect 651838 683576 651894 683632
rect 62118 676096 62174 676152
rect 652390 670384 652446 670440
rect 62118 663040 62174 663096
rect 651654 657056 651710 657112
rect 62118 649984 62174 650040
rect 651470 643728 651526 643784
rect 55862 643184 55918 643240
rect 62118 637064 62174 637120
rect 651562 630536 651618 630592
rect 62118 624008 62174 624064
rect 651470 617208 651526 617264
rect 62118 610952 62174 611008
rect 54482 600888 54538 600944
rect 47582 582392 47638 582448
rect 48962 557776 49018 557832
rect 50342 557504 50398 557560
rect 45650 556824 45706 556880
rect 45006 555600 45062 555656
rect 44638 555192 44694 555248
rect 44270 554376 44326 554432
rect 43810 548120 43866 548176
rect 43994 547032 44050 547088
rect 44454 552336 44510 552392
rect 44454 534248 44510 534304
rect 44914 551112 44970 551168
rect 45098 549480 45154 549536
rect 44822 548664 44878 548720
rect 44822 536832 44878 536888
rect 45282 549072 45338 549128
rect 45374 537376 45430 537432
rect 45282 533296 45338 533352
rect 45006 532616 45062 532672
rect 46018 556008 46074 556064
rect 45650 429664 45706 429720
rect 45834 429256 45890 429312
rect 45650 428440 45706 428496
rect 44638 428032 44694 428088
rect 44730 427624 44786 427680
rect 44270 427216 44326 427272
rect 44270 426808 44326 426864
rect 44454 423136 44510 423192
rect 44454 402872 44510 402928
rect 45098 423544 45154 423600
rect 44914 422320 44970 422376
rect 44914 405592 44970 405648
rect 45466 421504 45522 421560
rect 45282 421096 45338 421152
rect 45282 407768 45338 407824
rect 45466 406680 45522 406736
rect 45098 402464 45154 402520
rect 45282 386008 45338 386064
rect 45098 385192 45154 385248
rect 44730 384784 44786 384840
rect 44270 383968 44326 384024
rect 44546 379888 44602 379944
rect 44178 377440 44234 377496
rect 44362 376216 44418 376272
rect 44914 379480 44970 379536
rect 44730 379072 44786 379128
rect 46018 428848 46074 428904
rect 45834 387232 45890 387288
rect 45650 385600 45706 385656
rect 45834 384376 45890 384432
rect 45650 383560 45706 383616
rect 44822 365744 44878 365800
rect 44822 364248 44878 364304
rect 44178 356632 44234 356688
rect 44638 359896 44694 359952
rect 44454 356224 44510 356280
rect 43810 355272 43866 355328
rect 44638 355544 44694 355600
rect 44822 355272 44878 355328
rect 43258 353640 43314 353696
rect 28538 351192 28594 351248
rect 45190 356632 45246 356688
rect 45190 356224 45246 356280
rect 45144 353676 45146 353696
rect 45146 353676 45198 353696
rect 45198 353676 45200 353696
rect 45144 353640 45200 353676
rect 40222 345480 40278 345536
rect 28538 343848 28594 343904
rect 35806 343848 35862 343904
rect 45466 343304 45522 343360
rect 44822 342488 44878 342544
rect 45466 341264 45522 341320
rect 35806 339768 35862 339824
rect 35162 338952 35218 339008
rect 33782 338136 33838 338192
rect 37554 336504 37610 336560
rect 42798 334600 42854 334656
rect 43166 334600 43222 334656
rect 44178 334600 44234 334656
rect 44362 334600 44418 334656
rect 35162 329024 35218 329080
rect 33782 327664 33838 327720
rect 41786 325352 41842 325408
rect 41878 324672 41934 324728
rect 42246 324264 42302 324320
rect 42246 323584 42302 323640
rect 42062 322768 42118 322824
rect 42430 321408 42486 321464
rect 42430 321136 42486 321192
rect 42430 320048 42486 320104
rect 41786 319912 41842 319968
rect 42982 334328 43038 334384
rect 42982 323584 43038 323640
rect 43626 322904 43682 322960
rect 43166 322768 43222 322824
rect 41786 316784 41842 316840
rect 42154 315968 42210 316024
rect 41786 315560 41842 315616
rect 42154 313656 42210 313712
rect 42430 312704 42486 312760
rect 41970 312568 42026 312624
rect 41786 303048 41842 303104
rect 41786 300872 41842 300928
rect 42798 297200 42854 297256
rect 41786 296792 41842 296848
rect 41326 295976 41382 296032
rect 39302 294752 39358 294808
rect 41786 292848 41842 292904
rect 41786 292168 41842 292224
rect 41326 290264 41382 290320
rect 41970 281424 42026 281480
rect 42154 279792 42210 279848
rect 42430 278704 42486 278760
rect 42430 278160 42486 278216
rect 41786 277888 41842 277944
rect 42246 277616 42302 277672
rect 42062 277072 42118 277128
rect 42062 276664 42118 276720
rect 41786 274216 41842 274272
rect 42062 272992 42118 273048
rect 42062 272720 42118 272776
rect 41786 270408 41842 270464
rect 41786 269048 41842 269104
rect 42430 267688 42486 267744
rect 42982 295160 43038 295216
rect 43166 293120 43222 293176
rect 43442 291080 43498 291136
rect 43166 279792 43222 279848
rect 42982 276664 43038 276720
rect 35806 259936 35862 259992
rect 35806 258304 35862 258360
rect 42798 254768 42854 254824
rect 35622 253408 35678 253464
rect 35806 253000 35862 253056
rect 35806 252184 35862 252240
rect 34426 246880 34482 246936
rect 41694 242836 41696 242856
rect 41696 242836 41748 242856
rect 41748 242836 41750 242856
rect 41694 242800 41750 242836
rect 42430 242800 42486 242856
rect 40682 241440 40738 241496
rect 41786 240080 41842 240136
rect 42430 238040 42486 238096
rect 41786 235864 41842 235920
rect 42430 235864 42486 235920
rect 42246 234096 42302 234152
rect 42614 232464 42670 232520
rect 42430 232192 42486 232248
rect 42430 231784 42486 231840
rect 42154 230424 42210 230480
rect 41970 228928 42026 228984
rect 42430 227568 42486 227624
rect 42246 227296 42302 227352
rect 42430 226072 42486 226128
rect 42246 225528 42302 225584
rect 28538 222808 28594 222864
rect 42614 224848 42670 224904
rect 28538 214240 28594 214296
rect 41326 214240 41382 214296
rect 41142 212200 41198 212256
rect 43258 256400 43314 256456
rect 43166 255584 43222 255640
rect 42982 254360 43038 254416
rect 43258 213696 43314 213752
rect 42982 212880 43038 212936
rect 42798 212064 42854 212120
rect 41326 211792 41382 211848
rect 41326 210160 41382 210216
rect 41142 209752 41198 209808
rect 41326 209344 41382 209400
rect 41326 208936 41382 208992
rect 41142 207304 41198 207360
rect 40958 206896 41014 206952
rect 35806 204040 35862 204096
rect 41326 204448 41382 204504
rect 40958 203224 41014 203280
rect 35806 202136 35862 202192
rect 41694 208528 41750 208584
rect 42798 207576 42854 207632
rect 41510 200640 41566 200696
rect 41786 197104 41842 197160
rect 42154 195744 42210 195800
rect 41878 195200 41934 195256
rect 42430 193160 42486 193216
rect 42338 191664 42394 191720
rect 42430 191120 42486 191176
rect 42430 190440 42486 190496
rect 42430 189896 42486 189952
rect 42430 187584 42486 187640
rect 42430 186768 42486 186824
rect 42982 206352 43038 206408
rect 43258 203224 43314 203280
rect 42982 191120 43038 191176
rect 43258 186768 43314 186824
rect 41786 185816 41842 185872
rect 41786 184048 41842 184104
rect 42430 183096 42486 183152
rect 42430 180648 42486 180704
rect 44178 321136 44234 321192
rect 44362 320048 44418 320104
rect 44546 311344 44602 311400
rect 44362 311072 44418 311128
rect 44362 300056 44418 300112
rect 44178 299648 44234 299704
rect 43994 293528 44050 293584
rect 43810 291488 43866 291544
rect 43810 278160 43866 278216
rect 43994 272992 44050 273048
rect 43626 257624 43682 257680
rect 44546 299240 44602 299296
rect 45190 298832 45246 298888
rect 44362 298016 44418 298072
rect 44178 256808 44234 256864
rect 44822 294616 44878 294672
rect 44638 293936 44694 293992
rect 44546 272720 44602 272776
rect 44362 255176 44418 255232
rect 44178 253952 44234 254008
rect 43626 249056 43682 249112
rect 43810 241440 43866 241496
rect 43626 231784 43682 231840
rect 43810 227568 43866 227624
rect 44362 250280 44418 250336
rect 44546 248648 44602 248704
rect 44546 234096 44602 234152
rect 44362 230424 44418 230480
rect 45006 291760 45062 291816
rect 45006 277072 45062 277128
rect 47582 430072 47638 430128
rect 46938 426400 46994 426456
rect 46938 399744 46994 399800
rect 46938 380704 46994 380760
rect 46202 366968 46258 367024
rect 47122 380296 47178 380352
rect 47122 357312 47178 357368
rect 46938 355952 46994 356008
rect 45834 341672 45890 341728
rect 45650 340856 45706 340912
rect 45742 340040 45798 340096
rect 45926 338000 45982 338056
rect 45926 324264 45982 324320
rect 45742 313656 45798 313712
rect 45466 298424 45522 298480
rect 45466 294616 45522 294672
rect 45558 294344 45614 294400
rect 45558 267688 45614 267744
rect 47582 333104 47638 333160
rect 46202 257216 46258 257272
rect 45098 255992 45154 256048
rect 45558 252728 45614 252784
rect 45006 248240 45062 248296
rect 45006 235864 45062 235920
rect 47030 251912 47086 251968
rect 45834 251096 45890 251152
rect 45558 226072 45614 226128
rect 46018 249464 46074 249520
rect 46202 247832 46258 247888
rect 46018 232464 46074 232520
rect 45834 224848 45890 224904
rect 44822 214920 44878 214976
rect 44178 211248 44234 211304
rect 44178 207984 44234 208040
rect 43810 205536 43866 205592
rect 43626 202136 43682 202192
rect 43442 51720 43498 51776
rect 43994 205128 44050 205184
rect 43994 191664 44050 191720
rect 43810 190440 43866 190496
rect 44362 206760 44418 206816
rect 44638 205944 44694 206000
rect 44822 204720 44878 204776
rect 44546 203904 44602 203960
rect 44546 195744 44602 195800
rect 44362 193160 44418 193216
rect 44638 187584 44694 187640
rect 44178 183096 44234 183152
rect 47214 250688 47270 250744
rect 47030 232192 47086 232248
rect 47214 227296 47270 227352
rect 46938 209616 46994 209672
rect 46386 203496 46442 203552
rect 47122 208800 47178 208856
rect 47122 189896 47178 189952
rect 46938 180648 46994 180704
rect 50342 430888 50398 430944
rect 48962 386960 49018 387016
rect 48962 334056 49018 334112
rect 47766 300464 47822 300520
rect 47766 247424 47822 247480
rect 47950 213288 48006 213344
rect 48134 210840 48190 210896
rect 48134 194384 48190 194440
rect 47950 190440 48006 190496
rect 51722 386688 51778 386744
rect 51906 386416 51962 386472
rect 50526 351192 50582 351248
rect 50342 303048 50398 303104
rect 50342 290672 50398 290728
rect 49146 289856 49202 289912
rect 49330 208528 49386 208584
rect 49514 200640 49570 200696
rect 49330 196424 49386 196480
rect 49514 192344 49570 192400
rect 50526 246472 50582 246528
rect 54482 430480 54538 430536
rect 651470 603880 651526 603936
rect 62118 597896 62174 597952
rect 652390 590708 652446 590744
rect 652390 590688 652392 590708
rect 652392 590688 652444 590708
rect 652444 590688 652446 590708
rect 62118 584840 62174 584896
rect 664442 868672 664498 868728
rect 663062 760416 663118 760472
rect 661682 670656 661738 670712
rect 666466 879144 666522 879200
rect 666282 778368 666338 778424
rect 665822 761504 665878 761560
rect 664442 716488 664498 716544
rect 663062 689288 663118 689344
rect 661866 628496 661922 628552
rect 660302 625232 660358 625288
rect 660302 599528 660358 599584
rect 658922 579672 658978 579728
rect 651470 577360 651526 577416
rect 62118 571784 62174 571840
rect 62118 569200 62174 569256
rect 651654 564032 651710 564088
rect 62118 558728 62174 558784
rect 658922 553968 658978 554024
rect 651470 550840 651526 550896
rect 62118 545808 62174 545864
rect 56046 540232 56102 540288
rect 651470 537512 651526 537568
rect 62118 532772 62174 532808
rect 62118 532752 62120 532772
rect 62120 532752 62172 532772
rect 62172 532752 62174 532772
rect 651838 524184 651894 524240
rect 62118 519696 62174 519752
rect 651470 510992 651526 511048
rect 62118 506640 62174 506696
rect 652574 497664 652630 497720
rect 62118 493584 62174 493640
rect 651470 484492 651526 484528
rect 651470 484472 651472 484492
rect 651472 484472 651524 484492
rect 651524 484472 651526 484492
rect 62118 480528 62174 480584
rect 651470 471144 651526 471200
rect 62118 467472 62174 467528
rect 652390 457816 652446 457872
rect 62118 454552 62174 454608
rect 651470 444508 651526 444544
rect 651470 444488 651472 444508
rect 651472 444488 651524 444508
rect 651524 444488 651526 444508
rect 62118 441496 62174 441552
rect 651470 431296 651526 431352
rect 62118 428440 62174 428496
rect 651838 417968 651894 418024
rect 62762 415384 62818 415440
rect 55862 408448 55918 408504
rect 62118 402328 62174 402384
rect 54482 344256 54538 344312
rect 53102 321408 53158 321464
rect 51906 301280 51962 301336
rect 62118 389292 62174 389328
rect 62118 389272 62120 389292
rect 62120 389272 62172 389292
rect 62172 389272 62174 389292
rect 62118 376216 62174 376272
rect 62118 363296 62174 363352
rect 62118 350240 62174 350296
rect 651470 404640 651526 404696
rect 652574 391448 652630 391504
rect 652390 378156 652392 378176
rect 652392 378156 652444 378176
rect 652444 378156 652446 378176
rect 652390 378120 652446 378156
rect 651838 364792 651894 364848
rect 652390 351600 652446 351656
rect 62762 345616 62818 345672
rect 652022 338272 652078 338328
rect 62118 337184 62174 337240
rect 651470 324944 651526 325000
rect 651470 311752 651526 311808
rect 62118 311072 62174 311128
rect 62118 298172 62174 298208
rect 62118 298152 62120 298172
rect 62120 298152 62172 298172
rect 62172 298152 62174 298172
rect 651470 285232 651526 285288
rect 62762 285096 62818 285152
rect 55862 278704 55918 278760
rect 54482 259936 54538 259992
rect 51722 222808 51778 222864
rect 59266 224168 59322 224224
rect 102046 269728 102102 269784
rect 75918 267008 75974 267064
rect 138110 267008 138166 267064
rect 161294 269728 161350 269784
rect 467562 267008 467618 267064
rect 468758 269728 468814 269784
rect 470966 269184 471022 269240
rect 478602 271360 478658 271416
rect 497278 269456 497334 269512
rect 506110 268368 506166 268424
rect 507674 271088 507730 271144
rect 509698 267008 509754 267064
rect 513194 273808 513250 273864
rect 517150 267280 517206 267336
rect 519818 267552 519874 267608
rect 522394 274080 522450 274136
rect 521566 272720 521622 272776
rect 525154 275576 525210 275632
rect 525982 275596 526038 275632
rect 525982 275576 525984 275596
rect 525984 275576 526036 275596
rect 526036 275576 526038 275596
rect 529570 275168 529626 275224
rect 530950 270272 531006 270328
rect 533894 272448 533950 272504
rect 538034 270000 538090 270056
rect 537666 269728 537722 269784
rect 540518 269728 540574 269784
rect 539506 269184 539562 269240
rect 539690 267008 539746 267064
rect 551742 271360 551798 271416
rect 563702 267552 563758 267608
rect 568578 269456 568634 269512
rect 591026 268368 591082 268424
rect 593142 271088 593198 271144
rect 595442 274080 595498 274136
rect 602526 273808 602582 273864
rect 585782 267280 585838 267336
rect 614394 272720 614450 272776
rect 626170 275168 626226 275224
rect 626538 270272 626594 270328
rect 632150 272448 632206 272504
rect 625802 267008 625858 267064
rect 637578 270000 637634 270056
rect 640706 269728 640762 269784
rect 554410 262112 554466 262168
rect 554318 259936 554374 259992
rect 553950 257760 554006 257816
rect 553490 255584 553546 255640
rect 554410 253408 554466 253464
rect 554134 251252 554190 251288
rect 554134 251232 554136 251252
rect 554136 251232 554188 251252
rect 554188 251232 554190 251252
rect 553858 249056 553914 249112
rect 554410 246880 554466 246936
rect 553398 244704 553454 244760
rect 553950 242528 554006 242584
rect 554042 240352 554098 240408
rect 71042 230016 71098 230072
rect 65522 229744 65578 229800
rect 64142 228520 64198 228576
rect 62762 225528 62818 225584
rect 64786 222808 64842 222864
rect 66902 224440 66958 224496
rect 70858 218592 70914 218648
rect 73802 228248 73858 228304
rect 72422 224712 72478 224768
rect 71686 223080 71742 223136
rect 79966 226888 80022 226944
rect 77206 218864 77262 218920
rect 82542 225528 82598 225584
rect 89626 227160 89682 227216
rect 89166 225800 89222 225856
rect 92386 223352 92442 223408
rect 95698 221448 95754 221504
rect 97722 221720 97778 221776
rect 106922 230288 106978 230344
rect 108946 221992 109002 222048
rect 113086 228792 113142 228848
rect 118054 220088 118110 220144
rect 125506 226072 125562 226128
rect 124678 220360 124734 220416
rect 136362 227432 136418 227488
rect 143078 228520 143134 228576
rect 145010 224168 145066 224224
rect 148230 229744 148286 229800
rect 146850 223896 146906 223952
rect 146666 222808 146722 222864
rect 150806 230016 150862 230072
rect 149794 224440 149850 224496
rect 147586 220632 147642 220688
rect 151266 222808 151322 222864
rect 152738 224712 152794 224768
rect 152094 223080 152150 223136
rect 155314 228248 155370 228304
rect 153474 218592 153530 218648
rect 157522 218864 157578 218920
rect 160466 226888 160522 226944
rect 163042 225528 163098 225584
rect 166262 230288 166318 230344
rect 166906 227160 166962 227216
rect 169022 228248 169078 228304
rect 168194 225800 168250 225856
rect 167550 224168 167606 224224
rect 166906 218592 166962 218648
rect 170770 223352 170826 223408
rect 170586 221176 170642 221232
rect 172702 221720 172758 221776
rect 172978 221448 173034 221504
rect 176290 223896 176346 223952
rect 183650 221992 183706 222048
rect 184938 228792 184994 228848
rect 187882 220088 187938 220144
rect 193310 220360 193366 220416
rect 196530 226072 196586 226128
rect 199750 224168 199806 224224
rect 202970 227432 203026 227488
rect 206282 218592 206338 218648
rect 211342 220632 211398 220688
rect 213918 222808 213974 222864
rect 223578 228248 223634 228304
rect 229558 221176 229614 221232
rect 482742 222264 482798 222320
rect 485870 223624 485926 223680
rect 486606 223624 486662 223680
rect 488998 219408 489054 219464
rect 487802 218048 487858 218104
rect 490746 219136 490802 219192
rect 490562 218864 490618 218920
rect 491206 218864 491262 218920
rect 491942 218592 491998 218648
rect 492678 218320 492734 218376
rect 494794 219136 494850 219192
rect 493874 217640 493930 217696
rect 496818 223896 496874 223952
rect 497830 223896 497886 223952
rect 498842 217232 498898 217288
rect 501326 219680 501382 219736
rect 500222 219136 500278 219192
rect 500406 219136 500462 219192
rect 500038 218592 500094 218648
rect 500222 218592 500278 218648
rect 500222 217504 500278 217560
rect 503718 216960 503774 217016
rect 504546 219136 504602 219192
rect 504730 219156 504786 219192
rect 504730 219136 504732 219156
rect 504732 219136 504784 219156
rect 504784 219136 504786 219156
rect 504730 218864 504786 218920
rect 505282 218320 505338 218376
rect 505926 219952 505982 220008
rect 506294 219136 506350 219192
rect 507766 220224 507822 220280
rect 508870 217776 508926 217832
rect 508870 216960 508926 217016
rect 510710 220904 510766 220960
rect 512274 224168 512330 224224
rect 513470 221720 513526 221776
rect 514758 218592 514814 218648
rect 514942 218612 514998 218648
rect 514942 218592 514944 218612
rect 514944 218592 514996 218612
rect 514996 218592 514998 218612
rect 515770 221176 515826 221232
rect 518438 221448 518494 221504
rect 518806 220496 518862 220552
rect 519542 224440 519598 224496
rect 519542 223896 519598 223952
rect 523038 221992 523094 222048
rect 523406 221992 523462 222048
rect 524050 219172 524052 219192
rect 524052 219172 524104 219192
rect 524104 219172 524106 219192
rect 524050 219136 524106 219172
rect 524234 219136 524290 219192
rect 523774 218592 523830 218648
rect 524234 218592 524290 218648
rect 528558 220224 528614 220280
rect 528742 220224 528798 220280
rect 528282 219136 528338 219192
rect 528466 219172 528468 219192
rect 528468 219172 528520 219192
rect 528520 219172 528522 219192
rect 528466 219136 528522 219172
rect 528282 218628 528284 218648
rect 528284 218628 528336 218648
rect 528336 218628 528338 218648
rect 528282 218592 528338 218628
rect 528466 218592 528522 218648
rect 528650 218592 528706 218648
rect 529018 218592 529074 218648
rect 532698 221992 532754 222048
rect 532882 221992 532938 222048
rect 532882 221448 532938 221504
rect 533066 221448 533122 221504
rect 534078 220224 534134 220280
rect 534262 220224 534318 220280
rect 534262 219156 534318 219192
rect 534262 219136 534264 219156
rect 534264 219136 534316 219156
rect 534316 219136 534318 219156
rect 534446 219136 534502 219192
rect 534078 218592 534134 218648
rect 534262 218612 534318 218648
rect 534262 218592 534264 218612
rect 534264 218592 534316 218612
rect 534316 218592 534318 218612
rect 543738 220224 543794 220280
rect 543922 220224 543978 220280
rect 543462 219136 543518 219192
rect 543646 219136 543702 219192
rect 543922 219136 543978 219192
rect 544106 219136 544162 219192
rect 543462 218612 543518 218648
rect 543462 218592 543464 218612
rect 543464 218592 543516 218612
rect 543516 218592 543518 218612
rect 543922 218592 543978 218648
rect 554318 238176 554374 238232
rect 554502 236036 554504 236056
rect 554504 236036 554556 236056
rect 554556 236036 554558 236056
rect 554502 236000 554558 236036
rect 554410 233824 554466 233880
rect 552570 219136 552626 219192
rect 553122 220224 553178 220280
rect 553306 220224 553362 220280
rect 552938 219136 552994 219192
rect 553490 218864 553546 218920
rect 553122 218612 553178 218648
rect 553122 218592 553124 218612
rect 553124 218592 553176 218612
rect 553176 218592 553178 218612
rect 553306 218592 553362 218648
rect 553490 217776 553546 217832
rect 553214 217540 553216 217560
rect 553216 217540 553268 217560
rect 553268 217540 553270 217560
rect 553214 217504 553270 217540
rect 553490 216960 553546 217016
rect 553858 218900 553860 218920
rect 553860 218900 553912 218920
rect 553912 218900 553914 218920
rect 553858 218864 553914 218900
rect 553858 218612 553914 218648
rect 553858 218592 553860 218612
rect 553860 218592 553912 218612
rect 553912 218592 553914 218612
rect 554226 217540 554228 217560
rect 554228 217540 554280 217560
rect 554280 217540 554282 217560
rect 554226 217504 554282 217540
rect 562782 218864 562838 218920
rect 563058 218864 563114 218920
rect 563058 218320 563114 218376
rect 563242 218320 563298 218376
rect 562874 217812 562876 217832
rect 562876 217812 562928 217832
rect 562928 217812 562930 217832
rect 562874 217776 562930 217812
rect 563058 217252 563114 217288
rect 563058 217232 563060 217252
rect 563060 217232 563112 217252
rect 563112 217232 563114 217252
rect 563242 217232 563298 217288
rect 571706 216960 571762 217016
rect 572442 218320 572498 218376
rect 576582 218320 576638 218376
rect 576766 218320 576822 218376
rect 576582 217524 576638 217560
rect 576582 217504 576584 217524
rect 576584 217504 576636 217524
rect 576636 217504 576638 217524
rect 576766 217504 576822 217560
rect 572350 217232 572406 217288
rect 572534 217232 572590 217288
rect 575386 217232 575442 217288
rect 576950 216960 577006 217016
rect 577134 216688 577190 216744
rect 575386 216416 575442 216472
rect 578882 213968 578938 214024
rect 578514 211656 578570 211712
rect 578422 209788 578424 209808
rect 578424 209788 578476 209808
rect 578476 209788 578478 209808
rect 578422 209752 578478 209788
rect 579526 207440 579582 207496
rect 579526 205828 579582 205864
rect 579526 205808 579528 205828
rect 579528 205808 579580 205828
rect 579580 205808 579582 205828
rect 578514 203224 578570 203280
rect 578790 200776 578846 200832
rect 579526 198872 579582 198928
rect 578514 196424 578570 196480
rect 579526 194928 579582 194984
rect 579526 192208 579582 192264
rect 579526 190712 579582 190768
rect 579526 187992 579582 188048
rect 579526 186260 579528 186280
rect 579528 186260 579580 186280
rect 579580 186260 579582 186280
rect 579526 186224 579582 186260
rect 579526 184320 579582 184376
rect 579526 181872 579582 181928
rect 578790 180104 578846 180160
rect 579526 177656 579582 177712
rect 578790 175072 578846 175128
rect 578422 173440 578478 173496
rect 578238 170992 578294 171048
rect 578422 169224 578478 169280
rect 579526 166912 579582 166968
rect 579526 164464 579582 164520
rect 579342 162696 579398 162752
rect 578238 159840 578294 159896
rect 578422 158344 578478 158400
rect 578514 155896 578570 155952
rect 578698 153992 578754 154048
rect 578238 151680 578294 151736
rect 578330 149640 578386 149696
rect 579526 147464 579582 147520
rect 578606 138760 578662 138816
rect 579434 144644 579436 144664
rect 579436 144644 579488 144664
rect 579488 144644 579490 144664
rect 579434 144608 579490 144644
rect 579526 142976 579582 143032
rect 579526 140564 579528 140584
rect 579528 140564 579580 140584
rect 579580 140564 579582 140584
rect 579526 140528 579582 140564
rect 578882 136584 578938 136640
rect 579526 134408 579582 134464
rect 579066 132232 579122 132288
rect 578698 129648 578754 129704
rect 578514 127744 578570 127800
rect 578514 121080 578570 121136
rect 578514 114452 578516 114472
rect 578516 114452 578568 114472
rect 578568 114452 578570 114472
rect 578514 114416 578570 114452
rect 578882 110336 578938 110392
rect 578330 108296 578386 108352
rect 579526 125332 579528 125352
rect 579528 125332 579580 125352
rect 579580 125332 579582 125352
rect 579526 125296 579582 125332
rect 579250 123528 579306 123584
rect 579526 118396 579528 118416
rect 579528 118396 579580 118416
rect 579580 118396 579582 118416
rect 579526 118360 579582 118396
rect 579342 116864 579398 116920
rect 579526 112648 579582 112704
rect 579066 105848 579122 105904
rect 579250 103300 579252 103320
rect 579252 103300 579304 103320
rect 579304 103300 579306 103320
rect 579250 103264 579306 103300
rect 578330 101668 578332 101688
rect 578332 101668 578384 101688
rect 578384 101668 578386 101688
rect 578330 101632 578386 101668
rect 578606 99340 578662 99376
rect 578606 99320 578608 99340
rect 578608 99320 578660 99340
rect 578660 99320 578662 99340
rect 579250 97416 579306 97472
rect 129186 51720 129242 51776
rect 130474 44240 130530 44296
rect 308034 50224 308090 50280
rect 458086 48184 458142 48240
rect 457902 47912 457958 47968
rect 457718 47640 457774 47696
rect 458270 46824 458326 46880
rect 462594 52264 462650 52320
rect 461766 51992 461822 52048
rect 466642 52264 466698 52320
rect 466642 51584 466698 51640
rect 466458 48184 466514 48240
rect 466642 47912 466698 47968
rect 459006 47368 459062 47424
rect 458454 46552 458510 46608
rect 431222 44784 431278 44840
rect 132590 44276 132592 44296
rect 132592 44276 132644 44296
rect 132644 44276 132646 44296
rect 132590 44240 132646 44276
rect 142618 44240 142674 44296
rect 307298 44104 307354 44160
rect 194322 42064 194378 42120
rect 419722 43832 419778 43888
rect 415398 43560 415454 43616
rect 439594 43596 439596 43616
rect 439596 43596 439648 43616
rect 439648 43596 439650 43616
rect 439594 43560 439650 43596
rect 441618 43596 441620 43616
rect 441620 43596 441672 43616
rect 441672 43596 441674 43616
rect 441618 43560 441674 43596
rect 361946 41792 362002 41848
rect 365166 41792 365222 41848
rect 416686 42200 416742 42256
rect 446402 42200 446458 42256
rect 446402 41520 446458 41576
rect 460110 44784 460166 44840
rect 460754 43288 460810 43344
rect 462870 43832 462926 43888
rect 461582 43560 461638 43616
rect 462686 43560 462742 43616
rect 461398 42880 461454 42936
rect 463698 44376 463754 44432
rect 465078 46824 465134 46880
rect 466826 47640 466882 47696
rect 467010 47368 467066 47424
rect 545670 49408 545726 49464
rect 549994 48864 550050 48920
rect 579250 94968 579306 95024
rect 579342 93100 579344 93120
rect 579344 93100 579396 93120
rect 579396 93100 579398 93120
rect 579342 93064 579398 93100
rect 578238 90888 578294 90944
rect 579342 88032 579398 88088
rect 578790 86436 578792 86456
rect 578792 86436 578844 86456
rect 578844 86436 578846 86456
rect 578790 86400 578846 86436
rect 579342 83988 579344 84008
rect 579344 83988 579396 84008
rect 579396 83988 579398 84008
rect 579342 83952 579398 83988
rect 578698 82184 578754 82240
rect 578606 77832 578662 77888
rect 579526 80008 579582 80064
rect 593970 222264 594026 222320
rect 582378 219952 582434 220008
rect 582562 219988 582564 220008
rect 582564 219988 582616 220008
rect 582616 219988 582618 220008
rect 582562 219952 582618 219988
rect 582378 219680 582434 219736
rect 582378 216688 582434 216744
rect 582562 216724 582564 216744
rect 582564 216724 582616 216744
rect 582616 216724 582618 216744
rect 582562 216688 582618 216724
rect 583114 219408 583170 219464
rect 591762 217232 591818 217288
rect 591946 217252 592002 217288
rect 591946 217232 591948 217252
rect 591948 217232 592000 217252
rect 592000 217232 592002 217252
rect 591578 216960 591634 217016
rect 591946 216960 592002 217016
rect 591762 216416 591818 216472
rect 582930 216144 582986 216200
rect 594798 219680 594854 219736
rect 595902 218884 595958 218920
rect 595902 218864 595904 218884
rect 595904 218864 595956 218884
rect 595956 218864 595958 218884
rect 596086 218864 596142 218920
rect 596270 216552 596326 216608
rect 597558 217096 597614 217152
rect 597926 216280 597982 216336
rect 606758 224440 606814 224496
rect 617154 224168 617210 224224
rect 606758 223896 606814 223952
rect 611634 223624 611690 223680
rect 600686 221992 600742 222048
rect 599030 221720 599086 221776
rect 599214 220904 599270 220960
rect 601974 221448 602030 221504
rect 600870 221176 600926 221232
rect 604642 220224 604698 220280
rect 605102 218592 605158 218648
rect 608966 217776 609022 217832
rect 610070 217504 610126 217560
rect 612830 213152 612886 213208
rect 615682 220224 615738 220280
rect 617706 220496 617762 220552
rect 618810 219408 618866 219464
rect 623778 219136 623834 219192
rect 622950 218592 623006 218648
rect 630954 223896 631010 223952
rect 630678 218864 630734 218920
rect 629390 218048 629446 218104
rect 627826 216824 627882 216880
rect 639602 230016 639658 230072
rect 650642 225528 650698 225584
rect 649722 221448 649778 221504
rect 644754 220360 644810 220416
rect 643834 218864 643890 218920
rect 640614 218592 640670 218648
rect 639970 217776 640026 217832
rect 643006 215872 643062 215928
rect 644570 217504 644626 217560
rect 648618 219816 648674 219872
rect 646594 216144 646650 216200
rect 647146 213152 647202 213208
rect 651286 219136 651342 219192
rect 652206 298424 652262 298480
rect 668398 876288 668454 876344
rect 666466 755112 666522 755168
rect 666466 745456 666522 745512
rect 666282 711592 666338 711648
rect 666282 688608 666338 688664
rect 665822 626048 665878 626104
rect 667846 780680 667902 780736
rect 667662 742464 667718 742520
rect 667202 671064 667258 671120
rect 669042 872480 669098 872536
rect 668398 754160 668454 754216
rect 668398 735256 668454 735312
rect 668214 731448 668270 731504
rect 667846 710232 667902 710288
rect 667846 705064 667902 705120
rect 667662 665896 667718 665952
rect 666466 665352 666522 665408
rect 666282 621152 666338 621208
rect 667018 593408 667074 593464
rect 664442 580080 664498 580136
rect 663062 535472 663118 535528
rect 661682 491544 661738 491600
rect 660302 411848 660358 411904
rect 659106 360032 659162 360088
rect 661866 406272 661922 406328
rect 661682 313520 661738 313576
rect 660302 234096 660358 234152
rect 658922 233824 658978 233880
rect 664442 494672 664498 494728
rect 667662 603336 667718 603392
rect 667386 564440 667442 564496
rect 667202 535200 667258 535256
rect 667018 528536 667074 528592
rect 665822 492088 665878 492144
rect 667662 529896 667718 529952
rect 667386 485152 667442 485208
rect 663246 358536 663302 358592
rect 668030 693232 668086 693288
rect 669042 755384 669098 755440
rect 668858 738248 668914 738304
rect 669042 733760 669098 733816
rect 668766 730496 668822 730552
rect 668214 664128 668270 664184
rect 668582 669296 668638 669352
rect 668766 666168 668822 666224
rect 670606 928240 670662 928296
rect 669778 864184 669834 864240
rect 669778 750896 669834 750952
rect 669594 737024 669650 737080
rect 669226 728184 669282 728240
rect 668950 661680 669006 661736
rect 669778 730088 669834 730144
rect 669594 661952 669650 662008
rect 669134 661272 669190 661328
rect 670422 780000 670478 780056
rect 670330 779456 670386 779512
rect 670146 775648 670202 775704
rect 669962 715672 670018 715728
rect 670146 709960 670202 710016
rect 670330 707920 670386 707976
rect 670790 865272 670846 865328
rect 671986 935720 672042 935776
rect 671158 774968 671214 775024
rect 670974 758648 671030 758704
rect 670974 758240 671030 758296
rect 670790 754840 670846 754896
rect 670790 728592 670846 728648
rect 670790 714856 670846 714912
rect 670514 707104 670570 707160
rect 669778 659640 669834 659696
rect 669226 654200 669282 654256
rect 669042 645496 669098 645552
rect 668398 643864 668454 643920
rect 668030 619928 668086 619984
rect 668398 601704 668454 601760
rect 668858 638696 668914 638752
rect 669042 574776 669098 574832
rect 668858 574368 668914 574424
rect 669778 643456 669834 643512
rect 669594 623872 669650 623928
rect 669594 578992 669650 579048
rect 669594 577768 669650 577824
rect 669226 574096 669282 574152
rect 669042 557504 669098 557560
rect 668582 535880 668638 535936
rect 668398 527312 668454 527368
rect 669226 552608 669282 552664
rect 669042 485832 669098 485888
rect 669226 483928 669282 483984
rect 667846 456184 667902 456240
rect 667202 360848 667258 360904
rect 665822 315424 665878 315480
rect 664442 271088 664498 271144
rect 663062 268096 663118 268152
rect 663798 231784 663854 231840
rect 662050 231104 662106 231160
rect 660946 229744 661002 229800
rect 653402 229064 653458 229120
rect 652390 222808 652446 222864
rect 652942 221176 652998 221232
rect 653126 220632 653182 220688
rect 654782 226616 654838 226672
rect 658922 226344 658978 226400
rect 656714 224984 656770 225040
rect 656162 224440 656218 224496
rect 658186 223896 658242 223952
rect 656898 223624 656954 223680
rect 657542 223080 657598 223136
rect 656530 216960 656586 217016
rect 659382 214512 659438 214568
rect 660210 223352 660266 223408
rect 663062 230560 663118 230616
rect 664442 230832 664498 230888
rect 664810 213424 664866 213480
rect 665270 230288 665326 230344
rect 665822 225392 665878 225448
rect 665454 220904 665510 220960
rect 666282 215056 666338 215112
rect 589462 207984 589518 208040
rect 589462 206352 589518 206408
rect 589646 204720 589702 204776
rect 589462 203088 589518 203144
rect 589462 201456 589518 201512
rect 589462 199824 589518 199880
rect 590382 198192 590438 198248
rect 589462 196560 589518 196616
rect 589278 194928 589334 194984
rect 589462 193296 589518 193352
rect 589462 191664 589518 191720
rect 590566 190032 590622 190088
rect 589646 188400 589702 188456
rect 589462 186768 589518 186824
rect 589462 185136 589518 185192
rect 589462 183504 589518 183560
rect 590566 181872 590622 181928
rect 589646 180240 589702 180296
rect 589462 178608 589518 178664
rect 667018 218048 667074 218104
rect 667018 213152 667074 213208
rect 666650 178744 666706 178800
rect 666834 178472 666890 178528
rect 589646 176976 589702 177032
rect 589462 175364 589518 175400
rect 589462 175344 589464 175364
rect 589464 175344 589516 175364
rect 589516 175344 589518 175364
rect 589462 173712 589518 173768
rect 589462 172080 589518 172136
rect 589186 170448 589242 170504
rect 589830 168816 589886 168872
rect 589462 167184 589518 167240
rect 589646 165552 589702 165608
rect 589462 163920 589518 163976
rect 590566 162288 590622 162344
rect 589462 160656 589518 160712
rect 588542 159024 588598 159080
rect 589278 157412 589334 157448
rect 589278 157392 589280 157412
rect 589280 157392 589332 157412
rect 589332 157392 589334 157412
rect 589462 155760 589518 155816
rect 589462 154128 589518 154184
rect 589462 152496 589518 152552
rect 589922 150864 589978 150920
rect 589186 149232 589242 149288
rect 588726 145968 588782 146024
rect 578882 75656 578938 75712
rect 578514 61784 578570 61840
rect 579526 73108 579528 73128
rect 579528 73108 579580 73128
rect 579580 73108 579582 73128
rect 579526 73072 579582 73108
rect 579250 71168 579306 71224
rect 579526 66292 579582 66328
rect 579526 66272 579528 66292
rect 579528 66272 579580 66292
rect 579580 66272 579582 66292
rect 579066 64776 579122 64832
rect 579526 60288 579582 60344
rect 579526 57876 579528 57896
rect 579528 57876 579580 57896
rect 579580 57876 579582 57896
rect 579526 57840 579582 57876
rect 579526 56072 579582 56128
rect 588542 137808 588598 137864
rect 589462 147600 589518 147656
rect 589462 144336 589518 144392
rect 589646 142704 589702 142760
rect 589462 141072 589518 141128
rect 589462 139460 589518 139496
rect 589462 139440 589464 139460
rect 589464 139440 589516 139460
rect 589516 139440 589518 139460
rect 589462 136176 589518 136232
rect 590290 134544 590346 134600
rect 589922 132912 589978 132968
rect 589278 129648 589334 129704
rect 589462 128016 589518 128072
rect 589462 126384 589518 126440
rect 589738 124752 589794 124808
rect 589462 123120 589518 123176
rect 589278 121508 589334 121544
rect 589278 121488 589280 121508
rect 589280 121488 589332 121508
rect 589332 121488 589334 121508
rect 588726 119856 588782 119912
rect 589462 118224 589518 118280
rect 589462 116592 589518 116648
rect 589554 114960 589610 115016
rect 670422 684936 670478 684992
rect 670238 668208 670294 668264
rect 670974 713632 671030 713688
rect 671802 869216 671858 869272
rect 671342 763680 671398 763736
rect 671434 759872 671490 759928
rect 671618 759056 671674 759112
rect 671342 757424 671398 757480
rect 671434 715264 671490 715320
rect 675390 966456 675446 966512
rect 672998 966320 673054 966376
rect 675114 966320 675170 966376
rect 672722 947280 672778 947336
rect 672722 938032 672778 938088
rect 672538 933136 672594 933192
rect 672354 787344 672410 787400
rect 674378 962784 674434 962840
rect 673182 960744 673238 960800
rect 672998 932864 673054 932920
rect 674102 959248 674158 959304
rect 673366 937352 673422 937408
rect 673182 930688 673238 930744
rect 673182 872208 673238 872264
rect 672630 783808 672686 783864
rect 671986 757832 672042 757888
rect 671986 751712 672042 751768
rect 672354 750080 672410 750136
rect 671986 743416 672042 743472
rect 671802 735528 671858 735584
rect 671618 714448 671674 714504
rect 671710 714040 671766 714096
rect 671526 713224 671582 713280
rect 671342 712816 671398 712872
rect 671158 705472 671214 705528
rect 670974 689016 671030 689072
rect 670790 669840 670846 669896
rect 670606 666576 670662 666632
rect 670146 624280 670202 624336
rect 670790 647808 670846 647864
rect 670606 624688 670662 624744
rect 670422 622512 670478 622568
rect 670146 615712 670202 615768
rect 670606 614896 670662 614952
rect 669962 581032 670018 581088
rect 670146 580760 670202 580816
rect 670238 579400 670294 579456
rect 669962 578584 670018 578640
rect 669778 570288 669834 570344
rect 669778 569472 669834 569528
rect 669594 533024 669650 533080
rect 670422 553424 670478 553480
rect 670238 534928 670294 534984
rect 669962 534656 670018 534712
rect 670422 482296 670478 482352
rect 671250 670248 671306 670304
rect 672170 728184 672226 728240
rect 672170 712408 672226 712464
rect 672998 784216 673054 784272
rect 672814 759464 672870 759520
rect 672814 756200 672870 756256
rect 672814 755112 672870 755168
rect 672814 734032 672870 734088
rect 672538 710776 672594 710832
rect 672538 709416 672594 709472
rect 672538 698264 672594 698320
rect 672354 696904 672410 696960
rect 671802 680040 671858 680096
rect 671618 669432 671674 669488
rect 671434 668480 671490 668536
rect 671526 667936 671582 667992
rect 671250 625096 671306 625152
rect 671526 623464 671582 623520
rect 671158 622784 671214 622840
rect 670974 616528 671030 616584
rect 671618 622240 671674 622296
rect 671342 594768 671398 594824
rect 671158 578176 671214 578232
rect 670790 571920 670846 571976
rect 670790 570696 670846 570752
rect 671158 548392 671214 548448
rect 670974 532752 671030 532808
rect 670790 500928 670846 500984
rect 670974 489232 671030 489288
rect 672170 667392 672226 667448
rect 671986 664400 672042 664456
rect 671986 661000 672042 661056
rect 671802 620336 671858 620392
rect 671618 577360 671674 577416
rect 671802 576952 671858 577008
rect 671802 534248 671858 534304
rect 671618 531800 671674 531856
rect 671618 531392 671674 531448
rect 671342 524864 671398 524920
rect 671434 490456 671490 490512
rect 671158 485560 671214 485616
rect 670606 455368 670662 455424
rect 669778 455096 669834 455152
rect 669410 403688 669466 403744
rect 668582 311888 668638 311944
rect 667202 181328 667258 181384
rect 669226 302232 669282 302288
rect 667386 142704 667442 142760
rect 667938 231140 667940 231160
rect 667940 231140 667992 231160
rect 667992 231140 667994 231160
rect 667938 231104 667994 231140
rect 668490 234504 668546 234560
rect 668306 231512 668362 231568
rect 668306 230560 668362 230616
rect 667938 223080 667994 223136
rect 667938 221212 667940 221232
rect 667940 221212 667992 221232
rect 667992 221212 667994 221232
rect 667938 221176 667994 221212
rect 667846 219408 667902 219464
rect 668122 192616 668178 192672
rect 668030 187584 668086 187640
rect 667938 184492 667940 184512
rect 667940 184492 667992 184512
rect 667992 184492 667994 184512
rect 667938 184456 667994 184492
rect 668306 182824 668362 182880
rect 667754 174936 667810 174992
rect 667938 174664 667994 174720
rect 668030 169668 668032 169688
rect 668032 169668 668084 169688
rect 668084 169668 668086 169688
rect 668030 169632 668086 169668
rect 667938 164872 667994 164928
rect 667938 160012 667940 160032
rect 667940 160012 667992 160032
rect 667992 160012 667994 160032
rect 667938 159976 667994 160012
rect 668306 150220 668308 150240
rect 668308 150220 668360 150240
rect 668360 150220 668362 150240
rect 668306 150184 668362 150220
rect 668950 231784 669006 231840
rect 668950 231240 669006 231296
rect 669042 224304 669098 224360
rect 669042 221856 669098 221912
rect 671802 490864 671858 490920
rect 671802 489640 671858 489696
rect 671618 488416 671674 488472
rect 671434 402464 671490 402520
rect 672170 648624 672226 648680
rect 674746 958296 674802 958352
rect 674562 957072 674618 957128
rect 675298 964688 675354 964744
rect 675758 963328 675814 963384
rect 675482 962784 675538 962840
rect 675114 960744 675170 960800
rect 675114 959248 675170 959304
rect 675390 958296 675446 958352
rect 675206 957752 675262 957808
rect 675758 957752 675814 957808
rect 674102 933816 674158 933872
rect 674286 932592 674342 932648
rect 674838 953400 674894 953456
rect 674654 930416 674710 930472
rect 674470 930144 674526 930200
rect 675390 957072 675446 957128
rect 675758 956392 675814 956448
rect 675390 953400 675446 953456
rect 675390 952176 675446 952232
rect 675390 951496 675446 951552
rect 683302 950680 683358 950736
rect 679622 949456 679678 949512
rect 675206 937896 675262 937952
rect 675206 936944 675262 937000
rect 675390 935448 675446 935504
rect 676218 941704 676274 941760
rect 676218 939256 676274 939312
rect 675574 934632 675630 934688
rect 683118 947280 683174 947336
rect 683118 939664 683174 939720
rect 682382 935176 682438 935232
rect 679622 934360 679678 934416
rect 683302 932320 683358 932376
rect 683118 929056 683174 929112
rect 675298 879144 675354 879200
rect 675758 876560 675814 876616
rect 675114 876288 675170 876344
rect 675758 875880 675814 875936
rect 675390 873976 675446 874032
rect 675114 873160 675170 873216
rect 675114 872480 675170 872536
rect 675390 872208 675446 872264
rect 674562 868400 674618 868456
rect 674102 867176 674158 867232
rect 673734 864864 673790 864920
rect 673550 777416 673606 777472
rect 673366 760280 673422 760336
rect 673182 752528 673238 752584
rect 673182 751304 673238 751360
rect 673366 739880 673422 739936
rect 672998 709144 673054 709200
rect 673182 697176 673238 697232
rect 672998 665660 673000 665680
rect 673000 665660 673052 665680
rect 673052 665660 673054 665680
rect 672998 665624 673054 665660
rect 672814 662496 672870 662552
rect 672722 648896 672778 648952
rect 672538 621560 672594 621616
rect 672354 620608 672410 620664
rect 672446 608640 672502 608696
rect 672446 607280 672502 607336
rect 673918 779184 673974 779240
rect 673734 771976 673790 772032
rect 673734 734304 673790 734360
rect 673550 724240 673606 724296
rect 673550 693504 673606 693560
rect 673366 663312 673422 663368
rect 673366 659912 673422 659968
rect 673182 619656 673238 619712
rect 672814 604832 672870 604888
rect 672630 575048 672686 575104
rect 672262 532480 672318 532536
rect 672630 533432 672686 533488
rect 672446 528944 672502 529000
rect 672998 604288 673054 604344
rect 674930 868672 674986 868728
rect 675114 868672 675170 868728
rect 675298 868400 675354 868456
rect 674930 866768 674986 866824
rect 675298 867176 675354 867232
rect 675298 865272 675354 865328
rect 675482 864864 675538 864920
rect 675482 864184 675538 864240
rect 674286 788024 674342 788080
rect 674562 770616 674618 770672
rect 674102 753344 674158 753400
rect 675482 788024 675538 788080
rect 675482 787344 675538 787400
rect 674930 786664 674986 786720
rect 675390 786664 675446 786720
rect 675482 784216 675538 784272
rect 675482 783808 675538 783864
rect 675482 782992 675538 783048
rect 675482 780680 675538 780736
rect 675298 780408 675354 780464
rect 675482 780000 675538 780056
rect 675482 779456 675538 779512
rect 675482 779184 675538 779240
rect 675298 778912 675354 778968
rect 675022 777144 675078 777200
rect 675482 777416 675538 777472
rect 674930 775648 674986 775704
rect 674930 774560 674986 774616
rect 675482 776192 675538 776248
rect 675298 776056 675354 776112
rect 675022 766536 675078 766592
rect 675482 774968 675538 775024
rect 675482 774560 675538 774616
rect 675390 773336 675446 773392
rect 675206 765040 675262 765096
rect 674838 757152 674894 757208
rect 683210 772248 683266 772304
rect 681002 768712 681058 768768
rect 676770 761776 676826 761832
rect 676034 757172 676090 757208
rect 676034 757152 676036 757172
rect 676036 757152 676088 757172
rect 676088 757152 676090 757172
rect 675850 755792 675906 755848
rect 681002 757016 681058 757072
rect 676770 754568 676826 754624
rect 683854 771976 683910 772032
rect 683486 770616 683542 770672
rect 683394 763680 683450 763736
rect 683394 760688 683450 760744
rect 683210 753752 683266 753808
rect 683854 756608 683910 756664
rect 683578 752936 683634 752992
rect 683394 752120 683450 752176
rect 675298 745456 675354 745512
rect 675114 743416 675170 743472
rect 674930 742464 674986 742520
rect 675114 741512 675170 741568
rect 675298 739880 675354 739936
rect 675482 739336 675538 739392
rect 675206 738316 675262 738372
rect 675114 737024 675170 737080
rect 675390 735528 675446 735584
rect 674838 735256 674894 735312
rect 675114 734304 675170 734360
rect 674930 734032 674986 734088
rect 675114 733760 675170 733816
rect 675114 731448 675170 731504
rect 674378 728612 674434 728648
rect 674378 728592 674380 728612
rect 674380 728592 674432 728612
rect 674432 728592 674434 728612
rect 673918 726824 673974 726880
rect 675114 730496 675170 730552
rect 675114 730088 675170 730144
rect 683394 726824 683450 726880
rect 674746 726552 674802 726608
rect 681002 725736 681058 725792
rect 677322 724260 677378 724296
rect 677322 724240 677324 724260
rect 677324 724240 677376 724260
rect 677376 724240 677378 724260
rect 676034 710776 676090 710832
rect 681002 710776 681058 710832
rect 676034 709552 676090 709608
rect 675850 709416 675906 709472
rect 675850 708736 675906 708792
rect 683210 708328 683266 708384
rect 683762 726416 683818 726472
rect 683762 711184 683818 711240
rect 683394 706696 683450 706752
rect 674470 706288 674526 706344
rect 674102 690104 674158 690160
rect 673734 682624 673790 682680
rect 674286 687248 674342 687304
rect 673826 645088 673882 645144
rect 673550 618568 673606 618624
rect 673642 604016 673698 604072
rect 673458 592320 673514 592376
rect 675114 698264 675170 698320
rect 675114 697176 675170 697232
rect 675114 696904 675170 696960
rect 675390 696768 675446 696824
rect 675666 694320 675722 694376
rect 675114 693504 675170 693560
rect 674930 693232 674986 693288
rect 675114 692960 675170 693016
rect 675390 690104 675446 690160
rect 674194 642096 674250 642152
rect 674010 641688 674066 641744
rect 673826 598304 673882 598360
rect 673182 580760 673238 580816
rect 673182 579808 673238 579864
rect 673182 573280 673238 573336
rect 673182 560088 673238 560144
rect 672998 530576 673054 530632
rect 672814 530168 672870 530224
rect 672630 490048 672686 490104
rect 673182 484744 673238 484800
rect 674286 640736 674342 640792
rect 674470 636248 674526 636304
rect 674194 635704 674250 635760
rect 674194 597352 674250 597408
rect 674010 591232 674066 591288
rect 674010 558048 674066 558104
rect 673826 557912 673882 557968
rect 673642 545808 673698 545864
rect 673642 528264 673698 528320
rect 674930 689288 674986 689344
rect 675114 689016 675170 689072
rect 674930 688608 674986 688664
rect 675298 687248 675354 687304
rect 675114 685752 675170 685808
rect 675482 684936 675538 684992
rect 683118 682624 683174 682680
rect 675298 680040 675354 680096
rect 674838 668752 674894 668808
rect 674838 668208 674894 668264
rect 674838 664672 674894 664728
rect 674838 664128 674894 664184
rect 674838 662224 674894 662280
rect 674838 661680 674894 661736
rect 676494 670248 676550 670304
rect 676770 670248 676826 670304
rect 676494 669840 676550 669896
rect 676770 669024 676826 669080
rect 676494 665760 676550 665816
rect 676494 664944 676550 665000
rect 683302 682352 683358 682408
rect 683486 680992 683542 681048
rect 683302 666984 683358 667040
rect 683486 664128 683542 664184
rect 683118 662904 683174 662960
rect 675390 660184 675446 660240
rect 675390 659640 675446 659696
rect 675390 654200 675446 654256
rect 675574 652840 675630 652896
rect 675574 651480 675630 651536
rect 675390 648896 675446 648952
rect 675114 648624 675170 648680
rect 675390 647808 675446 647864
rect 675022 645768 675078 645824
rect 675114 645496 675170 645552
rect 675114 645088 675170 645144
rect 675758 644272 675814 644328
rect 675114 643864 675170 643920
rect 675298 643456 675354 643512
rect 675298 641688 675354 641744
rect 675114 640464 675170 640520
rect 675390 639784 675446 639840
rect 675482 638696 675538 638752
rect 674838 638152 674894 638208
rect 675758 638152 675814 638208
rect 674838 637880 674894 637936
rect 674930 637608 674986 637664
rect 674930 636152 674986 636208
rect 675298 637608 675354 637664
rect 676034 637880 676090 637936
rect 675482 636112 675538 636168
rect 675298 631352 675354 631408
rect 683394 636792 683450 636848
rect 683210 635432 683266 635488
rect 676034 631352 676090 631408
rect 674654 623192 674710 623248
rect 674838 608640 674894 608696
rect 674838 607008 674894 607064
rect 674838 601704 674894 601760
rect 674838 600480 674894 600536
rect 674654 599800 674710 599856
rect 674470 589872 674526 589928
rect 674378 554376 674434 554432
rect 674194 547032 674250 547088
rect 674194 529352 674250 529408
rect 674194 528536 674250 528592
rect 674010 487192 674066 487248
rect 673826 486104 673882 486160
rect 675574 623192 675630 623248
rect 675850 622820 675852 622840
rect 675852 622820 675904 622840
rect 675904 622820 675906 622840
rect 675850 622784 675906 622820
rect 676402 622784 676458 622840
rect 676678 622820 676680 622840
rect 676680 622820 676732 622840
rect 676732 622820 676734 622840
rect 676678 622784 676734 622820
rect 676034 622512 676090 622568
rect 683118 628496 683174 628552
rect 683118 625640 683174 625696
rect 682382 621968 682438 622024
rect 676494 621560 676550 621616
rect 676494 621152 676550 621208
rect 676494 620336 676550 620392
rect 676494 619928 676550 619984
rect 683302 618296 683358 618352
rect 675574 617752 675630 617808
rect 683486 617072 683542 617128
rect 675482 607824 675538 607880
rect 675298 607280 675354 607336
rect 675298 607008 675354 607064
rect 675298 604832 675354 604888
rect 675298 604288 675354 604344
rect 675390 604016 675446 604072
rect 675298 603336 675354 603392
rect 675482 602928 675538 602984
rect 675298 600480 675354 600536
rect 675482 599800 675538 599856
rect 674838 592592 674894 592648
rect 675298 599256 675354 599312
rect 675482 598440 675538 598496
rect 675482 597352 675538 597408
rect 675390 595312 675446 595368
rect 675482 594768 675538 594824
rect 675390 593408 675446 593464
rect 675574 593136 675630 593192
rect 675298 592048 675354 592104
rect 675114 575456 675170 575512
rect 676034 592864 676090 592920
rect 675850 592592 675906 592648
rect 675574 586200 675630 586256
rect 683394 592592 683450 592648
rect 681002 591640 681058 591696
rect 676034 576544 676090 576600
rect 681002 576000 681058 576056
rect 676034 575048 676090 575104
rect 676034 573688 676090 573744
rect 674838 571104 674894 571160
rect 674838 570288 674894 570344
rect 674838 559544 674894 559600
rect 675022 557504 675078 557560
rect 675022 555736 675078 555792
rect 683670 591232 683726 591288
rect 683854 589872 683910 589928
rect 683854 576408 683910 576464
rect 683670 573144 683726 573200
rect 683394 571920 683450 571976
rect 682382 570696 682438 570752
rect 675390 564440 675446 564496
rect 675482 562672 675538 562728
rect 675482 561176 675538 561232
rect 675390 560088 675446 560144
rect 675482 559544 675538 559600
rect 675390 558048 675446 558104
rect 675390 557776 675446 557832
rect 675482 557504 675538 557560
rect 675482 555736 675538 555792
rect 675390 554376 675446 554432
rect 675206 553968 675262 554024
rect 675390 553424 675446 553480
rect 675482 552608 675538 552664
rect 675758 550296 675814 550352
rect 675114 550160 675170 550216
rect 675482 548392 675538 548448
rect 674838 546352 674894 546408
rect 675850 547576 675906 547632
rect 678242 547576 678298 547632
rect 675666 546352 675722 546408
rect 674838 545536 674894 545592
rect 674654 526904 674710 526960
rect 674838 502560 674894 502616
rect 675298 546080 675354 546136
rect 674930 502152 674986 502208
rect 675114 487600 675170 487656
rect 675758 534656 675814 534712
rect 675758 534044 675814 534100
rect 675758 532480 675814 532536
rect 675758 531596 675814 531652
rect 683578 547304 683634 547360
rect 683302 545672 683358 545728
rect 681002 531392 681058 531448
rect 678242 530984 678298 531040
rect 676034 530576 676090 530632
rect 676034 528740 676090 528796
rect 683854 547032 683910 547088
rect 683854 528128 683910 528184
rect 683578 527312 683634 527368
rect 683302 526496 683358 526552
rect 683118 525680 683174 525736
rect 677874 524456 677930 524512
rect 675298 486376 675354 486432
rect 674378 483520 674434 483576
rect 672906 456456 672962 456512
rect 671986 455640 672042 455696
rect 672078 455116 672134 455152
rect 672078 455096 672080 455116
rect 672080 455096 672132 455116
rect 672132 455096 672134 455116
rect 673946 456204 674002 456240
rect 673946 456184 673948 456204
rect 673948 456184 674000 456204
rect 674000 456184 674002 456204
rect 673826 455948 673828 455968
rect 673828 455948 673880 455968
rect 673880 455948 673882 455968
rect 673826 455912 673882 455948
rect 673596 455660 673652 455696
rect 673596 455640 673598 455660
rect 673598 455640 673650 455660
rect 673650 455640 673652 455660
rect 673274 455388 673330 455424
rect 673274 455368 673276 455388
rect 673276 455368 673328 455388
rect 673328 455368 673330 455388
rect 673386 455252 673442 455288
rect 673386 455232 673388 455252
rect 673388 455232 673440 455252
rect 673440 455232 673442 455252
rect 676034 502560 676090 502616
rect 675850 502152 675906 502208
rect 676402 500928 676458 500984
rect 683118 503648 683174 503704
rect 676034 488008 676090 488064
rect 675850 487192 675906 487248
rect 675666 486104 675722 486160
rect 675850 484336 675906 484392
rect 675666 483112 675722 483168
rect 675666 481888 675722 481944
rect 673044 454844 673100 454880
rect 673044 454824 673046 454844
rect 673046 454824 673098 454844
rect 673098 454824 673100 454844
rect 675482 454824 675538 454880
rect 673162 454588 673164 454608
rect 673164 454588 673216 454608
rect 673216 454588 673218 454608
rect 673162 454552 673218 454588
rect 672814 454180 672816 454200
rect 672816 454180 672868 454200
rect 672868 454180 672870 454200
rect 672814 454144 672870 454180
rect 672722 453908 672724 453928
rect 672724 453908 672776 453928
rect 672776 453908 672778 453928
rect 672722 453872 672778 453908
rect 675206 453872 675262 453928
rect 675850 480664 675906 480720
rect 675850 454144 675906 454200
rect 676218 475360 676274 475416
rect 676218 455912 676274 455968
rect 677506 492768 677562 492824
rect 678242 486784 678298 486840
rect 683302 494672 683358 494728
rect 683302 491272 683358 491328
rect 683118 487192 683174 487248
rect 683302 482704 683358 482760
rect 683118 481516 683120 481536
rect 683120 481516 683172 481536
rect 683172 481516 683174 481536
rect 683118 481480 683174 481516
rect 676954 456456 677010 456512
rect 676770 454552 676826 454608
rect 676034 453736 676090 453792
rect 683302 411848 683358 411904
rect 676034 410488 676090 410544
rect 674194 402192 674250 402248
rect 671802 401648 671858 401704
rect 672814 400424 672870 400480
rect 672630 393896 672686 393952
rect 671986 393488 672042 393544
rect 671802 347656 671858 347712
rect 670606 347248 670662 347304
rect 669962 275304 670018 275360
rect 670422 261568 670478 261624
rect 670238 260344 670294 260400
rect 670422 247016 670478 247072
rect 670238 240216 670294 240272
rect 669962 237088 670018 237144
rect 669410 234912 669466 234968
rect 669226 206488 669282 206544
rect 669318 188400 669374 188456
rect 669410 177248 669466 177304
rect 669778 168272 669834 168328
rect 669226 168136 669282 168192
rect 669134 164192 669190 164248
rect 668950 163240 669006 163296
rect 668766 153448 668822 153504
rect 668766 153040 668822 153096
rect 668490 148552 668546 148608
rect 667938 137808 667994 137864
rect 667570 135904 667626 135960
rect 667938 135496 667994 135552
rect 667018 133048 667074 133104
rect 590106 131280 590162 131336
rect 669134 143656 669190 143712
rect 669226 141072 669282 141128
rect 669226 138760 669282 138816
rect 668950 128288 669006 128344
rect 668766 125704 668822 125760
rect 669226 122168 669282 122224
rect 668950 120808 669006 120864
rect 667938 119176 667994 119232
rect 667938 117544 667994 117600
rect 670238 236816 670294 236872
rect 671802 325624 671858 325680
rect 671710 261160 671766 261216
rect 671526 260888 671582 260944
rect 671342 256672 671398 256728
rect 671526 246608 671582 246664
rect 671710 245248 671766 245304
rect 670146 232736 670202 232792
rect 671342 237768 671398 237824
rect 671066 234504 671122 234560
rect 670606 232464 670662 232520
rect 670698 226208 670754 226264
rect 670698 225428 670700 225448
rect 670700 225428 670752 225448
rect 670752 225428 670754 225448
rect 670698 225392 670754 225428
rect 670698 225020 670700 225040
rect 670700 225020 670752 225040
rect 670752 225020 670754 225040
rect 670698 224984 670754 225020
rect 671158 225664 671214 225720
rect 671158 225392 671214 225448
rect 670514 223660 670516 223680
rect 670516 223660 670568 223680
rect 670568 223660 670570 223680
rect 670514 223624 670570 223660
rect 670882 224612 670884 224632
rect 670884 224612 670936 224632
rect 670936 224612 670938 224632
rect 670882 224576 670938 224612
rect 670928 223896 670984 223952
rect 670790 221992 670846 222048
rect 670606 220904 670662 220960
rect 670606 220632 670662 220688
rect 670790 220088 670846 220144
rect 670606 176432 670662 176488
rect 670974 199144 671030 199200
rect 671158 194248 671214 194304
rect 670790 175616 670846 175672
rect 670606 171944 670662 172000
rect 670422 169496 670478 169552
rect 670146 165008 670202 165064
rect 669962 121352 670018 121408
rect 669226 114280 669282 114336
rect 590290 113328 590346 113384
rect 589370 111696 589426 111752
rect 670422 154808 670478 154864
rect 671710 234504 671766 234560
rect 671710 229336 671766 229392
rect 671802 227024 671858 227080
rect 671618 226888 671674 226944
rect 671802 226636 671858 226672
rect 671802 226616 671804 226636
rect 671804 226616 671856 226636
rect 671856 226616 671858 226636
rect 671802 226092 671858 226128
rect 671802 226072 671804 226092
rect 671804 226072 671856 226092
rect 671856 226072 671858 226092
rect 671818 225700 671820 225720
rect 671820 225700 671872 225720
rect 671872 225700 671874 225720
rect 671818 225664 671874 225700
rect 671802 225120 671858 225176
rect 671710 224848 671766 224904
rect 672354 392264 672410 392320
rect 672170 357040 672226 357096
rect 672170 312432 672226 312488
rect 672630 376216 672686 376272
rect 672630 356224 672686 356280
rect 673182 399608 673238 399664
rect 672998 397160 673054 397216
rect 672998 377984 673054 378040
rect 673366 396344 673422 396400
rect 673826 396072 673882 396128
rect 673366 382200 673422 382256
rect 674010 395664 674066 395720
rect 673826 381384 673882 381440
rect 674010 375400 674066 375456
rect 672814 355816 672870 355872
rect 673182 355408 673238 355464
rect 672814 351328 672870 351384
rect 672998 348880 673054 348936
rect 672814 337184 672870 337240
rect 672998 331472 673054 331528
rect 674654 401376 674710 401432
rect 674470 394440 674526 394496
rect 674470 377712 674526 377768
rect 674194 357448 674250 357504
rect 683118 406272 683174 406328
rect 683302 403688 683358 403744
rect 683118 403280 683174 403336
rect 676034 400152 676090 400208
rect 676034 399336 676090 399392
rect 676218 398384 676274 398440
rect 676402 397976 676458 398032
rect 681002 397568 681058 397624
rect 683026 392672 683082 392728
rect 683026 389000 683082 389056
rect 681002 387640 681058 387696
rect 675758 384920 675814 384976
rect 675390 382200 675446 382256
rect 675114 381384 675170 381440
rect 675758 380568 675814 380624
rect 675758 378664 675814 378720
rect 675114 377712 675170 377768
rect 675758 377304 675814 377360
rect 675206 376896 675262 376952
rect 675390 376216 675446 376272
rect 675390 375400 675446 375456
rect 675666 372952 675722 373008
rect 675114 372544 675170 372600
rect 675850 360848 675906 360904
rect 676034 360032 676090 360088
rect 676034 358264 676090 358320
rect 675850 357856 675906 357912
rect 674654 356632 674710 356688
rect 673366 355000 673422 355056
rect 674654 354592 674710 354648
rect 673366 353368 673422 353424
rect 674470 352552 674526 352608
rect 674286 352144 674342 352200
rect 673734 350512 673790 350568
rect 673550 349424 673606 349480
rect 673366 340720 673422 340776
rect 673550 332696 673606 332752
rect 674102 349696 674158 349752
rect 673918 348472 673974 348528
rect 673734 331064 673790 331120
rect 672814 312704 672870 312760
rect 672630 311616 672686 311672
rect 672630 304272 672686 304328
rect 672630 287816 672686 287872
rect 673090 311208 673146 311264
rect 673274 310800 673330 310856
rect 673734 305496 673790 305552
rect 673550 304680 673606 304736
rect 673274 303456 673330 303512
rect 673090 267552 673146 267608
rect 672814 266872 672870 266928
rect 672814 266464 672870 266520
rect 672630 257896 672686 257952
rect 672630 257080 672686 257136
rect 672538 242800 672594 242856
rect 673090 266056 673146 266112
rect 673550 290536 673606 290592
rect 673734 285504 673790 285560
rect 673642 259664 673698 259720
rect 673642 258440 673698 258496
rect 673458 245792 673514 245848
rect 673526 237088 673582 237144
rect 673412 236852 673414 236872
rect 673414 236852 673466 236872
rect 673466 236852 673468 236872
rect 673412 236816 673468 236852
rect 673458 236272 673514 236328
rect 673366 232464 673422 232520
rect 672906 231784 672962 231840
rect 672262 228520 672318 228576
rect 672262 227044 672318 227080
rect 672262 227024 672264 227044
rect 672264 227024 672316 227044
rect 672316 227024 672318 227044
rect 672262 226480 672318 226536
rect 672170 225936 672226 225992
rect 672170 224576 672226 224632
rect 672170 216960 672226 217016
rect 672170 211384 672226 211440
rect 671986 211112 672042 211168
rect 672262 210160 672318 210216
rect 672078 209344 672134 209400
rect 672262 200776 672318 200832
rect 672170 197512 672226 197568
rect 671986 192344 672042 192400
rect 671710 189352 671766 189408
rect 673750 236000 673806 236056
rect 674286 336640 674342 336696
rect 674102 335824 674158 335880
rect 674470 333920 674526 333976
rect 676034 352960 676090 353016
rect 675942 349152 675998 349208
rect 675114 340720 675170 340776
rect 675758 340176 675814 340232
rect 675666 339360 675722 339416
rect 675574 337728 675630 337784
rect 675114 337184 675170 337240
rect 675482 335824 675538 335880
rect 675298 335280 675354 335336
rect 675114 333920 675170 333976
rect 675114 332696 675170 332752
rect 675758 332288 675814 332344
rect 675114 331472 675170 331528
rect 675114 331064 675170 331120
rect 675758 328344 675814 328400
rect 675390 326848 675446 326904
rect 675114 325624 675170 325680
rect 676034 315424 676090 315480
rect 676034 313248 676090 313304
rect 674654 312976 674710 313032
rect 674838 312704 674894 312760
rect 674838 312024 674894 312080
rect 674654 311888 674710 311944
rect 674654 310392 674710 310448
rect 674470 309984 674526 310040
rect 674194 309576 674250 309632
rect 674378 303864 674434 303920
rect 675114 309168 675170 309224
rect 676034 308352 676090 308408
rect 675390 307944 675446 308000
rect 674838 297064 674894 297120
rect 674378 286592 674434 286648
rect 681002 307536 681058 307592
rect 678242 307128 678298 307184
rect 675390 296656 675446 296712
rect 675942 297608 675998 297664
rect 678978 306312 679034 306368
rect 678242 297336 678298 297392
rect 676218 297084 676274 297120
rect 683026 302640 683082 302696
rect 683026 299376 683082 299432
rect 676218 297064 676220 297084
rect 676220 297064 676272 297084
rect 676272 297064 676274 297084
rect 675758 296248 675814 296304
rect 675758 295840 675814 295896
rect 675758 295160 675814 295216
rect 675390 292848 675446 292904
rect 675574 292032 675630 292088
rect 675758 291488 675814 291544
rect 675114 290536 675170 290592
rect 675114 287816 675170 287872
rect 675758 287000 675814 287056
rect 675390 286592 675446 286648
rect 675114 285504 675170 285560
rect 675758 283600 675814 283656
rect 675666 282784 675722 282840
rect 675666 281152 675722 281208
rect 683302 275304 683358 275360
rect 683118 271088 683174 271144
rect 683302 268504 683358 268560
rect 683118 268096 683174 268152
rect 675022 267552 675078 267608
rect 675022 266600 675078 266656
rect 674562 265784 674618 265840
rect 674562 265376 674618 265432
rect 674194 264968 674250 265024
rect 674378 264560 674434 264616
rect 674102 258848 674158 258904
rect 674102 241440 674158 241496
rect 673642 231784 673698 231840
rect 673458 230016 673514 230072
rect 673826 230016 673882 230072
rect 673274 229472 673330 229528
rect 675022 264152 675078 264208
rect 674838 261976 674894 262032
rect 674838 261160 674894 261216
rect 678242 263200 678298 263256
rect 676402 262792 676458 262848
rect 676218 262384 676274 262440
rect 676218 261160 676274 261216
rect 675666 259120 675722 259176
rect 675666 258168 675722 258224
rect 675298 257488 675354 257544
rect 675298 256672 675354 256728
rect 674838 249328 674894 249384
rect 675022 249328 675078 249384
rect 675022 248376 675078 248432
rect 675758 250280 675814 250336
rect 675390 249328 675446 249384
rect 675298 247016 675354 247072
rect 675298 246608 675354 246664
rect 675298 245792 675354 245848
rect 675022 245520 675078 245576
rect 674746 245248 674802 245304
rect 674930 245248 674986 245304
rect 674534 234948 674536 234968
rect 674536 234948 674588 234968
rect 674588 234948 674590 234968
rect 674534 234912 674590 234948
rect 675114 242800 675170 242856
rect 675114 241440 675170 241496
rect 675114 240216 675170 240272
rect 675390 238584 675446 238640
rect 675390 237768 675446 237824
rect 674746 234368 674802 234424
rect 675850 234388 675906 234424
rect 675850 234368 675852 234388
rect 675852 234368 675904 234388
rect 675904 234368 675906 234388
rect 674562 233416 674618 233472
rect 675850 233452 675852 233472
rect 675852 233452 675904 233472
rect 675904 233452 675906 233472
rect 675850 233416 675906 233452
rect 674470 231784 674526 231840
rect 675178 231512 675234 231568
rect 675068 231240 675124 231296
rect 675022 230968 675078 231024
rect 676034 230968 676090 231024
rect 674730 230868 674732 230888
rect 674732 230868 674784 230888
rect 674784 230868 674786 230888
rect 674730 230832 674786 230868
rect 674394 230308 674450 230344
rect 674394 230288 674396 230308
rect 674396 230288 674448 230308
rect 674448 230288 674450 230308
rect 674654 230288 674710 230344
rect 673458 229064 673514 229120
rect 673366 228828 673368 228848
rect 673368 228828 673420 228848
rect 673420 228828 673422 228848
rect 673366 228792 673422 228828
rect 673386 228540 673442 228576
rect 673386 228520 673388 228540
rect 673388 228520 673440 228540
rect 673440 228520 673442 228540
rect 672998 227024 673054 227080
rect 673162 226752 673218 226808
rect 673182 223896 673238 223952
rect 673366 221448 673422 221504
rect 673734 227024 673790 227080
rect 673734 226208 673790 226264
rect 673734 225664 673790 225720
rect 673734 225392 673790 225448
rect 673918 222808 673974 222864
rect 673734 221992 673790 222048
rect 673550 221176 673606 221232
rect 673458 220360 673514 220416
rect 673458 219816 673514 219872
rect 673182 219136 673238 219192
rect 672998 216144 673054 216200
rect 673366 215736 673422 215792
rect 672538 188400 672594 188456
rect 672078 183504 672134 183560
rect 671894 169904 671950 169960
rect 671710 166912 671766 166968
rect 671526 158344 671582 158400
rect 670606 148960 670662 149016
rect 671342 131688 671398 131744
rect 671526 130872 671582 130928
rect 667938 111016 667994 111072
rect 668582 111016 668638 111072
rect 590106 110064 590162 110120
rect 589462 108432 589518 108488
rect 589462 106800 589518 106856
rect 589830 105168 589886 105224
rect 589922 101904 589978 101960
rect 667938 109248 667994 109304
rect 590290 103536 590346 103592
rect 666650 102788 666706 102844
rect 666650 102312 666706 102368
rect 553674 49136 553730 49192
rect 603078 51856 603134 51912
rect 612002 95784 612058 95840
rect 617522 77288 617578 77344
rect 604458 51584 604514 51640
rect 635554 96328 635610 96384
rect 635738 96056 635794 96112
rect 637026 96872 637082 96928
rect 641994 96056 642050 96112
rect 647422 96328 647478 96384
rect 647146 94968 647202 95024
rect 626446 94424 626502 94480
rect 625986 93608 626042 93664
rect 626446 92792 626502 92848
rect 625802 91976 625858 92032
rect 625434 88712 625490 88768
rect 626446 91160 626502 91216
rect 626446 90344 626502 90400
rect 626446 89548 626502 89584
rect 626446 89528 626448 89548
rect 626448 89528 626500 89548
rect 626500 89528 626502 89548
rect 626262 87896 626318 87952
rect 626446 87080 626502 87136
rect 626446 86300 626448 86320
rect 626448 86300 626500 86320
rect 626500 86300 626502 86320
rect 626446 86264 626502 86300
rect 626446 85484 626448 85504
rect 626448 85484 626500 85504
rect 626500 85484 626502 85504
rect 626446 85448 626502 85484
rect 625250 84632 625306 84688
rect 648618 91976 648674 92032
rect 552018 47776 552074 47832
rect 547878 47504 547934 47560
rect 521106 46960 521162 47016
rect 465262 46552 465318 46608
rect 625802 83816 625858 83872
rect 628746 83272 628802 83328
rect 629206 81640 629262 81696
rect 625802 77696 625858 77752
rect 633898 78512 633954 78568
rect 633898 77288 633954 77344
rect 639602 77696 639658 77752
rect 646134 67088 646190 67144
rect 646502 74160 646558 74216
rect 646870 68924 646926 68980
rect 646318 59336 646374 59392
rect 650182 89528 650238 89584
rect 650550 87080 650606 87136
rect 655058 94152 655114 94208
rect 654690 91432 654746 91488
rect 655426 93336 655482 93392
rect 655426 90652 655428 90672
rect 655428 90652 655480 90672
rect 655480 90652 655482 90672
rect 655426 90616 655482 90652
rect 655794 89800 655850 89856
rect 663706 92792 663762 92848
rect 664166 90616 664222 90672
rect 664534 91704 664590 91760
rect 664350 89800 664406 89856
rect 665362 93336 665418 93392
rect 665178 88984 665234 89040
rect 649998 84632 650054 84688
rect 668122 106120 668178 106176
rect 668398 106156 668400 106176
rect 668400 106156 668452 106176
rect 668452 106156 668454 106176
rect 668398 106120 668454 106156
rect 671894 151816 671950 151872
rect 672446 177928 672502 177984
rect 672538 175208 672594 175264
rect 672078 140392 672134 140448
rect 673182 214104 673238 214160
rect 672906 209616 672962 209672
rect 672906 200776 672962 200832
rect 672722 153040 672778 153096
rect 672538 130464 672594 130520
rect 672354 125976 672410 126032
rect 671710 115776 671766 115832
rect 673642 215328 673698 215384
rect 673366 201320 673422 201376
rect 675114 230016 675170 230072
rect 674838 229744 674894 229800
rect 676862 230288 676918 230344
rect 675114 229472 675170 229528
rect 675114 228792 675170 228848
rect 674746 226480 674802 226536
rect 674378 225664 674434 225720
rect 674562 225120 674618 225176
rect 674378 220632 674434 220688
rect 674378 220360 674434 220416
rect 674954 225936 675010 225992
rect 674654 218048 674710 218104
rect 676218 227024 676274 227080
rect 675298 226752 675354 226808
rect 675114 223352 675170 223408
rect 675574 224304 675630 224360
rect 674838 217504 674894 217560
rect 674562 216552 674618 216608
rect 675574 218864 675630 218920
rect 676034 218320 676090 218376
rect 676034 217776 676090 217832
rect 675114 216008 675170 216064
rect 675574 216144 675630 216200
rect 673826 211112 673882 211168
rect 674010 208256 674066 208312
rect 673826 203904 673882 203960
rect 673642 200776 673698 200832
rect 673182 197648 673238 197704
rect 673366 174392 673422 174448
rect 673182 169088 673238 169144
rect 673182 152496 673238 152552
rect 673918 172896 673974 172952
rect 674838 214648 674894 214704
rect 674654 213696 674710 213752
rect 674562 209616 674618 209672
rect 675850 215092 675852 215112
rect 675852 215092 675904 215112
rect 675904 215092 675906 215112
rect 675850 215056 675906 215092
rect 675758 214648 675814 214704
rect 676034 214512 676090 214568
rect 675850 214412 675852 214432
rect 675852 214412 675904 214432
rect 675904 214412 675906 214432
rect 675850 214376 675906 214412
rect 675850 213424 675906 213480
rect 675022 207304 675078 207360
rect 676770 211384 676826 211440
rect 677046 211384 677102 211440
rect 676310 211112 676366 211168
rect 675482 209616 675538 209672
rect 677690 209344 677746 209400
rect 676770 208256 676826 208312
rect 683302 234096 683358 234152
rect 683670 233824 683726 233880
rect 683302 223488 683358 223544
rect 683670 223080 683726 223136
rect 683486 222672 683542 222728
rect 683118 221448 683174 221504
rect 681002 220632 681058 220688
rect 684498 219816 684554 219872
rect 679622 219000 679678 219056
rect 683302 213288 683358 213344
rect 683118 212472 683174 212528
rect 683118 211112 683174 211168
rect 683302 210296 683358 210352
rect 679622 207032 679678 207088
rect 677874 206352 677930 206408
rect 675758 205536 675814 205592
rect 675666 204176 675722 204232
rect 674930 202544 674986 202600
rect 675390 202544 675446 202600
rect 675114 201320 675170 201376
rect 674838 200776 674894 200832
rect 675758 200776 675814 200832
rect 674654 196016 674710 196072
rect 675390 198328 675446 198384
rect 675482 197648 675538 197704
rect 675758 197104 675814 197160
rect 675206 196016 675262 196072
rect 675666 193160 675722 193216
rect 675114 192344 675170 192400
rect 675758 191528 675814 191584
rect 675850 181328 675906 181384
rect 674286 179424 674342 179480
rect 676034 178744 676090 178800
rect 675850 178064 675906 178120
rect 676034 177656 676090 177712
rect 674286 176840 674342 176896
rect 674102 154536 674158 154592
rect 674654 176024 674710 176080
rect 674470 168680 674526 168736
rect 674470 151000 674526 151056
rect 674286 132096 674342 132152
rect 676034 173168 676090 173224
rect 674838 172760 674894 172816
rect 675022 171128 675078 171184
rect 681002 171536 681058 171592
rect 676586 170720 676642 170776
rect 676034 167864 676090 167920
rect 674838 157528 674894 157584
rect 675206 161336 675262 161392
rect 676586 166368 676642 166424
rect 676034 165008 676090 165064
rect 675850 161336 675906 161392
rect 675758 159296 675814 159352
rect 675482 157528 675538 157584
rect 675758 156304 675814 156360
rect 675114 154808 675170 154864
rect 675482 152496 675538 152552
rect 675482 151816 675538 151872
rect 675298 151544 675354 151600
rect 675114 151000 675170 151056
rect 675666 150320 675722 150376
rect 675298 148960 675354 149016
rect 675758 148416 675814 148472
rect 675666 147600 675722 147656
rect 683302 142704 683358 142760
rect 683118 135904 683174 135960
rect 683302 133048 683358 133104
rect 683118 132640 683174 132696
rect 674654 131280 674710 131336
rect 676218 130192 676274 130248
rect 673366 129648 673422 129704
rect 674102 129240 674158 129296
rect 673182 124344 673238 124400
rect 672906 124072 672962 124128
rect 672906 123800 672962 123856
rect 672722 123120 672778 123176
rect 672538 122712 672594 122768
rect 672722 122168 672778 122224
rect 672538 112648 672594 112704
rect 672354 111424 672410 111480
rect 671526 107752 671582 107808
rect 673366 123528 673422 123584
rect 673182 110336 673238 110392
rect 672814 106256 672870 106312
rect 674286 128152 674342 128208
rect 676218 128152 676274 128208
rect 676862 128152 676918 128208
rect 674102 111016 674158 111072
rect 673366 105576 673422 105632
rect 668582 104352 668638 104408
rect 674838 127608 674894 127664
rect 674654 125568 674710 125624
rect 674470 125160 674526 125216
rect 675022 126384 675078 126440
rect 679622 127744 679678 127800
rect 676862 117272 676918 117328
rect 675298 113056 675354 113112
rect 675114 111424 675170 111480
rect 675114 110336 675170 110392
rect 675758 108160 675814 108216
rect 675114 106256 675170 106312
rect 675758 106120 675814 106176
rect 675114 105576 675170 105632
rect 675666 103128 675722 103184
rect 675666 102448 675722 102504
rect 674286 102312 674342 102368
rect 675758 101360 675814 101416
rect 668306 95784 668362 95840
rect 648894 82184 648950 82240
rect 648986 71712 649042 71768
rect 649170 64368 649226 64424
rect 648618 62056 648674 62112
rect 647238 57296 647294 57352
rect 662418 48456 662474 48512
rect 661590 47733 661646 47789
rect 464710 44240 464766 44296
rect 463882 44104 463938 44160
rect 465814 43560 465870 43616
rect 463698 42880 463754 42936
rect 460938 42336 460994 42392
rect 471058 43288 471114 43344
rect 518806 42744 518862 42800
rect 662602 47368 662658 47424
rect 515402 42064 515458 42120
rect 520922 42064 520978 42120
rect 522118 42064 522174 42120
rect 526442 42064 526498 42120
rect 529570 42064 529626 42120
rect 141698 40432 141754 40488
<< metal3 >>
rect 202689 1007450 202755 1007453
rect 202492 1007448 202755 1007450
rect 202492 1007392 202694 1007448
rect 202750 1007392 202755 1007448
rect 202492 1007390 202755 1007392
rect 202689 1007387 202755 1007390
rect 505369 1007178 505435 1007181
rect 505369 1007176 505632 1007178
rect 505369 1007120 505374 1007176
rect 505430 1007120 505632 1007176
rect 505369 1007118 505632 1007120
rect 505369 1007115 505435 1007118
rect 357709 1006906 357775 1006909
rect 427997 1006906 428063 1006909
rect 505369 1006906 505435 1006909
rect 554773 1006906 554839 1006909
rect 357604 1006904 357775 1006906
rect 357604 1006848 357714 1006904
rect 357770 1006848 357775 1006904
rect 357604 1006846 357775 1006848
rect 427800 1006904 428063 1006906
rect 427800 1006848 428002 1006904
rect 428058 1006848 428063 1006904
rect 427800 1006846 428063 1006848
rect 505172 1006904 505435 1006906
rect 505172 1006848 505374 1006904
rect 505430 1006848 505435 1006904
rect 505172 1006846 505435 1006848
rect 554576 1006904 554839 1006906
rect 554576 1006848 554778 1006904
rect 554834 1006848 554839 1006904
rect 554576 1006846 554839 1006848
rect 357709 1006843 357775 1006846
rect 427997 1006843 428063 1006846
rect 505369 1006843 505435 1006846
rect 554773 1006843 554839 1006846
rect 360193 1006770 360259 1006773
rect 430849 1006770 430915 1006773
rect 506197 1006770 506263 1006773
rect 359996 1006768 360259 1006770
rect 359996 1006712 360198 1006768
rect 360254 1006712 360259 1006768
rect 359996 1006710 360259 1006712
rect 430652 1006768 430915 1006770
rect 430652 1006712 430854 1006768
rect 430910 1006712 430915 1006768
rect 430652 1006710 430915 1006712
rect 506000 1006768 506263 1006770
rect 506000 1006712 506202 1006768
rect 506258 1006712 506263 1006768
rect 506000 1006710 506263 1006712
rect 360193 1006707 360259 1006710
rect 430849 1006707 430915 1006710
rect 506197 1006707 506263 1006710
rect 555969 1006770 556035 1006773
rect 555969 1006768 556232 1006770
rect 555969 1006712 555974 1006768
rect 556030 1006712 556232 1006768
rect 555969 1006710 556232 1006712
rect 555969 1006707 556035 1006710
rect 153745 1006634 153811 1006637
rect 153548 1006632 153811 1006634
rect 153548 1006576 153750 1006632
rect 153806 1006576 153811 1006632
rect 153548 1006574 153811 1006576
rect 153745 1006571 153811 1006574
rect 102317 1006498 102383 1006501
rect 152089 1006498 152155 1006501
rect 157425 1006498 157491 1006501
rect 210049 1006498 210115 1006501
rect 306925 1006498 306991 1006501
rect 430021 1006498 430087 1006501
rect 102317 1006496 102580 1006498
rect 102317 1006440 102322 1006496
rect 102378 1006440 102580 1006496
rect 102317 1006438 102580 1006440
rect 152089 1006496 152352 1006498
rect 152089 1006440 152094 1006496
rect 152150 1006440 152352 1006496
rect 152089 1006438 152352 1006440
rect 157228 1006496 157491 1006498
rect 157228 1006440 157430 1006496
rect 157486 1006440 157491 1006496
rect 157228 1006438 157491 1006440
rect 209852 1006496 210115 1006498
rect 209852 1006440 210054 1006496
rect 210110 1006440 210115 1006496
rect 209852 1006438 210115 1006440
rect 306728 1006496 306991 1006498
rect 306728 1006440 306930 1006496
rect 306986 1006440 306991 1006496
rect 306728 1006438 306991 1006440
rect 429824 1006496 430087 1006498
rect 429824 1006440 430026 1006496
rect 430082 1006440 430087 1006496
rect 429824 1006438 430087 1006440
rect 102317 1006435 102383 1006438
rect 152089 1006435 152155 1006438
rect 157425 1006435 157491 1006438
rect 210049 1006435 210115 1006438
rect 306925 1006435 306991 1006438
rect 430021 1006435 430087 1006438
rect 431677 1006498 431743 1006501
rect 508221 1006498 508287 1006501
rect 559649 1006498 559715 1006501
rect 431677 1006496 431940 1006498
rect 431677 1006440 431682 1006496
rect 431738 1006440 431940 1006496
rect 431677 1006438 431940 1006440
rect 508221 1006496 508484 1006498
rect 508221 1006440 508226 1006496
rect 508282 1006440 508484 1006496
rect 508221 1006438 508484 1006440
rect 559452 1006496 559715 1006498
rect 559452 1006440 559654 1006496
rect 559710 1006440 559715 1006496
rect 559452 1006438 559715 1006440
rect 431677 1006435 431743 1006438
rect 508221 1006435 508287 1006438
rect 559649 1006435 559715 1006438
rect 101949 1006362 102015 1006365
rect 151721 1006362 151787 1006365
rect 158253 1006362 158319 1006365
rect 210417 1006362 210483 1006365
rect 256141 1006362 256207 1006365
rect 361389 1006362 361455 1006365
rect 101949 1006360 102212 1006362
rect 101949 1006304 101954 1006360
rect 102010 1006304 102212 1006360
rect 101949 1006302 102212 1006304
rect 151721 1006360 151892 1006362
rect 151721 1006304 151726 1006360
rect 151782 1006304 151892 1006360
rect 151721 1006302 151892 1006304
rect 158056 1006360 158319 1006362
rect 158056 1006304 158258 1006360
rect 158314 1006304 158319 1006360
rect 158056 1006302 158319 1006304
rect 210220 1006360 210483 1006362
rect 210220 1006304 210422 1006360
rect 210478 1006304 210483 1006360
rect 210220 1006302 210483 1006304
rect 255944 1006360 256207 1006362
rect 255944 1006304 256146 1006360
rect 256202 1006304 256207 1006360
rect 255944 1006302 256207 1006304
rect 361192 1006360 361455 1006362
rect 361192 1006304 361394 1006360
rect 361450 1006304 361455 1006360
rect 361192 1006302 361455 1006304
rect 101949 1006299 102015 1006302
rect 151721 1006299 151787 1006302
rect 158253 1006299 158319 1006302
rect 210417 1006299 210483 1006302
rect 256141 1006299 256207 1006302
rect 361389 1006299 361455 1006302
rect 429193 1006362 429259 1006365
rect 429193 1006360 429456 1006362
rect 429193 1006304 429198 1006360
rect 429254 1006304 429456 1006360
rect 429193 1006302 429456 1006304
rect 429193 1006299 429259 1006302
rect 103973 1006226 104039 1006229
rect 107653 1006226 107719 1006229
rect 103973 1006224 104236 1006226
rect 103973 1006168 103978 1006224
rect 104034 1006168 104236 1006224
rect 103973 1006166 104236 1006168
rect 107456 1006224 107719 1006226
rect 107456 1006168 107658 1006224
rect 107714 1006168 107719 1006224
rect 107456 1006166 107719 1006168
rect 103973 1006163 104039 1006166
rect 107653 1006163 107719 1006166
rect 150893 1006226 150959 1006229
rect 160277 1006226 160343 1006229
rect 150893 1006224 151156 1006226
rect 150893 1006168 150898 1006224
rect 150954 1006168 151156 1006224
rect 150893 1006166 151156 1006168
rect 160080 1006224 160343 1006226
rect 160080 1006168 160282 1006224
rect 160338 1006168 160343 1006224
rect 160080 1006166 160343 1006168
rect 150893 1006163 150959 1006166
rect 160277 1006163 160343 1006166
rect 208393 1006226 208459 1006229
rect 255313 1006226 255379 1006229
rect 261845 1006226 261911 1006229
rect 306097 1006226 306163 1006229
rect 357341 1006226 357407 1006229
rect 431677 1006226 431743 1006229
rect 507025 1006226 507091 1006229
rect 556797 1006226 556863 1006229
rect 208393 1006224 208656 1006226
rect 208393 1006168 208398 1006224
rect 208454 1006168 208656 1006224
rect 208393 1006166 208656 1006168
rect 255116 1006224 255379 1006226
rect 255116 1006168 255318 1006224
rect 255374 1006168 255379 1006224
rect 255116 1006166 255379 1006168
rect 261648 1006224 261911 1006226
rect 261648 1006168 261850 1006224
rect 261906 1006168 261911 1006224
rect 261648 1006166 261911 1006168
rect 305900 1006224 306163 1006226
rect 305900 1006168 306102 1006224
rect 306158 1006168 306163 1006224
rect 305900 1006166 306163 1006168
rect 357144 1006224 357407 1006226
rect 357144 1006168 357346 1006224
rect 357402 1006168 357407 1006224
rect 357144 1006166 357407 1006168
rect 431480 1006224 431743 1006226
rect 431480 1006168 431682 1006224
rect 431738 1006168 431743 1006224
rect 431480 1006166 431743 1006168
rect 506828 1006224 507091 1006226
rect 506828 1006168 507030 1006224
rect 507086 1006168 507091 1006224
rect 506828 1006166 507091 1006168
rect 556600 1006224 556863 1006226
rect 556600 1006168 556802 1006224
rect 556858 1006168 556863 1006224
rect 556600 1006166 556863 1006168
rect 208393 1006163 208459 1006166
rect 255313 1006163 255379 1006166
rect 261845 1006163 261911 1006166
rect 306097 1006163 306163 1006166
rect 357341 1006163 357407 1006166
rect 431677 1006163 431743 1006166
rect 507025 1006163 507091 1006166
rect 556797 1006163 556863 1006166
rect 98269 1006090 98335 1006093
rect 104801 1006090 104867 1006093
rect 108481 1006090 108547 1006093
rect 150065 1006090 150131 1006093
rect 159449 1006090 159515 1006093
rect 201033 1006090 201099 1006093
rect 209221 1006090 209287 1006093
rect 252461 1006090 252527 1006093
rect 260189 1006090 260255 1006093
rect 98269 1006088 98900 1006090
rect 98269 1006032 98274 1006088
rect 98330 1006032 98900 1006088
rect 98269 1006030 98900 1006032
rect 104801 1006088 104972 1006090
rect 104801 1006032 104806 1006088
rect 104862 1006032 104972 1006088
rect 104801 1006030 104972 1006032
rect 108284 1006088 108547 1006090
rect 108284 1006032 108486 1006088
rect 108542 1006032 108547 1006088
rect 108284 1006030 108547 1006032
rect 149868 1006088 150328 1006090
rect 149868 1006032 150070 1006088
rect 150126 1006032 150328 1006088
rect 149868 1006030 150328 1006032
rect 159449 1006088 159712 1006090
rect 159449 1006032 159454 1006088
rect 159510 1006032 159712 1006088
rect 159449 1006030 159712 1006032
rect 201033 1006088 201756 1006090
rect 201033 1006032 201038 1006088
rect 201094 1006032 201756 1006088
rect 201033 1006030 201756 1006032
rect 209221 1006088 209484 1006090
rect 209221 1006032 209226 1006088
rect 209282 1006032 209484 1006088
rect 209221 1006030 209484 1006032
rect 252461 1006088 253092 1006090
rect 252461 1006032 252466 1006088
rect 252522 1006032 253092 1006088
rect 252461 1006030 253092 1006032
rect 260084 1006088 260255 1006090
rect 260084 1006032 260194 1006088
rect 260250 1006032 260255 1006088
rect 260084 1006030 260255 1006032
rect 98269 1006027 98335 1006030
rect 104801 1006027 104867 1006030
rect 108481 1006027 108547 1006030
rect 150065 1006027 150131 1006030
rect 159449 1006027 159515 1006030
rect 201033 1006027 201099 1006030
rect 209221 1006027 209287 1006030
rect 252461 1006027 252527 1006030
rect 260189 1006027 260255 1006030
rect 301681 1006090 301747 1006093
rect 303245 1006090 303311 1006093
rect 301681 1006088 303311 1006090
rect 301681 1006032 301686 1006088
rect 301742 1006032 303250 1006088
rect 303306 1006032 303311 1006088
rect 301681 1006030 303311 1006032
rect 301681 1006027 301747 1006030
rect 303245 1006027 303311 1006030
rect 304073 1006090 304139 1006093
rect 311801 1006090 311867 1006093
rect 314653 1006090 314719 1006093
rect 354857 1006090 354923 1006093
rect 356881 1006090 356947 1006093
rect 363413 1006090 363479 1006093
rect 304073 1006088 304704 1006090
rect 304073 1006032 304078 1006088
rect 304134 1006032 304704 1006088
rect 304073 1006030 304704 1006032
rect 311801 1006088 312064 1006090
rect 311801 1006032 311806 1006088
rect 311862 1006032 312064 1006088
rect 311801 1006030 312064 1006032
rect 314653 1006088 314916 1006090
rect 314653 1006032 314658 1006088
rect 314714 1006032 314916 1006088
rect 314653 1006030 314916 1006032
rect 354660 1006088 355120 1006090
rect 354660 1006032 354862 1006088
rect 354918 1006032 355120 1006088
rect 354660 1006030 355120 1006032
rect 356684 1006088 356947 1006090
rect 356684 1006032 356886 1006088
rect 356942 1006032 356947 1006088
rect 356684 1006030 356947 1006032
rect 363308 1006088 363479 1006090
rect 363308 1006032 363418 1006088
rect 363474 1006032 363479 1006088
rect 363308 1006030 363479 1006032
rect 304073 1006027 304139 1006030
rect 311801 1006027 311867 1006030
rect 314653 1006027 314719 1006030
rect 354857 1006027 354923 1006030
rect 356881 1006027 356947 1006030
rect 363413 1006027 363479 1006030
rect 421833 1006090 421899 1006093
rect 428365 1006090 428431 1006093
rect 498837 1006090 498903 1006093
rect 502517 1006090 502583 1006093
rect 509049 1006090 509115 1006093
rect 551093 1006090 551159 1006093
rect 421833 1006088 422556 1006090
rect 421833 1006032 421838 1006088
rect 421894 1006032 422556 1006088
rect 421833 1006030 422556 1006032
rect 428365 1006088 428628 1006090
rect 428365 1006032 428370 1006088
rect 428426 1006032 428628 1006088
rect 428365 1006030 428628 1006032
rect 498837 1006088 499468 1006090
rect 498837 1006032 498842 1006088
rect 498898 1006032 499468 1006088
rect 498837 1006030 499468 1006032
rect 502517 1006088 502780 1006090
rect 502517 1006032 502522 1006088
rect 502578 1006032 502780 1006088
rect 502517 1006030 502780 1006032
rect 509049 1006088 509312 1006090
rect 509049 1006032 509054 1006088
rect 509110 1006032 509312 1006088
rect 509049 1006030 509312 1006032
rect 550436 1006088 551159 1006090
rect 550436 1006032 551098 1006088
rect 551154 1006032 551159 1006088
rect 550436 1006030 551159 1006032
rect 421833 1006027 421899 1006030
rect 428365 1006027 428431 1006030
rect 498837 1006027 498903 1006030
rect 502517 1006027 502583 1006030
rect 509049 1006027 509115 1006030
rect 551093 1006027 551159 1006030
rect 555141 1006090 555207 1006093
rect 557165 1006090 557231 1006093
rect 555141 1006088 555404 1006090
rect 555141 1006032 555146 1006088
rect 555202 1006032 555404 1006088
rect 555141 1006030 555404 1006032
rect 557060 1006088 557231 1006090
rect 557060 1006032 557170 1006088
rect 557226 1006032 557231 1006088
rect 557060 1006030 557231 1006032
rect 555141 1006027 555207 1006030
rect 557165 1006027 557231 1006030
rect 304073 1005818 304139 1005821
rect 303876 1005816 304139 1005818
rect 303876 1005760 304078 1005816
rect 304134 1005760 304139 1005816
rect 303876 1005758 304139 1005760
rect 304073 1005755 304139 1005758
rect 425513 1005682 425579 1005685
rect 505001 1005682 505067 1005685
rect 425316 1005680 425579 1005682
rect 425316 1005624 425518 1005680
rect 425574 1005624 425579 1005680
rect 425316 1005622 425579 1005624
rect 504804 1005680 505067 1005682
rect 504804 1005624 505006 1005680
rect 505062 1005624 505067 1005680
rect 504804 1005622 505067 1005624
rect 425513 1005619 425579 1005622
rect 505001 1005619 505067 1005622
rect 360561 1005546 360627 1005549
rect 427169 1005546 427235 1005549
rect 360364 1005544 360627 1005546
rect 360364 1005488 360566 1005544
rect 360622 1005488 360627 1005544
rect 360364 1005486 360627 1005488
rect 426972 1005544 427235 1005546
rect 426972 1005488 427174 1005544
rect 427230 1005488 427235 1005544
rect 426972 1005486 427235 1005488
rect 360561 1005483 360627 1005486
rect 427169 1005483 427235 1005486
rect 152917 1005410 152983 1005413
rect 152720 1005408 152983 1005410
rect 152720 1005352 152922 1005408
rect 152978 1005352 152983 1005408
rect 152720 1005350 152983 1005352
rect 152917 1005347 152983 1005350
rect 358537 1005410 358603 1005413
rect 428365 1005410 428431 1005413
rect 502149 1005410 502215 1005413
rect 553117 1005410 553183 1005413
rect 358537 1005408 358800 1005410
rect 358537 1005352 358542 1005408
rect 358598 1005352 358800 1005408
rect 358537 1005350 358800 1005352
rect 428260 1005408 428431 1005410
rect 428260 1005352 428370 1005408
rect 428426 1005352 428431 1005408
rect 428260 1005350 428431 1005352
rect 501952 1005408 502215 1005410
rect 501952 1005352 502154 1005408
rect 502210 1005352 502215 1005408
rect 501952 1005350 502215 1005352
rect 552920 1005408 553183 1005410
rect 552920 1005352 553122 1005408
rect 553178 1005352 553183 1005408
rect 552920 1005350 553183 1005352
rect 358537 1005347 358603 1005350
rect 428365 1005347 428431 1005350
rect 502149 1005347 502215 1005350
rect 553117 1005347 553183 1005350
rect 357709 1005274 357775 1005277
rect 423489 1005274 423555 1005277
rect 357709 1005272 357972 1005274
rect 357709 1005216 357714 1005272
rect 357770 1005216 357972 1005272
rect 357709 1005214 357972 1005216
rect 423292 1005272 423555 1005274
rect 423292 1005216 423494 1005272
rect 423550 1005216 423555 1005272
rect 423292 1005214 423555 1005216
rect 357709 1005211 357775 1005214
rect 423489 1005211 423555 1005214
rect 499665 1005274 499731 1005277
rect 551461 1005274 551527 1005277
rect 499665 1005272 499928 1005274
rect 499665 1005216 499670 1005272
rect 499726 1005216 499928 1005272
rect 499665 1005214 499928 1005216
rect 551356 1005272 551527 1005274
rect 551356 1005216 551466 1005272
rect 551522 1005216 551527 1005272
rect 551356 1005214 551527 1005216
rect 499665 1005211 499731 1005214
rect 551461 1005211 551527 1005214
rect 152917 1005138 152983 1005141
rect 208393 1005138 208459 1005141
rect 500493 1005138 500559 1005141
rect 152917 1005136 153180 1005138
rect 152917 1005080 152922 1005136
rect 152978 1005080 153180 1005136
rect 152917 1005078 153180 1005080
rect 208196 1005136 208459 1005138
rect 208196 1005080 208398 1005136
rect 208454 1005080 208459 1005136
rect 208196 1005078 208459 1005080
rect 500296 1005136 500559 1005138
rect 500296 1005080 500498 1005136
rect 500554 1005080 500559 1005136
rect 500296 1005078 500559 1005080
rect 152917 1005075 152983 1005078
rect 208393 1005075 208459 1005078
rect 500493 1005075 500559 1005078
rect 153745 1005002 153811 1005005
rect 158621 1005002 158687 1005005
rect 207565 1005002 207631 1005005
rect 263041 1005002 263107 1005005
rect 313825 1005002 313891 1005005
rect 153745 1005000 153916 1005002
rect 153745 1004944 153750 1005000
rect 153806 1004944 153916 1005000
rect 153745 1004942 153916 1004944
rect 158621 1005000 158884 1005002
rect 158621 1004944 158626 1005000
rect 158682 1004944 158884 1005000
rect 158621 1004942 158884 1004944
rect 207565 1005000 207828 1005002
rect 207565 1004944 207570 1005000
rect 207626 1004944 207828 1005000
rect 207565 1004942 207828 1004944
rect 262844 1005000 263107 1005002
rect 262844 1004944 263046 1005000
rect 263102 1004944 263107 1005000
rect 262844 1004942 263107 1004944
rect 313628 1005000 313891 1005002
rect 313628 1004944 313830 1005000
rect 313886 1004944 313891 1005000
rect 313628 1004942 313891 1004944
rect 153745 1004939 153811 1004942
rect 158621 1004939 158687 1004942
rect 207565 1004939 207631 1004942
rect 263041 1004939 263107 1004942
rect 313825 1004939 313891 1004942
rect 361389 1005002 361455 1005005
rect 431217 1005002 431283 1005005
rect 361389 1005000 361652 1005002
rect 361389 1004944 361394 1005000
rect 361450 1004944 361652 1005000
rect 361389 1004942 361652 1004944
rect 431020 1005000 431283 1005002
rect 431020 1004944 431222 1005000
rect 431278 1004944 431283 1005000
rect 431020 1004942 431283 1004944
rect 361389 1004939 361455 1004942
rect 431217 1004939 431283 1004942
rect 160645 1004866 160711 1004869
rect 209221 1004866 209287 1004869
rect 314653 1004866 314719 1004869
rect 355685 1004866 355751 1004869
rect 362585 1004866 362651 1004869
rect 160540 1004864 160711 1004866
rect 160540 1004808 160650 1004864
rect 160706 1004808 160711 1004864
rect 160540 1004806 160711 1004808
rect 209024 1004864 209287 1004866
rect 209024 1004808 209226 1004864
rect 209282 1004808 209287 1004864
rect 209024 1004806 209287 1004808
rect 314548 1004864 314719 1004866
rect 314548 1004808 314658 1004864
rect 314714 1004808 314719 1004864
rect 314548 1004806 314719 1004808
rect 355488 1004864 355751 1004866
rect 355488 1004808 355690 1004864
rect 355746 1004808 355751 1004864
rect 355488 1004806 355751 1004808
rect 362388 1004864 362651 1004866
rect 362388 1004808 362590 1004864
rect 362646 1004808 362651 1004864
rect 362388 1004806 362651 1004808
rect 160645 1004803 160711 1004806
rect 209221 1004803 209287 1004806
rect 314653 1004803 314719 1004806
rect 355685 1004803 355751 1004806
rect 362585 1004803 362651 1004806
rect 422661 1004866 422727 1004869
rect 432045 1004866 432111 1004869
rect 500493 1004866 500559 1004869
rect 507853 1004866 507919 1004869
rect 555969 1004866 556035 1004869
rect 422661 1004864 422924 1004866
rect 422661 1004808 422666 1004864
rect 422722 1004808 422924 1004864
rect 422661 1004806 422924 1004808
rect 432045 1004864 432308 1004866
rect 432045 1004808 432050 1004864
rect 432106 1004808 432308 1004864
rect 432045 1004806 432308 1004808
rect 500493 1004864 500756 1004866
rect 500493 1004808 500498 1004864
rect 500554 1004808 500756 1004864
rect 500493 1004806 500756 1004808
rect 507656 1004864 507919 1004866
rect 507656 1004808 507858 1004864
rect 507914 1004808 507919 1004864
rect 507656 1004806 507919 1004808
rect 555772 1004864 556035 1004866
rect 555772 1004808 555974 1004864
rect 556030 1004808 556035 1004864
rect 555772 1004806 556035 1004808
rect 422661 1004803 422727 1004806
rect 432045 1004803 432111 1004806
rect 500493 1004803 500559 1004806
rect 507853 1004803 507919 1004806
rect 555969 1004803 556035 1004806
rect 154113 1004730 154179 1004733
rect 161105 1004730 161171 1004733
rect 212533 1004730 212599 1004733
rect 315481 1004730 315547 1004733
rect 356513 1004730 356579 1004733
rect 364241 1004730 364307 1004733
rect 154113 1004728 154376 1004730
rect 154113 1004672 154118 1004728
rect 154174 1004672 154376 1004728
rect 154113 1004670 154376 1004672
rect 160908 1004728 161171 1004730
rect 160908 1004672 161110 1004728
rect 161166 1004672 161171 1004728
rect 160908 1004670 161171 1004672
rect 212336 1004728 212599 1004730
rect 212336 1004672 212538 1004728
rect 212594 1004672 212599 1004728
rect 212336 1004670 212599 1004672
rect 315284 1004728 315547 1004730
rect 315284 1004672 315486 1004728
rect 315542 1004672 315547 1004728
rect 315284 1004670 315547 1004672
rect 356316 1004728 356579 1004730
rect 356316 1004672 356518 1004728
rect 356574 1004672 356579 1004728
rect 356316 1004670 356579 1004672
rect 364044 1004728 364307 1004730
rect 364044 1004672 364246 1004728
rect 364302 1004672 364307 1004728
rect 364044 1004670 364307 1004672
rect 154113 1004667 154179 1004670
rect 161105 1004667 161171 1004670
rect 212533 1004667 212599 1004670
rect 315481 1004667 315547 1004670
rect 356513 1004667 356579 1004670
rect 364241 1004667 364307 1004670
rect 430021 1004730 430087 1004733
rect 501321 1004730 501387 1004733
rect 507393 1004730 507459 1004733
rect 557625 1004730 557691 1004733
rect 430021 1004728 430284 1004730
rect 430021 1004672 430026 1004728
rect 430082 1004672 430284 1004728
rect 430021 1004670 430284 1004672
rect 501124 1004728 501387 1004730
rect 501124 1004672 501326 1004728
rect 501382 1004672 501387 1004728
rect 501124 1004670 501387 1004672
rect 507196 1004728 507459 1004730
rect 507196 1004672 507398 1004728
rect 507454 1004672 507459 1004728
rect 507196 1004670 507459 1004672
rect 557428 1004728 557691 1004730
rect 557428 1004672 557630 1004728
rect 557686 1004672 557691 1004728
rect 557428 1004670 557691 1004672
rect 430021 1004667 430087 1004670
rect 501321 1004667 501387 1004670
rect 507393 1004667 507459 1004670
rect 557625 1004667 557691 1004670
rect 560845 1004730 560911 1004733
rect 560845 1004728 561108 1004730
rect 560845 1004672 560850 1004728
rect 560906 1004672 561108 1004728
rect 560845 1004670 561108 1004672
rect 560845 1004667 560911 1004670
rect 424685 1004050 424751 1004053
rect 424580 1004048 424751 1004050
rect 424580 1003992 424690 1004048
rect 424746 1003992 424751 1004048
rect 424580 1003990 424751 1003992
rect 424685 1003987 424751 1003990
rect 360561 1003914 360627 1003917
rect 426341 1003914 426407 1003917
rect 504541 1003914 504607 1003917
rect 360561 1003912 360824 1003914
rect 360561 1003856 360566 1003912
rect 360622 1003856 360824 1003912
rect 360561 1003854 360824 1003856
rect 426341 1003912 426604 1003914
rect 426341 1003856 426346 1003912
rect 426402 1003856 426604 1003912
rect 426341 1003854 426604 1003856
rect 504436 1003912 504607 1003914
rect 504436 1003856 504546 1003912
rect 504602 1003856 504607 1003912
rect 504436 1003854 504607 1003856
rect 360561 1003851 360627 1003854
rect 426341 1003851 426407 1003854
rect 504541 1003851 504607 1003854
rect 552289 1003914 552355 1003917
rect 552289 1003912 552552 1003914
rect 552289 1003856 552294 1003912
rect 552350 1003856 552552 1003912
rect 552289 1003854 552552 1003856
rect 552289 1003851 552355 1003854
rect 355685 1003370 355751 1003373
rect 355685 1003368 355948 1003370
rect 355685 1003312 355690 1003368
rect 355746 1003312 355948 1003368
rect 355685 1003310 355948 1003312
rect 355685 1003307 355751 1003310
rect 100293 1002690 100359 1002693
rect 106825 1002690 106891 1002693
rect 100293 1002688 100556 1002690
rect 100293 1002632 100298 1002688
rect 100354 1002632 100556 1002688
rect 100293 1002630 100556 1002632
rect 106628 1002688 106891 1002690
rect 106628 1002632 106830 1002688
rect 106886 1002632 106891 1002688
rect 106628 1002630 106891 1002632
rect 100293 1002627 100359 1002630
rect 106825 1002627 106891 1002630
rect 256141 1002690 256207 1002693
rect 558821 1002690 558887 1002693
rect 256141 1002688 256404 1002690
rect 256141 1002632 256146 1002688
rect 256202 1002632 256404 1002688
rect 256141 1002630 256404 1002632
rect 558821 1002688 559084 1002690
rect 558821 1002632 558826 1002688
rect 558882 1002632 559084 1002688
rect 558821 1002630 559084 1002632
rect 256141 1002627 256207 1002630
rect 558821 1002627 558887 1002630
rect 99465 1002554 99531 1002557
rect 103145 1002554 103211 1002557
rect 108021 1002554 108087 1002557
rect 99465 1002552 99728 1002554
rect 99465 1002496 99470 1002552
rect 99526 1002496 99728 1002552
rect 99465 1002494 99728 1002496
rect 103145 1002552 103408 1002554
rect 103145 1002496 103150 1002552
rect 103206 1002496 103408 1002552
rect 103145 1002494 103408 1002496
rect 107916 1002552 108087 1002554
rect 107916 1002496 108026 1002552
rect 108082 1002496 108087 1002552
rect 107916 1002494 108087 1002496
rect 99465 1002491 99531 1002494
rect 103145 1002491 103211 1002494
rect 108021 1002491 108087 1002494
rect 155769 1002554 155835 1002557
rect 207197 1002554 207263 1002557
rect 155769 1002552 156032 1002554
rect 155769 1002496 155774 1002552
rect 155830 1002496 156032 1002552
rect 155769 1002494 156032 1002496
rect 207000 1002552 207263 1002554
rect 207000 1002496 207202 1002552
rect 207258 1002496 207263 1002552
rect 207000 1002494 207263 1002496
rect 155769 1002491 155835 1002494
rect 207197 1002491 207263 1002494
rect 211245 1002554 211311 1002557
rect 254485 1002554 254551 1002557
rect 358537 1002554 358603 1002557
rect 211245 1002552 211508 1002554
rect 211245 1002496 211250 1002552
rect 211306 1002496 211508 1002552
rect 211245 1002494 211508 1002496
rect 254485 1002552 254748 1002554
rect 254485 1002496 254490 1002552
rect 254546 1002496 254748 1002552
rect 254485 1002494 254748 1002496
rect 358340 1002552 358603 1002554
rect 358340 1002496 358542 1002552
rect 358598 1002496 358603 1002552
rect 358340 1002494 358603 1002496
rect 211245 1002491 211311 1002494
rect 254485 1002491 254551 1002494
rect 358537 1002491 358603 1002494
rect 423489 1002554 423555 1002557
rect 560845 1002554 560911 1002557
rect 423489 1002552 423752 1002554
rect 423489 1002496 423494 1002552
rect 423550 1002496 423752 1002552
rect 423489 1002494 423752 1002496
rect 560740 1002552 560911 1002554
rect 560740 1002496 560850 1002552
rect 560906 1002496 560911 1002552
rect 560740 1002494 560911 1002496
rect 423489 1002491 423555 1002494
rect 560845 1002491 560911 1002494
rect 100293 1002418 100359 1002421
rect 105997 1002418 106063 1002421
rect 100096 1002416 100359 1002418
rect 100096 1002360 100298 1002416
rect 100354 1002360 100359 1002416
rect 100096 1002358 100359 1002360
rect 105892 1002416 106063 1002418
rect 105892 1002360 106002 1002416
rect 106058 1002360 106063 1002416
rect 105892 1002358 106063 1002360
rect 100293 1002355 100359 1002358
rect 105997 1002355 106063 1002358
rect 156597 1002418 156663 1002421
rect 261017 1002418 261083 1002421
rect 156597 1002416 156860 1002418
rect 156597 1002360 156602 1002416
rect 156658 1002360 156860 1002416
rect 156597 1002358 156860 1002360
rect 260820 1002416 261083 1002418
rect 260820 1002360 261022 1002416
rect 261078 1002360 261083 1002416
rect 260820 1002358 261083 1002360
rect 156597 1002355 156663 1002358
rect 261017 1002355 261083 1002358
rect 503345 1002418 503411 1002421
rect 557993 1002418 558059 1002421
rect 503345 1002416 503608 1002418
rect 503345 1002360 503350 1002416
rect 503406 1002360 503608 1002416
rect 503345 1002358 503608 1002360
rect 557993 1002416 558256 1002418
rect 557993 1002360 557998 1002416
rect 558054 1002360 558256 1002416
rect 557993 1002358 558256 1002360
rect 503345 1002355 503411 1002358
rect 557993 1002355 558059 1002358
rect 101121 1002282 101187 1002285
rect 105629 1002282 105695 1002285
rect 100924 1002280 101187 1002282
rect 100924 1002224 101126 1002280
rect 101182 1002224 101187 1002280
rect 100924 1002222 101187 1002224
rect 105432 1002280 105695 1002282
rect 105432 1002224 105634 1002280
rect 105690 1002224 105695 1002280
rect 105432 1002222 105695 1002224
rect 101121 1002219 101187 1002222
rect 105629 1002219 105695 1002222
rect 108849 1002282 108915 1002285
rect 151721 1002282 151787 1002285
rect 155769 1002282 155835 1002285
rect 108849 1002280 109112 1002282
rect 108849 1002224 108854 1002280
rect 108910 1002224 109112 1002280
rect 108849 1002222 109112 1002224
rect 151524 1002280 151787 1002282
rect 151524 1002224 151726 1002280
rect 151782 1002224 151787 1002280
rect 151524 1002222 151787 1002224
rect 155572 1002280 155835 1002282
rect 155572 1002224 155774 1002280
rect 155830 1002224 155835 1002280
rect 155572 1002222 155835 1002224
rect 108849 1002219 108915 1002222
rect 151721 1002219 151787 1002222
rect 155769 1002219 155835 1002222
rect 207197 1002282 207263 1002285
rect 211245 1002282 211311 1002285
rect 262673 1002282 262739 1002285
rect 207197 1002280 207460 1002282
rect 207197 1002224 207202 1002280
rect 207258 1002224 207460 1002280
rect 207197 1002222 207460 1002224
rect 211140 1002280 211311 1002282
rect 211140 1002224 211250 1002280
rect 211306 1002224 211311 1002280
rect 211140 1002222 211311 1002224
rect 262476 1002280 262739 1002282
rect 262476 1002224 262678 1002280
rect 262734 1002224 262739 1002280
rect 262476 1002222 262739 1002224
rect 207197 1002219 207263 1002222
rect 211245 1002219 211311 1002222
rect 262673 1002219 262739 1002222
rect 359365 1002282 359431 1002285
rect 365069 1002282 365135 1002285
rect 504173 1002282 504239 1002285
rect 553945 1002282 554011 1002285
rect 560477 1002282 560543 1002285
rect 359365 1002280 359628 1002282
rect 359365 1002224 359370 1002280
rect 359426 1002224 359628 1002280
rect 359365 1002222 359628 1002224
rect 364872 1002280 365135 1002282
rect 364872 1002224 365074 1002280
rect 365130 1002224 365135 1002280
rect 364872 1002222 365135 1002224
rect 503976 1002280 504239 1002282
rect 503976 1002224 504178 1002280
rect 504234 1002224 504239 1002280
rect 503976 1002222 504239 1002224
rect 553748 1002280 554011 1002282
rect 553748 1002224 553950 1002280
rect 554006 1002224 554011 1002280
rect 553748 1002222 554011 1002224
rect 560280 1002280 560543 1002282
rect 560280 1002224 560482 1002280
rect 560538 1002224 560543 1002280
rect 560280 1002222 560543 1002224
rect 359365 1002219 359431 1002222
rect 365069 1002219 365135 1002222
rect 504173 1002219 504239 1002222
rect 553945 1002219 554011 1002222
rect 560477 1002219 560543 1002222
rect 99097 1002146 99163 1002149
rect 101949 1002146 102015 1002149
rect 99097 1002144 99268 1002146
rect 99097 1002088 99102 1002144
rect 99158 1002088 99268 1002144
rect 99097 1002086 99268 1002088
rect 101752 1002144 102015 1002146
rect 101752 1002088 101954 1002144
rect 102010 1002088 102015 1002144
rect 101752 1002086 102015 1002088
rect 99097 1002083 99163 1002086
rect 101949 1002083 102015 1002086
rect 106825 1002146 106891 1002149
rect 109677 1002146 109743 1002149
rect 150893 1002146 150959 1002149
rect 156597 1002146 156663 1002149
rect 206369 1002146 206435 1002149
rect 210877 1002146 210943 1002149
rect 106825 1002144 107088 1002146
rect 106825 1002088 106830 1002144
rect 106886 1002088 107088 1002144
rect 106825 1002086 107088 1002088
rect 109480 1002144 109743 1002146
rect 109480 1002088 109682 1002144
rect 109738 1002088 109743 1002144
rect 109480 1002086 109743 1002088
rect 150696 1002144 150959 1002146
rect 150696 1002088 150898 1002144
rect 150954 1002088 150959 1002144
rect 150696 1002086 150959 1002088
rect 156400 1002144 156663 1002146
rect 156400 1002088 156602 1002144
rect 156658 1002088 156663 1002144
rect 156400 1002086 156663 1002088
rect 206172 1002144 206435 1002146
rect 206172 1002088 206374 1002144
rect 206430 1002088 206435 1002144
rect 206172 1002086 206435 1002088
rect 210680 1002144 210943 1002146
rect 210680 1002088 210882 1002144
rect 210938 1002088 210943 1002144
rect 210680 1002086 210943 1002088
rect 106825 1002083 106891 1002086
rect 109677 1002083 109743 1002086
rect 150893 1002083 150959 1002086
rect 156597 1002083 156663 1002086
rect 206369 1002083 206435 1002086
rect 210877 1002083 210943 1002086
rect 254117 1002146 254183 1002149
rect 263869 1002146 263935 1002149
rect 254117 1002144 254380 1002146
rect 254117 1002088 254122 1002144
rect 254178 1002088 254380 1002144
rect 254117 1002086 254380 1002088
rect 263764 1002144 263935 1002146
rect 263764 1002088 263874 1002144
rect 263930 1002088 263935 1002144
rect 263764 1002086 263935 1002088
rect 254117 1002083 254183 1002086
rect 263869 1002083 263935 1002086
rect 304901 1002146 304967 1002149
rect 310145 1002146 310211 1002149
rect 365897 1002146 365963 1002149
rect 304901 1002144 305164 1002146
rect 304901 1002088 304906 1002144
rect 304962 1002088 305164 1002144
rect 304901 1002086 305164 1002088
rect 309948 1002144 310211 1002146
rect 309948 1002088 310150 1002144
rect 310206 1002088 310211 1002144
rect 309948 1002086 310211 1002088
rect 365700 1002144 365963 1002146
rect 365700 1002088 365902 1002144
rect 365958 1002088 365963 1002144
rect 365700 1002086 365963 1002088
rect 304901 1002083 304967 1002086
rect 310145 1002083 310211 1002086
rect 365897 1002083 365963 1002086
rect 425513 1002146 425579 1002149
rect 427537 1002146 427603 1002149
rect 433333 1002146 433399 1002149
rect 502517 1002146 502583 1002149
rect 509877 1002146 509943 1002149
rect 560017 1002146 560083 1002149
rect 425513 1002144 425776 1002146
rect 425513 1002088 425518 1002144
rect 425574 1002088 425776 1002144
rect 425513 1002086 425776 1002088
rect 427340 1002144 427603 1002146
rect 427340 1002088 427542 1002144
rect 427598 1002088 427603 1002144
rect 427340 1002086 427603 1002088
rect 433136 1002144 433399 1002146
rect 433136 1002088 433338 1002144
rect 433394 1002088 433399 1002144
rect 433136 1002086 433399 1002088
rect 502412 1002144 502583 1002146
rect 502412 1002088 502522 1002144
rect 502578 1002088 502583 1002144
rect 502412 1002086 502583 1002088
rect 509680 1002144 509943 1002146
rect 509680 1002088 509882 1002144
rect 509938 1002088 509943 1002144
rect 509680 1002086 509943 1002088
rect 559820 1002144 560083 1002146
rect 559820 1002088 560022 1002144
rect 560078 1002088 560083 1002144
rect 559820 1002086 560083 1002088
rect 425513 1002083 425579 1002086
rect 427537 1002083 427603 1002086
rect 433333 1002083 433399 1002086
rect 502517 1002083 502583 1002086
rect 509877 1002083 509943 1002086
rect 560017 1002083 560083 1002086
rect 98269 1002010 98335 1002013
rect 98072 1002008 98335 1002010
rect 98072 1001952 98274 1002008
rect 98330 1001952 98335 1002008
rect 98072 1001950 98335 1001952
rect 98269 1001947 98335 1001950
rect 101121 1002010 101187 1002013
rect 103145 1002010 103211 1002013
rect 103973 1002010 104039 1002013
rect 101121 1002008 101292 1002010
rect 101121 1001952 101126 1002008
rect 101182 1001952 101292 1002008
rect 101121 1001950 101292 1001952
rect 102948 1002008 103211 1002010
rect 102948 1001952 103150 1002008
rect 103206 1001952 103211 1002008
rect 102948 1001950 103211 1001952
rect 103776 1002008 104039 1002010
rect 103776 1001952 103978 1002008
rect 104034 1001952 104039 1002008
rect 103776 1001950 104039 1001952
rect 101121 1001947 101187 1001950
rect 103145 1001947 103211 1001950
rect 103973 1001947 104039 1001950
rect 105997 1002010 106063 1002013
rect 108849 1002010 108915 1002013
rect 105997 1002008 106260 1002010
rect 105997 1001952 106002 1002008
rect 106058 1001952 106260 1002008
rect 105997 1001950 106260 1001952
rect 108652 1002008 108915 1002010
rect 108652 1001952 108854 1002008
rect 108910 1001952 108915 1002008
rect 108652 1001950 108915 1001952
rect 105997 1001947 106063 1001950
rect 108849 1001947 108915 1001950
rect 149237 1002010 149303 1002013
rect 154573 1002010 154639 1002013
rect 154941 1002010 155007 1002013
rect 157793 1002010 157859 1002013
rect 149237 1002008 149500 1002010
rect 149237 1001952 149242 1002008
rect 149298 1001952 149500 1002008
rect 149237 1001950 149500 1001952
rect 154573 1002008 154836 1002010
rect 154573 1001952 154578 1002008
rect 154634 1001952 154836 1002008
rect 154573 1001950 154836 1001952
rect 154941 1002008 155204 1002010
rect 154941 1001952 154946 1002008
rect 155002 1001952 155204 1002008
rect 154941 1001950 155204 1001952
rect 157596 1002008 157859 1002010
rect 157596 1001952 157798 1002008
rect 157854 1001952 157859 1002008
rect 157596 1001950 157859 1001952
rect 149237 1001947 149303 1001950
rect 154573 1001947 154639 1001950
rect 154941 1001947 155007 1001950
rect 157793 1001947 157859 1001950
rect 205541 1002010 205607 1002013
rect 206737 1002010 206803 1002013
rect 212073 1002010 212139 1002013
rect 205541 1002008 205804 1002010
rect 205541 1001952 205546 1002008
rect 205602 1001952 205804 1002008
rect 205541 1001950 205804 1001952
rect 206540 1002008 206803 1002010
rect 206540 1001952 206742 1002008
rect 206798 1001952 206803 1002008
rect 206540 1001950 206803 1001952
rect 211876 1002008 212139 1002010
rect 211876 1001952 212078 1002008
rect 212134 1001952 212139 1002008
rect 211876 1001950 212139 1001952
rect 205541 1001947 205607 1001950
rect 206737 1001947 206803 1001950
rect 212073 1001947 212139 1001950
rect 255313 1002010 255379 1002013
rect 263501 1002010 263567 1002013
rect 255313 1002008 255576 1002010
rect 255313 1001952 255318 1002008
rect 255374 1001952 255576 1002008
rect 255313 1001950 255576 1001952
rect 263304 1002008 263567 1002010
rect 263304 1001952 263506 1002008
rect 263562 1001952 263567 1002008
rect 263304 1001950 263567 1001952
rect 255313 1001947 255379 1001950
rect 263501 1001947 263567 1001950
rect 310973 1002010 311039 1002013
rect 354029 1002010 354095 1002013
rect 359365 1002010 359431 1002013
rect 310973 1002008 311236 1002010
rect 310973 1001952 310978 1002008
rect 311034 1001952 311236 1002008
rect 310973 1001950 311236 1001952
rect 354029 1002008 354292 1002010
rect 354029 1001952 354034 1002008
rect 354090 1001952 354292 1002008
rect 354029 1001950 354292 1001952
rect 359168 1002008 359431 1002010
rect 359168 1001952 359370 1002008
rect 359426 1001952 359431 1002008
rect 359168 1001950 359431 1001952
rect 310973 1001947 311039 1001950
rect 354029 1001947 354095 1001950
rect 359365 1001947 359431 1001950
rect 365069 1002010 365135 1002013
rect 421465 1002010 421531 1002013
rect 424317 1002010 424383 1002013
rect 425145 1002010 425211 1002013
rect 426341 1002010 426407 1002013
rect 429193 1002010 429259 1002013
rect 432873 1002010 432939 1002013
rect 365069 1002008 365332 1002010
rect 365069 1001952 365074 1002008
rect 365130 1001952 365332 1002008
rect 365069 1001950 365332 1001952
rect 421465 1002008 421636 1002010
rect 421465 1001952 421470 1002008
rect 421526 1001952 421636 1002008
rect 421465 1001950 421636 1001952
rect 424120 1002008 424383 1002010
rect 424120 1001952 424322 1002008
rect 424378 1001952 424383 1002008
rect 424120 1001950 424383 1001952
rect 424948 1002008 425211 1002010
rect 424948 1001952 425150 1002008
rect 425206 1001952 425211 1002008
rect 424948 1001950 425211 1001952
rect 426144 1002008 426407 1002010
rect 426144 1001952 426346 1002008
rect 426402 1001952 426407 1002008
rect 426144 1001950 426407 1001952
rect 428996 1002008 429259 1002010
rect 428996 1001952 429198 1002008
rect 429254 1001952 429259 1002008
rect 428996 1001950 429259 1001952
rect 432676 1002008 432939 1002010
rect 432676 1001952 432878 1002008
rect 432934 1001952 432939 1002008
rect 432676 1001950 432939 1001952
rect 365069 1001947 365135 1001950
rect 421465 1001947 421531 1001950
rect 424317 1001947 424383 1001950
rect 425145 1001947 425211 1001950
rect 426341 1001947 426407 1001950
rect 429193 1001947 429259 1001950
rect 432873 1001947 432939 1001950
rect 498469 1002010 498535 1002013
rect 501689 1002010 501755 1002013
rect 503345 1002010 503411 1002013
rect 498469 1002008 498732 1002010
rect 498469 1001952 498474 1002008
rect 498530 1001952 498732 1002008
rect 498469 1001950 498732 1001952
rect 501492 1002008 501755 1002010
rect 501492 1001952 501694 1002008
rect 501750 1001952 501755 1002008
rect 501492 1001950 501755 1001952
rect 503148 1002008 503411 1002010
rect 503148 1001952 503350 1002008
rect 503406 1001952 503411 1002008
rect 503148 1001950 503411 1001952
rect 498469 1001947 498535 1001950
rect 501689 1001947 501755 1001950
rect 503345 1001947 503411 1001950
rect 506197 1002010 506263 1002013
rect 510337 1002010 510403 1002013
rect 506197 1002008 506460 1002010
rect 506197 1001952 506202 1002008
rect 506258 1001952 506460 1002008
rect 506197 1001950 506460 1001952
rect 510140 1002008 510403 1002010
rect 510140 1001952 510342 1002008
rect 510398 1001952 510403 1002008
rect 510140 1001950 510403 1001952
rect 506197 1001947 506263 1001950
rect 510337 1001947 510403 1001950
rect 553945 1002010 554011 1002013
rect 554773 1002010 554839 1002013
rect 558821 1002010 558887 1002013
rect 561673 1002010 561739 1002013
rect 553945 1002008 554116 1002010
rect 553945 1001952 553950 1002008
rect 554006 1001952 554116 1002008
rect 553945 1001950 554116 1001952
rect 554773 1002008 555036 1002010
rect 554773 1001952 554778 1002008
rect 554834 1001952 555036 1002008
rect 554773 1001950 555036 1001952
rect 558624 1002008 558887 1002010
rect 558624 1001952 558826 1002008
rect 558882 1001952 558887 1002008
rect 558624 1001950 558887 1001952
rect 561476 1002008 561739 1002010
rect 561476 1001952 561678 1002008
rect 561734 1001952 561739 1002008
rect 561476 1001950 561739 1001952
rect 553945 1001947 554011 1001950
rect 554773 1001947 554839 1001950
rect 558821 1001947 558887 1001950
rect 561673 1001947 561739 1001950
rect 550265 1001194 550331 1001197
rect 550068 1001192 550331 1001194
rect 550068 1001136 550270 1001192
rect 550326 1001136 550331 1001192
rect 550068 1001134 550331 1001136
rect 550265 1001131 550331 1001134
rect 203885 998882 203951 998885
rect 203780 998880 203951 998882
rect 203780 998824 203890 998880
rect 203946 998824 203951 998880
rect 203780 998822 203951 998824
rect 203885 998819 203951 998822
rect 202689 998746 202755 998749
rect 202689 998744 202952 998746
rect 202689 998688 202694 998744
rect 202750 998688 202952 998744
rect 202689 998686 202952 998688
rect 202689 998683 202755 998686
rect 203885 998610 203951 998613
rect 308949 998610 309015 998613
rect 203885 998608 204148 998610
rect 203885 998552 203890 998608
rect 203946 998552 204148 998608
rect 203885 998550 204148 998552
rect 308752 998608 309015 998610
rect 308752 998552 308954 998608
rect 309010 998552 309015 998608
rect 308752 998550 309015 998552
rect 203885 998547 203951 998550
rect 308949 998547 309015 998550
rect 307293 998474 307359 998477
rect 552289 998474 552355 998477
rect 307293 998472 307556 998474
rect 307293 998416 307298 998472
rect 307354 998416 307556 998472
rect 307293 998414 307556 998416
rect 552092 998472 552355 998474
rect 552092 998416 552294 998472
rect 552350 998416 552355 998472
rect 552092 998414 552355 998416
rect 307293 998411 307359 998414
rect 552289 998411 552355 998414
rect 259361 998338 259427 998341
rect 259164 998336 259427 998338
rect 259164 998280 259366 998336
rect 259422 998280 259427 998336
rect 259164 998278 259427 998280
rect 259361 998275 259427 998278
rect 306097 998338 306163 998341
rect 373257 998338 373323 998341
rect 306097 998336 306360 998338
rect 306097 998280 306102 998336
rect 306158 998280 306360 998336
rect 306097 998278 306360 998280
rect 373257 998336 383670 998338
rect 373257 998280 373262 998336
rect 373318 998280 383670 998336
rect 373257 998278 383670 998280
rect 306097 998275 306163 998278
rect 373257 998275 373323 998278
rect 201861 998202 201927 998205
rect 253657 998202 253723 998205
rect 258165 998202 258231 998205
rect 201861 998200 202124 998202
rect 201861 998144 201866 998200
rect 201922 998144 202124 998200
rect 201861 998142 202124 998144
rect 253657 998200 253920 998202
rect 253657 998144 253662 998200
rect 253718 998144 253920 998200
rect 253657 998142 253920 998144
rect 257968 998200 258231 998202
rect 257968 998144 258170 998200
rect 258226 998144 258231 998200
rect 257968 998142 258231 998144
rect 201861 998139 201927 998142
rect 253657 998139 253723 998142
rect 258165 998139 258231 998142
rect 308121 998202 308187 998205
rect 308121 998200 308384 998202
rect 308121 998144 308126 998200
rect 308182 998144 308384 998200
rect 308121 998142 308384 998144
rect 308121 998139 308187 998142
rect 200665 998066 200731 998069
rect 205541 998066 205607 998069
rect 200665 998064 200836 998066
rect 200665 998008 200670 998064
rect 200726 998008 200836 998064
rect 200665 998006 200836 998008
rect 205344 998064 205607 998066
rect 205344 998008 205546 998064
rect 205602 998008 205607 998064
rect 205344 998006 205607 998008
rect 200665 998003 200731 998006
rect 205541 998003 205607 998006
rect 257337 998066 257403 998069
rect 259821 998066 259887 998069
rect 257337 998064 257600 998066
rect 257337 998008 257342 998064
rect 257398 998008 257600 998064
rect 257337 998006 257600 998008
rect 259624 998064 259887 998066
rect 259624 998008 259826 998064
rect 259882 998008 259887 998064
rect 259624 998006 259887 998008
rect 257337 998003 257403 998006
rect 259821 998003 259887 998006
rect 306925 998066 306991 998069
rect 310605 998066 310671 998069
rect 306925 998064 307188 998066
rect 306925 998008 306930 998064
rect 306986 998008 307188 998064
rect 306925 998006 307188 998008
rect 310605 998064 310868 998066
rect 310605 998008 310610 998064
rect 310666 998008 310868 998064
rect 310605 998006 310868 998008
rect 306925 998003 306991 998006
rect 310605 998003 310671 998006
rect 204713 997930 204779 997933
rect 253657 997930 253723 997933
rect 204713 997928 204976 997930
rect 204713 997872 204718 997928
rect 204774 997872 204976 997928
rect 204713 997870 204976 997872
rect 253460 997928 253723 997930
rect 253460 997872 253662 997928
rect 253718 997872 253723 997928
rect 253460 997870 253723 997872
rect 204713 997867 204779 997870
rect 253657 997867 253723 997870
rect 256509 997930 256575 997933
rect 258165 997930 258231 997933
rect 260189 997930 260255 997933
rect 298093 997930 298159 997933
rect 303245 997930 303311 997933
rect 256509 997928 256772 997930
rect 256509 997872 256514 997928
rect 256570 997872 256772 997928
rect 256509 997870 256772 997872
rect 258165 997928 258428 997930
rect 258165 997872 258170 997928
rect 258226 997872 258428 997928
rect 258165 997870 258428 997872
rect 260189 997928 260452 997930
rect 260189 997872 260194 997928
rect 260250 997872 260452 997928
rect 260189 997870 260452 997872
rect 298093 997928 303311 997930
rect 298093 997872 298098 997928
rect 298154 997872 303250 997928
rect 303306 997872 303311 997928
rect 298093 997870 303311 997872
rect 256509 997867 256575 997870
rect 258165 997867 258231 997870
rect 260189 997867 260255 997870
rect 298093 997867 298159 997870
rect 303245 997867 303311 997870
rect 305269 997930 305335 997933
rect 308949 997930 309015 997933
rect 305269 997928 305532 997930
rect 305269 997872 305274 997928
rect 305330 997872 305532 997928
rect 305269 997870 305532 997872
rect 308949 997928 309212 997930
rect 308949 997872 308954 997928
rect 309010 997872 309212 997928
rect 308949 997870 309212 997872
rect 305269 997867 305335 997870
rect 308949 997867 309015 997870
rect 252461 997794 252527 997797
rect 252264 997792 252527 997794
rect 252264 997736 252466 997792
rect 252522 997736 252527 997792
rect 252264 997734 252527 997736
rect 252461 997731 252527 997734
rect 256969 997794 257035 997797
rect 258993 997794 259059 997797
rect 256969 997792 257140 997794
rect 256969 997736 256974 997792
rect 257030 997736 257140 997792
rect 256969 997734 257140 997736
rect 258796 997792 259059 997794
rect 258796 997736 258998 997792
rect 259054 997736 259059 997792
rect 258796 997734 259059 997736
rect 256969 997731 257035 997734
rect 258993 997731 259059 997734
rect 261845 997794 261911 997797
rect 307753 997794 307819 997797
rect 310605 997794 310671 997797
rect 261845 997792 262108 997794
rect 261845 997736 261850 997792
rect 261906 997736 262108 997792
rect 261845 997734 262108 997736
rect 307753 997792 307924 997794
rect 307753 997736 307758 997792
rect 307814 997736 307924 997792
rect 307753 997734 307924 997736
rect 310408 997792 310671 997794
rect 310408 997736 310610 997792
rect 310666 997736 310671 997792
rect 310408 997734 310671 997736
rect 261845 997731 261911 997734
rect 307753 997731 307819 997734
rect 310605 997731 310671 997734
rect 84510 997188 84516 997252
rect 84580 997250 84586 997252
rect 92473 997250 92539 997253
rect 84580 997248 92539 997250
rect 84580 997192 92478 997248
rect 92534 997192 92539 997248
rect 84580 997190 92539 997192
rect 84580 997188 84586 997190
rect 92473 997187 92539 997190
rect 117221 997250 117287 997253
rect 143809 997250 143875 997253
rect 117221 997248 143875 997250
rect 117221 997192 117226 997248
rect 117282 997192 143814 997248
rect 143870 997192 143875 997248
rect 117221 997190 143875 997192
rect 117221 997187 117287 997190
rect 143809 997187 143875 997190
rect 170305 997250 170371 997253
rect 200205 997250 200271 997253
rect 170305 997248 200271 997250
rect 170305 997192 170310 997248
rect 170366 997192 200210 997248
rect 200266 997192 200271 997248
rect 170305 997190 200271 997192
rect 170305 997187 170371 997190
rect 200205 997187 200271 997190
rect 245694 997188 245700 997252
rect 245764 997250 245770 997252
rect 250621 997250 250687 997253
rect 245764 997248 250687 997250
rect 245764 997192 250626 997248
rect 250682 997192 250687 997248
rect 245764 997190 250687 997192
rect 245764 997188 245770 997190
rect 250621 997187 250687 997190
rect 293534 997188 293540 997252
rect 293604 997250 293610 997252
rect 303245 997250 303311 997253
rect 293604 997248 303311 997250
rect 293604 997192 303250 997248
rect 303306 997192 303311 997248
rect 293604 997190 303311 997192
rect 293604 997188 293610 997190
rect 303245 997187 303311 997190
rect 372337 997250 372403 997253
rect 383610 997250 383670 998278
rect 467097 998202 467163 998205
rect 467097 998200 470610 998202
rect 467097 998144 467102 998200
rect 467158 998144 470610 998200
rect 467097 998142 470610 998144
rect 467097 998139 467163 998142
rect 387926 997250 387932 997252
rect 372337 997248 374010 997250
rect 372337 997192 372342 997248
rect 372398 997192 374010 997248
rect 372337 997190 374010 997192
rect 383610 997190 387932 997250
rect 372337 997187 372403 997190
rect 86534 996916 86540 996980
rect 86604 996978 86610 996980
rect 92657 996978 92723 996981
rect 86604 996976 92723 996978
rect 86604 996920 92662 996976
rect 92718 996920 92723 996976
rect 86604 996918 92723 996920
rect 86604 996916 86610 996918
rect 92657 996915 92723 996918
rect 116301 996978 116367 996981
rect 144821 996978 144887 996981
rect 116301 996976 144887 996978
rect 116301 996920 116306 996976
rect 116362 996920 144826 996976
rect 144882 996920 144887 996976
rect 116301 996918 144887 996920
rect 116301 996915 116367 996918
rect 144821 996915 144887 996918
rect 293718 996916 293724 996980
rect 293788 996978 293794 996980
rect 298737 996978 298803 996981
rect 293788 996976 298803 996978
rect 293788 996920 298742 996976
rect 298798 996920 298803 996976
rect 293788 996918 298803 996920
rect 373950 996978 374010 997190
rect 387926 997188 387932 997190
rect 387996 997188 388002 997252
rect 470550 997250 470610 998142
rect 551461 998066 551527 998069
rect 551461 998064 551724 998066
rect 551461 998008 551466 998064
rect 551522 998008 551724 998064
rect 551461 998006 551724 998008
rect 551461 998003 551527 998006
rect 553117 997930 553183 997933
rect 553117 997928 553380 997930
rect 553117 997872 553122 997928
rect 553178 997872 553380 997928
rect 553117 997870 553380 997872
rect 553117 997867 553183 997870
rect 482686 997250 482692 997252
rect 470550 997190 482692 997250
rect 482686 997188 482692 997190
rect 482756 997188 482762 997252
rect 524045 997250 524111 997253
rect 530158 997250 530164 997252
rect 524045 997248 530164 997250
rect 524045 997192 524050 997248
rect 524106 997192 530164 997248
rect 524045 997190 530164 997192
rect 524045 997187 524111 997190
rect 530158 997188 530164 997190
rect 530228 997188 530234 997252
rect 399937 996978 400003 996981
rect 373950 996976 400003 996978
rect 373950 996920 399942 996976
rect 399998 996920 400003 996976
rect 373950 996918 400003 996920
rect 293788 996916 293794 996918
rect 298737 996915 298803 996918
rect 399937 996915 400003 996918
rect 439681 996978 439747 996981
rect 488993 996978 489059 996981
rect 439681 996976 489059 996978
rect 439681 996920 439686 996976
rect 439742 996920 488998 996976
rect 489054 996920 489059 996976
rect 439681 996918 489059 996920
rect 439681 996915 439747 996918
rect 488993 996915 489059 996918
rect 517329 996978 517395 996981
rect 540881 996978 540947 996981
rect 517329 996976 540947 996978
rect 517329 996920 517334 996976
rect 517390 996920 540886 996976
rect 540942 996920 540947 996976
rect 517329 996918 540947 996920
rect 517329 996915 517395 996918
rect 540881 996915 540947 996918
rect 590561 996978 590627 996981
rect 627126 996978 627132 996980
rect 590561 996976 627132 996978
rect 590561 996920 590566 996976
rect 590622 996920 627132 996976
rect 590561 996918 627132 996920
rect 590561 996915 590627 996918
rect 627126 996916 627132 996918
rect 627196 996916 627202 996980
rect 90214 996644 90220 996708
rect 90284 996706 90290 996708
rect 94497 996706 94563 996709
rect 90284 996704 94563 996706
rect 90284 996648 94502 996704
rect 94558 996648 94563 996704
rect 90284 996646 94563 996648
rect 90284 996644 90290 996646
rect 94497 996643 94563 996646
rect 141918 996644 141924 996708
rect 141988 996706 141994 996708
rect 143993 996706 144059 996709
rect 195421 996706 195487 996709
rect 141988 996704 144059 996706
rect 141988 996648 143998 996704
rect 144054 996648 144059 996704
rect 141988 996646 144059 996648
rect 141988 996644 141994 996646
rect 143993 996643 144059 996646
rect 190410 996704 195487 996706
rect 190410 996648 195426 996704
rect 195482 996648 195487 996704
rect 190410 996646 195487 996648
rect 87822 996372 87828 996436
rect 87892 996434 87898 996436
rect 92473 996434 92539 996437
rect 147673 996434 147739 996437
rect 87892 996432 92539 996434
rect 87892 996376 92478 996432
rect 92534 996376 92539 996432
rect 87892 996374 92539 996376
rect 87892 996372 87898 996374
rect 92473 996371 92539 996374
rect 140454 996432 147739 996434
rect 140454 996376 147678 996432
rect 147734 996376 147739 996432
rect 140454 996374 147739 996376
rect 98637 995890 98703 995893
rect 85438 995888 98703 995890
rect 85438 995832 98642 995888
rect 98698 995832 98703 995888
rect 85438 995830 98703 995832
rect 81249 995754 81315 995757
rect 85438 995754 85498 995830
rect 98637 995827 98703 995830
rect 81249 995752 85498 995754
rect 81249 995696 81254 995752
rect 81310 995696 85498 995752
rect 81249 995694 85498 995696
rect 81249 995691 81315 995694
rect 86493 995620 86559 995621
rect 87781 995620 87847 995621
rect 90173 995620 90239 995621
rect 86493 995618 86540 995620
rect 86448 995616 86540 995618
rect 86448 995560 86498 995616
rect 86448 995558 86540 995560
rect 86493 995556 86540 995558
rect 86604 995556 86610 995620
rect 87781 995618 87828 995620
rect 87736 995616 87828 995618
rect 87736 995560 87786 995616
rect 87736 995558 87828 995560
rect 87781 995556 87828 995558
rect 87892 995556 87898 995620
rect 90173 995618 90220 995620
rect 90128 995616 90220 995618
rect 90128 995560 90178 995616
rect 90128 995558 90220 995560
rect 90173 995556 90220 995558
rect 90284 995556 90290 995620
rect 86493 995555 86559 995556
rect 87781 995555 87847 995556
rect 90173 995555 90239 995556
rect 77201 995346 77267 995349
rect 101397 995346 101463 995349
rect 77201 995344 101463 995346
rect 77201 995288 77206 995344
rect 77262 995288 101402 995344
rect 101458 995288 101463 995344
rect 77201 995286 101463 995288
rect 77201 995283 77267 995286
rect 101397 995283 101463 995286
rect 84469 995076 84535 995077
rect 84469 995074 84516 995076
rect 84424 995072 84516 995074
rect 84424 995016 84474 995072
rect 84424 995014 84516 995016
rect 84469 995012 84516 995014
rect 84580 995012 84586 995076
rect 89345 995074 89411 995077
rect 104574 995074 104634 996132
rect 140454 995757 140514 996374
rect 147673 996371 147739 996374
rect 143993 996162 144059 996165
rect 140405 995752 140514 995757
rect 140405 995696 140410 995752
rect 140466 995696 140514 995752
rect 140405 995694 140514 995696
rect 140638 996160 144059 996162
rect 140638 996104 143998 996160
rect 144054 996104 144059 996160
rect 140638 996102 144059 996104
rect 140405 995691 140471 995694
rect 136265 995618 136331 995621
rect 136265 995616 140330 995618
rect 136265 995560 136270 995616
rect 136326 995584 140330 995616
rect 140638 995584 140698 996102
rect 143993 996099 144059 996102
rect 141049 995754 141115 995757
rect 143625 995754 143691 995757
rect 141049 995752 143691 995754
rect 141049 995696 141054 995752
rect 141110 995696 143630 995752
rect 143686 995696 143691 995752
rect 141049 995694 143691 995696
rect 141049 995691 141115 995694
rect 143625 995691 143691 995694
rect 136326 995560 140698 995584
rect 136265 995558 140698 995560
rect 136265 995555 136331 995558
rect 140270 995524 140698 995558
rect 155125 995618 155191 995621
rect 158486 995618 158546 996132
rect 155125 995616 158546 995618
rect 155125 995560 155130 995616
rect 155186 995560 158546 995616
rect 155125 995558 158546 995560
rect 155125 995555 155191 995558
rect 141693 995482 141759 995485
rect 141918 995482 141924 995484
rect 141693 995480 141924 995482
rect 141693 995424 141698 995480
rect 141754 995424 141924 995480
rect 141693 995422 141924 995424
rect 141693 995419 141759 995422
rect 141918 995420 141924 995422
rect 141988 995420 141994 995484
rect 126237 995346 126303 995349
rect 141509 995346 141575 995349
rect 126237 995344 141575 995346
rect 126237 995288 126242 995344
rect 126298 995288 141514 995344
rect 141570 995288 141575 995344
rect 126237 995286 141575 995288
rect 126237 995283 126303 995286
rect 141509 995283 141575 995286
rect 142061 995346 142127 995349
rect 159222 995346 159282 996132
rect 190410 996026 190470 996646
rect 195421 996643 195487 996646
rect 242014 996644 242020 996708
rect 242084 996706 242090 996708
rect 251633 996706 251699 996709
rect 242084 996704 251699 996706
rect 242084 996648 251638 996704
rect 251694 996648 251699 996704
rect 242084 996646 251699 996648
rect 242084 996644 242090 996646
rect 251633 996643 251699 996646
rect 288014 996644 288020 996708
rect 288084 996706 288090 996708
rect 383377 996706 383443 996709
rect 386638 996706 386644 996708
rect 288084 996646 293970 996706
rect 288084 996644 288090 996646
rect 195053 996434 195119 996437
rect 196801 996434 196867 996437
rect 195053 996432 196867 996434
rect 195053 996376 195058 996432
rect 195114 996376 196806 996432
rect 196862 996376 196867 996432
rect 195053 996374 196867 996376
rect 195053 996371 195119 996374
rect 196801 996371 196867 996374
rect 243854 996372 243860 996436
rect 243924 996434 243930 996436
rect 246941 996434 247007 996437
rect 293718 996434 293724 996436
rect 243924 996432 247007 996434
rect 243924 996376 246946 996432
rect 247002 996376 247007 996432
rect 243924 996374 247007 996376
rect 243924 996372 243930 996374
rect 246941 996371 247007 996374
rect 282686 996374 293724 996434
rect 203320 996102 203442 996162
rect 189950 995966 190470 996026
rect 203382 995992 203442 996102
rect 189441 995754 189507 995757
rect 189950 995754 190010 995966
rect 203290 995932 203442 995992
rect 202505 995890 202571 995893
rect 203290 995890 203350 995932
rect 202505 995888 203350 995890
rect 202505 995832 202510 995888
rect 202566 995832 203350 995888
rect 202505 995830 203350 995832
rect 202505 995827 202571 995830
rect 189441 995752 190010 995754
rect 189441 995696 189446 995752
rect 189502 995696 190010 995752
rect 189441 995694 190010 995696
rect 190453 995754 190519 995757
rect 200941 995754 201007 995757
rect 190453 995752 201007 995754
rect 190453 995696 190458 995752
rect 190514 995696 200946 995752
rect 201002 995696 201007 995752
rect 190453 995694 201007 995696
rect 189441 995691 189507 995694
rect 190453 995691 190519 995694
rect 200941 995691 201007 995694
rect 172421 995348 172487 995349
rect 172421 995346 172468 995348
rect 142061 995344 159282 995346
rect 142061 995288 142066 995344
rect 142122 995288 159282 995344
rect 142061 995286 159282 995288
rect 172376 995344 172468 995346
rect 172376 995288 172426 995344
rect 172376 995286 172468 995288
rect 142061 995283 142127 995286
rect 172421 995284 172468 995286
rect 172532 995284 172538 995348
rect 187601 995346 187667 995349
rect 203517 995346 203583 995349
rect 187601 995344 203583 995346
rect 187601 995288 187606 995344
rect 187662 995288 203522 995344
rect 203578 995288 203583 995344
rect 187601 995286 203583 995288
rect 172421 995283 172487 995284
rect 187601 995283 187667 995286
rect 203517 995283 203583 995286
rect 89345 995072 104634 995074
rect 89345 995016 89350 995072
rect 89406 995016 104634 995072
rect 89345 995014 104634 995016
rect 124857 995074 124923 995077
rect 155125 995074 155191 995077
rect 124857 995072 155191 995074
rect 124857 995016 124862 995072
rect 124918 995016 155130 995072
rect 155186 995016 155191 995072
rect 124857 995014 155191 995016
rect 84469 995011 84535 995012
rect 89345 995011 89411 995014
rect 124857 995011 124923 995014
rect 155125 995011 155191 995014
rect 184473 995074 184539 995077
rect 190361 995074 190427 995077
rect 184473 995072 190427 995074
rect 184473 995016 184478 995072
rect 184534 995016 190366 995072
rect 190422 995016 190427 995072
rect 184473 995014 190427 995016
rect 184473 995011 184539 995014
rect 190361 995011 190427 995014
rect 190545 995074 190611 995077
rect 204486 995074 204546 996132
rect 250437 996026 250503 996029
rect 243862 996024 250503 996026
rect 243862 995968 250442 996024
rect 250498 995968 250503 996024
rect 243862 995966 250503 995968
rect 240869 995754 240935 995757
rect 243862 995754 243922 995966
rect 250437 995963 250503 995966
rect 240869 995752 243922 995754
rect 240869 995696 240874 995752
rect 240930 995696 243922 995752
rect 240869 995694 243922 995696
rect 244089 995754 244155 995757
rect 246573 995754 246639 995757
rect 244089 995752 246639 995754
rect 244089 995696 244094 995752
rect 244150 995696 246578 995752
rect 246634 995696 246639 995752
rect 244089 995694 246639 995696
rect 240869 995691 240935 995694
rect 244089 995691 244155 995694
rect 246573 995691 246639 995694
rect 241973 995484 242039 995485
rect 243813 995484 243879 995485
rect 241973 995482 242020 995484
rect 241928 995480 242020 995482
rect 241928 995424 241978 995480
rect 241928 995422 242020 995424
rect 241973 995420 242020 995422
rect 242084 995420 242090 995484
rect 243813 995482 243860 995484
rect 243768 995480 243860 995482
rect 243768 995424 243818 995480
rect 243768 995422 243860 995424
rect 243813 995420 243860 995422
rect 243924 995420 243930 995484
rect 241973 995419 242039 995420
rect 243813 995419 243879 995420
rect 243997 995346 244063 995349
rect 247125 995346 247191 995349
rect 243997 995344 247191 995346
rect 243997 995288 244002 995344
rect 244058 995288 247130 995344
rect 247186 995288 247191 995344
rect 243997 995286 247191 995288
rect 243997 995283 244063 995286
rect 247125 995283 247191 995286
rect 190545 995072 204546 995074
rect 190545 995016 190550 995072
rect 190606 995016 204546 995072
rect 190545 995014 204546 995016
rect 228357 995074 228423 995077
rect 261250 995074 261310 996132
rect 282686 995757 282746 996374
rect 293718 996372 293724 996374
rect 293788 996372 293794 996436
rect 293910 996298 293970 996646
rect 383377 996704 386644 996706
rect 383377 996648 383382 996704
rect 383438 996648 386644 996704
rect 383377 996646 386644 996648
rect 383377 996643 383443 996646
rect 386638 996644 386644 996646
rect 386708 996644 386714 996708
rect 472249 996706 472315 996709
rect 476246 996706 476252 996708
rect 472249 996704 476252 996706
rect 472249 996648 472254 996704
rect 472310 996648 476252 996704
rect 472249 996646 476252 996648
rect 472249 996643 472315 996646
rect 476246 996644 476252 996646
rect 476316 996644 476322 996708
rect 516685 996706 516751 996709
rect 524045 996706 524111 996709
rect 516685 996704 524111 996706
rect 516685 996648 516690 996704
rect 516746 996648 524050 996704
rect 524106 996648 524111 996704
rect 516685 996646 524111 996648
rect 516685 996643 516751 996646
rect 524045 996643 524111 996646
rect 590561 996706 590627 996709
rect 626574 996706 626580 996708
rect 590561 996704 626580 996706
rect 590561 996648 590566 996704
rect 590622 996648 626580 996704
rect 590561 996646 626580 996648
rect 590561 996643 590627 996646
rect 626574 996644 626580 996646
rect 626644 996644 626650 996708
rect 295006 996508 295012 996572
rect 295076 996570 295082 996572
rect 299381 996570 299447 996573
rect 295076 996568 299447 996570
rect 295076 996512 299386 996568
rect 299442 996512 299447 996568
rect 295076 996510 299447 996512
rect 295076 996508 295082 996510
rect 299381 996507 299447 996510
rect 300301 996434 300367 996437
rect 299614 996432 300367 996434
rect 299614 996376 300306 996432
rect 300362 996376 300367 996432
rect 299614 996374 300367 996376
rect 299381 996298 299447 996301
rect 293910 996296 299447 996298
rect 293910 996240 299386 996296
rect 299442 996240 299447 996296
rect 293910 996238 299447 996240
rect 299381 996235 299447 996238
rect 299614 996026 299674 996374
rect 300301 996371 300367 996374
rect 372521 996434 372587 996437
rect 388110 996434 388116 996436
rect 372521 996432 388116 996434
rect 372521 996376 372526 996432
rect 372582 996376 388116 996432
rect 372521 996374 388116 996376
rect 372521 996371 372587 996374
rect 388110 996372 388116 996374
rect 388180 996372 388186 996436
rect 400121 996434 400187 996437
rect 396582 996432 400187 996434
rect 396582 996376 400126 996432
rect 400182 996376 400187 996432
rect 396582 996374 400187 996376
rect 292530 995966 299674 996026
rect 299841 996026 299907 996029
rect 301681 996026 301747 996029
rect 299841 996024 301747 996026
rect 299841 995968 299846 996024
rect 299902 995968 301686 996024
rect 301742 995968 301747 996024
rect 299841 995966 301747 995968
rect 282686 995752 282795 995757
rect 287973 995756 288039 995757
rect 287973 995754 288020 995756
rect 282686 995696 282734 995752
rect 282790 995696 282795 995752
rect 282686 995694 282795 995696
rect 287928 995752 288020 995754
rect 287928 995696 287978 995752
rect 287928 995694 288020 995696
rect 282729 995691 282795 995694
rect 287973 995692 288020 995694
rect 288084 995692 288090 995756
rect 291745 995754 291811 995757
rect 292530 995754 292590 995966
rect 299841 995963 299907 995966
rect 301681 995963 301747 995966
rect 293493 995756 293559 995757
rect 295057 995756 295123 995757
rect 293493 995754 293540 995756
rect 291745 995752 292590 995754
rect 291745 995696 291750 995752
rect 291806 995696 292590 995752
rect 291745 995694 292590 995696
rect 293448 995752 293540 995754
rect 293448 995696 293498 995752
rect 293448 995694 293540 995696
rect 287973 995691 288039 995692
rect 291745 995691 291811 995694
rect 293493 995692 293540 995694
rect 293604 995692 293610 995756
rect 295006 995692 295012 995756
rect 295076 995754 295123 995756
rect 299381 995754 299447 995757
rect 302877 995754 302943 995757
rect 295076 995752 295168 995754
rect 295118 995696 295168 995752
rect 295076 995694 295168 995696
rect 299381 995752 302943 995754
rect 299381 995696 299386 995752
rect 299442 995696 302882 995752
rect 302938 995696 302943 995752
rect 299381 995694 302943 995696
rect 295076 995692 295123 995694
rect 293493 995691 293559 995692
rect 295057 995691 295123 995692
rect 299381 995691 299447 995694
rect 302877 995691 302943 995694
rect 296161 995618 296227 995621
rect 299197 995618 299263 995621
rect 296161 995616 299263 995618
rect 296161 995560 296166 995616
rect 296222 995560 299202 995616
rect 299258 995560 299263 995616
rect 296161 995558 299263 995560
rect 296161 995555 296227 995558
rect 299197 995555 299263 995558
rect 286225 995346 286291 995349
rect 309550 995346 309610 996132
rect 286225 995344 309610 995346
rect 286225 995288 286230 995344
rect 286286 995288 309610 995344
rect 286225 995286 309610 995288
rect 286225 995283 286291 995286
rect 228357 995072 261310 995074
rect 228357 995016 228362 995072
rect 228418 995016 261310 995072
rect 228357 995014 261310 995016
rect 279417 995074 279483 995077
rect 312862 995074 312922 996132
rect 372337 996026 372403 996029
rect 372337 996024 388546 996026
rect 372337 995968 372342 996024
rect 372398 995968 388546 996024
rect 372337 995966 388546 995968
rect 372337 995963 372403 995966
rect 383193 995754 383259 995757
rect 385677 995754 385743 995757
rect 386689 995756 386755 995757
rect 383193 995752 385743 995754
rect 383193 995696 383198 995752
rect 383254 995696 385682 995752
rect 385738 995696 385743 995752
rect 383193 995694 385743 995696
rect 383193 995691 383259 995694
rect 385677 995691 385743 995694
rect 386638 995692 386644 995756
rect 386708 995754 386755 995756
rect 387885 995756 387951 995757
rect 388161 995756 388227 995757
rect 387885 995754 387932 995756
rect 386708 995752 386800 995754
rect 386750 995696 386800 995752
rect 386708 995694 386800 995696
rect 387840 995752 387932 995754
rect 387840 995696 387890 995752
rect 387840 995694 387932 995696
rect 386708 995692 386755 995694
rect 386689 995691 386755 995692
rect 387885 995692 387932 995694
rect 387996 995692 388002 995756
rect 388110 995692 388116 995756
rect 388180 995754 388227 995756
rect 388486 995754 388546 995966
rect 396582 995757 396642 996374
rect 400121 996371 400187 996374
rect 439865 996434 439931 996437
rect 474774 996434 474780 996436
rect 439865 996432 474780 996434
rect 439865 996376 439870 996432
rect 439926 996376 474780 996432
rect 439865 996374 474780 996376
rect 439865 996371 439931 996374
rect 474774 996372 474780 996374
rect 474844 996372 474850 996436
rect 494053 996434 494119 996437
rect 485638 996432 494119 996434
rect 485638 996376 494058 996432
rect 494114 996376 494119 996432
rect 485638 996374 494119 996376
rect 471237 996026 471303 996029
rect 471237 996024 477970 996026
rect 471237 995968 471242 996024
rect 471298 995968 477970 996024
rect 471237 995966 477970 995968
rect 471237 995963 471303 995966
rect 391933 995754 391999 995757
rect 388180 995752 388272 995754
rect 388222 995696 388272 995752
rect 388180 995694 388272 995696
rect 388486 995752 391999 995754
rect 388486 995696 391938 995752
rect 391994 995696 391999 995752
rect 388486 995694 391999 995696
rect 388180 995692 388227 995694
rect 387885 995691 387951 995692
rect 388161 995691 388227 995692
rect 391933 995691 391999 995694
rect 396533 995752 396642 995757
rect 416129 995754 416195 995757
rect 396533 995696 396538 995752
rect 396594 995696 396642 995752
rect 396533 995694 396642 995696
rect 398054 995752 416195 995754
rect 398054 995696 416134 995752
rect 416190 995696 416195 995752
rect 398054 995694 416195 995696
rect 396533 995691 396599 995694
rect 380893 995482 380959 995485
rect 398054 995482 398114 995694
rect 416129 995691 416195 995694
rect 472433 995754 472499 995757
rect 473997 995754 474063 995757
rect 474733 995756 474799 995757
rect 474733 995754 474780 995756
rect 472433 995752 474063 995754
rect 472433 995696 472438 995752
rect 472494 995696 474002 995752
rect 474058 995696 474063 995752
rect 472433 995694 474063 995696
rect 474688 995752 474780 995754
rect 474688 995696 474738 995752
rect 474688 995694 474780 995696
rect 472433 995691 472499 995694
rect 473997 995691 474063 995694
rect 474733 995692 474780 995694
rect 474844 995692 474850 995756
rect 476246 995692 476252 995756
rect 476316 995754 476322 995756
rect 477033 995754 477099 995757
rect 476316 995752 477099 995754
rect 476316 995696 477038 995752
rect 477094 995696 477099 995752
rect 476316 995694 477099 995696
rect 476316 995692 476322 995694
rect 474733 995691 474799 995692
rect 477033 995691 477099 995694
rect 460933 995618 460999 995621
rect 460933 995616 470610 995618
rect 460933 995560 460938 995616
rect 460994 995560 470610 995616
rect 460933 995558 470610 995560
rect 460933 995555 460999 995558
rect 415393 995482 415459 995485
rect 380893 995480 398114 995482
rect 380893 995424 380898 995480
rect 380954 995424 398114 995480
rect 380893 995422 398114 995424
rect 402930 995480 415459 995482
rect 402930 995424 415398 995480
rect 415454 995424 415459 995480
rect 402930 995422 415459 995424
rect 470550 995482 470610 995558
rect 477677 995482 477743 995485
rect 470550 995480 477743 995482
rect 470550 995424 477682 995480
rect 477738 995424 477743 995480
rect 470550 995422 477743 995424
rect 477910 995482 477970 995966
rect 485638 995757 485698 996374
rect 494053 996371 494119 996374
rect 516869 996434 516935 996437
rect 590745 996434 590811 996437
rect 627862 996434 627868 996436
rect 516869 996432 532802 996434
rect 516869 996376 516874 996432
rect 516930 996376 532802 996432
rect 516869 996374 532802 996376
rect 516869 996371 516935 996374
rect 518893 996162 518959 996165
rect 526294 996162 526300 996164
rect 518893 996160 526300 996162
rect 479926 995692 479932 995756
rect 479996 995754 480002 995756
rect 481449 995754 481515 995757
rect 482737 995756 482803 995757
rect 479996 995752 481515 995754
rect 479996 995696 481454 995752
rect 481510 995696 481515 995752
rect 479996 995694 481515 995696
rect 479996 995692 480002 995694
rect 481449 995691 481515 995694
rect 482686 995692 482692 995756
rect 482756 995754 482803 995756
rect 482756 995752 482848 995754
rect 482798 995696 482848 995752
rect 482756 995694 482848 995696
rect 485589 995752 485698 995757
rect 485589 995696 485594 995752
rect 485650 995696 485698 995752
rect 485589 995694 485698 995696
rect 487981 995754 488047 995757
rect 488901 995754 488967 995757
rect 487981 995752 488967 995754
rect 487981 995696 487986 995752
rect 488042 995696 488906 995752
rect 488962 995696 488967 995752
rect 487981 995694 488967 995696
rect 482756 995692 482803 995694
rect 482737 995691 482803 995692
rect 485589 995691 485655 995694
rect 487981 995691 488047 995694
rect 488901 995691 488967 995694
rect 502057 995618 502123 995621
rect 508086 995618 508146 996132
rect 502057 995616 508146 995618
rect 502057 995560 502062 995616
rect 502118 995560 508146 995616
rect 502057 995558 508146 995560
rect 502057 995555 502123 995558
rect 477910 995422 480270 995482
rect 380893 995419 380959 995422
rect 382273 995210 382339 995213
rect 402930 995210 402990 995422
rect 415393 995419 415459 995422
rect 477677 995419 477743 995422
rect 480210 995346 480270 995422
rect 508822 995346 508882 996132
rect 518893 996104 518898 996160
rect 518954 996104 526300 996160
rect 518893 996102 526300 996104
rect 518893 996099 518959 996102
rect 526294 996100 526300 996102
rect 526364 996100 526370 996164
rect 517145 995890 517211 995893
rect 517145 995888 524522 995890
rect 517145 995832 517150 995888
rect 517206 995832 524522 995888
rect 517145 995830 524522 995832
rect 517145 995827 517211 995830
rect 524462 995754 524522 995830
rect 525006 995828 525012 995892
rect 525076 995890 525082 995892
rect 525076 995830 525442 995890
rect 525076 995828 525082 995830
rect 524781 995754 524847 995757
rect 524462 995752 524847 995754
rect 524462 995696 524786 995752
rect 524842 995696 524847 995752
rect 524462 995694 524847 995696
rect 525382 995754 525442 995830
rect 532742 995757 532802 996374
rect 590745 996432 626274 996434
rect 590745 996376 590750 996432
rect 590806 996376 626274 996432
rect 590745 996374 626274 996376
rect 590745 996371 590811 996374
rect 626214 996298 626274 996374
rect 626766 996374 627868 996434
rect 626766 996298 626826 996374
rect 627862 996372 627868 996374
rect 627932 996372 627938 996436
rect 626214 996238 626826 996298
rect 532141 995754 532207 995757
rect 525382 995752 532207 995754
rect 525382 995696 532146 995752
rect 532202 995696 532207 995752
rect 525382 995694 532207 995696
rect 532742 995752 532851 995757
rect 532742 995696 532790 995752
rect 532846 995696 532851 995752
rect 532742 995694 532851 995696
rect 524781 995691 524847 995694
rect 532141 995691 532207 995694
rect 532785 995691 532851 995694
rect 535913 995754 535979 995757
rect 538213 995754 538279 995757
rect 535913 995752 538279 995754
rect 535913 995696 535918 995752
rect 535974 995696 538218 995752
rect 538274 995696 538279 995752
rect 535913 995694 538279 995696
rect 535913 995691 535979 995694
rect 538213 995691 538279 995694
rect 516961 995618 517027 995621
rect 516961 995616 524430 995618
rect 516961 995560 516966 995616
rect 517022 995584 524430 995616
rect 517022 995560 525258 995584
rect 516961 995558 525258 995560
rect 516961 995555 517027 995558
rect 524370 995524 525258 995558
rect 525198 995482 525258 995524
rect 529841 995482 529907 995485
rect 530209 995484 530275 995485
rect 525198 995480 529907 995482
rect 525198 995424 529846 995480
rect 529902 995424 529907 995480
rect 525198 995422 529907 995424
rect 529841 995419 529907 995422
rect 530158 995420 530164 995484
rect 530228 995482 530275 995484
rect 530228 995480 530320 995482
rect 530270 995424 530320 995480
rect 530228 995422 530320 995424
rect 530228 995420 530275 995422
rect 530209 995419 530275 995420
rect 480210 995286 508882 995346
rect 516685 995346 516751 995349
rect 525006 995346 525012 995348
rect 516685 995344 525012 995346
rect 516685 995288 516690 995344
rect 516746 995288 525012 995344
rect 516685 995286 525012 995288
rect 516685 995283 516751 995286
rect 525006 995284 525012 995286
rect 525076 995284 525082 995348
rect 382273 995208 402990 995210
rect 382273 995152 382278 995208
rect 382334 995152 402990 995208
rect 382273 995150 402990 995152
rect 382273 995147 382339 995150
rect 279417 995072 312922 995074
rect 279417 995016 279422 995072
rect 279478 995016 312922 995072
rect 279417 995014 312922 995016
rect 469857 995074 469923 995077
rect 502057 995074 502123 995077
rect 469857 995072 502123 995074
rect 469857 995016 469862 995072
rect 469918 995016 502062 995072
rect 502118 995016 502123 995072
rect 469857 995014 502123 995016
rect 190545 995011 190611 995014
rect 228357 995011 228423 995014
rect 279417 995011 279483 995014
rect 469857 995011 469923 995014
rect 502057 995011 502123 995014
rect 520917 995074 520983 995077
rect 557766 995074 557826 996132
rect 627686 996102 629770 996162
rect 622393 996026 622459 996029
rect 627686 996026 627746 996102
rect 622393 996024 627746 996026
rect 622393 995968 622398 996024
rect 622454 995968 627746 996024
rect 622393 995966 627746 995968
rect 622393 995963 622459 995966
rect 626625 995756 626691 995757
rect 627177 995756 627243 995757
rect 627913 995756 627979 995757
rect 626574 995692 626580 995756
rect 626644 995754 626691 995756
rect 626644 995752 626736 995754
rect 626686 995696 626736 995752
rect 626644 995694 626736 995696
rect 626644 995692 626691 995694
rect 627126 995692 627132 995756
rect 627196 995754 627243 995756
rect 627196 995752 627288 995754
rect 627238 995696 627288 995752
rect 627196 995694 627288 995696
rect 627196 995692 627243 995694
rect 627862 995692 627868 995756
rect 627932 995754 627979 995756
rect 629710 995754 629770 996102
rect 633985 995754 634051 995757
rect 627932 995752 628024 995754
rect 627974 995696 628024 995752
rect 627932 995694 628024 995696
rect 629710 995752 634051 995754
rect 629710 995696 633990 995752
rect 634046 995696 634051 995752
rect 629710 995694 634051 995696
rect 627932 995692 627979 995694
rect 626625 995691 626691 995692
rect 627177 995691 627243 995692
rect 627913 995691 627979 995692
rect 633985 995691 634051 995694
rect 635825 995754 635891 995757
rect 642081 995754 642147 995757
rect 635825 995752 642147 995754
rect 635825 995696 635830 995752
rect 635886 995696 642086 995752
rect 642142 995696 642147 995752
rect 635825 995694 642147 995696
rect 635825 995691 635891 995694
rect 642081 995691 642147 995694
rect 620277 995482 620343 995485
rect 631501 995482 631567 995485
rect 620277 995480 631567 995482
rect 620277 995424 620282 995480
rect 620338 995424 631506 995480
rect 631562 995424 631567 995480
rect 620277 995422 631567 995424
rect 620277 995419 620343 995422
rect 631501 995419 631567 995422
rect 520917 995072 557826 995074
rect 520917 995016 520922 995072
rect 520978 995016 557826 995072
rect 520917 995014 557826 995016
rect 590561 995074 590627 995077
rect 660573 995074 660639 995077
rect 590561 995072 660639 995074
rect 590561 995016 590566 995072
rect 590622 995016 660578 995072
rect 660634 995016 660639 995072
rect 590561 995014 660639 995016
rect 520917 995011 520983 995014
rect 590561 995011 590627 995014
rect 660573 995011 660639 995014
rect 374637 994938 374703 994941
rect 395153 994938 395219 994941
rect 374637 994936 395219 994938
rect 374637 994880 374642 994936
rect 374698 994880 395158 994936
rect 395214 994880 395219 994936
rect 374637 994878 395219 994880
rect 374637 994875 374703 994878
rect 395153 994875 395219 994878
rect 81985 994802 82051 994805
rect 97441 994802 97507 994805
rect 81985 994800 97507 994802
rect 81985 994744 81990 994800
rect 82046 994744 97446 994800
rect 97502 994744 97507 994800
rect 81985 994742 97507 994744
rect 81985 994739 82051 994742
rect 97441 994739 97507 994742
rect 129089 994802 129155 994805
rect 151077 994802 151143 994805
rect 129089 994800 151143 994802
rect 129089 994744 129094 994800
rect 129150 994744 151082 994800
rect 151138 994744 151143 994800
rect 129089 994742 151143 994744
rect 129089 994739 129155 994742
rect 151077 994739 151143 994742
rect 184841 994802 184907 994805
rect 200757 994802 200823 994805
rect 184841 994800 200823 994802
rect 184841 994744 184846 994800
rect 184902 994744 200762 994800
rect 200818 994744 200823 994800
rect 184841 994742 200823 994744
rect 184841 994739 184907 994742
rect 200757 994739 200823 994742
rect 236545 994802 236611 994805
rect 251817 994802 251883 994805
rect 236545 994800 251883 994802
rect 236545 994744 236550 994800
rect 236606 994744 251822 994800
rect 251878 994744 251883 994800
rect 236545 994742 251883 994744
rect 236545 994739 236611 994742
rect 251817 994739 251883 994742
rect 290273 994802 290339 994805
rect 307017 994802 307083 994805
rect 290273 994800 307083 994802
rect 290273 994744 290278 994800
rect 290334 994744 307022 994800
rect 307078 994744 307083 994800
rect 290273 994742 307083 994744
rect 290273 994739 290339 994742
rect 307017 994739 307083 994742
rect 469213 994802 469279 994805
rect 482277 994802 482343 994805
rect 469213 994800 482343 994802
rect 469213 994744 469218 994800
rect 469274 994744 482282 994800
rect 482338 994744 482343 994800
rect 469213 994742 482343 994744
rect 469213 994739 469279 994742
rect 482277 994739 482343 994742
rect 520181 994802 520247 994805
rect 526345 994804 526411 994805
rect 520181 994800 524430 994802
rect 520181 994744 520186 994800
rect 520242 994744 524430 994800
rect 520181 994742 524430 994744
rect 520181 994739 520247 994742
rect 85021 994530 85087 994533
rect 97257 994530 97323 994533
rect 85021 994528 97323 994530
rect 85021 994472 85026 994528
rect 85082 994472 97262 994528
rect 97318 994472 97323 994528
rect 85021 994470 97323 994472
rect 85021 994467 85087 994470
rect 97257 994467 97323 994470
rect 137093 994530 137159 994533
rect 142061 994530 142127 994533
rect 137093 994528 142127 994530
rect 137093 994472 137098 994528
rect 137154 994472 142066 994528
rect 142122 994472 142127 994528
rect 137093 994470 142127 994472
rect 137093 994467 137159 994470
rect 142061 994467 142127 994470
rect 142286 994468 142292 994532
rect 142356 994530 142362 994532
rect 149697 994530 149763 994533
rect 142356 994528 149763 994530
rect 142356 994472 149702 994528
rect 149758 994472 149763 994528
rect 142356 994470 149763 994472
rect 142356 994468 142362 994470
rect 149697 994467 149763 994470
rect 188153 994530 188219 994533
rect 197997 994530 198063 994533
rect 188153 994528 198063 994530
rect 188153 994472 188158 994528
rect 188214 994472 198002 994528
rect 198058 994472 198063 994528
rect 188153 994470 198063 994472
rect 188153 994467 188219 994470
rect 197997 994467 198063 994470
rect 239581 994530 239647 994533
rect 246941 994530 247007 994533
rect 239581 994528 247007 994530
rect 239581 994472 239586 994528
rect 239642 994472 246946 994528
rect 247002 994472 247007 994528
rect 239581 994470 247007 994472
rect 239581 994467 239647 994470
rect 246941 994467 247007 994470
rect 458817 994530 458883 994533
rect 524370 994530 524430 994742
rect 526294 994740 526300 994804
rect 526364 994802 526411 994804
rect 536741 994804 536807 994805
rect 526364 994800 526456 994802
rect 526406 994744 526456 994800
rect 526364 994742 526456 994744
rect 536741 994800 536788 994804
rect 536852 994802 536858 994804
rect 570781 994802 570847 994805
rect 634537 994802 634603 994805
rect 536741 994744 536746 994800
rect 526364 994740 526411 994742
rect 526345 994739 526411 994740
rect 536741 994740 536788 994744
rect 536852 994742 536898 994802
rect 570781 994800 634603 994802
rect 570781 994744 570786 994800
rect 570842 994744 634542 994800
rect 634598 994744 634603 994800
rect 570781 994742 634603 994744
rect 536852 994740 536858 994742
rect 536741 994739 536807 994740
rect 570781 994739 570847 994742
rect 634537 994739 634603 994742
rect 538029 994530 538095 994533
rect 458817 994528 480270 994530
rect 458817 994472 458822 994528
rect 458878 994472 480270 994528
rect 458817 994470 480270 994472
rect 524370 994528 538095 994530
rect 524370 994472 538034 994528
rect 538090 994472 538095 994528
rect 524370 994470 538095 994472
rect 458817 994467 458883 994470
rect 85665 994258 85731 994261
rect 95141 994258 95207 994261
rect 85665 994256 95207 994258
rect 85665 994200 85670 994256
rect 85726 994200 95146 994256
rect 95202 994200 95207 994256
rect 85665 994198 95207 994200
rect 85665 994195 85731 994198
rect 95141 994195 95207 994198
rect 132769 994258 132835 994261
rect 149881 994258 149947 994261
rect 132769 994256 149947 994258
rect 132769 994200 132774 994256
rect 132830 994200 149886 994256
rect 149942 994200 149947 994256
rect 132769 994198 149947 994200
rect 132769 994195 132835 994198
rect 149881 994195 149947 994198
rect 189073 994258 189139 994261
rect 196617 994258 196683 994261
rect 189073 994256 196683 994258
rect 189073 994200 189078 994256
rect 189134 994200 196622 994256
rect 196678 994200 196683 994256
rect 189073 994198 196683 994200
rect 189073 994195 189139 994198
rect 196617 994195 196683 994198
rect 238661 994258 238727 994261
rect 254761 994258 254827 994261
rect 238661 994256 254827 994258
rect 238661 994200 238666 994256
rect 238722 994200 254766 994256
rect 254822 994200 254827 994256
rect 238661 994198 254827 994200
rect 238661 994195 238727 994198
rect 254761 994195 254827 994198
rect 290825 994258 290891 994261
rect 300117 994258 300183 994261
rect 290825 994256 300183 994258
rect 290825 994200 290830 994256
rect 290886 994200 300122 994256
rect 300178 994200 300183 994256
rect 290825 994198 300183 994200
rect 290825 994195 290891 994198
rect 300117 994195 300183 994198
rect 471881 994258 471947 994261
rect 476757 994258 476823 994261
rect 471881 994256 476823 994258
rect 471881 994200 471886 994256
rect 471942 994200 476762 994256
rect 476818 994200 476823 994256
rect 471881 994198 476823 994200
rect 471881 994195 471947 994198
rect 476757 994195 476823 994198
rect 139393 993986 139459 993989
rect 142102 993986 142108 993988
rect 139393 993984 142108 993986
rect 139393 993928 139398 993984
rect 139454 993928 142108 993984
rect 139393 993926 142108 993928
rect 139393 993923 139459 993926
rect 142102 993924 142108 993926
rect 142172 993924 142178 993988
rect 142337 993986 142403 993989
rect 145557 993986 145623 993989
rect 142337 993984 145623 993986
rect 142337 993928 142342 993984
rect 142398 993928 145562 993984
rect 145618 993928 145623 993984
rect 142337 993926 145623 993928
rect 142337 993923 142403 993926
rect 145557 993923 145623 993926
rect 240041 993986 240107 993989
rect 249057 993986 249123 993989
rect 240041 993984 249123 993986
rect 240041 993928 240046 993984
rect 240102 993928 249062 993984
rect 249118 993928 249123 993984
rect 240041 993926 249123 993928
rect 240041 993923 240107 993926
rect 249057 993923 249123 993926
rect 468477 993986 468543 993989
rect 479926 993986 479932 993988
rect 468477 993984 479932 993986
rect 468477 993928 468482 993984
rect 468538 993928 479932 993984
rect 468477 993926 479932 993928
rect 468477 993923 468543 993926
rect 479926 993924 479932 993926
rect 479996 993924 480002 993988
rect 480210 993986 480270 994470
rect 538029 994467 538095 994470
rect 481081 993986 481147 993989
rect 480210 993984 481147 993986
rect 480210 993928 481086 993984
rect 481142 993928 481147 993984
rect 480210 993926 481147 993928
rect 481081 993923 481147 993926
rect 133873 993714 133939 993717
rect 142061 993714 142127 993717
rect 133873 993712 142127 993714
rect 133873 993656 133878 993712
rect 133934 993656 142066 993712
rect 142122 993656 142127 993712
rect 133873 993654 142127 993656
rect 133873 993651 133939 993654
rect 142061 993651 142127 993654
rect 142245 993714 142311 993717
rect 144361 993714 144427 993717
rect 142245 993712 144427 993714
rect 142245 993656 142250 993712
rect 142306 993656 144366 993712
rect 144422 993656 144427 993712
rect 142245 993654 144427 993656
rect 142245 993651 142311 993654
rect 144361 993651 144427 993654
rect 183829 993578 183895 993581
rect 202137 993578 202203 993581
rect 183829 993576 202203 993578
rect 183829 993520 183834 993576
rect 183890 993520 202142 993576
rect 202198 993520 202203 993576
rect 183829 993518 202203 993520
rect 183829 993515 183895 993518
rect 202137 993515 202203 993518
rect 191833 992898 191899 992901
rect 251449 992898 251515 992901
rect 191833 992896 251515 992898
rect 191833 992840 191838 992896
rect 191894 992840 251454 992896
rect 251510 992840 251515 992896
rect 191833 992838 251515 992840
rect 191833 992835 191899 992838
rect 251449 992835 251515 992838
rect 572662 990932 572668 990996
rect 572732 990994 572738 990996
rect 576301 990994 576367 990997
rect 572732 990992 576367 990994
rect 572732 990936 576306 990992
rect 576362 990936 576367 990992
rect 572732 990934 576367 990936
rect 572732 990932 572738 990934
rect 576301 990931 576367 990934
rect 62113 976034 62179 976037
rect 62113 976032 64492 976034
rect 62113 975976 62118 976032
rect 62174 975976 64492 976032
rect 62113 975974 64492 975976
rect 62113 975971 62179 975974
rect 651649 975898 651715 975901
rect 650164 975896 651715 975898
rect 650164 975840 651654 975896
rect 651710 975840 651715 975896
rect 650164 975838 651715 975840
rect 651649 975835 651715 975838
rect 42149 968826 42215 968829
rect 44541 968826 44607 968829
rect 42149 968824 44607 968826
rect 42149 968768 42154 968824
rect 42210 968768 44546 968824
rect 44602 968768 44607 968824
rect 42149 968766 44607 968768
rect 42149 968763 42215 968766
rect 44541 968763 44607 968766
rect 42149 967602 42215 967605
rect 42793 967602 42859 967605
rect 42149 967600 42859 967602
rect 42149 967544 42154 967600
rect 42210 967544 42798 967600
rect 42854 967544 42859 967600
rect 42149 967542 42859 967544
rect 42149 967539 42215 967542
rect 42793 967539 42859 967542
rect 41965 967196 42031 967197
rect 41965 967192 42012 967196
rect 42076 967194 42082 967196
rect 41965 967136 41970 967192
rect 41965 967132 42012 967136
rect 42076 967134 42122 967194
rect 42076 967132 42082 967134
rect 41965 967131 42031 967132
rect 42425 966786 42491 966789
rect 43437 966786 43503 966789
rect 42425 966784 43503 966786
rect 42425 966728 42430 966784
rect 42486 966728 43442 966784
rect 43498 966728 43503 966784
rect 42425 966726 43503 966728
rect 42425 966723 42491 966726
rect 43437 966723 43503 966726
rect 675385 966516 675451 966517
rect 675334 966452 675340 966516
rect 675404 966514 675451 966516
rect 675404 966512 675496 966514
rect 675446 966456 675496 966512
rect 675404 966454 675496 966456
rect 675404 966452 675451 966454
rect 675385 966451 675451 966452
rect 672993 966378 673059 966381
rect 675109 966378 675175 966381
rect 672993 966376 675175 966378
rect 672993 966320 672998 966376
rect 673054 966320 675114 966376
rect 675170 966320 675175 966376
rect 672993 966318 675175 966320
rect 672993 966315 673059 966318
rect 675109 966315 675175 966318
rect 42425 964746 42491 964749
rect 44357 964746 44423 964749
rect 42425 964744 44423 964746
rect 42425 964688 42430 964744
rect 42486 964688 44362 964744
rect 44418 964688 44423 964744
rect 42425 964686 44423 964688
rect 42425 964683 42491 964686
rect 44357 964683 44423 964686
rect 675293 964746 675359 964749
rect 676806 964746 676812 964748
rect 675293 964744 676812 964746
rect 675293 964688 675298 964744
rect 675354 964688 676812 964744
rect 675293 964686 676812 964688
rect 675293 964683 675359 964686
rect 676806 964684 676812 964686
rect 676876 964684 676882 964748
rect 42425 963930 42491 963933
rect 44173 963930 44239 963933
rect 42425 963928 44239 963930
rect 42425 963872 42430 963928
rect 42486 963872 44178 963928
rect 44234 963872 44239 963928
rect 42425 963870 44239 963872
rect 42425 963867 42491 963870
rect 44173 963867 44239 963870
rect 42425 963386 42491 963389
rect 43161 963386 43227 963389
rect 42425 963384 43227 963386
rect 42425 963328 42430 963384
rect 42486 963328 43166 963384
rect 43222 963328 43227 963384
rect 42425 963326 43227 963328
rect 42425 963323 42491 963326
rect 43161 963323 43227 963326
rect 675753 963386 675819 963389
rect 676070 963386 676076 963388
rect 675753 963384 676076 963386
rect 675753 963328 675758 963384
rect 675814 963328 676076 963384
rect 675753 963326 676076 963328
rect 675753 963323 675819 963326
rect 676070 963324 676076 963326
rect 676140 963324 676146 963388
rect 42425 963114 42491 963117
rect 42977 963114 43043 963117
rect 42425 963112 43043 963114
rect 42425 963056 42430 963112
rect 42486 963056 42982 963112
rect 43038 963056 43043 963112
rect 42425 963054 43043 963056
rect 42425 963051 42491 963054
rect 42977 963051 43043 963054
rect 62113 962978 62179 962981
rect 62113 962976 64492 962978
rect 62113 962920 62118 962976
rect 62174 962920 64492 962976
rect 62113 962918 64492 962920
rect 62113 962915 62179 962918
rect 674373 962842 674439 962845
rect 675477 962842 675543 962845
rect 674373 962840 675543 962842
rect 674373 962784 674378 962840
rect 674434 962784 675482 962840
rect 675538 962784 675543 962840
rect 674373 962782 675543 962784
rect 674373 962779 674439 962782
rect 675477 962779 675543 962782
rect 651465 962570 651531 962573
rect 650164 962568 651531 962570
rect 650164 962512 651470 962568
rect 651526 962512 651531 962568
rect 650164 962510 651531 962512
rect 651465 962507 651531 962510
rect 41454 962100 41460 962164
rect 41524 962162 41530 962164
rect 41781 962162 41847 962165
rect 41524 962160 41847 962162
rect 41524 962104 41786 962160
rect 41842 962104 41847 962160
rect 41524 962102 41847 962104
rect 41524 962100 41530 962102
rect 41781 962099 41847 962102
rect 673177 960802 673243 960805
rect 675109 960802 675175 960805
rect 673177 960800 675175 960802
rect 673177 960744 673182 960800
rect 673238 960744 675114 960800
rect 675170 960744 675175 960800
rect 673177 960742 675175 960744
rect 673177 960739 673243 960742
rect 675109 960739 675175 960742
rect 41270 959788 41276 959852
rect 41340 959850 41346 959852
rect 41781 959850 41847 959853
rect 41340 959848 41847 959850
rect 41340 959792 41786 959848
rect 41842 959792 41847 959848
rect 41340 959790 41847 959792
rect 41340 959788 41346 959790
rect 41781 959787 41847 959790
rect 674097 959306 674163 959309
rect 675109 959306 675175 959309
rect 674097 959304 675175 959306
rect 674097 959248 674102 959304
rect 674158 959248 675114 959304
rect 675170 959248 675175 959304
rect 674097 959246 675175 959248
rect 674097 959243 674163 959246
rect 675109 959243 675175 959246
rect 40534 959108 40540 959172
rect 40604 959170 40610 959172
rect 41781 959170 41847 959173
rect 40604 959168 41847 959170
rect 40604 959112 41786 959168
rect 41842 959112 41847 959168
rect 40604 959110 41847 959112
rect 40604 959108 40610 959110
rect 41781 959107 41847 959110
rect 42425 958762 42491 958765
rect 43713 958762 43779 958765
rect 42425 958760 43779 958762
rect 42425 958704 42430 958760
rect 42486 958704 43718 958760
rect 43774 958704 43779 958760
rect 42425 958702 43779 958704
rect 42425 958699 42491 958702
rect 43713 958699 43779 958702
rect 674741 958354 674807 958357
rect 675385 958354 675451 958357
rect 674741 958352 675451 958354
rect 674741 958296 674746 958352
rect 674802 958296 675390 958352
rect 675446 958296 675451 958352
rect 674741 958294 675451 958296
rect 674741 958291 674807 958294
rect 675385 958291 675451 958294
rect 42057 957946 42123 957949
rect 42558 957946 42564 957948
rect 42057 957944 42564 957946
rect 42057 957888 42062 957944
rect 42118 957888 42564 957944
rect 42057 957886 42564 957888
rect 42057 957883 42123 957886
rect 42558 957884 42564 957886
rect 42628 957884 42634 957948
rect 661677 957810 661743 957813
rect 675201 957810 675267 957813
rect 661677 957808 675267 957810
rect 661677 957752 661682 957808
rect 661738 957752 675206 957808
rect 675262 957752 675267 957808
rect 661677 957750 675267 957752
rect 661677 957747 661743 957750
rect 675201 957747 675267 957750
rect 675753 957810 675819 957813
rect 676990 957810 676996 957812
rect 675753 957808 676996 957810
rect 675753 957752 675758 957808
rect 675814 957752 676996 957808
rect 675753 957750 676996 957752
rect 675753 957747 675819 957750
rect 676990 957748 676996 957750
rect 677060 957748 677066 957812
rect 674557 957130 674623 957133
rect 675385 957130 675451 957133
rect 674557 957128 675451 957130
rect 674557 957072 674562 957128
rect 674618 957072 675390 957128
rect 675446 957072 675451 957128
rect 674557 957070 675451 957072
rect 674557 957067 674623 957070
rect 675385 957067 675451 957070
rect 675753 956450 675819 956453
rect 676622 956450 676628 956452
rect 675753 956448 676628 956450
rect 675753 956392 675758 956448
rect 675814 956392 676628 956448
rect 675753 956390 676628 956392
rect 675753 956387 675819 956390
rect 676622 956388 676628 956390
rect 676692 956388 676698 956452
rect 40718 955436 40724 955500
rect 40788 955498 40794 955500
rect 41781 955498 41847 955501
rect 40788 955496 41847 955498
rect 40788 955440 41786 955496
rect 41842 955440 41847 955496
rect 40788 955438 41847 955440
rect 40788 955436 40794 955438
rect 41781 955435 41847 955438
rect 674833 953458 674899 953461
rect 675385 953458 675451 953461
rect 674833 953456 675451 953458
rect 674833 953400 674838 953456
rect 674894 953400 675390 953456
rect 675446 953400 675451 953456
rect 674833 953398 675451 953400
rect 674833 953395 674899 953398
rect 675385 953395 675451 953398
rect 28533 952914 28599 952917
rect 43437 952914 43503 952917
rect 28533 952912 43503 952914
rect 28533 952856 28538 952912
rect 28594 952856 43442 952912
rect 43498 952856 43503 952912
rect 28533 952854 43503 952856
rect 28533 952851 28599 952854
rect 43437 952851 43503 952854
rect 39297 952234 39363 952237
rect 41454 952234 41460 952236
rect 39297 952232 41460 952234
rect 39297 952176 39302 952232
rect 39358 952176 41460 952232
rect 39297 952174 41460 952176
rect 39297 952171 39363 952174
rect 41454 952172 41460 952174
rect 41524 952172 41530 952236
rect 672533 952234 672599 952237
rect 675385 952234 675451 952237
rect 672533 952232 675451 952234
rect 672533 952176 672538 952232
rect 672594 952176 675390 952232
rect 675446 952176 675451 952232
rect 672533 952174 675451 952176
rect 672533 952171 672599 952174
rect 675385 952171 675451 952174
rect 42057 951962 42123 951965
rect 42558 951962 42564 951964
rect 42057 951960 42564 951962
rect 42057 951904 42062 951960
rect 42118 951904 42564 951960
rect 42057 951902 42564 951904
rect 42057 951899 42123 951902
rect 42558 951900 42564 951902
rect 42628 951900 42634 951964
rect 40033 951826 40099 951829
rect 41270 951826 41276 951828
rect 40033 951824 41276 951826
rect 40033 951768 40038 951824
rect 40094 951768 41276 951824
rect 40033 951766 41276 951768
rect 40033 951763 40099 951766
rect 41270 951764 41276 951766
rect 41340 951764 41346 951828
rect 41413 951690 41479 951693
rect 42006 951690 42012 951692
rect 41413 951688 42012 951690
rect 41413 951632 41418 951688
rect 41474 951632 42012 951688
rect 41413 951630 42012 951632
rect 41413 951627 41479 951630
rect 42006 951628 42012 951630
rect 42076 951628 42082 951692
rect 675385 951556 675451 951557
rect 675334 951554 675340 951556
rect 675294 951494 675340 951554
rect 675404 951552 675451 951556
rect 675446 951496 675451 951552
rect 675334 951492 675340 951494
rect 675404 951492 675451 951496
rect 675385 951491 675451 951492
rect 676806 950676 676812 950740
rect 676876 950738 676882 950740
rect 683297 950738 683363 950741
rect 676876 950736 683363 950738
rect 676876 950680 683302 950736
rect 683358 950680 683363 950736
rect 676876 950678 683363 950680
rect 676876 950676 676882 950678
rect 683297 950675 683363 950678
rect 62113 949922 62179 949925
rect 62113 949920 64492 949922
rect 62113 949864 62118 949920
rect 62174 949864 64492 949920
rect 62113 949862 64492 949864
rect 62113 949859 62179 949862
rect 676070 949452 676076 949516
rect 676140 949514 676146 949516
rect 679617 949514 679683 949517
rect 676140 949512 679683 949514
rect 676140 949456 679622 949512
rect 679678 949456 679683 949512
rect 676140 949454 679683 949456
rect 676140 949452 676146 949454
rect 679617 949451 679683 949454
rect 652201 949378 652267 949381
rect 650164 949376 652267 949378
rect 650164 949320 652206 949376
rect 652262 949320 652267 949376
rect 650164 949318 652267 949320
rect 652201 949315 652267 949318
rect 672717 947338 672783 947341
rect 683113 947338 683179 947341
rect 672717 947336 683179 947338
rect 672717 947280 672722 947336
rect 672778 947280 683118 947336
rect 683174 947280 683179 947336
rect 672717 947278 683179 947280
rect 672717 947275 672783 947278
rect 683113 947275 683179 947278
rect 45553 943530 45619 943533
rect 41492 943528 45619 943530
rect 41492 943472 45558 943528
rect 45614 943472 45619 943528
rect 41492 943470 45619 943472
rect 45553 943467 45619 943470
rect 41229 943122 41295 943125
rect 41229 943120 41308 943122
rect 41229 943064 41234 943120
rect 41290 943064 41308 943120
rect 41229 943062 41308 943064
rect 41229 943059 41295 943062
rect 28533 942714 28599 942717
rect 28533 942712 28612 942714
rect 28533 942656 28538 942712
rect 28594 942656 28612 942712
rect 28533 942654 28612 942656
rect 28533 942651 28599 942654
rect 48957 942306 49023 942309
rect 41492 942304 49023 942306
rect 41492 942248 48962 942304
rect 49018 942248 49023 942304
rect 41492 942246 49023 942248
rect 48957 942243 49023 942246
rect 41229 941898 41295 941901
rect 41229 941896 41308 941898
rect 41229 941840 41234 941896
rect 41290 941840 41308 941896
rect 41229 941838 41308 941840
rect 41229 941835 41295 941838
rect 660297 941762 660363 941765
rect 676213 941762 676279 941765
rect 660297 941760 676279 941762
rect 660297 941704 660302 941760
rect 660358 941704 676218 941760
rect 676274 941704 676279 941760
rect 660297 941702 676279 941704
rect 660297 941699 660363 941702
rect 676213 941699 676279 941702
rect 44817 941490 44883 941493
rect 41492 941488 44883 941490
rect 41492 941432 44822 941488
rect 44878 941432 44883 941488
rect 41492 941430 44883 941432
rect 44817 941427 44883 941430
rect 41822 941082 41828 941084
rect 41492 941022 41828 941082
rect 41822 941020 41828 941022
rect 41892 941020 41898 941084
rect 50337 940674 50403 940677
rect 41492 940672 50403 940674
rect 41492 940616 50342 940672
rect 50398 940616 50403 940672
rect 41492 940614 50403 940616
rect 50337 940611 50403 940614
rect 43529 940266 43595 940269
rect 41492 940264 43595 940266
rect 41492 940208 43534 940264
rect 43590 940208 43595 940264
rect 41492 940206 43595 940208
rect 43529 940203 43595 940206
rect 51717 939858 51783 939861
rect 41492 939856 51783 939858
rect 41492 939800 51722 939856
rect 51778 939800 51783 939856
rect 41492 939798 51783 939800
rect 51717 939795 51783 939798
rect 665817 939858 665883 939861
rect 676262 939858 676322 939964
rect 665817 939856 676322 939858
rect 665817 939800 665822 939856
rect 665878 939800 676322 939856
rect 665817 939798 676322 939800
rect 665817 939795 665883 939798
rect 683113 939722 683179 939725
rect 683070 939720 683179 939722
rect 683070 939664 683118 939720
rect 683174 939664 683179 939720
rect 683070 939659 683179 939664
rect 683070 939556 683130 939659
rect 41137 939450 41203 939453
rect 41124 939448 41203 939450
rect 41124 939392 41142 939448
rect 41198 939392 41203 939448
rect 41124 939390 41203 939392
rect 41137 939387 41203 939390
rect 676213 939314 676279 939317
rect 676213 939312 676322 939314
rect 676213 939256 676218 939312
rect 676274 939256 676322 939312
rect 676213 939251 676322 939256
rect 676262 939148 676322 939251
rect 37917 939042 37983 939045
rect 37917 939040 37996 939042
rect 37917 938984 37922 939040
rect 37978 938984 37996 939040
rect 37917 938982 37996 938984
rect 37917 938979 37983 938982
rect 40910 938467 40970 938604
rect 669957 938498 670023 938501
rect 676262 938498 676322 938740
rect 669957 938496 676322 938498
rect 36537 938464 36603 938467
rect 36494 938462 36603 938464
rect 36494 938406 36542 938462
rect 36598 938406 36603 938462
rect 36494 938401 36603 938406
rect 40910 938462 41019 938467
rect 40910 938406 40958 938462
rect 41014 938406 41019 938462
rect 669957 938440 669962 938496
rect 670018 938440 676322 938496
rect 669957 938438 676322 938440
rect 669957 938435 670023 938438
rect 40910 938404 41019 938406
rect 40953 938401 41019 938404
rect 36494 938196 36554 938401
rect 675150 938164 675156 938228
rect 675220 938226 675226 938228
rect 676262 938226 676322 938332
rect 675220 938166 676322 938226
rect 675220 938164 675226 938166
rect 672717 938090 672783 938093
rect 672717 938088 675034 938090
rect 672717 938032 672722 938088
rect 672778 938032 675034 938088
rect 672717 938030 675034 938032
rect 672717 938027 672783 938030
rect 42057 937818 42123 937821
rect 41492 937816 42123 937818
rect 41492 937760 42062 937816
rect 42118 937760 42123 937816
rect 41492 937758 42123 937760
rect 42057 937755 42123 937758
rect 668577 937682 668643 937685
rect 674974 937682 675034 938030
rect 675201 937954 675267 937957
rect 675201 937952 676292 937954
rect 675201 937896 675206 937952
rect 675262 937896 676292 937952
rect 675201 937894 676292 937896
rect 675201 937891 675267 937894
rect 668577 937680 674850 937682
rect 668577 937624 668582 937680
rect 668638 937624 674850 937680
rect 668577 937622 674850 937624
rect 674974 937622 676322 937682
rect 668577 937619 668643 937622
rect 39297 937410 39363 937413
rect 39284 937408 39363 937410
rect 39284 937352 39302 937408
rect 39358 937352 39363 937408
rect 39284 937350 39363 937352
rect 39297 937347 39363 937350
rect 673361 937410 673427 937413
rect 674598 937410 674604 937412
rect 673361 937408 674604 937410
rect 673361 937352 673366 937408
rect 673422 937352 674604 937408
rect 673361 937350 674604 937352
rect 673361 937347 673427 937350
rect 674598 937348 674604 937350
rect 674668 937348 674674 937412
rect 40166 937178 40172 937242
rect 40236 937240 40242 937242
rect 41822 937240 41828 937276
rect 40236 937212 41828 937240
rect 41892 937212 41898 937276
rect 674790 937274 674850 937622
rect 676262 937516 676322 937622
rect 674790 937214 676322 937274
rect 40236 937180 41890 937212
rect 40236 937178 40242 937180
rect 667197 937138 667263 937141
rect 667197 937136 673470 937138
rect 667197 937080 667202 937136
rect 667258 937080 673470 937136
rect 676262 937108 676322 937214
rect 667197 937078 673470 937080
rect 667197 937075 667263 937078
rect 44541 937002 44607 937005
rect 41492 937000 44607 937002
rect 41492 936944 44546 937000
rect 44602 936944 44607 937000
rect 41492 936942 44607 936944
rect 673410 937002 673470 937078
rect 675201 937002 675267 937005
rect 673410 937000 675267 937002
rect 673410 936944 675206 937000
rect 675262 936944 675267 937000
rect 673410 936942 675267 936944
rect 44541 936939 44607 936942
rect 675201 936939 675267 936942
rect 41822 936594 41828 936596
rect 41492 936534 41828 936594
rect 41822 936532 41828 936534
rect 41892 936532 41898 936596
rect 43713 936186 43779 936189
rect 41492 936184 43779 936186
rect 41492 936128 43718 936184
rect 43774 936128 43779 936184
rect 41492 936126 43779 936128
rect 43713 936123 43779 936126
rect 41822 935778 41828 935780
rect 41492 935718 41828 935778
rect 41822 935716 41828 935718
rect 41892 935716 41898 935780
rect 42057 935778 42123 935781
rect 64462 935778 64522 936836
rect 670969 936458 671035 936461
rect 676262 936458 676322 936700
rect 670969 936456 676322 936458
rect 670969 936400 670974 936456
rect 671030 936400 676322 936456
rect 670969 936398 676322 936400
rect 670969 936395 671035 936398
rect 651465 936186 651531 936189
rect 650164 936184 651531 936186
rect 650164 936128 651470 936184
rect 651526 936128 651531 936184
rect 650164 936126 651531 936128
rect 651465 936123 651531 936126
rect 658917 936050 658983 936053
rect 676262 936050 676322 936292
rect 658917 936048 676322 936050
rect 658917 935992 658922 936048
rect 658978 935992 676322 936048
rect 658917 935990 676322 935992
rect 658917 935987 658983 935990
rect 42057 935776 64522 935778
rect 42057 935720 42062 935776
rect 42118 935720 64522 935776
rect 42057 935718 64522 935720
rect 671981 935778 672047 935781
rect 676262 935778 676322 935884
rect 671981 935776 676322 935778
rect 671981 935720 671986 935776
rect 672042 935720 676322 935776
rect 671981 935718 676322 935720
rect 42057 935715 42123 935718
rect 671981 935715 672047 935718
rect 675385 935506 675451 935509
rect 675385 935504 676292 935506
rect 675385 935448 675390 935504
rect 675446 935448 676292 935504
rect 675385 935446 676292 935448
rect 675385 935443 675451 935446
rect 44357 935370 44423 935373
rect 41492 935368 44423 935370
rect 41492 935312 44362 935368
rect 44418 935312 44423 935368
rect 41492 935310 44423 935312
rect 44357 935307 44423 935310
rect 682377 935234 682443 935237
rect 682334 935232 682443 935234
rect 682334 935176 682382 935232
rect 682438 935176 682443 935232
rect 682334 935171 682443 935176
rect 682334 935068 682394 935171
rect 43161 934962 43227 934965
rect 41492 934960 43227 934962
rect 41492 934904 43166 934960
rect 43222 934904 43227 934960
rect 41492 934902 43227 934904
rect 43161 934899 43227 934902
rect 675569 934690 675635 934693
rect 675569 934688 676292 934690
rect 675569 934632 675574 934688
rect 675630 934632 676292 934688
rect 675569 934630 676292 934632
rect 675569 934627 675635 934630
rect 40033 934554 40099 934557
rect 40020 934552 40099 934554
rect 40020 934496 40038 934552
rect 40094 934496 40099 934552
rect 40020 934494 40099 934496
rect 40033 934491 40099 934494
rect 679617 934418 679683 934421
rect 679574 934416 679683 934418
rect 679574 934360 679622 934416
rect 679678 934360 679683 934416
rect 679574 934355 679683 934360
rect 679574 934252 679634 934355
rect 42977 934146 43043 934149
rect 41492 934144 43043 934146
rect 41492 934088 42982 934144
rect 43038 934088 43043 934144
rect 41492 934086 43043 934088
rect 42977 934083 43043 934086
rect 674097 933874 674163 933877
rect 674097 933872 676292 933874
rect 674097 933816 674102 933872
rect 674158 933816 676292 933872
rect 674097 933814 676292 933816
rect 674097 933811 674163 933814
rect 44173 933738 44239 933741
rect 41492 933736 44239 933738
rect 41492 933680 44178 933736
rect 44234 933680 44239 933736
rect 41492 933678 44239 933680
rect 44173 933675 44239 933678
rect 46933 933330 46999 933333
rect 41492 933328 46999 933330
rect 41492 933272 46938 933328
rect 46994 933272 46999 933328
rect 41492 933270 46999 933272
rect 46933 933267 46999 933270
rect 672533 933194 672599 933197
rect 676262 933194 676322 933436
rect 672533 933192 676322 933194
rect 672533 933136 672538 933192
rect 672594 933136 676322 933192
rect 672533 933134 676322 933136
rect 672533 933131 672599 933134
rect 42241 932922 42307 932925
rect 41492 932920 42307 932922
rect 41492 932864 42246 932920
rect 42302 932864 42307 932920
rect 41492 932862 42307 932864
rect 42241 932859 42307 932862
rect 672993 932922 673059 932925
rect 676262 932922 676322 933028
rect 672993 932920 676322 932922
rect 672993 932864 672998 932920
rect 673054 932864 676322 932920
rect 672993 932862 676322 932864
rect 672993 932859 673059 932862
rect 674281 932650 674347 932653
rect 674281 932648 676292 932650
rect 674281 932592 674286 932648
rect 674342 932592 676292 932648
rect 674281 932590 676292 932592
rect 674281 932587 674347 932590
rect 683297 932378 683363 932381
rect 683254 932376 683363 932378
rect 683254 932320 683302 932376
rect 683358 932320 683363 932376
rect 683254 932315 683363 932320
rect 683254 932212 683314 932315
rect 43345 932106 43411 932109
rect 41492 932104 43411 932106
rect 41492 932048 43350 932104
rect 43406 932048 43411 932104
rect 41492 932046 43411 932048
rect 43345 932043 43411 932046
rect 676622 931908 676628 931972
rect 676692 931908 676698 931972
rect 676630 931804 676690 931908
rect 676990 931500 676996 931564
rect 677060 931500 677066 931564
rect 676998 931396 677058 931500
rect 673177 930746 673243 930749
rect 676262 930746 676322 930988
rect 673177 930744 676322 930746
rect 673177 930688 673182 930744
rect 673238 930688 676322 930744
rect 673177 930686 676322 930688
rect 673177 930683 673243 930686
rect 674649 930474 674715 930477
rect 676262 930474 676322 930580
rect 674649 930472 676322 930474
rect 674649 930416 674654 930472
rect 674710 930416 676322 930472
rect 674649 930414 676322 930416
rect 674649 930411 674715 930414
rect 674465 930202 674531 930205
rect 674465 930200 676292 930202
rect 674465 930144 674470 930200
rect 674526 930144 676292 930200
rect 674465 930142 676292 930144
rect 674465 930139 674531 930142
rect 669221 929522 669287 929525
rect 676262 929522 676322 929764
rect 669221 929520 676322 929522
rect 669221 929464 669226 929520
rect 669282 929464 676322 929520
rect 669221 929462 676322 929464
rect 669221 929459 669287 929462
rect 682886 929114 682946 929356
rect 683113 929114 683179 929117
rect 682886 929112 683179 929114
rect 682886 929056 683118 929112
rect 683174 929056 683179 929112
rect 682886 929054 683179 929056
rect 682886 928948 682946 929054
rect 683113 929051 683179 929054
rect 670601 928298 670667 928301
rect 676262 928298 676322 928540
rect 670601 928296 676322 928298
rect 670601 928240 670606 928296
rect 670662 928240 676322 928296
rect 670601 928238 676322 928240
rect 670601 928235 670667 928238
rect 62113 923810 62179 923813
rect 62113 923808 64492 923810
rect 62113 923752 62118 923808
rect 62174 923752 64492 923808
rect 62113 923750 64492 923752
rect 62113 923747 62179 923750
rect 651465 922722 651531 922725
rect 650164 922720 651531 922722
rect 650164 922664 651470 922720
rect 651526 922664 651531 922720
rect 650164 922662 651531 922664
rect 651465 922659 651531 922662
rect 41689 911978 41755 911981
rect 42006 911978 42012 911980
rect 41689 911976 42012 911978
rect 41689 911920 41694 911976
rect 41750 911920 42012 911976
rect 41689 911918 42012 911920
rect 41689 911915 41755 911918
rect 42006 911916 42012 911918
rect 42076 911916 42082 911980
rect 41505 911706 41571 911709
rect 42190 911706 42196 911708
rect 41505 911704 42196 911706
rect 41505 911648 41510 911704
rect 41566 911648 42196 911704
rect 41505 911646 42196 911648
rect 41505 911643 41571 911646
rect 42190 911644 42196 911646
rect 42260 911644 42266 911708
rect 62113 910754 62179 910757
rect 62113 910752 64492 910754
rect 62113 910696 62118 910752
rect 62174 910696 64492 910752
rect 62113 910694 64492 910696
rect 62113 910691 62179 910694
rect 652385 909530 652451 909533
rect 650164 909528 652451 909530
rect 650164 909472 652390 909528
rect 652446 909472 652451 909528
rect 650164 909470 652451 909472
rect 652385 909467 652451 909470
rect 62113 897834 62179 897837
rect 62113 897832 64492 897834
rect 62113 897776 62118 897832
rect 62174 897776 64492 897832
rect 62113 897774 64492 897776
rect 62113 897771 62179 897774
rect 651465 896202 651531 896205
rect 650164 896200 651531 896202
rect 650164 896144 651470 896200
rect 651526 896144 651531 896200
rect 650164 896142 651531 896144
rect 651465 896139 651531 896142
rect 44081 892802 44147 892805
rect 55857 892802 55923 892805
rect 44081 892800 55923 892802
rect 44081 892744 44086 892800
rect 44142 892744 55862 892800
rect 55918 892744 55923 892800
rect 44081 892742 55923 892744
rect 44081 892739 44147 892742
rect 55857 892739 55923 892742
rect 42931 892530 42997 892533
rect 54477 892530 54543 892533
rect 42931 892528 54543 892530
rect 42931 892472 42936 892528
rect 42992 892472 54482 892528
rect 54538 892472 54543 892528
rect 42931 892470 54543 892472
rect 42931 892467 42997 892470
rect 54477 892467 54543 892470
rect 44081 892258 44147 892261
rect 53281 892258 53347 892261
rect 44081 892256 53347 892258
rect 44081 892200 44086 892256
rect 44142 892200 53286 892256
rect 53342 892200 53347 892256
rect 44081 892198 53347 892200
rect 44081 892195 44147 892198
rect 53281 892195 53347 892198
rect 43069 891986 43135 891989
rect 47577 891986 47643 891989
rect 43069 891984 47643 891986
rect 43069 891928 43074 891984
rect 43130 891928 47582 891984
rect 47638 891928 47643 891984
rect 43069 891926 47643 891928
rect 43069 891923 43135 891926
rect 47577 891923 47643 891926
rect 41597 885458 41663 885461
rect 42006 885458 42012 885460
rect 41597 885456 42012 885458
rect 41597 885400 41602 885456
rect 41658 885400 42012 885456
rect 41597 885398 42012 885400
rect 41597 885395 41663 885398
rect 42006 885396 42012 885398
rect 42076 885396 42082 885460
rect 41413 885186 41479 885189
rect 42190 885186 42196 885188
rect 41413 885184 42196 885186
rect 41413 885128 41418 885184
rect 41474 885128 42196 885184
rect 41413 885126 42196 885128
rect 41413 885123 41479 885126
rect 42190 885124 42196 885126
rect 42260 885124 42266 885188
rect 45510 884718 64492 884778
rect 42057 884642 42123 884645
rect 45510 884642 45570 884718
rect 42057 884640 45570 884642
rect 42057 884584 42062 884640
rect 42118 884584 45570 884640
rect 42057 884582 45570 884584
rect 42057 884579 42123 884582
rect 651649 882874 651715 882877
rect 650164 882872 651715 882874
rect 650164 882816 651654 882872
rect 651710 882816 651715 882872
rect 650164 882814 651715 882816
rect 651649 882811 651715 882814
rect 666461 879202 666527 879205
rect 675293 879202 675359 879205
rect 666461 879200 675359 879202
rect 666461 879144 666466 879200
rect 666522 879144 675298 879200
rect 675354 879144 675359 879200
rect 666461 879142 675359 879144
rect 666461 879139 666527 879142
rect 675293 879139 675359 879142
rect 675753 876618 675819 876621
rect 676806 876618 676812 876620
rect 675753 876616 676812 876618
rect 675753 876560 675758 876616
rect 675814 876560 676812 876616
rect 675753 876558 676812 876560
rect 675753 876555 675819 876558
rect 676806 876556 676812 876558
rect 676876 876556 676882 876620
rect 668393 876346 668459 876349
rect 675109 876346 675175 876349
rect 668393 876344 675175 876346
rect 668393 876288 668398 876344
rect 668454 876288 675114 876344
rect 675170 876288 675175 876344
rect 668393 876286 675175 876288
rect 668393 876283 668459 876286
rect 675109 876283 675175 876286
rect 675753 875938 675819 875941
rect 676070 875938 676076 875940
rect 675753 875936 676076 875938
rect 675753 875880 675758 875936
rect 675814 875880 676076 875936
rect 675753 875878 676076 875880
rect 675753 875875 675819 875878
rect 676070 875876 676076 875878
rect 676140 875876 676146 875940
rect 675150 873972 675156 874036
rect 675220 874034 675226 874036
rect 675385 874034 675451 874037
rect 675220 874032 675451 874034
rect 675220 873976 675390 874032
rect 675446 873976 675451 874032
rect 675220 873974 675451 873976
rect 675220 873972 675226 873974
rect 675385 873971 675451 873974
rect 673862 873156 673868 873220
rect 673932 873218 673938 873220
rect 675109 873218 675175 873221
rect 673932 873216 675175 873218
rect 673932 873160 675114 873216
rect 675170 873160 675175 873216
rect 673932 873158 675175 873160
rect 673932 873156 673938 873158
rect 675109 873155 675175 873158
rect 669037 872538 669103 872541
rect 675109 872538 675175 872541
rect 669037 872536 675175 872538
rect 669037 872480 669042 872536
rect 669098 872480 675114 872536
rect 675170 872480 675175 872536
rect 669037 872478 675175 872480
rect 669037 872475 669103 872478
rect 675109 872475 675175 872478
rect 673177 872266 673243 872269
rect 675385 872266 675451 872269
rect 673177 872264 675451 872266
rect 673177 872208 673182 872264
rect 673238 872208 675390 872264
rect 675446 872208 675451 872264
rect 673177 872206 675451 872208
rect 673177 872203 673243 872206
rect 675385 872203 675451 872206
rect 62113 871722 62179 871725
rect 62113 871720 64492 871722
rect 62113 871664 62118 871720
rect 62174 871664 64492 871720
rect 62113 871662 64492 871664
rect 62113 871659 62179 871662
rect 651465 869682 651531 869685
rect 650164 869680 651531 869682
rect 650164 869624 651470 869680
rect 651526 869624 651531 869680
rect 650164 869622 651531 869624
rect 651465 869619 651531 869622
rect 671797 869274 671863 869277
rect 671797 869272 675172 869274
rect 671797 869216 671802 869272
rect 671858 869216 675172 869272
rect 671797 869214 675172 869216
rect 671797 869211 671863 869214
rect 675112 868733 675172 869214
rect 664437 868730 664503 868733
rect 674925 868730 674991 868733
rect 664437 868728 674991 868730
rect 664437 868672 664442 868728
rect 664498 868672 674930 868728
rect 674986 868672 674991 868728
rect 664437 868670 674991 868672
rect 664437 868667 664503 868670
rect 674925 868667 674991 868670
rect 675109 868728 675175 868733
rect 675109 868672 675114 868728
rect 675170 868672 675175 868728
rect 675109 868667 675175 868672
rect 674557 868458 674623 868461
rect 675293 868458 675359 868461
rect 674557 868456 675359 868458
rect 674557 868400 674562 868456
rect 674618 868400 675298 868456
rect 675354 868400 675359 868456
rect 674557 868398 675359 868400
rect 674557 868395 674623 868398
rect 675293 868395 675359 868398
rect 674097 867234 674163 867237
rect 675293 867234 675359 867237
rect 674097 867232 675359 867234
rect 674097 867176 674102 867232
rect 674158 867176 675298 867232
rect 675354 867176 675359 867232
rect 674097 867174 675359 867176
rect 674097 867171 674163 867174
rect 675293 867171 675359 867174
rect 674925 866826 674991 866829
rect 675150 866826 675156 866828
rect 674925 866824 675156 866826
rect 674925 866768 674930 866824
rect 674986 866768 675156 866824
rect 674925 866766 675156 866768
rect 674925 866763 674991 866766
rect 675150 866764 675156 866766
rect 675220 866764 675226 866828
rect 670785 865330 670851 865333
rect 675293 865330 675359 865333
rect 670785 865328 675359 865330
rect 670785 865272 670790 865328
rect 670846 865272 675298 865328
rect 675354 865272 675359 865328
rect 670785 865270 675359 865272
rect 670785 865267 670851 865270
rect 675293 865267 675359 865270
rect 673729 864922 673795 864925
rect 675477 864922 675543 864925
rect 673729 864920 675543 864922
rect 673729 864864 673734 864920
rect 673790 864864 675482 864920
rect 675538 864864 675543 864920
rect 673729 864862 675543 864864
rect 673729 864859 673795 864862
rect 675477 864859 675543 864862
rect 669773 864242 669839 864245
rect 675477 864242 675543 864245
rect 669773 864240 675543 864242
rect 669773 864184 669778 864240
rect 669834 864184 675482 864240
rect 675538 864184 675543 864240
rect 669773 864182 675543 864184
rect 669773 864179 669839 864182
rect 675477 864179 675543 864182
rect 62113 858666 62179 858669
rect 62113 858664 64492 858666
rect 62113 858608 62118 858664
rect 62174 858608 64492 858664
rect 62113 858606 64492 858608
rect 62113 858603 62179 858606
rect 651465 856354 651531 856357
rect 650164 856352 651531 856354
rect 650164 856296 651470 856352
rect 651526 856296 651531 856352
rect 650164 856294 651531 856296
rect 651465 856291 651531 856294
rect 62113 845610 62179 845613
rect 62113 845608 64492 845610
rect 62113 845552 62118 845608
rect 62174 845552 64492 845608
rect 62113 845550 64492 845552
rect 62113 845547 62179 845550
rect 651833 843026 651899 843029
rect 650164 843024 651899 843026
rect 650164 842968 651838 843024
rect 651894 842968 651899 843024
rect 650164 842966 651899 842968
rect 651833 842963 651899 842966
rect 62757 832554 62823 832557
rect 62757 832552 64492 832554
rect 62757 832496 62762 832552
rect 62818 832496 64492 832552
rect 62757 832494 64492 832496
rect 62757 832491 62823 832494
rect 651465 829834 651531 829837
rect 650164 829832 651531 829834
rect 650164 829776 651470 829832
rect 651526 829776 651531 829832
rect 650164 829774 651531 829776
rect 651465 829771 651531 829774
rect 62113 819498 62179 819501
rect 62113 819496 64492 819498
rect 62113 819440 62118 819496
rect 62174 819440 64492 819496
rect 62113 819438 64492 819440
rect 62113 819435 62179 819438
rect 47761 817730 47827 817733
rect 41492 817728 47827 817730
rect 41492 817672 47766 817728
rect 47822 817672 47827 817728
rect 41492 817670 47827 817672
rect 47761 817667 47827 817670
rect 41229 817322 41295 817325
rect 41229 817320 41308 817322
rect 41229 817264 41234 817320
rect 41290 817264 41308 817320
rect 41229 817262 41308 817264
rect 41229 817259 41295 817262
rect 50337 816914 50403 816917
rect 41492 816912 50403 816914
rect 41492 816856 50342 816912
rect 50398 816856 50403 816912
rect 41492 816854 50403 816856
rect 50337 816851 50403 816854
rect 41229 816506 41295 816509
rect 651465 816506 651531 816509
rect 41229 816504 41308 816506
rect 41229 816448 41234 816504
rect 41290 816448 41308 816504
rect 41229 816446 41308 816448
rect 650164 816504 651531 816506
rect 650164 816448 651470 816504
rect 651526 816448 651531 816504
rect 650164 816446 651531 816448
rect 41229 816443 41295 816446
rect 651465 816443 651531 816446
rect 44173 816098 44239 816101
rect 41492 816096 44239 816098
rect 41492 816040 44178 816096
rect 44234 816040 44239 816096
rect 41492 816038 44239 816040
rect 44173 816035 44239 816038
rect 40174 815658 40234 815660
rect 40166 815594 40172 815658
rect 40236 815594 40242 815658
rect 45001 815282 45067 815285
rect 41492 815280 45067 815282
rect 41492 815224 45006 815280
rect 45062 815224 45067 815280
rect 41492 815222 45067 815224
rect 45001 815219 45067 815222
rect 43529 814874 43595 814877
rect 41492 814872 43595 814874
rect 41492 814816 43534 814872
rect 43590 814816 43595 814872
rect 41492 814814 43595 814816
rect 43529 814811 43595 814814
rect 44357 814466 44423 814469
rect 41492 814464 44423 814466
rect 41492 814408 44362 814464
rect 44418 814408 44423 814464
rect 41492 814406 44423 814408
rect 44357 814403 44423 814406
rect 41781 814058 41847 814061
rect 41492 814056 41847 814058
rect 41492 814000 41786 814056
rect 41842 814000 41847 814056
rect 41492 813998 41847 814000
rect 41781 813995 41847 813998
rect 44633 813650 44699 813653
rect 41492 813648 44699 813650
rect 41492 813592 44638 813648
rect 44694 813592 44699 813648
rect 41492 813590 44699 813592
rect 44633 813587 44699 813590
rect 40953 813242 41019 813245
rect 40940 813240 41019 813242
rect 40940 813184 40958 813240
rect 41014 813184 41019 813240
rect 40940 813182 41019 813184
rect 40953 813179 41019 813182
rect 40769 812834 40835 812837
rect 40756 812832 40835 812834
rect 40756 812776 40774 812832
rect 40830 812776 40835 812832
rect 40756 812774 40835 812776
rect 40769 812771 40835 812774
rect 41137 812426 41203 812429
rect 41124 812424 41203 812426
rect 41124 812368 41142 812424
rect 41198 812368 41203 812424
rect 41124 812366 41203 812368
rect 41137 812363 41203 812366
rect 42006 812018 42012 812020
rect 41492 811958 42012 812018
rect 42006 811956 42012 811958
rect 42076 811956 42082 812020
rect 39297 811610 39363 811613
rect 39284 811608 39363 811610
rect 39284 811552 39302 811608
rect 39358 811552 39363 811608
rect 39284 811550 39363 811552
rect 39297 811547 39363 811550
rect 33041 811202 33107 811205
rect 33028 811200 33107 811202
rect 33028 811144 33046 811200
rect 33102 811144 33107 811200
rect 33028 811142 33107 811144
rect 33041 811139 33107 811142
rect 45185 810794 45251 810797
rect 41492 810792 45251 810794
rect 41492 810736 45190 810792
rect 45246 810736 45251 810792
rect 41492 810734 45251 810736
rect 45185 810731 45251 810734
rect 42977 810386 43043 810389
rect 41492 810384 43043 810386
rect 41492 810328 42982 810384
rect 43038 810328 43043 810384
rect 41492 810326 43043 810328
rect 42977 810323 43043 810326
rect 44817 809978 44883 809981
rect 41492 809976 44883 809978
rect 41492 809920 44822 809976
rect 44878 809920 44883 809976
rect 41492 809918 44883 809920
rect 44817 809915 44883 809918
rect 43161 809570 43227 809573
rect 41492 809568 43227 809570
rect 41492 809512 43166 809568
rect 43222 809512 43227 809568
rect 41492 809510 43227 809512
rect 43161 809507 43227 809510
rect 41822 809162 41828 809164
rect 41492 809102 41828 809162
rect 41822 809100 41828 809102
rect 41892 809100 41898 809164
rect 40542 808712 40602 808724
rect 40534 808648 40540 808712
rect 40604 808648 40610 808712
rect 41965 808346 42031 808349
rect 41492 808344 42031 808346
rect 41492 808288 41970 808344
rect 42026 808288 42031 808344
rect 41492 808286 42031 808288
rect 41965 808283 42031 808286
rect 42793 807938 42859 807941
rect 41492 807936 42859 807938
rect 41492 807880 42798 807936
rect 42854 807880 42859 807936
rect 41492 807878 42859 807880
rect 42793 807875 42859 807878
rect 43529 807666 43595 807669
rect 41830 807664 43595 807666
rect 41830 807608 43534 807664
rect 43590 807608 43595 807664
rect 41830 807606 43595 807608
rect 41830 807530 41890 807606
rect 43529 807603 43595 807606
rect 41492 807470 41890 807530
rect 41781 807260 41847 807261
rect 41781 807256 41828 807260
rect 41892 807258 41898 807260
rect 41781 807200 41786 807256
rect 41781 807196 41828 807200
rect 41892 807198 41938 807258
rect 41892 807196 41898 807198
rect 41781 807195 41847 807196
rect 41462 806714 41522 807092
rect 42241 806714 42307 806717
rect 41462 806712 42307 806714
rect 41462 806684 42246 806712
rect 41492 806656 42246 806684
rect 42302 806656 42307 806712
rect 41492 806654 42307 806656
rect 42241 806651 42307 806654
rect 62113 806578 62179 806581
rect 62113 806576 64492 806578
rect 62113 806520 62118 806576
rect 62174 806520 64492 806576
rect 62113 806518 64492 806520
rect 62113 806515 62179 806518
rect 43713 806306 43779 806309
rect 41492 806304 43779 806306
rect 41492 806248 43718 806304
rect 43774 806248 43779 806304
rect 41492 806246 43779 806248
rect 43713 806243 43779 806246
rect 40953 805626 41019 805629
rect 41454 805626 41460 805628
rect 40953 805624 41460 805626
rect 40953 805568 40958 805624
rect 41014 805568 41460 805624
rect 40953 805566 41460 805568
rect 40953 805563 41019 805566
rect 41454 805564 41460 805566
rect 41524 805564 41530 805628
rect 40718 805020 40724 805084
rect 40788 805082 40794 805084
rect 41965 805082 42031 805085
rect 40788 805080 42031 805082
rect 40788 805024 41970 805080
rect 42026 805024 42031 805080
rect 40788 805022 42031 805024
rect 40788 805020 40794 805022
rect 41965 805019 42031 805022
rect 651465 803314 651531 803317
rect 650164 803312 651531 803314
rect 650164 803256 651470 803312
rect 651526 803256 651531 803312
rect 650164 803254 651531 803256
rect 651465 803251 651531 803254
rect 41597 801682 41663 801685
rect 42609 801682 42675 801685
rect 41597 801680 42675 801682
rect 41597 801624 41602 801680
rect 41658 801624 42614 801680
rect 42670 801624 42675 801680
rect 41597 801622 42675 801624
rect 41597 801619 41663 801622
rect 42609 801619 42675 801622
rect 41781 800322 41847 800325
rect 41781 800320 41890 800322
rect 41781 800264 41786 800320
rect 41842 800264 41890 800320
rect 41781 800259 41890 800264
rect 41830 799917 41890 800259
rect 41781 799912 41890 799917
rect 41781 799856 41786 799912
rect 41842 799856 41890 799912
rect 41781 799854 41890 799856
rect 41781 799851 41847 799854
rect 45369 799098 45435 799101
rect 53097 799098 53163 799101
rect 45369 799096 53163 799098
rect 45369 799040 45374 799096
rect 45430 799040 53102 799096
rect 53158 799040 53163 799096
rect 45369 799038 53163 799040
rect 45369 799035 45435 799038
rect 53097 799035 53163 799038
rect 42149 797330 42215 797333
rect 45369 797330 45435 797333
rect 42149 797328 45435 797330
rect 42149 797272 42154 797328
rect 42210 797272 45374 797328
rect 45430 797272 45435 797328
rect 42149 797270 45435 797272
rect 42149 797267 42215 797270
rect 45369 797267 45435 797270
rect 42149 796242 42215 796245
rect 43161 796242 43227 796245
rect 42149 796240 43227 796242
rect 42149 796184 42154 796240
rect 42210 796184 43166 796240
rect 43222 796184 43227 796240
rect 42149 796182 43227 796184
rect 42149 796179 42215 796182
rect 43161 796179 43227 796182
rect 42057 795018 42123 795021
rect 42701 795018 42767 795021
rect 42057 795016 42767 795018
rect 42057 794960 42062 795016
rect 42118 794960 42706 795016
rect 42762 794960 42767 795016
rect 42057 794958 42767 794960
rect 42057 794955 42123 794958
rect 42701 794955 42767 794958
rect 40902 794412 40908 794476
rect 40972 794474 40978 794476
rect 41781 794474 41847 794477
rect 40972 794472 41847 794474
rect 40972 794416 41786 794472
rect 41842 794416 41847 794472
rect 40972 794414 41847 794416
rect 40972 794412 40978 794414
rect 41781 794411 41847 794414
rect 40718 793732 40724 793796
rect 40788 793794 40794 793796
rect 41781 793794 41847 793797
rect 40788 793792 41847 793794
rect 40788 793736 41786 793792
rect 41842 793736 41847 793792
rect 40788 793734 41847 793736
rect 40788 793732 40794 793734
rect 41781 793731 41847 793734
rect 62113 793658 62179 793661
rect 62113 793656 64492 793658
rect 62113 793600 62118 793656
rect 62174 793600 64492 793656
rect 62113 793598 64492 793600
rect 62113 793595 62179 793598
rect 40534 792508 40540 792572
rect 40604 792570 40610 792572
rect 42241 792570 42307 792573
rect 40604 792568 42307 792570
rect 40604 792512 42246 792568
rect 42302 792512 42307 792568
rect 40604 792510 42307 792512
rect 40604 792508 40610 792510
rect 42241 792507 42307 792510
rect 42425 792298 42491 792301
rect 44817 792298 44883 792301
rect 42425 792296 44883 792298
rect 42425 792240 42430 792296
rect 42486 792240 44822 792296
rect 44878 792240 44883 792296
rect 42425 792238 44883 792240
rect 42425 792235 42491 792238
rect 44817 792235 44883 792238
rect 651465 789986 651531 789989
rect 650164 789984 651531 789986
rect 650164 789928 651470 789984
rect 651526 789928 651531 789984
rect 650164 789926 651531 789928
rect 651465 789923 651531 789926
rect 42149 789442 42215 789445
rect 42793 789442 42859 789445
rect 42149 789440 42859 789442
rect 42149 789384 42154 789440
rect 42210 789384 42798 789440
rect 42854 789384 42859 789440
rect 42149 789382 42859 789384
rect 42149 789379 42215 789382
rect 42793 789379 42859 789382
rect 41638 789108 41644 789172
rect 41708 789170 41714 789172
rect 42333 789170 42399 789173
rect 41708 789168 42399 789170
rect 41708 789112 42338 789168
rect 42394 789112 42399 789168
rect 41708 789110 42399 789112
rect 41708 789108 41714 789110
rect 42333 789107 42399 789110
rect 41822 788700 41828 788764
rect 41892 788762 41898 788764
rect 42609 788762 42675 788765
rect 41892 788760 42675 788762
rect 41892 788704 42614 788760
rect 42670 788704 42675 788760
rect 41892 788702 42675 788704
rect 41892 788700 41898 788702
rect 42609 788699 42675 788702
rect 42793 788626 42859 788629
rect 62757 788626 62823 788629
rect 42793 788624 62823 788626
rect 42793 788568 42798 788624
rect 42854 788568 62762 788624
rect 62818 788568 62823 788624
rect 42793 788566 62823 788568
rect 42793 788563 42859 788566
rect 62757 788563 62823 788566
rect 41454 788156 41460 788220
rect 41524 788218 41530 788220
rect 42241 788218 42307 788221
rect 41524 788216 42307 788218
rect 41524 788160 42246 788216
rect 42302 788160 42307 788216
rect 41524 788158 42307 788160
rect 41524 788156 41530 788158
rect 42241 788155 42307 788158
rect 42425 788218 42491 788221
rect 45185 788218 45251 788221
rect 42425 788216 45251 788218
rect 42425 788160 42430 788216
rect 42486 788160 45190 788216
rect 45246 788160 45251 788216
rect 42425 788158 45251 788160
rect 42425 788155 42491 788158
rect 45185 788155 45251 788158
rect 674281 788082 674347 788085
rect 675477 788082 675543 788085
rect 674281 788080 675543 788082
rect 674281 788024 674286 788080
rect 674342 788024 675482 788080
rect 675538 788024 675543 788080
rect 674281 788022 675543 788024
rect 674281 788019 674347 788022
rect 675477 788019 675543 788022
rect 672349 787402 672415 787405
rect 675477 787402 675543 787405
rect 672349 787400 675543 787402
rect 672349 787344 672354 787400
rect 672410 787344 675482 787400
rect 675538 787344 675543 787400
rect 672349 787342 675543 787344
rect 672349 787339 672415 787342
rect 675477 787339 675543 787342
rect 674925 786722 674991 786725
rect 675385 786722 675451 786725
rect 674925 786720 675451 786722
rect 674925 786664 674930 786720
rect 674986 786664 675390 786720
rect 675446 786664 675451 786720
rect 674925 786662 675451 786664
rect 674925 786659 674991 786662
rect 675385 786659 675451 786662
rect 672993 784274 673059 784277
rect 675477 784274 675543 784277
rect 672993 784272 675543 784274
rect 672993 784216 672998 784272
rect 673054 784216 675482 784272
rect 675538 784216 675543 784272
rect 672993 784214 675543 784216
rect 672993 784211 673059 784214
rect 675477 784211 675543 784214
rect 672625 783866 672691 783869
rect 675477 783866 675543 783869
rect 672625 783864 675543 783866
rect 672625 783808 672630 783864
rect 672686 783808 675482 783864
rect 675538 783808 675543 783864
rect 672625 783806 675543 783808
rect 672625 783803 672691 783806
rect 675477 783803 675543 783806
rect 674414 782988 674420 783052
rect 674484 783050 674490 783052
rect 675477 783050 675543 783053
rect 674484 783048 675543 783050
rect 674484 782992 675482 783048
rect 675538 782992 675543 783048
rect 674484 782990 675543 782992
rect 674484 782988 674490 782990
rect 675477 782987 675543 782990
rect 667841 780738 667907 780741
rect 675477 780738 675543 780741
rect 667841 780736 675543 780738
rect 667841 780680 667846 780736
rect 667902 780680 675482 780736
rect 675538 780680 675543 780736
rect 667841 780678 675543 780680
rect 667841 780675 667907 780678
rect 675477 780675 675543 780678
rect 62757 780466 62823 780469
rect 675293 780468 675359 780469
rect 62757 780464 64492 780466
rect 62757 780408 62762 780464
rect 62818 780408 64492 780464
rect 62757 780406 64492 780408
rect 675293 780464 675340 780468
rect 675404 780466 675410 780468
rect 675293 780408 675298 780464
rect 62757 780403 62823 780406
rect 675293 780404 675340 780408
rect 675404 780406 675450 780466
rect 675404 780404 675410 780406
rect 675293 780403 675359 780404
rect 670417 780058 670483 780061
rect 675477 780058 675543 780061
rect 670417 780056 675543 780058
rect 670417 780000 670422 780056
rect 670478 780000 675482 780056
rect 675538 780000 675543 780056
rect 670417 779998 675543 780000
rect 670417 779995 670483 779998
rect 675477 779995 675543 779998
rect 670325 779514 670391 779517
rect 675477 779514 675543 779517
rect 670325 779512 675543 779514
rect 670325 779456 670330 779512
rect 670386 779456 675482 779512
rect 675538 779456 675543 779512
rect 670325 779454 675543 779456
rect 670325 779451 670391 779454
rect 675477 779451 675543 779454
rect 673913 779242 673979 779245
rect 675477 779242 675543 779245
rect 673913 779240 675543 779242
rect 673913 779184 673918 779240
rect 673974 779184 675482 779240
rect 675538 779184 675543 779240
rect 673913 779182 675543 779184
rect 673913 779179 673979 779182
rect 675477 779179 675543 779182
rect 660297 778970 660363 778973
rect 675293 778970 675359 778973
rect 660297 778968 675359 778970
rect 660297 778912 660302 778968
rect 660358 778912 675298 778968
rect 675354 778912 675359 778968
rect 660297 778910 675359 778912
rect 660297 778907 660363 778910
rect 675293 778907 675359 778910
rect 666277 778426 666343 778429
rect 675518 778426 675524 778428
rect 666277 778424 675524 778426
rect 666277 778368 666282 778424
rect 666338 778368 675524 778424
rect 666277 778366 675524 778368
rect 666277 778363 666343 778366
rect 675518 778364 675524 778366
rect 675588 778364 675594 778428
rect 673545 777474 673611 777477
rect 675477 777474 675543 777477
rect 673545 777472 675543 777474
rect 673545 777416 673550 777472
rect 673606 777416 675482 777472
rect 675538 777416 675543 777472
rect 673545 777414 675543 777416
rect 673545 777411 673611 777414
rect 675477 777411 675543 777414
rect 675017 777204 675083 777205
rect 674966 777140 674972 777204
rect 675036 777202 675083 777204
rect 675036 777200 675128 777202
rect 675078 777144 675128 777200
rect 675036 777142 675128 777144
rect 675036 777140 675083 777142
rect 675017 777139 675083 777140
rect 652385 776658 652451 776661
rect 650164 776656 652451 776658
rect 650164 776600 652390 776656
rect 652446 776600 652451 776656
rect 650164 776598 652451 776600
rect 652385 776595 652451 776598
rect 675477 776252 675543 776253
rect 675477 776248 675524 776252
rect 675588 776250 675594 776252
rect 675477 776192 675482 776248
rect 675477 776188 675524 776192
rect 675588 776190 675634 776250
rect 675588 776188 675594 776190
rect 675477 776187 675543 776188
rect 675293 776116 675359 776117
rect 675293 776114 675340 776116
rect 675248 776112 675340 776114
rect 675248 776056 675298 776112
rect 675248 776054 675340 776056
rect 675293 776052 675340 776054
rect 675404 776052 675410 776116
rect 675293 776051 675359 776052
rect 670141 775706 670207 775709
rect 674925 775706 674991 775709
rect 670141 775704 674991 775706
rect 670141 775648 670146 775704
rect 670202 775648 674930 775704
rect 674986 775648 674991 775704
rect 670141 775646 674991 775648
rect 670141 775643 670207 775646
rect 674925 775643 674991 775646
rect 671153 775026 671219 775029
rect 675477 775026 675543 775029
rect 671153 775024 675543 775026
rect 671153 774968 671158 775024
rect 671214 774968 675482 775024
rect 675538 774968 675543 775024
rect 671153 774966 675543 774968
rect 671153 774963 671219 774966
rect 675477 774963 675543 774966
rect 674925 774618 674991 774621
rect 675477 774618 675543 774621
rect 674925 774616 675543 774618
rect 674925 774560 674930 774616
rect 674986 774560 675482 774616
rect 675538 774560 675543 774616
rect 674925 774558 675543 774560
rect 674925 774555 674991 774558
rect 675477 774555 675543 774558
rect 41462 774346 41522 774452
rect 54477 774346 54543 774349
rect 41462 774344 54543 774346
rect 41462 774288 54482 774344
rect 54538 774288 54543 774344
rect 41462 774286 54543 774288
rect 54477 774283 54543 774286
rect 35758 773941 35818 774044
rect 35758 773936 35867 773941
rect 35758 773880 35806 773936
rect 35862 773880 35867 773936
rect 35758 773878 35867 773880
rect 35801 773875 35867 773878
rect 41462 773530 41522 773636
rect 51717 773530 51783 773533
rect 41462 773528 51783 773530
rect 41462 773472 51722 773528
rect 51778 773472 51783 773528
rect 41462 773470 51783 773472
rect 51717 773467 51783 773470
rect 674966 773332 674972 773396
rect 675036 773394 675042 773396
rect 675385 773394 675451 773397
rect 675036 773392 675451 773394
rect 675036 773336 675390 773392
rect 675446 773336 675451 773392
rect 675036 773334 675451 773336
rect 675036 773332 675042 773334
rect 675385 773331 675451 773334
rect 44173 773258 44239 773261
rect 41492 773256 44239 773258
rect 41492 773200 44178 773256
rect 44234 773200 44239 773256
rect 41492 773198 44239 773200
rect 44173 773195 44239 773198
rect 44817 772850 44883 772853
rect 41492 772848 44883 772850
rect 41492 772792 44822 772848
rect 44878 772792 44883 772848
rect 41492 772790 44883 772792
rect 44817 772787 44883 772790
rect 45001 772442 45067 772445
rect 41492 772440 45067 772442
rect 41492 772384 45006 772440
rect 45062 772384 45067 772440
rect 41492 772382 45067 772384
rect 45001 772379 45067 772382
rect 673862 772244 673868 772308
rect 673932 772306 673938 772308
rect 683205 772306 683271 772309
rect 673932 772304 683271 772306
rect 673932 772248 683210 772304
rect 683266 772248 683271 772304
rect 673932 772246 683271 772248
rect 673932 772244 673938 772246
rect 683205 772243 683271 772246
rect 44449 772034 44515 772037
rect 41492 772032 44515 772034
rect 41492 771976 44454 772032
rect 44510 771976 44515 772032
rect 41492 771974 44515 771976
rect 44449 771971 44515 771974
rect 673729 772034 673795 772037
rect 683849 772034 683915 772037
rect 673729 772032 683915 772034
rect 673729 771976 673734 772032
rect 673790 771976 683854 772032
rect 683910 771976 683915 772032
rect 673729 771974 683915 771976
rect 673729 771971 673795 771974
rect 683849 771971 683915 771974
rect 44265 771626 44331 771629
rect 41492 771624 44331 771626
rect 41492 771568 44270 771624
rect 44326 771568 44331 771624
rect 41492 771566 44331 771568
rect 44265 771563 44331 771566
rect 45001 771218 45067 771221
rect 41492 771216 45067 771218
rect 41492 771160 45006 771216
rect 45062 771160 45067 771216
rect 41492 771158 45067 771160
rect 45001 771155 45067 771158
rect 44633 770810 44699 770813
rect 41492 770808 44699 770810
rect 41492 770752 44638 770808
rect 44694 770752 44699 770808
rect 41492 770750 44699 770752
rect 44633 770747 44699 770750
rect 674557 770674 674623 770677
rect 683481 770674 683547 770677
rect 674557 770672 683547 770674
rect 674557 770616 674562 770672
rect 674618 770616 683486 770672
rect 683542 770616 683547 770672
rect 674557 770614 683547 770616
rect 674557 770611 674623 770614
rect 683481 770611 683547 770614
rect 44265 770402 44331 770405
rect 41492 770400 44331 770402
rect 41492 770344 44270 770400
rect 44326 770344 44331 770400
rect 41492 770342 44331 770344
rect 44265 770339 44331 770342
rect 41462 769860 41522 769964
rect 41454 769796 41460 769860
rect 41524 769796 41530 769860
rect 35390 769453 35450 769556
rect 35341 769448 35450 769453
rect 35341 769392 35346 769448
rect 35402 769392 35450 769448
rect 35341 769390 35450 769392
rect 35341 769387 35407 769390
rect 35574 769045 35634 769148
rect 35525 769040 35634 769045
rect 35801 769042 35867 769045
rect 35525 768984 35530 769040
rect 35586 768984 35634 769040
rect 35525 768982 35634 768984
rect 35758 769040 35867 769042
rect 35758 768984 35806 769040
rect 35862 768984 35867 769040
rect 35525 768979 35591 768982
rect 35758 768979 35867 768984
rect 35758 768740 35818 768979
rect 676070 768708 676076 768772
rect 676140 768770 676146 768772
rect 680997 768770 681063 768773
rect 676140 768768 681063 768770
rect 676140 768712 681002 768768
rect 681058 768712 681063 768768
rect 676140 768710 681063 768712
rect 676140 768708 676146 768710
rect 680997 768707 681063 768710
rect 35574 768229 35634 768332
rect 35574 768224 35683 768229
rect 35574 768168 35622 768224
rect 35678 768168 35683 768224
rect 35574 768166 35683 768168
rect 35617 768163 35683 768166
rect 30974 767821 31034 767924
rect 30974 767816 31083 767821
rect 35801 767818 35867 767821
rect 30974 767760 31022 767816
rect 31078 767760 31083 767816
rect 30974 767758 31083 767760
rect 31017 767755 31083 767758
rect 35758 767816 35867 767818
rect 35758 767760 35806 767816
rect 35862 767760 35867 767816
rect 35758 767755 35867 767760
rect 35758 767516 35818 767755
rect 62113 767410 62179 767413
rect 62113 767408 64492 767410
rect 62113 767352 62118 767408
rect 62174 767352 64492 767408
rect 62113 767350 64492 767352
rect 62113 767347 62179 767350
rect 35206 767005 35266 767108
rect 35157 767000 35266 767005
rect 35157 766944 35162 767000
rect 35218 766944 35266 767000
rect 35157 766942 35266 766944
rect 35157 766939 35223 766942
rect 43069 766730 43135 766733
rect 41492 766728 43135 766730
rect 41492 766672 43074 766728
rect 43130 766672 43135 766728
rect 41492 766670 43135 766672
rect 43069 766667 43135 766670
rect 675017 766594 675083 766597
rect 675886 766594 675892 766596
rect 675017 766592 675892 766594
rect 675017 766536 675022 766592
rect 675078 766536 675892 766592
rect 675017 766534 675892 766536
rect 675017 766531 675083 766534
rect 675886 766532 675892 766534
rect 675956 766532 675962 766596
rect 44633 766322 44699 766325
rect 41492 766320 44699 766322
rect 41492 766264 44638 766320
rect 44694 766264 44699 766320
rect 41492 766262 44699 766264
rect 44633 766259 44699 766262
rect 40910 765780 40970 765884
rect 40902 765716 40908 765780
rect 40972 765716 40978 765780
rect 40542 765372 40602 765476
rect 40534 765308 40540 765372
rect 40604 765308 40610 765372
rect 41321 765370 41387 765373
rect 42517 765370 42583 765373
rect 41321 765368 42583 765370
rect 41321 765312 41326 765368
rect 41382 765312 42522 765368
rect 42578 765312 42583 765368
rect 41321 765310 42583 765312
rect 41321 765307 41387 765310
rect 42517 765307 42583 765310
rect 675201 765098 675267 765101
rect 676070 765098 676076 765100
rect 675201 765096 676076 765098
rect 40726 764964 40786 765068
rect 675201 765040 675206 765096
rect 675262 765040 676076 765096
rect 675201 765038 676076 765040
rect 675201 765035 675267 765038
rect 676070 765036 676076 765038
rect 676140 765036 676146 765100
rect 40718 764900 40724 764964
rect 40788 764900 40794 764964
rect 42793 764690 42859 764693
rect 41492 764688 42859 764690
rect 41492 764632 42798 764688
rect 42854 764632 42859 764688
rect 41492 764630 42859 764632
rect 42793 764627 42859 764630
rect 45553 764282 45619 764285
rect 41492 764280 45619 764282
rect 41492 764224 45558 764280
rect 45614 764224 45619 764280
rect 41492 764222 45619 764224
rect 45553 764219 45619 764222
rect 35758 763333 35818 763844
rect 671337 763738 671403 763741
rect 683389 763738 683455 763741
rect 671337 763736 683455 763738
rect 671337 763680 671342 763736
rect 671398 763680 683394 763736
rect 683450 763680 683455 763736
rect 671337 763678 683455 763680
rect 671337 763675 671403 763678
rect 683389 763675 683455 763678
rect 35758 763328 35867 763333
rect 651465 763330 651531 763333
rect 35758 763272 35806 763328
rect 35862 763272 35867 763328
rect 35758 763270 35867 763272
rect 650164 763328 651531 763330
rect 650164 763272 651470 763328
rect 651526 763272 651531 763328
rect 650164 763270 651531 763272
rect 35801 763267 35867 763270
rect 651465 763267 651531 763270
rect 43897 763058 43963 763061
rect 41492 763056 43963 763058
rect 41492 763000 43902 763056
rect 43958 763000 43963 763056
rect 41492 762998 43963 763000
rect 43897 762995 43963 762998
rect 676765 761836 676831 761837
rect 676765 761832 676812 761836
rect 676876 761834 676882 761836
rect 676765 761776 676770 761832
rect 676765 761772 676812 761776
rect 676876 761774 676922 761834
rect 676876 761772 676882 761774
rect 676765 761771 676831 761772
rect 665817 761562 665883 761565
rect 665817 761560 676292 761562
rect 665817 761504 665822 761560
rect 665878 761504 676292 761560
rect 665817 761502 676292 761504
rect 665817 761499 665883 761502
rect 669270 761094 676292 761154
rect 663057 760474 663123 760477
rect 669270 760474 669330 761094
rect 683389 760746 683455 760749
rect 683389 760744 683468 760746
rect 683389 760688 683394 760744
rect 683450 760688 683468 760744
rect 683389 760686 683468 760688
rect 683389 760683 683455 760686
rect 663057 760472 669330 760474
rect 663057 760416 663062 760472
rect 663118 760416 669330 760472
rect 663057 760414 669330 760416
rect 663057 760411 663123 760414
rect 673361 760338 673427 760341
rect 673361 760336 676292 760338
rect 673361 760280 673366 760336
rect 673422 760280 676292 760336
rect 673361 760278 676292 760280
rect 673361 760275 673427 760278
rect 671429 759930 671495 759933
rect 671429 759928 676292 759930
rect 671429 759872 671434 759928
rect 671490 759872 676292 759928
rect 671429 759870 676292 759872
rect 671429 759867 671495 759870
rect 672809 759522 672875 759525
rect 672809 759520 676292 759522
rect 672809 759464 672814 759520
rect 672870 759464 676292 759520
rect 672809 759462 676292 759464
rect 672809 759459 672875 759462
rect 36537 759114 36603 759117
rect 41638 759114 41644 759116
rect 36537 759112 41644 759114
rect 36537 759056 36542 759112
rect 36598 759056 41644 759112
rect 36537 759054 41644 759056
rect 36537 759051 36603 759054
rect 41638 759052 41644 759054
rect 41708 759052 41714 759116
rect 671613 759114 671679 759117
rect 671613 759112 676292 759114
rect 671613 759056 671618 759112
rect 671674 759056 676292 759112
rect 671613 759054 676292 759056
rect 671613 759051 671679 759054
rect 670969 758706 671035 758709
rect 670969 758704 676292 758706
rect 670969 758648 670974 758704
rect 671030 758648 676292 758704
rect 670969 758646 676292 758648
rect 670969 758643 671035 758646
rect 670969 758298 671035 758301
rect 670969 758296 676292 758298
rect 670969 758240 670974 758296
rect 671030 758240 676292 758296
rect 670969 758238 676292 758240
rect 670969 758235 671035 758238
rect 40309 758026 40375 758029
rect 41086 758026 41092 758028
rect 40309 758024 41092 758026
rect 40309 757968 40314 758024
rect 40370 757968 41092 758024
rect 40309 757966 41092 757968
rect 40309 757963 40375 757966
rect 41086 757964 41092 757966
rect 41156 757964 41162 758028
rect 42149 757890 42215 757893
rect 42374 757890 42380 757892
rect 42149 757888 42380 757890
rect 42149 757832 42154 757888
rect 42210 757832 42380 757888
rect 42149 757830 42380 757832
rect 42149 757827 42215 757830
rect 42374 757828 42380 757830
rect 42444 757828 42450 757892
rect 671981 757890 672047 757893
rect 671981 757888 676292 757890
rect 671981 757832 671986 757888
rect 672042 757832 676292 757888
rect 671981 757830 676292 757832
rect 671981 757827 672047 757830
rect 39297 757754 39363 757757
rect 42006 757754 42012 757756
rect 39297 757752 42012 757754
rect 39297 757696 39302 757752
rect 39358 757696 42012 757752
rect 39297 757694 42012 757696
rect 39297 757691 39363 757694
rect 42006 757692 42012 757694
rect 42076 757692 42082 757756
rect 40309 757484 40375 757485
rect 40309 757482 40356 757484
rect 40264 757480 40356 757482
rect 40264 757424 40314 757480
rect 40264 757422 40356 757424
rect 40309 757420 40356 757422
rect 40420 757420 40426 757484
rect 671337 757482 671403 757485
rect 671337 757480 676292 757482
rect 671337 757424 671342 757480
rect 671398 757424 676292 757480
rect 671337 757422 676292 757424
rect 40309 757419 40375 757420
rect 671337 757419 671403 757422
rect 674833 757210 674899 757213
rect 676029 757210 676095 757213
rect 674833 757208 676095 757210
rect 674833 757152 674838 757208
rect 674894 757152 676034 757208
rect 676090 757152 676095 757208
rect 674833 757150 676095 757152
rect 674833 757147 674899 757150
rect 676029 757147 676095 757150
rect 680997 757074 681063 757077
rect 680997 757072 681076 757074
rect 680997 757016 681002 757072
rect 681058 757016 681076 757072
rect 680997 757014 681076 757016
rect 680997 757011 681063 757014
rect 683849 756666 683915 756669
rect 683836 756664 683915 756666
rect 683836 756608 683854 756664
rect 683910 756608 683915 756664
rect 683836 756606 683915 756608
rect 683849 756603 683915 756606
rect 672809 756258 672875 756261
rect 672809 756256 676292 756258
rect 672809 756200 672814 756256
rect 672870 756200 676292 756256
rect 672809 756198 676292 756200
rect 672809 756195 672875 756198
rect 675845 755850 675911 755853
rect 675845 755848 676292 755850
rect 675845 755792 675850 755848
rect 675906 755792 676292 755848
rect 675845 755790 676292 755792
rect 675845 755787 675911 755790
rect 40350 755380 40356 755444
rect 40420 755442 40426 755444
rect 41781 755442 41847 755445
rect 40420 755440 41847 755442
rect 40420 755384 41786 755440
rect 41842 755384 41847 755440
rect 40420 755382 41847 755384
rect 40420 755380 40426 755382
rect 41781 755379 41847 755382
rect 669037 755442 669103 755445
rect 669037 755440 676292 755442
rect 669037 755384 669042 755440
rect 669098 755384 676292 755440
rect 669037 755382 676292 755384
rect 669037 755379 669103 755382
rect 666461 755170 666527 755173
rect 672809 755170 672875 755173
rect 666461 755168 672875 755170
rect 666461 755112 666466 755168
rect 666522 755112 672814 755168
rect 672870 755112 672875 755168
rect 666461 755110 672875 755112
rect 666461 755107 666527 755110
rect 672809 755107 672875 755110
rect 672950 754974 676292 755034
rect 42190 754836 42196 754900
rect 42260 754898 42266 754900
rect 44633 754898 44699 754901
rect 42260 754896 44699 754898
rect 42260 754840 44638 754896
rect 44694 754840 44699 754896
rect 42260 754838 44699 754840
rect 42260 754836 42266 754838
rect 44633 754835 44699 754838
rect 670785 754898 670851 754901
rect 672950 754898 673010 754974
rect 670785 754896 673010 754898
rect 670785 754840 670790 754896
rect 670846 754840 673010 754896
rect 670785 754838 673010 754840
rect 670785 754835 670851 754838
rect 676765 754626 676831 754629
rect 676765 754624 676844 754626
rect 676765 754568 676770 754624
rect 676826 754568 676844 754624
rect 676765 754566 676844 754568
rect 676765 754563 676831 754566
rect 62113 754354 62179 754357
rect 62113 754352 64492 754354
rect 62113 754296 62118 754352
rect 62174 754296 64492 754352
rect 62113 754294 64492 754296
rect 62113 754291 62179 754294
rect 668393 754218 668459 754221
rect 668393 754216 676292 754218
rect 668393 754160 668398 754216
rect 668454 754160 676292 754216
rect 668393 754158 676292 754160
rect 668393 754155 668459 754158
rect 42057 754082 42123 754085
rect 46197 754082 46263 754085
rect 42057 754080 46263 754082
rect 42057 754024 42062 754080
rect 42118 754024 46202 754080
rect 46258 754024 46263 754080
rect 42057 754022 46263 754024
rect 42057 754019 42123 754022
rect 46197 754019 46263 754022
rect 683205 753810 683271 753813
rect 683205 753808 683284 753810
rect 683205 753752 683210 753808
rect 683266 753752 683284 753808
rect 683205 753750 683284 753752
rect 683205 753747 683271 753750
rect 41086 753612 41092 753676
rect 41156 753674 41162 753676
rect 42241 753674 42307 753677
rect 41156 753672 42307 753674
rect 41156 753616 42246 753672
rect 42302 753616 42307 753672
rect 41156 753614 42307 753616
rect 41156 753612 41162 753614
rect 42241 753611 42307 753614
rect 42374 753340 42380 753404
rect 42444 753402 42450 753404
rect 42609 753402 42675 753405
rect 42444 753400 42675 753402
rect 42444 753344 42614 753400
rect 42670 753344 42675 753400
rect 42444 753342 42675 753344
rect 42444 753340 42450 753342
rect 42609 753339 42675 753342
rect 674097 753402 674163 753405
rect 674097 753400 676292 753402
rect 674097 753344 674102 753400
rect 674158 753344 676292 753400
rect 674097 753342 676292 753344
rect 674097 753339 674163 753342
rect 41965 752994 42031 752997
rect 42190 752994 42196 752996
rect 41965 752992 42196 752994
rect 41965 752936 41970 752992
rect 42026 752936 42196 752992
rect 41965 752934 42196 752936
rect 41965 752931 42031 752934
rect 42190 752932 42196 752934
rect 42260 752932 42266 752996
rect 683573 752994 683639 752997
rect 683573 752992 683652 752994
rect 683573 752936 683578 752992
rect 683634 752936 683652 752992
rect 683573 752934 683652 752936
rect 683573 752931 683639 752934
rect 673177 752586 673243 752589
rect 673177 752584 676292 752586
rect 673177 752528 673182 752584
rect 673238 752528 676292 752584
rect 673177 752526 676292 752528
rect 673177 752523 673243 752526
rect 683389 752178 683455 752181
rect 683389 752176 683468 752178
rect 683389 752120 683394 752176
rect 683450 752120 683468 752176
rect 683389 752118 683468 752120
rect 683389 752115 683455 752118
rect 42241 752044 42307 752045
rect 42190 752042 42196 752044
rect 42150 751982 42196 752042
rect 42260 752040 42307 752044
rect 42302 751984 42307 752040
rect 42190 751980 42196 751982
rect 42260 751980 42307 751984
rect 42241 751979 42307 751980
rect 42057 751770 42123 751773
rect 42793 751770 42859 751773
rect 42057 751768 42859 751770
rect 42057 751712 42062 751768
rect 42118 751712 42798 751768
rect 42854 751712 42859 751768
rect 42057 751710 42859 751712
rect 42057 751707 42123 751710
rect 42793 751707 42859 751710
rect 671981 751770 672047 751773
rect 671981 751768 676292 751770
rect 671981 751712 671986 751768
rect 672042 751712 676292 751768
rect 671981 751710 676292 751712
rect 671981 751707 672047 751710
rect 673177 751362 673243 751365
rect 673177 751360 676292 751362
rect 673177 751304 673182 751360
rect 673238 751304 676292 751360
rect 673177 751302 676292 751304
rect 673177 751299 673243 751302
rect 40902 751028 40908 751092
rect 40972 751090 40978 751092
rect 41781 751090 41847 751093
rect 40972 751088 41847 751090
rect 40972 751032 41786 751088
rect 41842 751032 41847 751088
rect 40972 751030 41847 751032
rect 40972 751028 40978 751030
rect 41781 751027 41847 751030
rect 669773 750954 669839 750957
rect 669773 750952 676292 750954
rect 669773 750896 669778 750952
rect 669834 750924 676292 750952
rect 669834 750896 676322 750924
rect 669773 750894 676322 750896
rect 669773 750891 669839 750894
rect 676262 750516 676322 750894
rect 40718 750348 40724 750412
rect 40788 750410 40794 750412
rect 41781 750410 41847 750413
rect 40788 750408 41847 750410
rect 40788 750352 41786 750408
rect 41842 750352 41847 750408
rect 40788 750350 41847 750352
rect 40788 750348 40794 750350
rect 41781 750347 41847 750350
rect 651465 750138 651531 750141
rect 650164 750136 651531 750138
rect 650164 750080 651470 750136
rect 651526 750080 651531 750136
rect 650164 750078 651531 750080
rect 651465 750075 651531 750078
rect 672349 750138 672415 750141
rect 672349 750136 676292 750138
rect 672349 750080 672354 750136
rect 672410 750080 676292 750136
rect 672349 750078 676292 750080
rect 672349 750075 672415 750078
rect 40534 749396 40540 749460
rect 40604 749458 40610 749460
rect 42241 749458 42307 749461
rect 40604 749456 42307 749458
rect 40604 749400 42246 749456
rect 42302 749400 42307 749456
rect 40604 749398 42307 749400
rect 40604 749396 40610 749398
rect 42241 749395 42307 749398
rect 42425 749322 42491 749325
rect 43069 749322 43135 749325
rect 42425 749320 43135 749322
rect 42425 749264 42430 749320
rect 42486 749264 43074 749320
rect 43130 749264 43135 749320
rect 42425 749262 43135 749264
rect 42425 749259 42491 749262
rect 43069 749259 43135 749262
rect 41454 746540 41460 746604
rect 41524 746602 41530 746604
rect 42241 746602 42307 746605
rect 41524 746600 42307 746602
rect 41524 746544 42246 746600
rect 42302 746544 42307 746600
rect 41524 746542 42307 746544
rect 41524 746540 41530 746542
rect 42241 746539 42307 746542
rect 41638 746268 41644 746332
rect 41708 746330 41714 746332
rect 42425 746330 42491 746333
rect 41708 746328 42491 746330
rect 41708 746272 42430 746328
rect 42486 746272 42491 746328
rect 41708 746270 42491 746272
rect 41708 746268 41714 746270
rect 42425 746267 42491 746270
rect 41965 746058 42031 746061
rect 42190 746058 42196 746060
rect 41965 746056 42196 746058
rect 41965 746000 41970 746056
rect 42026 746000 42196 746056
rect 41965 745998 42196 746000
rect 41965 745995 42031 745998
rect 42190 745996 42196 745998
rect 42260 745996 42266 746060
rect 42057 745514 42123 745517
rect 42609 745514 42675 745517
rect 42057 745512 42675 745514
rect 42057 745456 42062 745512
rect 42118 745456 42614 745512
rect 42670 745456 42675 745512
rect 42057 745454 42675 745456
rect 42057 745451 42123 745454
rect 42609 745451 42675 745454
rect 666461 745514 666527 745517
rect 675293 745514 675359 745517
rect 666461 745512 675359 745514
rect 666461 745456 666466 745512
rect 666522 745456 675298 745512
rect 675354 745456 675359 745512
rect 666461 745454 675359 745456
rect 666461 745451 666527 745454
rect 675293 745451 675359 745454
rect 41822 745044 41828 745108
rect 41892 745106 41898 745108
rect 42701 745106 42767 745109
rect 41892 745104 42767 745106
rect 41892 745048 42706 745104
rect 42762 745048 42767 745104
rect 41892 745046 42767 745048
rect 41892 745044 41898 745046
rect 42701 745043 42767 745046
rect 671981 743474 672047 743477
rect 675109 743474 675175 743477
rect 671981 743472 675175 743474
rect 671981 743416 671986 743472
rect 672042 743416 675114 743472
rect 675170 743416 675175 743472
rect 671981 743414 675175 743416
rect 671981 743411 672047 743414
rect 675109 743411 675175 743414
rect 42701 743066 42767 743069
rect 62757 743066 62823 743069
rect 42701 743064 62823 743066
rect 42701 743008 42706 743064
rect 42762 743008 62762 743064
rect 62818 743008 62823 743064
rect 42701 743006 62823 743008
rect 42701 743003 42767 743006
rect 62757 743003 62823 743006
rect 667657 742522 667723 742525
rect 674925 742522 674991 742525
rect 667657 742520 674991 742522
rect 667657 742464 667662 742520
rect 667718 742464 674930 742520
rect 674986 742464 674991 742520
rect 667657 742462 674991 742464
rect 667657 742459 667723 742462
rect 674925 742459 674991 742462
rect 674598 741508 674604 741572
rect 674668 741570 674674 741572
rect 675109 741570 675175 741573
rect 674668 741568 675175 741570
rect 674668 741512 675114 741568
rect 675170 741512 675175 741568
rect 674668 741510 675175 741512
rect 674668 741508 674674 741510
rect 675109 741507 675175 741510
rect 62113 741298 62179 741301
rect 62113 741296 64492 741298
rect 62113 741240 62118 741296
rect 62174 741240 64492 741296
rect 62113 741238 64492 741240
rect 62113 741235 62179 741238
rect 673361 739938 673427 739941
rect 675293 739938 675359 739941
rect 673361 739936 675359 739938
rect 673361 739880 673366 739936
rect 673422 739880 675298 739936
rect 675354 739880 675359 739936
rect 673361 739878 675359 739880
rect 673361 739875 673427 739878
rect 675293 739875 675359 739878
rect 674230 739332 674236 739396
rect 674300 739394 674306 739396
rect 675477 739394 675543 739397
rect 674300 739392 675543 739394
rect 674300 739336 675482 739392
rect 675538 739336 675543 739392
rect 674300 739334 675543 739336
rect 674300 739332 674306 739334
rect 675477 739331 675543 739334
rect 675201 738374 675267 738377
rect 675158 738372 675267 738374
rect 675158 738316 675206 738372
rect 675262 738316 675267 738372
rect 675158 738311 675267 738316
rect 668853 738306 668919 738309
rect 675158 738306 675218 738311
rect 668853 738304 675218 738306
rect 668853 738248 668858 738304
rect 668914 738248 675218 738304
rect 668853 738246 675218 738248
rect 668853 738243 668919 738246
rect 669589 737082 669655 737085
rect 675109 737082 675175 737085
rect 669589 737080 675175 737082
rect 669589 737024 669594 737080
rect 669650 737024 675114 737080
rect 675170 737024 675175 737080
rect 669589 737022 675175 737024
rect 669589 737019 669655 737022
rect 675109 737019 675175 737022
rect 651833 736810 651899 736813
rect 650164 736808 651899 736810
rect 650164 736752 651838 736808
rect 651894 736752 651899 736808
rect 650164 736750 651899 736752
rect 651833 736747 651899 736750
rect 671797 735586 671863 735589
rect 675385 735586 675451 735589
rect 671797 735584 675451 735586
rect 671797 735528 671802 735584
rect 671858 735528 675390 735584
rect 675446 735528 675451 735584
rect 671797 735526 675451 735528
rect 671797 735523 671863 735526
rect 675385 735523 675451 735526
rect 668393 735314 668459 735317
rect 674833 735314 674899 735317
rect 668393 735312 674899 735314
rect 668393 735256 668398 735312
rect 668454 735256 674838 735312
rect 674894 735256 674899 735312
rect 668393 735254 674899 735256
rect 668393 735251 668459 735254
rect 674833 735251 674899 735254
rect 673729 734362 673795 734365
rect 675109 734362 675175 734365
rect 673729 734360 675175 734362
rect 673729 734304 673734 734360
rect 673790 734304 675114 734360
rect 675170 734304 675175 734360
rect 673729 734302 675175 734304
rect 673729 734299 673795 734302
rect 675109 734299 675175 734302
rect 672809 734090 672875 734093
rect 674925 734090 674991 734093
rect 672809 734088 674991 734090
rect 672809 734032 672814 734088
rect 672870 734032 674930 734088
rect 674986 734032 674991 734088
rect 672809 734030 674991 734032
rect 672809 734027 672875 734030
rect 674925 734027 674991 734030
rect 669037 733818 669103 733821
rect 675109 733818 675175 733821
rect 669037 733816 675175 733818
rect 669037 733760 669042 733816
rect 669098 733760 675114 733816
rect 675170 733760 675175 733816
rect 669037 733758 675175 733760
rect 669037 733755 669103 733758
rect 675109 733755 675175 733758
rect 668209 731506 668275 731509
rect 675109 731506 675175 731509
rect 668209 731504 675175 731506
rect 668209 731448 668214 731504
rect 668270 731448 675114 731504
rect 675170 731448 675175 731504
rect 668209 731446 675175 731448
rect 668209 731443 668275 731446
rect 675109 731443 675175 731446
rect 41492 731310 51090 731370
rect 35801 730962 35867 730965
rect 35788 730960 35867 730962
rect 35788 730904 35806 730960
rect 35862 730904 35867 730960
rect 35788 730902 35867 730904
rect 35801 730899 35867 730902
rect 50337 730554 50403 730557
rect 41492 730552 50403 730554
rect 41492 730496 50342 730552
rect 50398 730496 50403 730552
rect 41492 730494 50403 730496
rect 50337 730491 50403 730494
rect 44817 730146 44883 730149
rect 41492 730144 44883 730146
rect 41492 730088 44822 730144
rect 44878 730088 44883 730144
rect 41492 730086 44883 730088
rect 51030 730146 51090 731310
rect 668761 730554 668827 730557
rect 675109 730554 675175 730557
rect 668761 730552 675175 730554
rect 668761 730496 668766 730552
rect 668822 730496 675114 730552
rect 675170 730496 675175 730552
rect 668761 730494 675175 730496
rect 668761 730491 668827 730494
rect 675109 730491 675175 730494
rect 55857 730146 55923 730149
rect 51030 730144 55923 730146
rect 51030 730088 55862 730144
rect 55918 730088 55923 730144
rect 51030 730086 55923 730088
rect 44817 730083 44883 730086
rect 55857 730083 55923 730086
rect 669773 730146 669839 730149
rect 675109 730146 675175 730149
rect 669773 730144 675175 730146
rect 669773 730088 669778 730144
rect 669834 730088 675114 730144
rect 675170 730088 675175 730144
rect 669773 730086 675175 730088
rect 669773 730083 669839 730086
rect 675109 730083 675175 730086
rect 44633 729738 44699 729741
rect 41492 729736 44699 729738
rect 41492 729680 44638 729736
rect 44694 729680 44699 729736
rect 41492 729678 44699 729680
rect 44633 729675 44699 729678
rect 44449 729330 44515 729333
rect 41492 729328 44515 729330
rect 41492 729272 44454 729328
rect 44510 729272 44515 729328
rect 41492 729270 44515 729272
rect 44449 729267 44515 729270
rect 45185 728922 45251 728925
rect 41492 728920 45251 728922
rect 41492 728864 45190 728920
rect 45246 728864 45251 728920
rect 41492 728862 45251 728864
rect 45185 728859 45251 728862
rect 675886 728724 675892 728788
rect 675956 728786 675962 728788
rect 676806 728786 676812 728788
rect 675956 728726 676812 728786
rect 675956 728724 675962 728726
rect 676806 728724 676812 728726
rect 676876 728724 676882 728788
rect 670785 728650 670851 728653
rect 674373 728650 674439 728653
rect 670785 728648 674439 728650
rect 670785 728592 670790 728648
rect 670846 728592 674378 728648
rect 674434 728592 674439 728648
rect 670785 728590 674439 728592
rect 670785 728587 670851 728590
rect 674373 728587 674439 728590
rect 45001 728514 45067 728517
rect 41492 728512 45067 728514
rect 41492 728456 45006 728512
rect 45062 728456 45067 728512
rect 41492 728454 45067 728456
rect 45001 728451 45067 728454
rect 62757 728242 62823 728245
rect 669221 728242 669287 728245
rect 672165 728242 672231 728245
rect 62757 728240 64492 728242
rect 62757 728184 62762 728240
rect 62818 728184 64492 728240
rect 62757 728182 64492 728184
rect 669221 728240 672231 728242
rect 669221 728184 669226 728240
rect 669282 728184 672170 728240
rect 672226 728184 672231 728240
rect 669221 728182 672231 728184
rect 62757 728179 62823 728182
rect 669221 728179 669287 728182
rect 672165 728179 672231 728182
rect 45737 728106 45803 728109
rect 41492 728104 45803 728106
rect 41492 728048 45742 728104
rect 45798 728048 45803 728104
rect 41492 728046 45803 728048
rect 45737 728043 45803 728046
rect 44265 727698 44331 727701
rect 41492 727696 44331 727698
rect 41492 727640 44270 727696
rect 44326 727640 44331 727696
rect 41492 727638 44331 727640
rect 44265 727635 44331 727638
rect 46105 727426 46171 727429
rect 41830 727424 46171 727426
rect 41830 727368 46110 727424
rect 46166 727368 46171 727424
rect 41830 727366 46171 727368
rect 41830 727290 41890 727366
rect 46105 727363 46171 727366
rect 41492 727230 41890 727290
rect 41822 726882 41828 726884
rect 41492 726822 41828 726882
rect 41822 726820 41828 726822
rect 41892 726820 41898 726884
rect 673913 726882 673979 726885
rect 683389 726882 683455 726885
rect 673913 726880 683455 726882
rect 673913 726824 673918 726880
rect 673974 726824 683394 726880
rect 683450 726824 683455 726880
rect 673913 726822 683455 726824
rect 673913 726819 673979 726822
rect 683389 726819 683455 726822
rect 674741 726610 674807 726613
rect 674741 726608 674850 726610
rect 674741 726552 674746 726608
rect 674802 726552 674850 726608
rect 674741 726547 674850 726552
rect 41321 726474 41387 726477
rect 41308 726472 41387 726474
rect 41308 726416 41326 726472
rect 41382 726416 41387 726472
rect 41308 726414 41387 726416
rect 674790 726474 674850 726547
rect 683757 726474 683823 726477
rect 674790 726472 683823 726474
rect 674790 726416 683762 726472
rect 683818 726416 683823 726472
rect 674790 726414 683823 726416
rect 41321 726411 41387 726414
rect 683757 726411 683823 726414
rect 41137 726066 41203 726069
rect 41124 726064 41203 726066
rect 41124 726008 41142 726064
rect 41198 726008 41203 726064
rect 41124 726006 41203 726008
rect 41137 726003 41203 726006
rect 676070 725732 676076 725796
rect 676140 725794 676146 725796
rect 680997 725794 681063 725797
rect 676140 725792 681063 725794
rect 676140 725736 681002 725792
rect 681058 725736 681063 725792
rect 676140 725734 681063 725736
rect 676140 725732 676146 725734
rect 680997 725731 681063 725734
rect 41321 725658 41387 725661
rect 41308 725656 41387 725658
rect 41308 725600 41326 725656
rect 41382 725600 41387 725656
rect 41308 725598 41387 725600
rect 41321 725595 41387 725598
rect 39297 725250 39363 725253
rect 39284 725248 39363 725250
rect 39284 725192 39302 725248
rect 39358 725192 39363 725248
rect 39284 725190 39363 725192
rect 39297 725187 39363 725190
rect 36537 724842 36603 724845
rect 36524 724840 36603 724842
rect 36524 724784 36542 724840
rect 36598 724784 36603 724840
rect 36524 724782 36603 724784
rect 36537 724779 36603 724782
rect 31661 724434 31727 724437
rect 31661 724432 31740 724434
rect 31661 724376 31666 724432
rect 31722 724376 31740 724432
rect 31661 724374 31740 724376
rect 31661 724371 31727 724374
rect 673545 724298 673611 724301
rect 677317 724298 677383 724301
rect 673545 724296 677383 724298
rect 673545 724240 673550 724296
rect 673606 724240 677322 724296
rect 677378 724240 677383 724296
rect 673545 724238 677383 724240
rect 673545 724235 673611 724238
rect 677317 724235 677383 724238
rect 34513 724026 34579 724029
rect 34500 724024 34579 724026
rect 34500 723968 34518 724024
rect 34574 723968 34579 724024
rect 34500 723966 34579 723968
rect 34513 723963 34579 723966
rect 44449 723618 44515 723621
rect 41492 723616 44515 723618
rect 41492 723560 44454 723616
rect 44510 723560 44515 723616
rect 41492 723558 44515 723560
rect 44449 723555 44515 723558
rect 651465 723482 651531 723485
rect 650164 723480 651531 723482
rect 650164 723424 651470 723480
rect 651526 723424 651531 723480
rect 650164 723422 651531 723424
rect 651465 723419 651531 723422
rect 40677 723210 40743 723213
rect 40677 723208 40756 723210
rect 40677 723152 40682 723208
rect 40738 723152 40756 723208
rect 40677 723150 40756 723152
rect 40677 723147 40743 723150
rect 44173 722802 44239 722805
rect 41492 722800 44239 722802
rect 41492 722744 44178 722800
rect 44234 722744 44239 722800
rect 41492 722742 44239 722744
rect 44173 722739 44239 722742
rect 41822 722394 41828 722396
rect 41492 722334 41828 722394
rect 41822 722332 41828 722334
rect 41892 722332 41898 722396
rect 40726 721772 40786 721956
rect 40718 721708 40724 721772
rect 40788 721708 40794 721772
rect 41137 721770 41203 721773
rect 41638 721770 41644 721772
rect 41137 721768 41644 721770
rect 41137 721712 41142 721768
rect 41198 721712 41644 721768
rect 41137 721710 41644 721712
rect 41137 721707 41203 721710
rect 41638 721708 41644 721710
rect 41708 721708 41714 721772
rect 45369 721578 45435 721581
rect 41492 721576 45435 721578
rect 41492 721520 45374 721576
rect 45430 721520 45435 721576
rect 41492 721518 45435 721520
rect 45369 721515 45435 721518
rect 44909 721170 44975 721173
rect 41492 721168 44975 721170
rect 41492 721112 44914 721168
rect 44970 721112 44975 721168
rect 41492 721110 44975 721112
rect 44909 721107 44975 721110
rect 34102 720357 34162 720732
rect 34102 720352 34211 720357
rect 34102 720324 34150 720352
rect 34132 720296 34150 720324
rect 34206 720296 34211 720352
rect 34132 720294 34211 720296
rect 34145 720291 34211 720294
rect 41492 719886 41890 719946
rect 41830 719810 41890 719886
rect 43069 719810 43135 719813
rect 41830 719808 43135 719810
rect 41830 719752 43074 719808
rect 43130 719752 43135 719808
rect 41830 719750 43135 719752
rect 43069 719747 43135 719750
rect 41873 719538 41939 719541
rect 42517 719538 42583 719541
rect 41873 719536 42583 719538
rect 41873 719480 41878 719536
rect 41934 719480 42522 719536
rect 42578 719480 42583 719536
rect 41873 719478 42583 719480
rect 41873 719475 41939 719478
rect 42517 719475 42583 719478
rect 41689 719130 41755 719133
rect 42701 719130 42767 719133
rect 41689 719128 42767 719130
rect 41689 719072 41694 719128
rect 41750 719072 42706 719128
rect 42762 719072 42767 719128
rect 41689 719070 42767 719072
rect 41689 719067 41755 719070
rect 42701 719067 42767 719070
rect 40534 717980 40540 718044
rect 40604 718042 40610 718044
rect 41822 718042 41828 718044
rect 40604 717982 41828 718042
rect 40604 717980 40610 717982
rect 41822 717980 41828 717982
rect 41892 717980 41898 718044
rect 664437 716546 664503 716549
rect 664437 716544 676292 716546
rect 664437 716488 664442 716544
rect 664498 716488 676292 716544
rect 664437 716486 676292 716488
rect 664437 716483 664503 716486
rect 663750 716078 676292 716138
rect 658917 716002 658983 716005
rect 663750 716002 663810 716078
rect 658917 716000 663810 716002
rect 658917 715944 658922 716000
rect 658978 715944 663810 716000
rect 658917 715942 663810 715944
rect 658917 715939 658983 715942
rect 669957 715730 670023 715733
rect 669957 715728 676292 715730
rect 669957 715672 669962 715728
rect 670018 715672 676292 715728
rect 669957 715670 676292 715672
rect 669957 715667 670023 715670
rect 31661 715458 31727 715461
rect 41822 715458 41828 715460
rect 31661 715456 41828 715458
rect 31661 715400 31666 715456
rect 31722 715400 41828 715456
rect 31661 715398 41828 715400
rect 31661 715395 31727 715398
rect 41822 715396 41828 715398
rect 41892 715396 41898 715460
rect 62113 715322 62179 715325
rect 671429 715322 671495 715325
rect 62113 715320 64492 715322
rect 62113 715264 62118 715320
rect 62174 715264 64492 715320
rect 62113 715262 64492 715264
rect 671429 715320 676292 715322
rect 671429 715264 671434 715320
rect 671490 715264 676292 715320
rect 671429 715262 676292 715264
rect 62113 715259 62179 715262
rect 671429 715259 671495 715262
rect 40309 715186 40375 715189
rect 42333 715186 42399 715189
rect 40309 715184 42399 715186
rect 40309 715128 40314 715184
rect 40370 715128 42338 715184
rect 42394 715128 42399 715184
rect 40309 715126 42399 715128
rect 40309 715123 40375 715126
rect 42333 715123 42399 715126
rect 670785 714914 670851 714917
rect 670785 714912 676292 714914
rect 670785 714856 670790 714912
rect 670846 714856 676292 714912
rect 670785 714854 676292 714856
rect 670785 714851 670851 714854
rect 38653 714506 38719 714509
rect 42057 714506 42123 714509
rect 38653 714504 42123 714506
rect 38653 714448 38658 714504
rect 38714 714448 42062 714504
rect 42118 714448 42123 714504
rect 38653 714446 42123 714448
rect 38653 714443 38719 714446
rect 42057 714443 42123 714446
rect 671613 714506 671679 714509
rect 671613 714504 676292 714506
rect 671613 714448 671618 714504
rect 671674 714448 676292 714504
rect 671613 714446 676292 714448
rect 671613 714443 671679 714446
rect 40677 714234 40743 714237
rect 40902 714234 40908 714236
rect 40677 714232 40908 714234
rect 40677 714176 40682 714232
rect 40738 714176 40908 714232
rect 40677 714174 40908 714176
rect 40677 714171 40743 714174
rect 40902 714172 40908 714174
rect 40972 714172 40978 714236
rect 41505 714234 41571 714237
rect 42006 714234 42012 714236
rect 41505 714232 42012 714234
rect 41505 714176 41510 714232
rect 41566 714176 42012 714232
rect 41505 714174 42012 714176
rect 41505 714171 41571 714174
rect 42006 714172 42012 714174
rect 42076 714172 42082 714236
rect 671705 714098 671771 714101
rect 671705 714096 676292 714098
rect 671705 714040 671710 714096
rect 671766 714040 676292 714096
rect 671705 714038 676292 714040
rect 671705 714035 671771 714038
rect 41781 713960 41847 713965
rect 41781 713904 41786 713960
rect 41842 713904 41847 713960
rect 41781 713899 41847 713904
rect 41784 713557 41844 713899
rect 670969 713690 671035 713693
rect 670969 713688 676292 713690
rect 670969 713632 670974 713688
rect 671030 713632 676292 713688
rect 670969 713630 676292 713632
rect 670969 713627 671035 713630
rect 41781 713552 41847 713557
rect 41781 713496 41786 713552
rect 41842 713496 41847 713552
rect 41781 713491 41847 713496
rect 671521 713282 671587 713285
rect 671521 713280 676292 713282
rect 671521 713224 671526 713280
rect 671582 713224 676292 713280
rect 671521 713222 676292 713224
rect 671521 713219 671587 713222
rect 671337 712874 671403 712877
rect 671337 712872 676292 712874
rect 671337 712816 671342 712872
rect 671398 712816 676292 712872
rect 671337 712814 676292 712816
rect 671337 712811 671403 712814
rect 672165 712466 672231 712469
rect 672165 712464 676292 712466
rect 672165 712408 672170 712464
rect 672226 712408 676292 712464
rect 672165 712406 676292 712408
rect 672165 712403 672231 712406
rect 675886 711996 675892 712060
rect 675956 712058 675962 712060
rect 675956 711998 676292 712058
rect 675956 711996 675962 711998
rect 666277 711650 666343 711653
rect 666277 711648 676292 711650
rect 666277 711592 666282 711648
rect 666338 711592 676292 711648
rect 666277 711590 676292 711592
rect 666277 711587 666343 711590
rect 42149 711378 42215 711381
rect 42609 711378 42675 711381
rect 42149 711376 42675 711378
rect 42149 711320 42154 711376
rect 42210 711320 42614 711376
rect 42670 711320 42675 711376
rect 42149 711318 42675 711320
rect 42149 711315 42215 711318
rect 42609 711315 42675 711318
rect 683757 711242 683823 711245
rect 683757 711240 683836 711242
rect 683757 711184 683762 711240
rect 683818 711184 683836 711240
rect 683757 711182 683836 711184
rect 683757 711179 683823 711182
rect 42149 711106 42215 711109
rect 47577 711106 47643 711109
rect 42149 711104 47643 711106
rect 42149 711048 42154 711104
rect 42210 711048 47582 711104
rect 47638 711048 47643 711104
rect 42149 711046 47643 711048
rect 42149 711043 42215 711046
rect 47577 711043 47643 711046
rect 42885 710834 42951 710837
rect 45369 710834 45435 710837
rect 42885 710832 45435 710834
rect 42885 710776 42890 710832
rect 42946 710776 45374 710832
rect 45430 710776 45435 710832
rect 42885 710774 45435 710776
rect 42885 710771 42951 710774
rect 45369 710771 45435 710774
rect 672533 710834 672599 710837
rect 676029 710834 676095 710837
rect 672533 710832 676095 710834
rect 672533 710776 672538 710832
rect 672594 710776 676034 710832
rect 676090 710776 676095 710832
rect 672533 710774 676095 710776
rect 672533 710771 672599 710774
rect 676029 710771 676095 710774
rect 680997 710834 681063 710837
rect 680997 710832 681076 710834
rect 680997 710776 681002 710832
rect 681058 710776 681076 710832
rect 680997 710774 681076 710776
rect 680997 710771 681063 710774
rect 669270 710366 676292 710426
rect 652569 710290 652635 710293
rect 650164 710288 652635 710290
rect 650164 710232 652574 710288
rect 652630 710232 652635 710288
rect 650164 710230 652635 710232
rect 652569 710227 652635 710230
rect 667841 710290 667907 710293
rect 669270 710290 669330 710366
rect 667841 710288 669330 710290
rect 667841 710232 667846 710288
rect 667902 710232 669330 710288
rect 667841 710230 669330 710232
rect 667841 710227 667907 710230
rect 670141 710018 670207 710021
rect 670141 710016 676292 710018
rect 670141 709960 670146 710016
rect 670202 709960 676292 710016
rect 670141 709958 676292 709960
rect 670141 709955 670207 709958
rect 40902 709820 40908 709884
rect 40972 709882 40978 709884
rect 41781 709882 41847 709885
rect 40972 709880 41847 709882
rect 40972 709824 41786 709880
rect 41842 709824 41847 709880
rect 40972 709822 41847 709824
rect 40972 709820 40978 709822
rect 41781 709819 41847 709822
rect 676029 709610 676095 709613
rect 676029 709608 676292 709610
rect 676029 709552 676034 709608
rect 676090 709552 676292 709608
rect 676029 709550 676292 709552
rect 676029 709547 676095 709550
rect 40718 709412 40724 709476
rect 40788 709474 40794 709476
rect 672533 709474 672599 709477
rect 675845 709474 675911 709477
rect 40788 709414 42258 709474
rect 40788 709412 40794 709414
rect 42198 709205 42258 709414
rect 672533 709472 675911 709474
rect 672533 709416 672538 709472
rect 672594 709416 675850 709472
rect 675906 709416 675911 709472
rect 672533 709414 675911 709416
rect 672533 709411 672599 709414
rect 675845 709411 675911 709414
rect 42198 709200 42307 709205
rect 42198 709144 42246 709200
rect 42302 709144 42307 709200
rect 42198 709142 42307 709144
rect 42241 709139 42307 709142
rect 672993 709202 673059 709205
rect 672993 709200 676292 709202
rect 672993 709144 672998 709200
rect 673054 709144 676292 709200
rect 672993 709142 676292 709144
rect 672993 709139 673059 709142
rect 675845 708794 675911 708797
rect 675845 708792 676292 708794
rect 675845 708736 675850 708792
rect 675906 708736 676292 708792
rect 675845 708734 676292 708736
rect 675845 708731 675911 708734
rect 42057 708522 42123 708525
rect 42885 708522 42951 708525
rect 42057 708520 42951 708522
rect 42057 708464 42062 708520
rect 42118 708464 42890 708520
rect 42946 708464 42951 708520
rect 42057 708462 42951 708464
rect 42057 708459 42123 708462
rect 42885 708459 42951 708462
rect 683205 708386 683271 708389
rect 683205 708384 683284 708386
rect 683205 708328 683210 708384
rect 683266 708328 683284 708384
rect 683205 708326 683284 708328
rect 683205 708323 683271 708326
rect 670325 707978 670391 707981
rect 670325 707976 676292 707978
rect 670325 707920 670330 707976
rect 670386 707920 676292 707976
rect 670325 707918 676292 707920
rect 670325 707915 670391 707918
rect 42057 707842 42123 707845
rect 44173 707842 44239 707845
rect 42057 707840 44239 707842
rect 42057 707784 42062 707840
rect 42118 707784 44178 707840
rect 44234 707784 44239 707840
rect 42057 707782 44239 707784
rect 42057 707779 42123 707782
rect 44173 707779 44239 707782
rect 674414 707508 674420 707572
rect 674484 707570 674490 707572
rect 674484 707510 676292 707570
rect 674484 707508 674490 707510
rect 670509 707162 670575 707165
rect 670509 707160 676292 707162
rect 670509 707104 670514 707160
rect 670570 707104 676292 707160
rect 670509 707102 676292 707104
rect 670509 707099 670575 707102
rect 42057 706756 42123 706757
rect 42006 706754 42012 706756
rect 41966 706694 42012 706754
rect 42076 706752 42123 706756
rect 42118 706696 42123 706752
rect 42006 706692 42012 706694
rect 42076 706692 42123 706696
rect 42057 706691 42123 706692
rect 683389 706754 683455 706757
rect 683389 706752 683468 706754
rect 683389 706696 683394 706752
rect 683450 706696 683468 706752
rect 683389 706694 683468 706696
rect 683389 706691 683455 706694
rect 674465 706346 674531 706349
rect 674465 706344 676292 706346
rect 674465 706288 674470 706344
rect 674526 706288 676292 706344
rect 674465 706286 676292 706288
rect 674465 706283 674531 706286
rect 42241 705530 42307 705533
rect 44449 705530 44515 705533
rect 42241 705528 44515 705530
rect 42241 705472 42246 705528
rect 42302 705472 44454 705528
rect 44510 705472 44515 705528
rect 42241 705470 44515 705472
rect 42241 705467 42307 705470
rect 44449 705467 44515 705470
rect 671153 705530 671219 705533
rect 676262 705530 676322 705908
rect 671153 705528 676322 705530
rect 671153 705472 671158 705528
rect 671214 705500 676322 705528
rect 671214 705472 676292 705500
rect 671153 705470 676292 705472
rect 671153 705467 671219 705470
rect 667841 705122 667907 705125
rect 667841 705120 676292 705122
rect 667841 705064 667846 705120
rect 667902 705064 676292 705120
rect 667841 705062 676292 705064
rect 667841 705059 667907 705062
rect 40534 704244 40540 704308
rect 40604 704306 40610 704308
rect 41781 704306 41847 704309
rect 40604 704304 41847 704306
rect 40604 704248 41786 704304
rect 41842 704248 41847 704304
rect 40604 704246 41847 704248
rect 40604 704244 40610 704246
rect 41781 704243 41847 704246
rect 41454 702476 41460 702540
rect 41524 702538 41530 702540
rect 41524 702478 41706 702538
rect 41524 702476 41530 702478
rect 41646 702130 41706 702478
rect 41822 702340 41828 702404
rect 41892 702402 41898 702404
rect 42425 702402 42491 702405
rect 41892 702400 42491 702402
rect 41892 702344 42430 702400
rect 42486 702344 42491 702400
rect 41892 702342 42491 702344
rect 41892 702340 41898 702342
rect 42425 702339 42491 702342
rect 62113 702266 62179 702269
rect 62113 702264 64492 702266
rect 62113 702208 62118 702264
rect 62174 702208 64492 702264
rect 62113 702206 64492 702208
rect 62113 702203 62179 702206
rect 42241 702130 42307 702133
rect 41646 702128 42307 702130
rect 41646 702072 42246 702128
rect 42302 702072 42307 702128
rect 41646 702070 42307 702072
rect 42241 702067 42307 702070
rect 42057 701858 42123 701861
rect 42701 701858 42767 701861
rect 42057 701856 42767 701858
rect 42057 701800 42062 701856
rect 42118 701800 42706 701856
rect 42762 701800 42767 701856
rect 42057 701798 42767 701800
rect 42057 701795 42123 701798
rect 42701 701795 42767 701798
rect 41638 701524 41644 701588
rect 41708 701586 41714 701588
rect 42609 701586 42675 701589
rect 41708 701584 42675 701586
rect 41708 701528 42614 701584
rect 42670 701528 42675 701584
rect 41708 701526 42675 701528
rect 41708 701524 41714 701526
rect 42609 701523 42675 701526
rect 672533 698322 672599 698325
rect 675109 698322 675175 698325
rect 672533 698320 675175 698322
rect 672533 698264 672538 698320
rect 672594 698264 675114 698320
rect 675170 698264 675175 698320
rect 672533 698262 675175 698264
rect 672533 698259 672599 698262
rect 675109 698259 675175 698262
rect 673177 697234 673243 697237
rect 675109 697234 675175 697237
rect 673177 697232 675175 697234
rect 673177 697176 673182 697232
rect 673238 697176 675114 697232
rect 675170 697176 675175 697232
rect 673177 697174 675175 697176
rect 673177 697171 673243 697174
rect 675109 697171 675175 697174
rect 652385 696962 652451 696965
rect 650164 696960 652451 696962
rect 650164 696904 652390 696960
rect 652446 696904 652451 696960
rect 650164 696902 652451 696904
rect 652385 696899 652451 696902
rect 672349 696962 672415 696965
rect 675109 696962 675175 696965
rect 672349 696960 675175 696962
rect 672349 696904 672354 696960
rect 672410 696904 675114 696960
rect 675170 696904 675175 696960
rect 672349 696902 675175 696904
rect 672349 696899 672415 696902
rect 675109 696899 675175 696902
rect 675385 696828 675451 696829
rect 675334 696764 675340 696828
rect 675404 696826 675451 696828
rect 675404 696824 675496 696826
rect 675446 696768 675496 696824
rect 675404 696766 675496 696768
rect 675404 696764 675451 696766
rect 675385 696763 675451 696764
rect 675661 694378 675727 694381
rect 675661 694376 675954 694378
rect 675661 694320 675666 694376
rect 675722 694320 675954 694376
rect 675661 694318 675954 694320
rect 675661 694315 675727 694318
rect 675894 694106 675954 694318
rect 676806 694106 676812 694108
rect 675894 694046 676812 694106
rect 676806 694044 676812 694046
rect 676876 694044 676882 694108
rect 673545 693562 673611 693565
rect 675109 693562 675175 693565
rect 673545 693560 675175 693562
rect 673545 693504 673550 693560
rect 673606 693504 675114 693560
rect 675170 693504 675175 693560
rect 673545 693502 675175 693504
rect 673545 693499 673611 693502
rect 675109 693499 675175 693502
rect 668025 693290 668091 693293
rect 674925 693290 674991 693293
rect 668025 693288 674991 693290
rect 668025 693232 668030 693288
rect 668086 693232 674930 693288
rect 674986 693232 674991 693288
rect 668025 693230 674991 693232
rect 668025 693227 668091 693230
rect 674925 693227 674991 693230
rect 674414 692956 674420 693020
rect 674484 693018 674490 693020
rect 675109 693018 675175 693021
rect 674484 693016 675175 693018
rect 674484 692960 675114 693016
rect 675170 692960 675175 693016
rect 674484 692958 675175 692960
rect 674484 692956 674490 692958
rect 675109 692955 675175 692958
rect 35617 691386 35683 691389
rect 51717 691386 51783 691389
rect 35617 691384 51783 691386
rect 35617 691328 35622 691384
rect 35678 691328 51722 691384
rect 51778 691328 51783 691384
rect 35617 691326 51783 691328
rect 35617 691323 35683 691326
rect 51717 691323 51783 691326
rect 674097 690162 674163 690165
rect 675385 690162 675451 690165
rect 674097 690160 675451 690162
rect 674097 690104 674102 690160
rect 674158 690104 675390 690160
rect 675446 690104 675451 690160
rect 674097 690102 675451 690104
rect 674097 690099 674163 690102
rect 675385 690099 675451 690102
rect 62757 689482 62823 689485
rect 45510 689480 62823 689482
rect 45510 689424 62762 689480
rect 62818 689424 62823 689480
rect 45510 689422 62823 689424
rect 41413 689346 41479 689349
rect 45510 689346 45570 689422
rect 62757 689419 62823 689422
rect 41413 689344 45570 689346
rect 41413 689288 41418 689344
rect 41474 689288 45570 689344
rect 41413 689286 45570 689288
rect 663057 689346 663123 689349
rect 674925 689346 674991 689349
rect 663057 689344 674991 689346
rect 663057 689288 663062 689344
rect 663118 689288 674930 689344
rect 674986 689288 674991 689344
rect 663057 689286 674991 689288
rect 41413 689283 41479 689286
rect 663057 689283 663123 689286
rect 674925 689283 674991 689286
rect 62113 689210 62179 689213
rect 62113 689208 64492 689210
rect 62113 689152 62118 689208
rect 62174 689152 64492 689208
rect 62113 689150 64492 689152
rect 62113 689147 62179 689150
rect 670969 689074 671035 689077
rect 675109 689074 675175 689077
rect 670969 689072 675175 689074
rect 670969 689016 670974 689072
rect 671030 689016 675114 689072
rect 675170 689016 675175 689072
rect 670969 689014 675175 689016
rect 670969 689011 671035 689014
rect 675109 689011 675175 689014
rect 666277 688666 666343 688669
rect 674925 688666 674991 688669
rect 666277 688664 674991 688666
rect 666277 688608 666282 688664
rect 666338 688608 674930 688664
rect 674986 688608 674991 688664
rect 666277 688606 674991 688608
rect 666277 688603 666343 688606
rect 674925 688603 674991 688606
rect 54477 688122 54543 688125
rect 41492 688120 54543 688122
rect 41492 688064 54482 688120
rect 54538 688064 54543 688120
rect 41492 688062 54543 688064
rect 54477 688059 54543 688062
rect 35801 687714 35867 687717
rect 35788 687712 35867 687714
rect 35788 687656 35806 687712
rect 35862 687656 35867 687712
rect 35788 687654 35867 687656
rect 35801 687651 35867 687654
rect 35617 687306 35683 687309
rect 35604 687304 35683 687306
rect 35604 687248 35622 687304
rect 35678 687248 35683 687304
rect 35604 687246 35683 687248
rect 35617 687243 35683 687246
rect 674281 687306 674347 687309
rect 675293 687306 675359 687309
rect 674281 687304 675359 687306
rect 674281 687248 674286 687304
rect 674342 687248 675298 687304
rect 675354 687248 675359 687304
rect 674281 687246 675359 687248
rect 674281 687243 674347 687246
rect 675293 687243 675359 687246
rect 44633 686898 44699 686901
rect 41492 686896 44699 686898
rect 41492 686840 44638 686896
rect 44694 686840 44699 686896
rect 41492 686838 44699 686840
rect 44633 686835 44699 686838
rect 44357 686490 44423 686493
rect 41492 686488 44423 686490
rect 41492 686432 44362 686488
rect 44418 686432 44423 686488
rect 41492 686430 44423 686432
rect 44357 686427 44423 686430
rect 45185 686082 45251 686085
rect 41492 686080 45251 686082
rect 41492 686024 45190 686080
rect 45246 686024 45251 686080
rect 41492 686022 45251 686024
rect 45185 686019 45251 686022
rect 675334 685890 675340 685948
rect 675296 685884 675340 685890
rect 675404 685884 675410 685948
rect 675296 685830 675402 685884
rect 675109 685810 675175 685813
rect 675296 685810 675356 685830
rect 675109 685808 675356 685810
rect 675109 685752 675114 685808
rect 675170 685752 675356 685808
rect 675109 685750 675356 685752
rect 675109 685747 675175 685750
rect 45277 685674 45343 685677
rect 41492 685672 45343 685674
rect 41492 685616 45282 685672
rect 45338 685616 45343 685672
rect 41492 685614 45343 685616
rect 45277 685611 45343 685614
rect 45737 685266 45803 685269
rect 41492 685264 45803 685266
rect 41492 685208 45742 685264
rect 45798 685208 45803 685264
rect 41492 685206 45803 685208
rect 45737 685203 45803 685206
rect 670417 684994 670483 684997
rect 675477 684994 675543 684997
rect 670417 684992 675543 684994
rect 670417 684936 670422 684992
rect 670478 684936 675482 684992
rect 675538 684936 675543 684992
rect 670417 684934 675543 684936
rect 670417 684931 670483 684934
rect 675477 684931 675543 684934
rect 45921 684858 45987 684861
rect 41492 684856 45987 684858
rect 41492 684800 45926 684856
rect 45982 684800 45987 684856
rect 41492 684798 45987 684800
rect 45921 684795 45987 684798
rect 46105 684450 46171 684453
rect 41492 684448 46171 684450
rect 41492 684392 46110 684448
rect 46166 684392 46171 684448
rect 41492 684390 46171 684392
rect 46105 684387 46171 684390
rect 45737 684042 45803 684045
rect 41492 684040 45803 684042
rect 41492 683984 45742 684040
rect 45798 683984 45803 684040
rect 41492 683982 45803 683984
rect 45737 683979 45803 683982
rect 41822 683634 41828 683636
rect 41492 683574 41828 683634
rect 41822 683572 41828 683574
rect 41892 683572 41898 683636
rect 651833 683634 651899 683637
rect 650164 683632 651899 683634
rect 650164 683576 651838 683632
rect 651894 683576 651899 683632
rect 650164 683574 651899 683576
rect 651833 683571 651899 683574
rect 35801 683226 35867 683229
rect 35788 683224 35867 683226
rect 35788 683168 35806 683224
rect 35862 683168 35867 683224
rect 35788 683166 35867 683168
rect 35801 683163 35867 683166
rect 35433 682818 35499 682821
rect 35420 682816 35499 682818
rect 35420 682760 35438 682816
rect 35494 682760 35499 682816
rect 35420 682758 35499 682760
rect 35433 682755 35499 682758
rect 673729 682682 673795 682685
rect 683113 682682 683179 682685
rect 673729 682680 683179 682682
rect 673729 682624 673734 682680
rect 673790 682624 683118 682680
rect 683174 682624 683179 682680
rect 673729 682622 683179 682624
rect 673729 682619 673795 682622
rect 683113 682619 683179 682622
rect 35617 682410 35683 682413
rect 35604 682408 35683 682410
rect 35604 682352 35622 682408
rect 35678 682352 35683 682408
rect 35604 682350 35683 682352
rect 35617 682347 35683 682350
rect 674598 682348 674604 682412
rect 674668 682410 674674 682412
rect 683297 682410 683363 682413
rect 674668 682408 683363 682410
rect 674668 682352 683302 682408
rect 683358 682352 683363 682408
rect 674668 682350 683363 682352
rect 674668 682348 674674 682350
rect 683297 682347 683363 682350
rect 35801 682002 35867 682005
rect 35788 682000 35867 682002
rect 35788 681944 35806 682000
rect 35862 681944 35867 682000
rect 35788 681942 35867 681944
rect 35801 681939 35867 681942
rect 41689 681866 41755 681869
rect 42517 681866 42583 681869
rect 41689 681864 42583 681866
rect 41689 681808 41694 681864
rect 41750 681808 42522 681864
rect 42578 681808 42583 681864
rect 41689 681806 42583 681808
rect 41689 681803 41755 681806
rect 42517 681803 42583 681806
rect 32397 681594 32463 681597
rect 32397 681592 32476 681594
rect 32397 681536 32402 681592
rect 32458 681536 32476 681592
rect 32397 681534 32476 681536
rect 32397 681531 32463 681534
rect 31017 681186 31083 681189
rect 31004 681184 31083 681186
rect 31004 681128 31022 681184
rect 31078 681128 31083 681184
rect 31004 681126 31083 681128
rect 31017 681123 31083 681126
rect 674230 680988 674236 681052
rect 674300 681050 674306 681052
rect 683481 681050 683547 681053
rect 674300 681048 683547 681050
rect 674300 680992 683486 681048
rect 683542 680992 683547 681048
rect 674300 680990 683547 680992
rect 674300 680988 674306 680990
rect 683481 680987 683547 680990
rect 35157 680778 35223 680781
rect 35157 680776 35236 680778
rect 35157 680720 35162 680776
rect 35218 680720 35236 680776
rect 35157 680718 35236 680720
rect 35157 680715 35223 680718
rect 46105 680370 46171 680373
rect 41492 680368 46171 680370
rect 41492 680312 46110 680368
rect 46166 680312 46171 680368
rect 41492 680310 46171 680312
rect 46105 680307 46171 680310
rect 671797 680098 671863 680101
rect 675293 680098 675359 680101
rect 671797 680096 675359 680098
rect 671797 680040 671802 680096
rect 671858 680040 675298 680096
rect 675354 680040 675359 680096
rect 671797 680038 675359 680040
rect 671797 680035 671863 680038
rect 675293 680035 675359 680038
rect 42793 679962 42859 679965
rect 41492 679960 42859 679962
rect 41492 679904 42798 679960
rect 42854 679904 42859 679960
rect 41492 679902 42859 679904
rect 42793 679899 42859 679902
rect 44173 679554 44239 679557
rect 41492 679552 44239 679554
rect 41492 679496 44178 679552
rect 44234 679496 44239 679552
rect 41492 679494 44239 679496
rect 44173 679491 44239 679494
rect 44541 679146 44607 679149
rect 41492 679144 44607 679146
rect 41492 679088 44546 679144
rect 44602 679088 44607 679144
rect 41492 679086 44607 679088
rect 44541 679083 44607 679086
rect 40718 678928 40724 678992
rect 40788 678928 40794 678992
rect 40902 678928 40908 678992
rect 40972 678990 40978 678992
rect 40972 678930 41844 678990
rect 40972 678928 40978 678930
rect 40726 678708 40786 678928
rect 41784 678874 41844 678930
rect 41784 678814 42074 678874
rect 41781 678604 41847 678605
rect 41781 678602 41828 678604
rect 41736 678600 41828 678602
rect 41736 678544 41786 678600
rect 41736 678542 41828 678544
rect 41781 678540 41828 678542
rect 41892 678540 41898 678604
rect 41781 678539 41847 678540
rect 42014 678330 42074 678814
rect 41492 678270 42074 678330
rect 44725 677922 44791 677925
rect 41492 677920 44791 677922
rect 41492 677864 44730 677920
rect 44786 677864 44791 677920
rect 41492 677862 44791 677864
rect 44725 677859 44791 677862
rect 41278 677109 41338 677484
rect 41278 677104 41387 677109
rect 41278 677076 41326 677104
rect 41308 677048 41326 677076
rect 41382 677048 41387 677104
rect 41308 677046 41387 677048
rect 41321 677043 41387 677046
rect 43069 676698 43135 676701
rect 41492 676696 43135 676698
rect 41492 676640 43074 676696
rect 43130 676640 43135 676696
rect 41492 676638 43135 676640
rect 43069 676635 43135 676638
rect 62113 676154 62179 676157
rect 62113 676152 64492 676154
rect 62113 676096 62118 676152
rect 62174 676096 64492 676152
rect 62113 676094 64492 676096
rect 62113 676091 62179 676094
rect 31017 672754 31083 672757
rect 41822 672754 41828 672756
rect 31017 672752 41828 672754
rect 31017 672696 31022 672752
rect 31078 672696 41828 672752
rect 31017 672694 41828 672696
rect 31017 672691 31083 672694
rect 41822 672692 41828 672694
rect 41892 672692 41898 672756
rect 41321 672484 41387 672485
rect 41270 672420 41276 672484
rect 41340 672482 41387 672484
rect 41340 672480 41432 672482
rect 41382 672424 41432 672480
rect 41340 672422 41432 672424
rect 41340 672420 41387 672422
rect 41321 672419 41387 672420
rect 42149 672212 42215 672213
rect 42149 672210 42196 672212
rect 42104 672208 42196 672210
rect 42104 672152 42154 672208
rect 42104 672150 42196 672152
rect 42149 672148 42196 672150
rect 42260 672148 42266 672212
rect 42149 672147 42215 672148
rect 41321 671122 41387 671125
rect 42609 671122 42675 671125
rect 41321 671120 42675 671122
rect 41321 671064 41326 671120
rect 41382 671064 42614 671120
rect 42670 671064 42675 671120
rect 41321 671062 42675 671064
rect 41321 671059 41387 671062
rect 42609 671059 42675 671062
rect 667197 671122 667263 671125
rect 676262 671122 676322 671364
rect 667197 671120 676322 671122
rect 667197 671064 667202 671120
rect 667258 671064 676322 671120
rect 667197 671062 676322 671064
rect 667197 671059 667263 671062
rect 39665 670986 39731 670989
rect 40350 670986 40356 670988
rect 39665 670984 40356 670986
rect 39665 670928 39670 670984
rect 39726 670928 40356 670984
rect 39665 670926 40356 670928
rect 39665 670923 39731 670926
rect 40350 670924 40356 670926
rect 40420 670924 40426 670988
rect 41781 670714 41847 670717
rect 661677 670714 661743 670717
rect 676262 670714 676322 670956
rect 41781 670712 41890 670714
rect 41781 670656 41786 670712
rect 41842 670656 41890 670712
rect 41781 670651 41890 670656
rect 661677 670712 676322 670714
rect 661677 670656 661682 670712
rect 661738 670656 676322 670712
rect 661677 670654 676322 670656
rect 661677 670651 661743 670654
rect 41830 670309 41890 670651
rect 652385 670442 652451 670445
rect 650164 670440 652451 670442
rect 650164 670384 652390 670440
rect 652446 670384 652451 670440
rect 650164 670382 652451 670384
rect 652385 670379 652451 670382
rect 676814 670309 676874 670548
rect 41781 670304 41890 670309
rect 41781 670248 41786 670304
rect 41842 670248 41890 670304
rect 41781 670246 41890 670248
rect 671245 670306 671311 670309
rect 676489 670306 676555 670309
rect 671245 670304 676555 670306
rect 671245 670248 671250 670304
rect 671306 670248 676494 670304
rect 676550 670248 676555 670304
rect 671245 670246 676555 670248
rect 41781 670243 41847 670246
rect 671245 670243 671311 670246
rect 676489 670243 676555 670246
rect 676765 670304 676874 670309
rect 676765 670248 676770 670304
rect 676826 670248 676874 670304
rect 676765 670246 676874 670248
rect 676765 670243 676831 670246
rect 670785 669898 670851 669901
rect 676262 669898 676322 670140
rect 676489 669898 676555 669901
rect 670785 669896 676322 669898
rect 670785 669840 670790 669896
rect 670846 669840 676322 669896
rect 670785 669838 676322 669840
rect 676446 669896 676555 669898
rect 676446 669840 676494 669896
rect 676550 669840 676555 669896
rect 670785 669835 670851 669838
rect 676446 669835 676555 669840
rect 676446 669732 676506 669835
rect 671613 669490 671679 669493
rect 671613 669488 676322 669490
rect 671613 669432 671618 669488
rect 671674 669432 676322 669488
rect 671613 669430 676322 669432
rect 671613 669427 671679 669430
rect 42006 669292 42012 669356
rect 42076 669354 42082 669356
rect 48957 669354 49023 669357
rect 42076 669352 49023 669354
rect 42076 669296 48962 669352
rect 49018 669296 49023 669352
rect 42076 669294 49023 669296
rect 42076 669292 42082 669294
rect 48957 669291 49023 669294
rect 668577 669354 668643 669357
rect 668577 669352 671538 669354
rect 668577 669296 668582 669352
rect 668638 669296 671538 669352
rect 676262 669324 676322 669430
rect 668577 669294 671538 669296
rect 668577 669291 668643 669294
rect 671478 669218 671538 669294
rect 671478 669158 673470 669218
rect 41270 669020 41276 669084
rect 41340 669082 41346 669084
rect 41781 669082 41847 669085
rect 41340 669080 41847 669082
rect 41340 669024 41786 669080
rect 41842 669024 41847 669080
rect 41340 669022 41847 669024
rect 673410 669082 673470 669158
rect 676765 669082 676831 669085
rect 673410 669080 676831 669082
rect 673410 669024 676770 669080
rect 676826 669024 676831 669080
rect 673410 669022 676831 669024
rect 41340 669020 41346 669022
rect 41781 669019 41847 669022
rect 676765 669019 676831 669022
rect 42241 668948 42307 668949
rect 42190 668946 42196 668948
rect 42150 668886 42196 668946
rect 42260 668944 42307 668948
rect 42302 668888 42307 668944
rect 42190 668884 42196 668886
rect 42260 668884 42307 668888
rect 42241 668883 42307 668884
rect 674833 668810 674899 668813
rect 676262 668810 676322 668916
rect 674833 668808 676322 668810
rect 674833 668752 674838 668808
rect 674894 668752 676322 668808
rect 674833 668750 676322 668752
rect 674833 668747 674899 668750
rect 671429 668538 671495 668541
rect 671429 668536 676292 668538
rect 671429 668480 671434 668536
rect 671490 668480 676292 668536
rect 671429 668478 676292 668480
rect 671429 668475 671495 668478
rect 670233 668266 670299 668269
rect 674833 668266 674899 668269
rect 670233 668264 674899 668266
rect 670233 668208 670238 668264
rect 670294 668208 674838 668264
rect 674894 668208 674899 668264
rect 670233 668206 674899 668208
rect 670233 668203 670299 668206
rect 674833 668203 674899 668206
rect 40350 668068 40356 668132
rect 40420 668130 40426 668132
rect 40420 668070 42304 668130
rect 40420 668068 40426 668070
rect 42244 667861 42304 668070
rect 671521 667994 671587 667997
rect 676262 667994 676322 668100
rect 671521 667992 676322 667994
rect 671521 667936 671526 667992
rect 671582 667936 676322 667992
rect 671521 667934 676322 667936
rect 671521 667931 671587 667934
rect 42241 667856 42307 667861
rect 42241 667800 42246 667856
rect 42302 667800 42307 667856
rect 42241 667795 42307 667800
rect 41965 667724 42031 667725
rect 41965 667720 42012 667724
rect 42076 667722 42082 667724
rect 41965 667664 41970 667720
rect 41965 667660 42012 667664
rect 42076 667662 42122 667722
rect 42076 667660 42082 667662
rect 41965 667659 42031 667660
rect 42241 667586 42307 667589
rect 44173 667586 44239 667589
rect 42241 667584 44239 667586
rect 42241 667528 42246 667584
rect 42302 667528 44178 667584
rect 44234 667528 44239 667584
rect 42241 667526 44239 667528
rect 42241 667523 42307 667526
rect 44173 667523 44239 667526
rect 672165 667450 672231 667453
rect 676262 667450 676322 667692
rect 672165 667448 676322 667450
rect 672165 667392 672170 667448
rect 672226 667392 676322 667448
rect 672165 667390 676322 667392
rect 672165 667387 672231 667390
rect 40718 666980 40724 667044
rect 40788 667042 40794 667044
rect 42057 667042 42123 667045
rect 676262 667042 676322 667284
rect 683297 667042 683363 667045
rect 40788 667040 42123 667042
rect 40788 666984 42062 667040
rect 42118 666984 42123 667040
rect 40788 666982 42123 666984
rect 40788 666980 40794 666982
rect 42057 666979 42123 666982
rect 674790 666982 676322 667042
rect 683254 667040 683363 667042
rect 683254 666984 683302 667040
rect 683358 666984 683363 667040
rect 42057 666634 42123 666637
rect 42885 666634 42951 666637
rect 42057 666632 42951 666634
rect 42057 666576 42062 666632
rect 42118 666576 42890 666632
rect 42946 666576 42951 666632
rect 42057 666574 42951 666576
rect 42057 666571 42123 666574
rect 42885 666571 42951 666574
rect 670601 666634 670667 666637
rect 674790 666634 674850 666982
rect 683254 666979 683363 666984
rect 683254 666876 683314 666979
rect 670601 666632 674850 666634
rect 670601 666576 670606 666632
rect 670662 666576 674850 666632
rect 670601 666574 674850 666576
rect 670601 666571 670667 666574
rect 668761 666226 668827 666229
rect 676262 666226 676322 666468
rect 668761 666224 676322 666226
rect 668761 666168 668766 666224
rect 668822 666168 676322 666224
rect 668761 666166 676322 666168
rect 668761 666163 668827 666166
rect 667657 665954 667723 665957
rect 667657 665952 674850 665954
rect 667657 665896 667662 665952
rect 667718 665896 674850 665952
rect 667657 665894 674850 665896
rect 667657 665891 667723 665894
rect 674790 665818 674850 665894
rect 676446 665821 676506 666060
rect 674790 665758 676322 665818
rect 676446 665816 676555 665821
rect 676446 665760 676494 665816
rect 676550 665760 676555 665816
rect 676446 665758 676555 665760
rect 42057 665684 42123 665685
rect 42006 665682 42012 665684
rect 41966 665622 42012 665682
rect 42076 665680 42123 665684
rect 42118 665624 42123 665680
rect 42006 665620 42012 665622
rect 42076 665620 42123 665624
rect 42057 665619 42123 665620
rect 672993 665682 673059 665685
rect 672993 665680 674666 665682
rect 672993 665624 672998 665680
rect 673054 665624 674666 665680
rect 676262 665652 676322 665758
rect 676489 665755 676555 665758
rect 672993 665622 674666 665624
rect 672993 665619 673059 665622
rect 40534 665348 40540 665412
rect 40604 665410 40610 665412
rect 41781 665410 41847 665413
rect 40604 665408 41847 665410
rect 40604 665352 41786 665408
rect 41842 665352 41847 665408
rect 40604 665350 41847 665352
rect 40604 665348 40610 665350
rect 41781 665347 41847 665350
rect 666461 665410 666527 665413
rect 674606 665410 674666 665622
rect 666461 665408 674482 665410
rect 666461 665352 666466 665408
rect 666522 665352 674482 665408
rect 666461 665350 674482 665352
rect 674606 665350 676322 665410
rect 666461 665347 666527 665350
rect 42149 665136 42215 665141
rect 42149 665080 42154 665136
rect 42210 665080 42215 665136
rect 42149 665075 42215 665080
rect 42152 664869 42212 665075
rect 674422 665002 674482 665350
rect 676262 665244 676322 665350
rect 676489 665002 676555 665005
rect 674422 665000 676555 665002
rect 674422 664944 676494 665000
rect 676550 664944 676555 665000
rect 674422 664942 676555 664944
rect 676489 664939 676555 664942
rect 42149 664864 42215 664869
rect 42149 664808 42154 664864
rect 42210 664808 42215 664864
rect 42149 664803 42215 664808
rect 674833 664730 674899 664733
rect 676262 664730 676322 664836
rect 674833 664728 676322 664730
rect 674833 664672 674838 664728
rect 674894 664672 676322 664728
rect 674833 664670 676322 664672
rect 674833 664667 674899 664670
rect 671981 664458 672047 664461
rect 671981 664456 676292 664458
rect 671981 664400 671986 664456
rect 672042 664400 676292 664456
rect 671981 664398 676292 664400
rect 671981 664395 672047 664398
rect 668209 664186 668275 664189
rect 674833 664186 674899 664189
rect 683481 664186 683547 664189
rect 668209 664184 674899 664186
rect 668209 664128 668214 664184
rect 668270 664128 674838 664184
rect 674894 664128 674899 664184
rect 668209 664126 674899 664128
rect 668209 664123 668275 664126
rect 674833 664123 674899 664126
rect 683438 664184 683547 664186
rect 683438 664128 683486 664184
rect 683542 664128 683547 664184
rect 683438 664123 683547 664128
rect 41965 664052 42031 664053
rect 41965 664050 42012 664052
rect 41920 664048 42012 664050
rect 41920 663992 41970 664048
rect 41920 663990 42012 663992
rect 41965 663988 42012 663990
rect 42076 663988 42082 664052
rect 683438 664020 683498 664123
rect 41965 663987 42031 663988
rect 673361 663370 673427 663373
rect 676262 663370 676322 663612
rect 673361 663368 676322 663370
rect 673361 663312 673366 663368
rect 673422 663312 676322 663368
rect 673361 663310 676322 663312
rect 673361 663307 673427 663310
rect 62113 663098 62179 663101
rect 62113 663096 64492 663098
rect 62113 663040 62118 663096
rect 62174 663040 64492 663096
rect 62113 663038 64492 663040
rect 62113 663035 62179 663038
rect 42190 662900 42196 662964
rect 42260 662962 42266 662964
rect 42517 662962 42583 662965
rect 676262 662962 676322 663204
rect 683113 662962 683179 662965
rect 42260 662960 42583 662962
rect 42260 662904 42522 662960
rect 42578 662904 42583 662960
rect 42260 662902 42583 662904
rect 42260 662900 42266 662902
rect 42517 662899 42583 662902
rect 674422 662902 676322 662962
rect 683070 662960 683179 662962
rect 683070 662904 683118 662960
rect 683174 662904 683179 662960
rect 42701 662824 42767 662829
rect 42701 662768 42706 662824
rect 42762 662768 42767 662824
rect 42701 662763 42767 662768
rect 42333 662554 42399 662557
rect 42704 662554 42764 662763
rect 42333 662552 42764 662554
rect 42333 662496 42338 662552
rect 42394 662496 42764 662552
rect 42333 662494 42764 662496
rect 672809 662554 672875 662557
rect 674422 662554 674482 662902
rect 683070 662899 683179 662904
rect 683070 662796 683130 662899
rect 672809 662552 674482 662554
rect 672809 662496 672814 662552
rect 672870 662496 674482 662552
rect 672809 662494 674482 662496
rect 42333 662491 42399 662494
rect 672809 662491 672875 662494
rect 674833 662282 674899 662285
rect 676262 662282 676322 662388
rect 674833 662280 676322 662282
rect 674833 662224 674838 662280
rect 674894 662224 676322 662280
rect 674833 662222 676322 662224
rect 674833 662219 674899 662222
rect 669589 662010 669655 662013
rect 669589 662008 676292 662010
rect 669589 661952 669594 662008
rect 669650 661952 676292 662008
rect 669589 661950 676292 661952
rect 669589 661947 669655 661950
rect 668945 661738 669011 661741
rect 674833 661738 674899 661741
rect 668945 661736 674899 661738
rect 668945 661680 668950 661736
rect 669006 661680 674838 661736
rect 674894 661680 674899 661736
rect 668945 661678 674899 661680
rect 668945 661675 669011 661678
rect 674833 661675 674899 661678
rect 669129 661330 669195 661333
rect 676262 661330 676322 661572
rect 669129 661328 676322 661330
rect 669129 661272 669134 661328
rect 669190 661272 676322 661328
rect 669129 661270 676322 661272
rect 669129 661267 669195 661270
rect 42149 661058 42215 661061
rect 44541 661058 44607 661061
rect 42149 661056 44607 661058
rect 42149 661000 42154 661056
rect 42210 661000 44546 661056
rect 44602 661000 44607 661056
rect 42149 660998 44607 661000
rect 42149 660995 42215 660998
rect 44541 660995 44607 660998
rect 671981 661058 672047 661061
rect 676262 661058 676322 661164
rect 671981 661056 676322 661058
rect 671981 661000 671986 661056
rect 672042 661000 676322 661056
rect 671981 660998 676322 661000
rect 671981 660995 672047 660998
rect 42149 660514 42215 660517
rect 46105 660514 46171 660517
rect 42149 660512 46171 660514
rect 42149 660456 42154 660512
rect 42210 660456 46110 660512
rect 46166 660456 46171 660512
rect 42149 660454 46171 660456
rect 42149 660451 42215 660454
rect 46105 660451 46171 660454
rect 675385 660242 675451 660245
rect 676262 660242 676322 660756
rect 675385 660240 676322 660242
rect 675385 660184 675390 660240
rect 675446 660184 676322 660240
rect 675385 660182 676322 660184
rect 675385 660179 675451 660182
rect 673361 659970 673427 659973
rect 673361 659968 676292 659970
rect 673361 659912 673366 659968
rect 673422 659912 676292 659968
rect 673361 659910 676292 659912
rect 673361 659907 673427 659910
rect 41454 659772 41460 659836
rect 41524 659834 41530 659836
rect 42701 659834 42767 659837
rect 41524 659832 42767 659834
rect 41524 659776 42706 659832
rect 42762 659776 42767 659832
rect 41524 659774 42767 659776
rect 41524 659772 41530 659774
rect 42701 659771 42767 659774
rect 669773 659698 669839 659701
rect 675385 659698 675451 659701
rect 669773 659696 675451 659698
rect 669773 659640 669778 659696
rect 669834 659640 675390 659696
rect 675446 659640 675451 659696
rect 669773 659638 675451 659640
rect 669773 659635 669839 659638
rect 675385 659635 675451 659638
rect 42149 659020 42215 659021
rect 42149 659018 42196 659020
rect 42104 659016 42196 659018
rect 42104 658960 42154 659016
rect 42104 658958 42196 658960
rect 42149 658956 42196 658958
rect 42260 658956 42266 659020
rect 42149 658955 42215 658956
rect 41822 658548 41828 658612
rect 41892 658610 41898 658612
rect 42333 658610 42399 658613
rect 41892 658608 42399 658610
rect 41892 658552 42338 658608
rect 42394 658552 42399 658608
rect 41892 658550 42399 658552
rect 41892 658548 41898 658550
rect 42333 658547 42399 658550
rect 41638 658276 41644 658340
rect 41708 658338 41714 658340
rect 42517 658338 42583 658341
rect 41708 658336 42583 658338
rect 41708 658280 42522 658336
rect 42578 658280 42583 658336
rect 41708 658278 42583 658280
rect 41708 658276 41714 658278
rect 42517 658275 42583 658278
rect 42149 657386 42215 657389
rect 42701 657386 42767 657389
rect 42149 657384 42767 657386
rect 42149 657328 42154 657384
rect 42210 657328 42706 657384
rect 42762 657328 42767 657384
rect 42149 657326 42767 657328
rect 42149 657323 42215 657326
rect 42701 657323 42767 657326
rect 651649 657114 651715 657117
rect 650164 657112 651715 657114
rect 650164 657056 651654 657112
rect 651710 657056 651715 657112
rect 650164 657054 651715 657056
rect 651649 657051 651715 657054
rect 669221 654258 669287 654261
rect 675385 654258 675451 654261
rect 669221 654256 675451 654258
rect 669221 654200 669226 654256
rect 669282 654200 675390 654256
rect 675446 654200 675451 654256
rect 669221 654198 675451 654200
rect 669221 654195 669287 654198
rect 675385 654195 675451 654198
rect 675334 652836 675340 652900
rect 675404 652898 675410 652900
rect 675569 652898 675635 652901
rect 675404 652896 675635 652898
rect 675404 652840 675574 652896
rect 675630 652840 675635 652896
rect 675404 652838 675635 652840
rect 675404 652836 675410 652838
rect 675569 652835 675635 652838
rect 675569 651540 675635 651541
rect 675518 651538 675524 651540
rect 675478 651478 675524 651538
rect 675588 651536 675635 651540
rect 675630 651480 675635 651536
rect 675518 651476 675524 651478
rect 675588 651476 675635 651480
rect 675569 651475 675635 651476
rect 62113 650042 62179 650045
rect 62113 650040 64492 650042
rect 62113 649984 62118 650040
rect 62174 649984 64492 650040
rect 62113 649982 64492 649984
rect 62113 649979 62179 649982
rect 672717 648954 672783 648957
rect 675385 648954 675451 648957
rect 672717 648952 675451 648954
rect 672717 648896 672722 648952
rect 672778 648896 675390 648952
rect 675446 648896 675451 648952
rect 672717 648894 675451 648896
rect 672717 648891 672783 648894
rect 675385 648891 675451 648894
rect 672165 648682 672231 648685
rect 675109 648682 675175 648685
rect 672165 648680 675175 648682
rect 672165 648624 672170 648680
rect 672226 648624 675114 648680
rect 675170 648624 675175 648680
rect 672165 648622 675175 648624
rect 672165 648619 672231 648622
rect 675109 648619 675175 648622
rect 670785 647866 670851 647869
rect 675385 647866 675451 647869
rect 670785 647864 675451 647866
rect 670785 647808 670790 647864
rect 670846 647808 675390 647864
rect 675446 647808 675451 647864
rect 670785 647806 675451 647808
rect 670785 647803 670851 647806
rect 675385 647803 675451 647806
rect 35801 646778 35867 646781
rect 35801 646776 35910 646778
rect 35801 646720 35806 646776
rect 35862 646720 35910 646776
rect 35801 646715 35910 646720
rect 35850 646642 35910 646715
rect 51717 646642 51783 646645
rect 35850 646640 51783 646642
rect 35850 646584 51722 646640
rect 51778 646584 51783 646640
rect 35850 646582 51783 646584
rect 51717 646579 51783 646582
rect 675017 645828 675083 645829
rect 674966 645826 674972 645828
rect 674926 645766 674972 645826
rect 675036 645824 675083 645828
rect 675078 645768 675083 645824
rect 674966 645764 674972 645766
rect 675036 645764 675083 645768
rect 675017 645763 675083 645764
rect 669037 645554 669103 645557
rect 675109 645554 675175 645557
rect 669037 645552 675175 645554
rect 669037 645496 669042 645552
rect 669098 645496 675114 645552
rect 675170 645496 675175 645552
rect 669037 645494 675175 645496
rect 669037 645491 669103 645494
rect 675109 645491 675175 645494
rect 673821 645146 673887 645149
rect 675109 645146 675175 645149
rect 673821 645144 675175 645146
rect 673821 645088 673826 645144
rect 673882 645088 675114 645144
rect 675170 645088 675175 645144
rect 673821 645086 675175 645088
rect 673821 645083 673887 645086
rect 675109 645083 675175 645086
rect 35801 644738 35867 644741
rect 35758 644736 35867 644738
rect 35758 644680 35806 644736
rect 35862 644680 35867 644736
rect 35758 644675 35867 644680
rect 41462 644738 41522 644912
rect 53097 644738 53163 644741
rect 41462 644736 53163 644738
rect 41462 644680 53102 644736
rect 53158 644680 53163 644736
rect 41462 644678 53163 644680
rect 53097 644675 53163 644678
rect 35758 644504 35818 644675
rect 675753 644330 675819 644333
rect 676990 644330 676996 644332
rect 675753 644328 676996 644330
rect 675753 644272 675758 644328
rect 675814 644272 676996 644328
rect 675753 644270 676996 644272
rect 675753 644267 675819 644270
rect 676990 644268 676996 644270
rect 677060 644268 677066 644332
rect 41462 643922 41522 644096
rect 668393 643922 668459 643925
rect 675109 643922 675175 643925
rect 41462 643862 45570 643922
rect 41462 643650 41522 643688
rect 44357 643650 44423 643653
rect 41462 643648 44423 643650
rect 41462 643592 44362 643648
rect 44418 643592 44423 643648
rect 41462 643590 44423 643592
rect 44357 643587 44423 643590
rect 45093 643378 45159 643381
rect 41462 643376 45159 643378
rect 41462 643320 45098 643376
rect 45154 643320 45159 643376
rect 41462 643318 45159 643320
rect 41462 643280 41522 643318
rect 45093 643315 45159 643318
rect 45510 643242 45570 643862
rect 668393 643920 675175 643922
rect 668393 643864 668398 643920
rect 668454 643864 675114 643920
rect 675170 643864 675175 643920
rect 668393 643862 675175 643864
rect 668393 643859 668459 643862
rect 675109 643859 675175 643862
rect 651465 643786 651531 643789
rect 650164 643784 651531 643786
rect 650164 643728 651470 643784
rect 651526 643728 651531 643784
rect 650164 643726 651531 643728
rect 651465 643723 651531 643726
rect 669773 643514 669839 643517
rect 675293 643514 675359 643517
rect 669773 643512 675359 643514
rect 669773 643456 669778 643512
rect 669834 643456 675298 643512
rect 675354 643456 675359 643512
rect 669773 643454 675359 643456
rect 669773 643451 669839 643454
rect 675293 643451 675359 643454
rect 55857 643242 55923 643245
rect 45510 643240 55923 643242
rect 45510 643184 55862 643240
rect 55918 643184 55923 643240
rect 45510 643182 55923 643184
rect 55857 643179 55923 643182
rect 45277 643106 45343 643109
rect 41462 643104 45343 643106
rect 41462 643048 45282 643104
rect 45338 643048 45343 643104
rect 41462 643046 45343 643048
rect 41462 642872 41522 643046
rect 45277 643043 45343 643046
rect 45369 642562 45435 642565
rect 41462 642560 45435 642562
rect 41462 642504 45374 642560
rect 45430 642504 45435 642560
rect 41462 642502 45435 642504
rect 41462 642464 41522 642502
rect 45369 642499 45435 642502
rect 45921 642290 45987 642293
rect 41462 642288 45987 642290
rect 41462 642232 45926 642288
rect 45982 642232 45987 642288
rect 41462 642230 45987 642232
rect 41462 642056 41522 642230
rect 45921 642227 45987 642230
rect 674189 642156 674255 642157
rect 674189 642154 674236 642156
rect 674144 642152 674236 642154
rect 674144 642096 674194 642152
rect 674144 642094 674236 642096
rect 674189 642092 674236 642094
rect 674300 642092 674306 642156
rect 674189 642091 674255 642092
rect 674005 641746 674071 641749
rect 675293 641746 675359 641749
rect 674005 641744 675359 641746
rect 674005 641688 674010 641744
rect 674066 641688 675298 641744
rect 675354 641688 675359 641744
rect 674005 641686 675359 641688
rect 674005 641683 674071 641686
rect 675293 641683 675359 641686
rect 41781 641678 41847 641681
rect 41492 641676 41847 641678
rect 41492 641620 41786 641676
rect 41842 641620 41847 641676
rect 41492 641618 41847 641620
rect 41781 641615 41847 641618
rect 45737 641474 45803 641477
rect 41462 641472 45803 641474
rect 41462 641416 45742 641472
rect 45798 641416 45803 641472
rect 41462 641414 45803 641416
rect 41462 641240 41522 641414
rect 45737 641411 45803 641414
rect 41781 641202 41847 641205
rect 45921 641202 45987 641205
rect 41781 641200 45987 641202
rect 41781 641144 41786 641200
rect 41842 641144 45926 641200
rect 45982 641144 45987 641200
rect 41781 641142 45987 641144
rect 41781 641139 41847 641142
rect 45921 641139 45987 641142
rect 46105 640930 46171 640933
rect 41462 640928 46171 640930
rect 41462 640872 46110 640928
rect 46166 640872 46171 640928
rect 41462 640870 46171 640872
rect 41462 640832 41522 640870
rect 46105 640867 46171 640870
rect 674281 640794 674347 640797
rect 674598 640794 674604 640796
rect 674281 640792 674604 640794
rect 674281 640736 674286 640792
rect 674342 640736 674604 640792
rect 674281 640734 674604 640736
rect 674281 640731 674347 640734
rect 674598 640732 674604 640734
rect 674668 640732 674674 640796
rect 41454 640596 41460 640660
rect 41524 640596 41530 640660
rect 41462 640424 41522 640596
rect 674046 640460 674052 640524
rect 674116 640522 674122 640524
rect 675109 640522 675175 640525
rect 674116 640520 675175 640522
rect 674116 640464 675114 640520
rect 675170 640464 675175 640520
rect 674116 640462 675175 640464
rect 674116 640460 674122 640462
rect 675109 640459 675175 640462
rect 35574 639845 35634 640016
rect 35574 639840 35683 639845
rect 35574 639784 35622 639840
rect 35678 639784 35683 639840
rect 35574 639782 35683 639784
rect 35617 639779 35683 639782
rect 675150 639780 675156 639844
rect 675220 639842 675226 639844
rect 675385 639842 675451 639845
rect 675220 639840 675451 639842
rect 675220 639784 675390 639840
rect 675446 639784 675451 639840
rect 675220 639782 675451 639784
rect 675220 639780 675226 639782
rect 675385 639779 675451 639782
rect 35758 639437 35818 639608
rect 35758 639432 35867 639437
rect 35758 639376 35806 639432
rect 35862 639376 35867 639432
rect 35758 639374 35867 639376
rect 35801 639371 35867 639374
rect 41462 639026 41522 639200
rect 41638 639026 41644 639028
rect 41462 638966 41644 639026
rect 41638 638964 41644 638966
rect 41708 638964 41714 639028
rect 35758 638621 35818 638792
rect 668853 638754 668919 638757
rect 675477 638754 675543 638757
rect 668853 638752 675543 638754
rect 668853 638696 668858 638752
rect 668914 638696 675482 638752
rect 675538 638696 675543 638752
rect 668853 638694 675543 638696
rect 668853 638691 668919 638694
rect 675477 638691 675543 638694
rect 35758 638616 35867 638621
rect 35758 638560 35806 638616
rect 35862 638560 35867 638616
rect 35758 638558 35867 638560
rect 35801 638555 35867 638558
rect 32446 638213 32506 638384
rect 32397 638208 32506 638213
rect 32397 638152 32402 638208
rect 32458 638152 32506 638208
rect 32397 638150 32506 638152
rect 674833 638210 674899 638213
rect 675753 638210 675819 638213
rect 674833 638208 675819 638210
rect 674833 638152 674838 638208
rect 674894 638152 675758 638208
rect 675814 638152 675819 638208
rect 674833 638150 675819 638152
rect 32397 638147 32463 638150
rect 674833 638147 674899 638150
rect 675753 638147 675819 638150
rect 41462 637938 41522 637976
rect 47301 637938 47367 637941
rect 41462 637936 47367 637938
rect 41462 637880 47306 637936
rect 47362 637880 47367 637936
rect 41462 637878 47367 637880
rect 47301 637875 47367 637878
rect 674833 637938 674899 637941
rect 675150 637938 675156 637940
rect 674833 637936 675156 637938
rect 674833 637880 674838 637936
rect 674894 637880 675156 637936
rect 674833 637878 675156 637880
rect 674833 637875 674899 637878
rect 675150 637876 675156 637878
rect 675220 637876 675226 637940
rect 675334 637876 675340 637940
rect 675404 637938 675410 637940
rect 676029 637938 676095 637941
rect 675404 637936 676095 637938
rect 675404 637880 676034 637936
rect 676090 637880 676095 637936
rect 675404 637878 676095 637880
rect 675404 637876 675410 637878
rect 676029 637875 676095 637878
rect 47117 637666 47183 637669
rect 674925 637668 674991 637669
rect 674925 637666 674972 637668
rect 41462 637664 47183 637666
rect 41462 637608 47122 637664
rect 47178 637608 47183 637664
rect 41462 637606 47183 637608
rect 674880 637664 674972 637666
rect 674880 637608 674930 637664
rect 674880 637606 674972 637608
rect 41462 637568 41522 637606
rect 47117 637603 47183 637606
rect 674925 637604 674972 637606
rect 675036 637604 675042 637668
rect 675293 637666 675359 637669
rect 675518 637666 675524 637668
rect 675293 637664 675524 637666
rect 675293 637608 675298 637664
rect 675354 637608 675524 637664
rect 675293 637606 675524 637608
rect 674925 637603 674991 637604
rect 675293 637603 675359 637606
rect 675518 637604 675524 637606
rect 675588 637604 675594 637668
rect 41462 636986 41522 637160
rect 62113 637122 62179 637125
rect 62113 637120 64492 637122
rect 62113 637064 62118 637120
rect 62174 637064 64492 637120
rect 62113 637062 64492 637064
rect 62113 637059 62179 637062
rect 47761 636986 47827 636989
rect 41462 636984 47827 636986
rect 41462 636928 47766 636984
rect 47822 636928 47827 636984
rect 41462 636926 47827 636928
rect 47761 636923 47827 636926
rect 674230 636788 674236 636852
rect 674300 636850 674306 636852
rect 683389 636850 683455 636853
rect 674300 636848 683455 636850
rect 674300 636792 683394 636848
rect 683450 636792 683455 636848
rect 674300 636790 683455 636792
rect 674300 636788 674306 636790
rect 683389 636787 683455 636790
rect 41462 636578 41522 636752
rect 44173 636578 44239 636581
rect 41462 636576 44239 636578
rect 41462 636520 44178 636576
rect 44234 636520 44239 636576
rect 41462 636518 44239 636520
rect 44173 636515 44239 636518
rect 41462 636306 41522 636344
rect 44357 636306 44423 636309
rect 41462 636304 44423 636306
rect 41462 636248 44362 636304
rect 44418 636248 44423 636304
rect 41462 636246 44423 636248
rect 44357 636243 44423 636246
rect 674046 636244 674052 636308
rect 674116 636306 674122 636308
rect 674465 636306 674531 636309
rect 674116 636304 674531 636306
rect 674116 636248 674470 636304
rect 674526 636248 674531 636304
rect 674116 636246 674531 636248
rect 674116 636244 674122 636246
rect 674465 636243 674531 636246
rect 674925 636210 674991 636213
rect 674925 636208 675034 636210
rect 674925 636152 674930 636208
rect 674986 636170 675034 636208
rect 675477 636170 675543 636173
rect 674986 636168 675543 636170
rect 674986 636152 675482 636168
rect 674925 636147 675482 636152
rect 674974 636112 675482 636147
rect 675538 636112 675543 636168
rect 674974 636110 675543 636112
rect 675477 636107 675543 636110
rect 41462 635762 41522 635936
rect 44541 635762 44607 635765
rect 41462 635760 44607 635762
rect 41462 635704 44546 635760
rect 44602 635704 44607 635760
rect 41462 635702 44607 635704
rect 44541 635699 44607 635702
rect 674189 635762 674255 635765
rect 674189 635760 678990 635762
rect 674189 635704 674194 635760
rect 674250 635704 678990 635760
rect 674189 635702 678990 635704
rect 674189 635699 674255 635702
rect 41462 635354 41522 635528
rect 678930 635490 678990 635702
rect 683205 635490 683271 635493
rect 678930 635488 683271 635490
rect 678930 635432 683210 635488
rect 683266 635432 683271 635488
rect 678930 635430 683271 635432
rect 683205 635427 683271 635430
rect 44173 635354 44239 635357
rect 41462 635352 44239 635354
rect 41462 635296 44178 635352
rect 44234 635296 44239 635352
rect 41462 635294 44239 635296
rect 44173 635291 44239 635294
rect 40726 634948 40786 635120
rect 40718 634884 40724 634948
rect 40788 634884 40794 634948
rect 40542 634540 40602 634712
rect 40534 634476 40540 634540
rect 40604 634476 40610 634540
rect 41462 633858 41522 634304
rect 42333 633858 42399 633861
rect 41462 633856 42399 633858
rect 41462 633800 42338 633856
rect 42394 633800 42399 633856
rect 41462 633798 42399 633800
rect 42333 633795 42399 633798
rect 41462 633450 41522 633488
rect 45737 633450 45803 633453
rect 41462 633448 45803 633450
rect 41462 633392 45742 633448
rect 45798 633392 45803 633448
rect 41462 633390 45803 633392
rect 45737 633387 45803 633390
rect 674966 631348 674972 631412
rect 675036 631410 675042 631412
rect 675293 631410 675359 631413
rect 676029 631412 676095 631413
rect 676029 631410 676076 631412
rect 675036 631408 675359 631410
rect 675036 631352 675298 631408
rect 675354 631352 675359 631408
rect 675036 631350 675359 631352
rect 675984 631408 676076 631410
rect 675984 631352 676034 631408
rect 675984 631350 676076 631352
rect 675036 631348 675042 631350
rect 675293 631347 675359 631350
rect 676029 631348 676076 631350
rect 676140 631348 676146 631412
rect 676029 631347 676095 631348
rect 36537 630730 36603 630733
rect 41822 630730 41828 630732
rect 36537 630728 41828 630730
rect 36537 630672 36542 630728
rect 36598 630672 41828 630728
rect 36537 630670 41828 630672
rect 36537 630667 36603 630670
rect 41822 630668 41828 630670
rect 41892 630668 41898 630732
rect 651557 630594 651623 630597
rect 650164 630592 651623 630594
rect 650164 630536 651562 630592
rect 651618 630536 651623 630592
rect 650164 630534 651623 630536
rect 651557 630531 651623 630534
rect 661861 628554 661927 628557
rect 683113 628554 683179 628557
rect 661861 628552 683179 628554
rect 661861 628496 661866 628552
rect 661922 628496 683118 628552
rect 683174 628496 683179 628552
rect 661861 628494 683179 628496
rect 661861 628491 661927 628494
rect 683113 628491 683179 628494
rect 42190 626588 42196 626652
rect 42260 626650 42266 626652
rect 50337 626650 50403 626653
rect 42260 626648 50403 626650
rect 42260 626592 50342 626648
rect 50398 626592 50403 626648
rect 42260 626590 50403 626592
rect 42260 626588 42266 626590
rect 50337 626587 50403 626590
rect 665817 626106 665883 626109
rect 676262 626106 676322 626348
rect 665817 626104 676322 626106
rect 665817 626048 665822 626104
rect 665878 626048 676322 626104
rect 665817 626046 676322 626048
rect 665817 626043 665883 626046
rect 676262 625698 676322 625940
rect 683113 625698 683179 625701
rect 669270 625638 676322 625698
rect 683070 625696 683179 625698
rect 683070 625640 683118 625696
rect 683174 625640 683179 625696
rect 42006 625228 42012 625292
rect 42076 625290 42082 625292
rect 44081 625290 44147 625293
rect 42076 625288 44147 625290
rect 42076 625232 44086 625288
rect 44142 625232 44147 625288
rect 42076 625230 44147 625232
rect 42076 625228 42082 625230
rect 44081 625227 44147 625230
rect 660297 625290 660363 625293
rect 669270 625290 669330 625638
rect 683070 625635 683179 625640
rect 683070 625532 683130 625635
rect 660297 625288 669330 625290
rect 660297 625232 660302 625288
rect 660358 625232 669330 625288
rect 660297 625230 669330 625232
rect 660297 625227 660363 625230
rect 671245 625154 671311 625157
rect 671245 625152 676292 625154
rect 671245 625096 671250 625152
rect 671306 625096 676292 625152
rect 671245 625094 676292 625096
rect 671245 625091 671311 625094
rect 670601 624746 670667 624749
rect 670601 624744 676292 624746
rect 670601 624688 670606 624744
rect 670662 624688 676292 624744
rect 670601 624686 676292 624688
rect 670601 624683 670667 624686
rect 42149 624476 42215 624477
rect 42149 624474 42196 624476
rect 42104 624472 42196 624474
rect 42104 624416 42154 624472
rect 42104 624414 42196 624416
rect 42149 624412 42196 624414
rect 42260 624412 42266 624476
rect 42425 624474 42491 624477
rect 44357 624474 44423 624477
rect 42425 624472 44423 624474
rect 42425 624416 42430 624472
rect 42486 624416 44362 624472
rect 44418 624416 44423 624472
rect 42425 624414 44423 624416
rect 42149 624411 42215 624412
rect 42425 624411 42491 624414
rect 44357 624411 44423 624414
rect 670141 624338 670207 624341
rect 670141 624336 676292 624338
rect 670141 624280 670146 624336
rect 670202 624280 676292 624336
rect 670141 624278 676292 624280
rect 670141 624275 670207 624278
rect 62113 624066 62179 624069
rect 62113 624064 64492 624066
rect 62113 624008 62118 624064
rect 62174 624008 64492 624064
rect 62113 624006 64492 624008
rect 62113 624003 62179 624006
rect 669589 623930 669655 623933
rect 669589 623928 676292 623930
rect 669589 623872 669594 623928
rect 669650 623872 676292 623928
rect 669589 623870 676292 623872
rect 669589 623867 669655 623870
rect 40718 623732 40724 623796
rect 40788 623794 40794 623796
rect 42241 623794 42307 623797
rect 40788 623792 42307 623794
rect 40788 623736 42246 623792
rect 42302 623736 42307 623792
rect 40788 623734 42307 623736
rect 40788 623732 40794 623734
rect 42241 623731 42307 623734
rect 671521 623522 671587 623525
rect 671521 623520 676292 623522
rect 671521 623464 671526 623520
rect 671582 623464 676292 623520
rect 671521 623462 676292 623464
rect 671521 623459 671587 623462
rect 42057 623388 42123 623389
rect 42006 623324 42012 623388
rect 42076 623386 42123 623388
rect 42076 623384 42168 623386
rect 42118 623328 42168 623384
rect 42076 623326 42168 623328
rect 42076 623324 42123 623326
rect 42057 623323 42123 623324
rect 674649 623250 674715 623253
rect 675569 623250 675635 623253
rect 674649 623248 675635 623250
rect 674649 623192 674654 623248
rect 674710 623192 675574 623248
rect 675630 623192 675635 623248
rect 674649 623190 675635 623192
rect 674649 623187 674715 623190
rect 675569 623187 675635 623190
rect 676630 622845 676690 623084
rect 671153 622842 671219 622845
rect 675845 622842 675911 622845
rect 671153 622840 675911 622842
rect 671153 622784 671158 622840
rect 671214 622784 675850 622840
rect 675906 622784 675911 622840
rect 671153 622782 675911 622784
rect 671153 622779 671219 622782
rect 675845 622779 675911 622782
rect 676397 622842 676463 622845
rect 676397 622840 676506 622842
rect 676397 622784 676402 622840
rect 676458 622784 676506 622840
rect 676397 622779 676506 622784
rect 676630 622840 676739 622845
rect 676630 622784 676678 622840
rect 676734 622784 676739 622840
rect 676630 622782 676739 622784
rect 676673 622779 676739 622782
rect 676446 622676 676506 622779
rect 670417 622570 670483 622573
rect 676029 622570 676095 622573
rect 670417 622568 676095 622570
rect 670417 622512 670422 622568
rect 670478 622512 676034 622568
rect 676090 622512 676095 622568
rect 670417 622510 676095 622512
rect 670417 622507 670483 622510
rect 676029 622507 676095 622510
rect 671613 622298 671679 622301
rect 671613 622296 676292 622298
rect 671613 622240 671618 622296
rect 671674 622240 676292 622296
rect 671613 622238 676292 622240
rect 671613 622235 671679 622238
rect 682377 622026 682443 622029
rect 682334 622024 682443 622026
rect 682334 621968 682382 622024
rect 682438 621968 682443 622024
rect 682334 621963 682443 621968
rect 682334 621860 682394 621963
rect 672533 621618 672599 621621
rect 676489 621618 676555 621621
rect 672533 621616 676555 621618
rect 672533 621560 672538 621616
rect 672594 621560 676494 621616
rect 676550 621560 676555 621616
rect 672533 621558 676555 621560
rect 672533 621555 672599 621558
rect 676489 621555 676555 621558
rect 666277 621210 666343 621213
rect 676262 621210 676322 621452
rect 676489 621210 676555 621213
rect 666277 621208 676322 621210
rect 666277 621152 666282 621208
rect 666338 621152 676322 621208
rect 666277 621150 676322 621152
rect 676446 621208 676555 621210
rect 676446 621152 676494 621208
rect 676550 621152 676555 621208
rect 666277 621147 666343 621150
rect 676446 621147 676555 621152
rect 676446 621044 676506 621147
rect 42057 620938 42123 620941
rect 44173 620938 44239 620941
rect 42057 620936 44239 620938
rect 42057 620880 42062 620936
rect 42118 620880 44178 620936
rect 44234 620880 44239 620936
rect 42057 620878 44239 620880
rect 42057 620875 42123 620878
rect 44173 620875 44239 620878
rect 672349 620666 672415 620669
rect 672349 620664 676292 620666
rect 672349 620608 672354 620664
rect 672410 620608 676292 620664
rect 672349 620606 676292 620608
rect 672349 620603 672415 620606
rect 40534 620332 40540 620396
rect 40604 620394 40610 620396
rect 42701 620394 42767 620397
rect 40604 620392 42767 620394
rect 40604 620336 42706 620392
rect 42762 620336 42767 620392
rect 40604 620334 42767 620336
rect 40604 620332 40610 620334
rect 42701 620331 42767 620334
rect 671797 620394 671863 620397
rect 676489 620394 676555 620397
rect 671797 620392 676555 620394
rect 671797 620336 671802 620392
rect 671858 620336 676494 620392
rect 676550 620336 676555 620392
rect 671797 620334 676555 620336
rect 671797 620331 671863 620334
rect 676489 620331 676555 620334
rect 668025 619986 668091 619989
rect 676262 619986 676322 620228
rect 676489 619986 676555 619989
rect 668025 619984 676322 619986
rect 668025 619928 668030 619984
rect 668086 619928 676322 619984
rect 668025 619926 676322 619928
rect 676446 619984 676555 619986
rect 676446 619928 676494 619984
rect 676550 619928 676555 619984
rect 668025 619923 668091 619926
rect 676446 619923 676555 619928
rect 676446 619820 676506 619923
rect 42241 619714 42307 619717
rect 44541 619714 44607 619717
rect 42241 619712 44607 619714
rect 42241 619656 42246 619712
rect 42302 619656 44546 619712
rect 44602 619656 44607 619712
rect 42241 619654 44607 619656
rect 42241 619651 42307 619654
rect 44541 619651 44607 619654
rect 673177 619714 673243 619717
rect 673177 619712 675954 619714
rect 673177 619656 673182 619712
rect 673238 619656 675954 619712
rect 673177 619654 675954 619656
rect 673177 619651 673243 619654
rect 675894 619578 675954 619654
rect 675894 619518 676322 619578
rect 676262 619412 676322 619518
rect 676806 619108 676812 619172
rect 676876 619108 676882 619172
rect 676814 619004 676874 619108
rect 42517 618626 42583 618629
rect 47117 618626 47183 618629
rect 42517 618624 47183 618626
rect 42517 618568 42522 618624
rect 42578 618568 47122 618624
rect 47178 618568 47183 618624
rect 42517 618566 47183 618568
rect 42517 618563 42583 618566
rect 47117 618563 47183 618566
rect 673545 618626 673611 618629
rect 673545 618624 676292 618626
rect 673545 618568 673550 618624
rect 673606 618568 676292 618624
rect 673545 618566 676292 618568
rect 673545 618563 673611 618566
rect 41638 618292 41644 618356
rect 41708 618354 41714 618356
rect 42057 618354 42123 618357
rect 47761 618354 47827 618357
rect 683297 618354 683363 618357
rect 41708 618352 42123 618354
rect 41708 618296 42062 618352
rect 42118 618296 42123 618352
rect 41708 618294 42123 618296
rect 41708 618292 41714 618294
rect 42057 618291 42123 618294
rect 42520 618352 47827 618354
rect 42520 618296 47766 618352
rect 47822 618296 47827 618352
rect 42520 618294 47827 618296
rect 42241 617676 42307 617677
rect 42190 617674 42196 617676
rect 42150 617614 42196 617674
rect 42260 617672 42307 617676
rect 42302 617616 42307 617672
rect 42190 617612 42196 617614
rect 42260 617612 42307 617616
rect 42241 617611 42307 617612
rect 42057 617130 42123 617133
rect 42520 617130 42580 618294
rect 47761 618291 47827 618294
rect 683254 618352 683363 618354
rect 683254 618296 683302 618352
rect 683358 618296 683363 618352
rect 683254 618291 683363 618296
rect 683254 618188 683314 618291
rect 675569 617810 675635 617813
rect 675569 617808 676292 617810
rect 675569 617752 675574 617808
rect 675630 617752 676292 617808
rect 675569 617750 676292 617752
rect 675569 617747 675635 617750
rect 674414 617340 674420 617404
rect 674484 617402 674490 617404
rect 674484 617342 676292 617402
rect 674484 617340 674490 617342
rect 651465 617266 651531 617269
rect 650164 617264 651531 617266
rect 650164 617208 651470 617264
rect 651526 617208 651531 617264
rect 650164 617206 651531 617208
rect 651465 617203 651531 617206
rect 683481 617130 683547 617133
rect 42057 617128 42580 617130
rect 42057 617072 42062 617128
rect 42118 617072 42580 617128
rect 42057 617070 42580 617072
rect 683438 617128 683547 617130
rect 683438 617072 683486 617128
rect 683542 617072 683547 617128
rect 42057 617067 42123 617070
rect 683438 617067 683547 617072
rect 683438 616964 683498 617067
rect 42057 616586 42123 616589
rect 42517 616586 42583 616589
rect 42057 616584 42583 616586
rect 42057 616528 42062 616584
rect 42118 616528 42522 616584
rect 42578 616528 42583 616584
rect 42057 616526 42583 616528
rect 42057 616523 42123 616526
rect 42517 616523 42583 616526
rect 670969 616586 671035 616589
rect 670969 616584 676292 616586
rect 670969 616528 670974 616584
rect 671030 616528 676292 616584
rect 670969 616526 676292 616528
rect 670969 616523 671035 616526
rect 42885 616178 42951 616181
rect 44081 616178 44147 616181
rect 42885 616176 44147 616178
rect 42885 616120 42890 616176
rect 42946 616120 44086 616176
rect 44142 616120 44147 616176
rect 42885 616118 44147 616120
rect 42885 616115 42951 616118
rect 44081 616115 44147 616118
rect 673862 616116 673868 616180
rect 673932 616178 673938 616180
rect 673932 616118 676292 616178
rect 673932 616116 673938 616118
rect 42149 615908 42215 615909
rect 42149 615906 42196 615908
rect 42104 615904 42196 615906
rect 42104 615848 42154 615904
rect 42104 615846 42196 615848
rect 42149 615844 42196 615846
rect 42260 615844 42266 615908
rect 42149 615843 42215 615844
rect 670141 615770 670207 615773
rect 670141 615768 676292 615770
rect 670141 615712 670146 615768
rect 670202 615740 676292 615768
rect 670202 615712 676322 615740
rect 670141 615710 676322 615712
rect 670141 615707 670207 615710
rect 47301 615634 47367 615637
rect 42934 615632 47367 615634
rect 42934 615576 47306 615632
rect 47362 615576 47367 615632
rect 42934 615574 47367 615576
rect 41822 615436 41828 615500
rect 41892 615498 41898 615500
rect 42609 615498 42675 615501
rect 41892 615496 42675 615498
rect 41892 615440 42614 615496
rect 42670 615440 42675 615496
rect 41892 615438 42675 615440
rect 41892 615436 41898 615438
rect 42609 615435 42675 615438
rect 42241 615226 42307 615229
rect 42934 615226 42994 615574
rect 47301 615571 47367 615574
rect 676262 615332 676322 615710
rect 42241 615224 42994 615226
rect 42241 615168 42246 615224
rect 42302 615168 42994 615224
rect 42241 615166 42994 615168
rect 42241 615163 42307 615166
rect 670601 614954 670667 614957
rect 670601 614952 676292 614954
rect 670601 614896 670606 614952
rect 670662 614896 676292 614952
rect 670601 614894 676292 614896
rect 670601 614891 670667 614894
rect 41454 614076 41460 614140
rect 41524 614138 41530 614140
rect 41781 614138 41847 614141
rect 41524 614136 41847 614138
rect 41524 614080 41786 614136
rect 41842 614080 41847 614136
rect 41524 614078 41847 614080
rect 41524 614076 41530 614078
rect 41781 614075 41847 614078
rect 43069 611962 43135 611965
rect 43924 611962 43990 611965
rect 43069 611960 43990 611962
rect 43069 611904 43074 611960
rect 43130 611904 43929 611960
rect 43985 611904 43990 611960
rect 43069 611902 43990 611904
rect 43069 611899 43135 611902
rect 43924 611899 43990 611902
rect 42517 611010 42583 611013
rect 44495 611010 44561 611013
rect 42517 611008 44561 611010
rect 42517 610952 42522 611008
rect 42578 610952 44500 611008
rect 44556 610952 44561 611008
rect 42517 610950 44561 610952
rect 42517 610947 42583 610950
rect 44495 610947 44561 610950
rect 62113 611010 62179 611013
rect 62113 611008 64492 611010
rect 62113 610952 62118 611008
rect 62174 610952 64492 611008
rect 62113 610950 64492 610952
rect 62113 610947 62179 610950
rect 672441 608698 672507 608701
rect 674833 608698 674899 608701
rect 672441 608696 674899 608698
rect 672441 608640 672446 608696
rect 672502 608640 674838 608696
rect 674894 608640 674899 608696
rect 672441 608638 674899 608640
rect 672441 608635 672507 608638
rect 674833 608635 674899 608638
rect 675477 607884 675543 607885
rect 675477 607880 675524 607884
rect 675588 607882 675594 607884
rect 675477 607824 675482 607880
rect 675477 607820 675524 607824
rect 675588 607822 675634 607882
rect 675588 607820 675594 607822
rect 675477 607819 675543 607820
rect 672441 607338 672507 607341
rect 675293 607338 675359 607341
rect 672441 607336 675359 607338
rect 672441 607280 672446 607336
rect 672502 607280 675298 607336
rect 675354 607280 675359 607336
rect 672441 607278 675359 607280
rect 672441 607275 672507 607278
rect 675293 607275 675359 607278
rect 674833 607066 674899 607069
rect 675293 607066 675359 607069
rect 674833 607064 675359 607066
rect 674833 607008 674838 607064
rect 674894 607008 675298 607064
rect 675354 607008 675359 607064
rect 674833 607006 675359 607008
rect 674833 607003 674899 607006
rect 675293 607003 675359 607006
rect 672809 604890 672875 604893
rect 675293 604890 675359 604893
rect 672809 604888 675359 604890
rect 672809 604832 672814 604888
rect 672870 604832 675298 604888
rect 675354 604832 675359 604888
rect 672809 604830 675359 604832
rect 672809 604827 672875 604830
rect 675293 604827 675359 604830
rect 672993 604346 673059 604349
rect 675293 604346 675359 604349
rect 672993 604344 675359 604346
rect 672993 604288 672998 604344
rect 673054 604288 675298 604344
rect 675354 604288 675359 604344
rect 672993 604286 675359 604288
rect 672993 604283 673059 604286
rect 675293 604283 675359 604286
rect 673637 604074 673703 604077
rect 675385 604074 675451 604077
rect 673637 604072 675451 604074
rect 673637 604016 673642 604072
rect 673698 604016 675390 604072
rect 675446 604016 675451 604072
rect 673637 604014 675451 604016
rect 673637 604011 673703 604014
rect 675385 604011 675451 604014
rect 651465 603938 651531 603941
rect 650164 603936 651531 603938
rect 650164 603880 651470 603936
rect 651526 603880 651531 603936
rect 650164 603878 651531 603880
rect 651465 603875 651531 603878
rect 667657 603394 667723 603397
rect 675293 603394 675359 603397
rect 667657 603392 675359 603394
rect 667657 603336 667662 603392
rect 667718 603336 675298 603392
rect 675354 603336 675359 603392
rect 667657 603334 675359 603336
rect 667657 603331 667723 603334
rect 675293 603331 675359 603334
rect 674230 602924 674236 602988
rect 674300 602986 674306 602988
rect 675477 602986 675543 602989
rect 674300 602984 675543 602986
rect 674300 602928 675482 602984
rect 675538 602928 675543 602984
rect 674300 602926 675543 602928
rect 674300 602924 674306 602926
rect 675477 602923 675543 602926
rect 51717 601762 51783 601765
rect 41492 601760 51783 601762
rect 41492 601704 51722 601760
rect 51778 601704 51783 601760
rect 41492 601702 51783 601704
rect 51717 601699 51783 601702
rect 668393 601762 668459 601765
rect 674833 601762 674899 601765
rect 668393 601760 674899 601762
rect 668393 601704 668398 601760
rect 668454 601704 674838 601760
rect 674894 601704 674899 601760
rect 668393 601702 674899 601704
rect 668393 601699 668459 601702
rect 674833 601699 674899 601702
rect 48957 601354 49023 601357
rect 41492 601352 49023 601354
rect 41492 601296 48962 601352
rect 49018 601296 49023 601352
rect 41492 601294 49023 601296
rect 48957 601291 49023 601294
rect 54477 600946 54543 600949
rect 41492 600944 54543 600946
rect 41492 600888 54482 600944
rect 54538 600888 54543 600944
rect 41492 600886 54543 600888
rect 54477 600883 54543 600886
rect 45093 600538 45159 600541
rect 41492 600536 45159 600538
rect 41492 600480 45098 600536
rect 45154 600480 45159 600536
rect 41492 600478 45159 600480
rect 45093 600475 45159 600478
rect 674833 600538 674899 600541
rect 675293 600538 675359 600541
rect 674833 600536 675359 600538
rect 674833 600480 674838 600536
rect 674894 600480 675298 600536
rect 675354 600480 675359 600536
rect 674833 600478 675359 600480
rect 674833 600475 674899 600478
rect 675293 600475 675359 600478
rect 44633 600130 44699 600133
rect 41492 600128 44699 600130
rect 41492 600072 44638 600128
rect 44694 600072 44699 600128
rect 41492 600070 44699 600072
rect 44633 600067 44699 600070
rect 674649 599858 674715 599861
rect 675477 599858 675543 599861
rect 674649 599856 675543 599858
rect 674649 599800 674654 599856
rect 674710 599800 675482 599856
rect 675538 599800 675543 599856
rect 674649 599798 675543 599800
rect 674649 599795 674715 599798
rect 675477 599795 675543 599798
rect 45369 599722 45435 599725
rect 41492 599720 45435 599722
rect 41492 599664 45374 599720
rect 45430 599664 45435 599720
rect 41492 599662 45435 599664
rect 45369 599659 45435 599662
rect 660297 599586 660363 599589
rect 660297 599584 663810 599586
rect 660297 599528 660302 599584
rect 660358 599528 663810 599584
rect 660297 599526 663810 599528
rect 660297 599523 660363 599526
rect 44817 599314 44883 599317
rect 41492 599312 44883 599314
rect 41492 599256 44822 599312
rect 44878 599256 44883 599312
rect 41492 599254 44883 599256
rect 663750 599314 663810 599526
rect 675293 599314 675359 599317
rect 663750 599312 675359 599314
rect 663750 599256 675298 599312
rect 675354 599256 675359 599312
rect 663750 599254 675359 599256
rect 44817 599251 44883 599254
rect 675293 599251 675359 599254
rect 45921 598906 45987 598909
rect 41492 598904 45987 598906
rect 41492 598848 45926 598904
rect 45982 598848 45987 598904
rect 41492 598846 45987 598848
rect 45921 598843 45987 598846
rect 45001 598498 45067 598501
rect 675477 598498 675543 598501
rect 41492 598496 45067 598498
rect 41492 598440 45006 598496
rect 45062 598440 45067 598496
rect 41492 598438 45067 598440
rect 45001 598435 45067 598438
rect 673870 598496 675543 598498
rect 673870 598440 675482 598496
rect 675538 598440 675543 598496
rect 673870 598438 675543 598440
rect 673870 598365 673930 598438
rect 675477 598435 675543 598438
rect 673821 598360 673930 598365
rect 673821 598304 673826 598360
rect 673882 598304 673930 598360
rect 673821 598302 673930 598304
rect 673821 598299 673887 598302
rect 46105 598090 46171 598093
rect 41492 598088 46171 598090
rect 41492 598032 46110 598088
rect 46166 598032 46171 598088
rect 41492 598030 46171 598032
rect 46105 598027 46171 598030
rect 62113 597954 62179 597957
rect 62113 597952 64492 597954
rect 62113 597896 62118 597952
rect 62174 597896 64492 597952
rect 62113 597894 64492 597896
rect 62113 597891 62179 597894
rect 41492 597622 42994 597682
rect 41822 597274 41828 597276
rect 41492 597214 41828 597274
rect 41822 597212 41828 597214
rect 41892 597212 41898 597276
rect 42934 597005 42994 597622
rect 674189 597410 674255 597413
rect 675477 597410 675543 597413
rect 674189 597408 675543 597410
rect 674189 597352 674194 597408
rect 674250 597352 675482 597408
rect 675538 597352 675543 597408
rect 674189 597350 675543 597352
rect 674189 597347 674255 597350
rect 675477 597347 675543 597350
rect 42934 597000 43043 597005
rect 42934 596944 42982 597000
rect 43038 596944 43043 597000
rect 42934 596942 43043 596944
rect 42977 596939 43043 596942
rect 42149 596866 42215 596869
rect 41492 596864 42215 596866
rect 41492 596808 42154 596864
rect 42210 596808 42215 596864
rect 41492 596806 42215 596808
rect 42149 596803 42215 596806
rect 41822 596458 41828 596460
rect 41492 596398 41828 596458
rect 41822 596396 41828 596398
rect 41892 596396 41898 596460
rect 41229 596050 41295 596053
rect 41229 596048 41308 596050
rect 41229 595992 41234 596048
rect 41290 595992 41308 596048
rect 41229 595990 41308 595992
rect 41229 595987 41295 595990
rect 33041 595642 33107 595645
rect 33028 595640 33107 595642
rect 33028 595584 33046 595640
rect 33102 595584 33107 595640
rect 33028 595582 33107 595584
rect 33041 595579 33107 595582
rect 675385 595372 675451 595373
rect 675334 595370 675340 595372
rect 675294 595310 675340 595370
rect 675404 595368 675451 595372
rect 675446 595312 675451 595368
rect 675334 595308 675340 595310
rect 675404 595308 675451 595312
rect 675385 595307 675451 595308
rect 35157 595234 35223 595237
rect 35157 595232 35236 595234
rect 35157 595176 35162 595232
rect 35218 595176 35236 595232
rect 35157 595174 35236 595176
rect 35157 595171 35223 595174
rect 40677 594826 40743 594829
rect 671337 594826 671403 594829
rect 675477 594826 675543 594829
rect 40677 594824 40756 594826
rect 40677 594768 40682 594824
rect 40738 594768 40756 594824
rect 40677 594766 40756 594768
rect 671337 594824 675543 594826
rect 671337 594768 671342 594824
rect 671398 594768 675482 594824
rect 675538 594768 675543 594824
rect 671337 594766 675543 594768
rect 40677 594763 40743 594766
rect 671337 594763 671403 594766
rect 675477 594763 675543 594766
rect 41689 594554 41755 594557
rect 42609 594554 42675 594557
rect 41689 594552 42675 594554
rect 41689 594496 41694 594552
rect 41750 594496 42614 594552
rect 42670 594496 42675 594552
rect 41689 594494 42675 594496
rect 41689 594491 41755 594494
rect 42609 594491 42675 594494
rect 31017 594418 31083 594421
rect 31004 594416 31083 594418
rect 31004 594360 31022 594416
rect 31078 594360 31083 594416
rect 31004 594358 31083 594360
rect 31017 594355 31083 594358
rect 42793 594010 42859 594013
rect 41492 594008 42859 594010
rect 41492 593952 42798 594008
rect 42854 593952 42859 594008
rect 41492 593950 42859 593952
rect 42793 593947 42859 593950
rect 41781 593602 41847 593605
rect 41492 593600 41847 593602
rect 41492 593544 41786 593600
rect 41842 593544 41847 593600
rect 41492 593542 41847 593544
rect 41781 593539 41847 593542
rect 667013 593466 667079 593469
rect 675385 593466 675451 593469
rect 667013 593464 675451 593466
rect 667013 593408 667018 593464
rect 667074 593408 675390 593464
rect 675446 593408 675451 593464
rect 667013 593406 675451 593408
rect 667013 593403 667079 593406
rect 675385 593403 675451 593406
rect 40493 593194 40559 593197
rect 675569 593196 675635 593197
rect 675518 593194 675524 593196
rect 40493 593192 40572 593194
rect 40493 593136 40498 593192
rect 40554 593136 40572 593192
rect 40493 593134 40572 593136
rect 675478 593134 675524 593194
rect 675588 593192 675635 593196
rect 675630 593136 675635 593192
rect 40493 593131 40559 593134
rect 675518 593132 675524 593134
rect 675588 593132 675635 593136
rect 675569 593131 675635 593132
rect 675150 592860 675156 592924
rect 675220 592922 675226 592924
rect 676029 592922 676095 592925
rect 675220 592920 676095 592922
rect 675220 592864 676034 592920
rect 676090 592864 676095 592920
rect 675220 592862 676095 592864
rect 675220 592860 675226 592862
rect 676029 592859 676095 592862
rect 41781 592786 41847 592789
rect 41492 592784 41847 592786
rect 41492 592728 41786 592784
rect 41842 592728 41847 592784
rect 41492 592726 41847 592728
rect 41781 592723 41847 592726
rect 674833 592650 674899 592653
rect 675845 592650 675911 592653
rect 683389 592650 683455 592653
rect 674833 592648 675911 592650
rect 674833 592592 674838 592648
rect 674894 592592 675850 592648
rect 675906 592592 675911 592648
rect 674833 592590 675911 592592
rect 674833 592587 674899 592590
rect 675845 592587 675911 592590
rect 678930 592648 683455 592650
rect 678930 592592 683394 592648
rect 683450 592592 683455 592648
rect 678930 592590 683455 592592
rect 41781 592378 41847 592381
rect 41492 592376 41847 592378
rect 41492 592320 41786 592376
rect 41842 592320 41847 592376
rect 41492 592318 41847 592320
rect 41781 592315 41847 592318
rect 673453 592378 673519 592381
rect 678930 592378 678990 592590
rect 683389 592587 683455 592590
rect 673453 592376 678990 592378
rect 673453 592320 673458 592376
rect 673514 592320 678990 592376
rect 673453 592318 678990 592320
rect 673453 592315 673519 592318
rect 675293 592108 675359 592109
rect 675293 592106 675340 592108
rect 675248 592104 675340 592106
rect 675248 592048 675298 592104
rect 675248 592046 675340 592048
rect 675293 592044 675340 592046
rect 675404 592044 675410 592108
rect 675293 592043 675359 592044
rect 44449 591970 44515 591973
rect 41492 591968 44515 591970
rect 41492 591912 44454 591968
rect 44510 591912 44515 591968
rect 41492 591910 44515 591912
rect 44449 591907 44515 591910
rect 676070 591636 676076 591700
rect 676140 591698 676146 591700
rect 680997 591698 681063 591701
rect 676140 591696 681063 591698
rect 676140 591640 681002 591696
rect 681058 591640 681063 591696
rect 676140 591638 681063 591640
rect 676140 591636 676146 591638
rect 680997 591635 681063 591638
rect 43437 591562 43503 591565
rect 41492 591560 43503 591562
rect 41492 591504 43442 591560
rect 43498 591504 43503 591560
rect 41492 591502 43503 591504
rect 43437 591499 43503 591502
rect 674005 591290 674071 591293
rect 683665 591290 683731 591293
rect 674005 591288 683731 591290
rect 674005 591232 674010 591288
rect 674066 591232 683670 591288
rect 683726 591232 683731 591288
rect 674005 591230 683731 591232
rect 674005 591227 674071 591230
rect 683665 591227 683731 591230
rect 39990 590749 40050 591124
rect 39941 590744 40050 590749
rect 652385 590746 652451 590749
rect 39941 590688 39946 590744
rect 40002 590716 40050 590744
rect 650164 590744 652451 590746
rect 40002 590688 40020 590716
rect 39941 590686 40020 590688
rect 650164 590688 652390 590744
rect 652446 590688 652451 590744
rect 650164 590686 652451 590688
rect 39941 590683 40007 590686
rect 652385 590683 652451 590686
rect 43621 590338 43687 590341
rect 41492 590336 43687 590338
rect 41492 590280 43626 590336
rect 43682 590280 43687 590336
rect 41492 590278 43687 590280
rect 43621 590275 43687 590278
rect 674465 589930 674531 589933
rect 683849 589930 683915 589933
rect 674465 589928 683915 589930
rect 674465 589872 674470 589928
rect 674526 589872 683854 589928
rect 683910 589872 683915 589928
rect 674465 589870 683915 589872
rect 674465 589867 674531 589870
rect 683849 589867 683915 589870
rect 40493 589658 40559 589661
rect 40718 589658 40724 589660
rect 40493 589656 40724 589658
rect 40493 589600 40498 589656
rect 40554 589600 40724 589656
rect 40493 589598 40724 589600
rect 40493 589595 40559 589598
rect 40718 589596 40724 589598
rect 40788 589596 40794 589660
rect 40902 589460 40908 589524
rect 40972 589522 40978 589524
rect 41781 589522 41847 589525
rect 40972 589520 41847 589522
rect 40972 589464 41786 589520
rect 41842 589464 41847 589520
rect 40972 589462 41847 589464
rect 40972 589460 40978 589462
rect 41781 589459 41847 589462
rect 40309 589386 40375 589389
rect 40534 589386 40540 589388
rect 40309 589384 40540 589386
rect 40309 589328 40314 589384
rect 40370 589328 40540 589384
rect 40309 589326 40540 589328
rect 40309 589323 40375 589326
rect 40534 589324 40540 589326
rect 40604 589324 40610 589388
rect 42057 586804 42123 586805
rect 42006 586802 42012 586804
rect 41966 586742 42012 586802
rect 42076 586800 42123 586804
rect 42118 586744 42123 586800
rect 42006 586740 42012 586742
rect 42076 586740 42123 586744
rect 42057 586739 42123 586740
rect 40401 586530 40467 586533
rect 42517 586530 42583 586533
rect 40401 586528 42583 586530
rect 40401 586472 40406 586528
rect 40462 586472 42522 586528
rect 42578 586472 42583 586528
rect 40401 586470 42583 586472
rect 40401 586467 40467 586470
rect 42517 586467 42583 586470
rect 675569 586258 675635 586261
rect 676070 586258 676076 586260
rect 675569 586256 676076 586258
rect 675569 586200 675574 586256
rect 675630 586200 676076 586256
rect 675569 586198 676076 586200
rect 675569 586195 675635 586198
rect 676070 586196 676076 586198
rect 676140 586196 676146 586260
rect 41689 584898 41755 584901
rect 43161 584898 43227 584901
rect 41689 584896 43227 584898
rect 41689 584840 41694 584896
rect 41750 584840 43166 584896
rect 43222 584840 43227 584896
rect 41689 584838 43227 584840
rect 41689 584835 41755 584838
rect 43161 584835 43227 584838
rect 62113 584898 62179 584901
rect 62113 584896 64492 584898
rect 62113 584840 62118 584896
rect 62174 584840 64492 584896
rect 62113 584838 64492 584840
rect 62113 584835 62179 584838
rect 40677 584626 40743 584629
rect 41822 584626 41828 584628
rect 40677 584624 41828 584626
rect 40677 584568 40682 584624
rect 40738 584568 41828 584624
rect 40677 584566 41828 584568
rect 40677 584563 40743 584566
rect 41822 584564 41828 584566
rect 41892 584564 41898 584628
rect 41781 584354 41847 584357
rect 42190 584354 42196 584356
rect 41781 584352 42196 584354
rect 41781 584296 41786 584352
rect 41842 584296 42196 584352
rect 41781 584294 42196 584296
rect 41781 584291 41847 584294
rect 42190 584292 42196 584294
rect 42260 584292 42266 584356
rect 47577 582450 47643 582453
rect 42014 582448 47643 582450
rect 42014 582392 47582 582448
rect 47638 582392 47643 582448
rect 42014 582390 47643 582392
rect 42014 581770 42074 582390
rect 47577 582387 47643 582390
rect 42333 581770 42399 581773
rect 42014 581768 42399 581770
rect 42014 581712 42338 581768
rect 42394 581712 42399 581768
rect 42014 581710 42399 581712
rect 42333 581707 42399 581710
rect 41965 581500 42031 581501
rect 41965 581498 42012 581500
rect 41920 581496 42012 581498
rect 41920 581440 41970 581496
rect 41920 581438 42012 581440
rect 41965 581436 42012 581438
rect 42076 581436 42082 581500
rect 41965 581435 42031 581436
rect 44449 581090 44515 581093
rect 42198 581088 44515 581090
rect 42198 581032 44454 581088
rect 44510 581032 44515 581088
rect 42198 581030 44515 581032
rect 42198 580821 42258 581030
rect 44449 581027 44515 581030
rect 669957 581090 670023 581093
rect 669957 581088 676292 581090
rect 669957 581032 669962 581088
rect 670018 581032 676292 581088
rect 669957 581030 676292 581032
rect 669957 581027 670023 581030
rect 42198 580816 42307 580821
rect 42198 580760 42246 580816
rect 42302 580760 42307 580816
rect 42198 580758 42307 580760
rect 42241 580755 42307 580758
rect 42425 580818 42491 580821
rect 43161 580818 43227 580821
rect 42425 580816 43227 580818
rect 42425 580760 42430 580816
rect 42486 580760 43166 580816
rect 43222 580760 43227 580816
rect 42425 580758 43227 580760
rect 42425 580755 42491 580758
rect 43161 580755 43227 580758
rect 670141 580818 670207 580821
rect 673177 580818 673243 580821
rect 670141 580816 673243 580818
rect 670141 580760 670146 580816
rect 670202 580760 673182 580816
rect 673238 580760 673243 580816
rect 670141 580758 673243 580760
rect 670141 580755 670207 580758
rect 673177 580755 673243 580758
rect 676262 580546 676322 580652
rect 669270 580486 676322 580546
rect 41965 580274 42031 580277
rect 42190 580274 42196 580276
rect 41965 580272 42196 580274
rect 41965 580216 41970 580272
rect 42026 580216 42196 580272
rect 41965 580214 42196 580216
rect 41965 580211 42031 580214
rect 42190 580212 42196 580214
rect 42260 580212 42266 580276
rect 664437 580138 664503 580141
rect 669270 580138 669330 580486
rect 676262 580138 676322 580244
rect 664437 580136 669330 580138
rect 664437 580080 664442 580136
rect 664498 580080 669330 580136
rect 664437 580078 669330 580080
rect 672766 580078 676322 580138
rect 664437 580075 664503 580078
rect 658917 579730 658983 579733
rect 672766 579730 672826 580078
rect 673177 579866 673243 579869
rect 673177 579864 676292 579866
rect 673177 579808 673182 579864
rect 673238 579808 676292 579864
rect 673177 579806 676292 579808
rect 673177 579803 673243 579806
rect 658917 579728 672826 579730
rect 658917 579672 658922 579728
rect 658978 579672 672826 579728
rect 658917 579670 672826 579672
rect 658917 579667 658983 579670
rect 670233 579458 670299 579461
rect 670233 579456 676292 579458
rect 670233 579400 670238 579456
rect 670294 579400 676292 579456
rect 670233 579398 676292 579400
rect 670233 579395 670299 579398
rect 669589 579050 669655 579053
rect 669589 579048 676292 579050
rect 669589 578992 669594 579048
rect 669650 578992 676292 579048
rect 669589 578990 676292 578992
rect 669589 578987 669655 578990
rect 669957 578642 670023 578645
rect 669957 578640 676292 578642
rect 669957 578584 669962 578640
rect 670018 578584 676292 578640
rect 669957 578582 676292 578584
rect 669957 578579 670023 578582
rect 40718 578172 40724 578236
rect 40788 578234 40794 578236
rect 41781 578234 41847 578237
rect 40788 578232 41847 578234
rect 40788 578176 41786 578232
rect 41842 578176 41847 578232
rect 40788 578174 41847 578176
rect 40788 578172 40794 578174
rect 41781 578171 41847 578174
rect 671153 578234 671219 578237
rect 671153 578232 676292 578234
rect 671153 578176 671158 578232
rect 671214 578176 676292 578232
rect 671153 578174 676292 578176
rect 671153 578171 671219 578174
rect 42558 577900 42564 577964
rect 42628 577962 42634 577964
rect 42885 577962 42951 577965
rect 42628 577960 42951 577962
rect 42628 577904 42890 577960
rect 42946 577904 42951 577960
rect 42628 577902 42951 577904
rect 42628 577900 42634 577902
rect 42885 577899 42951 577902
rect 669589 577826 669655 577829
rect 669589 577824 676292 577826
rect 669589 577768 669594 577824
rect 669650 577768 676292 577824
rect 669589 577766 676292 577768
rect 669589 577763 669655 577766
rect 40902 577492 40908 577556
rect 40972 577554 40978 577556
rect 41781 577554 41847 577557
rect 42701 577554 42767 577557
rect 40972 577552 41847 577554
rect 40972 577496 41786 577552
rect 41842 577496 41847 577552
rect 40972 577494 41847 577496
rect 40972 577492 40978 577494
rect 41781 577491 41847 577494
rect 42152 577552 42767 577554
rect 42152 577496 42706 577552
rect 42762 577496 42767 577552
rect 42152 577494 42767 577496
rect 42152 577149 42212 577494
rect 42701 577491 42767 577494
rect 651465 577418 651531 577421
rect 650164 577416 651531 577418
rect 650164 577360 651470 577416
rect 651526 577360 651531 577416
rect 650164 577358 651531 577360
rect 651465 577355 651531 577358
rect 671613 577418 671679 577421
rect 671613 577416 676292 577418
rect 671613 577360 671618 577416
rect 671674 577360 676292 577416
rect 671613 577358 676292 577360
rect 671613 577355 671679 577358
rect 42149 577144 42215 577149
rect 42149 577088 42154 577144
rect 42210 577088 42215 577144
rect 42149 577083 42215 577088
rect 671797 577010 671863 577013
rect 671797 577008 676292 577010
rect 671797 576952 671802 577008
rect 671858 576952 676292 577008
rect 671797 576950 676292 576952
rect 671797 576947 671863 576950
rect 40534 576812 40540 576876
rect 40604 576874 40610 576876
rect 40604 576814 42074 576874
rect 40604 576812 40610 576814
rect 42014 576605 42074 576814
rect 41965 576600 42074 576605
rect 41965 576544 41970 576600
rect 42026 576544 42074 576600
rect 41965 576542 42074 576544
rect 676029 576602 676095 576605
rect 676029 576600 676292 576602
rect 676029 576544 676034 576600
rect 676090 576544 676292 576600
rect 676029 576542 676292 576544
rect 41965 576539 42031 576542
rect 676029 576539 676095 576542
rect 683849 576466 683915 576469
rect 683806 576464 683915 576466
rect 683806 576408 683854 576464
rect 683910 576408 683915 576464
rect 683806 576403 683915 576408
rect 683806 576164 683866 576403
rect 680997 576058 681063 576061
rect 680997 576056 681106 576058
rect 680997 576000 681002 576056
rect 681058 576000 681106 576056
rect 680997 575995 681106 576000
rect 681046 575756 681106 575995
rect 675109 575514 675175 575517
rect 675109 575512 676322 575514
rect 675109 575456 675114 575512
rect 675170 575456 676322 575512
rect 675109 575454 676322 575456
rect 675109 575451 675175 575454
rect 676262 575348 676322 575454
rect 672625 575106 672691 575109
rect 676029 575106 676095 575109
rect 672625 575104 676095 575106
rect 672625 575048 672630 575104
rect 672686 575048 676034 575104
rect 676090 575048 676095 575104
rect 672625 575046 676095 575048
rect 672625 575043 672691 575046
rect 676029 575043 676095 575046
rect 669037 574834 669103 574837
rect 676262 574834 676322 574940
rect 669037 574832 676322 574834
rect 669037 574776 669042 574832
rect 669098 574776 676322 574832
rect 669037 574774 676322 574776
rect 669037 574771 669103 574774
rect 668853 574426 668919 574429
rect 676262 574426 676322 574532
rect 668853 574424 676322 574426
rect 668853 574368 668858 574424
rect 668914 574368 676322 574424
rect 668853 574366 676322 574368
rect 668853 574363 668919 574366
rect 42149 574154 42215 574157
rect 42558 574154 42564 574156
rect 42149 574152 42564 574154
rect 42149 574096 42154 574152
rect 42210 574096 42564 574152
rect 42149 574094 42564 574096
rect 42149 574091 42215 574094
rect 42558 574092 42564 574094
rect 42628 574092 42634 574156
rect 669221 574154 669287 574157
rect 669221 574152 676292 574154
rect 669221 574096 669226 574152
rect 669282 574096 676292 574152
rect 669221 574094 676292 574096
rect 669221 574091 669287 574094
rect 676029 573746 676095 573749
rect 676029 573744 676292 573746
rect 676029 573688 676034 573744
rect 676090 573688 676292 573744
rect 676029 573686 676292 573688
rect 676029 573683 676095 573686
rect 41454 573276 41460 573340
rect 41524 573338 41530 573340
rect 42609 573338 42675 573341
rect 41524 573336 42675 573338
rect 41524 573280 42614 573336
rect 42670 573280 42675 573336
rect 41524 573278 42675 573280
rect 41524 573276 41530 573278
rect 42609 573275 42675 573278
rect 673177 573338 673243 573341
rect 673177 573336 676292 573338
rect 673177 573280 673182 573336
rect 673238 573280 676292 573336
rect 673177 573278 676292 573280
rect 673177 573275 673243 573278
rect 683665 573202 683731 573205
rect 683622 573200 683731 573202
rect 683622 573144 683670 573200
rect 683726 573144 683731 573200
rect 683622 573139 683731 573144
rect 683622 572900 683682 573139
rect 676990 572732 676996 572796
rect 677060 572732 677066 572796
rect 676998 572492 677058 572732
rect 41638 572052 41644 572116
rect 41708 572114 41714 572116
rect 42517 572114 42583 572117
rect 41708 572112 42583 572114
rect 41708 572056 42522 572112
rect 42578 572056 42583 572112
rect 41708 572054 42583 572056
rect 41708 572052 41714 572054
rect 42517 572051 42583 572054
rect 670785 571978 670851 571981
rect 676262 571978 676322 572084
rect 670785 571976 676322 571978
rect 670785 571920 670790 571976
rect 670846 571920 676322 571976
rect 670785 571918 676322 571920
rect 683389 571978 683455 571981
rect 683389 571976 683498 571978
rect 683389 571920 683394 571976
rect 683450 571920 683498 571976
rect 670785 571915 670851 571918
rect 683389 571915 683498 571920
rect 62113 571842 62179 571845
rect 62113 571840 64492 571842
rect 62113 571784 62118 571840
rect 62174 571784 64492 571840
rect 62113 571782 64492 571784
rect 62113 571779 62179 571782
rect 683438 571676 683498 571915
rect 674833 571162 674899 571165
rect 676262 571162 676322 571268
rect 674833 571160 676322 571162
rect 674833 571104 674838 571160
rect 674894 571104 676322 571160
rect 674833 571102 676322 571104
rect 674833 571099 674899 571102
rect 670785 570754 670851 570757
rect 676262 570754 676322 570860
rect 682377 570754 682443 570757
rect 670785 570752 676322 570754
rect 670785 570696 670790 570752
rect 670846 570696 676322 570752
rect 670785 570694 676322 570696
rect 682334 570752 682443 570754
rect 682334 570696 682382 570752
rect 682438 570696 682443 570752
rect 670785 570691 670851 570694
rect 682334 570691 682443 570696
rect 669773 570346 669839 570349
rect 674833 570346 674899 570349
rect 669773 570344 674899 570346
rect 669773 570288 669778 570344
rect 669834 570288 674838 570344
rect 674894 570288 674899 570344
rect 669773 570286 674899 570288
rect 669773 570283 669839 570286
rect 674833 570283 674899 570286
rect 41781 570212 41847 570213
rect 41781 570208 41828 570212
rect 41892 570210 41898 570212
rect 41781 570152 41786 570208
rect 41781 570148 41828 570152
rect 41892 570150 41938 570210
rect 41892 570148 41898 570150
rect 41781 570147 41847 570148
rect 682334 570044 682394 570691
rect 669773 569530 669839 569533
rect 676262 569530 676322 569636
rect 669773 569528 676322 569530
rect 669773 569472 669778 569528
rect 669834 569472 676322 569528
rect 669773 569470 676322 569472
rect 669773 569467 669839 569470
rect 42333 569258 42399 569261
rect 62113 569258 62179 569261
rect 42333 569256 62179 569258
rect 42333 569200 42338 569256
rect 42394 569200 62118 569256
rect 62174 569200 62179 569256
rect 42333 569198 62179 569200
rect 42333 569195 42399 569198
rect 62113 569195 62179 569198
rect 667381 564498 667447 564501
rect 675385 564498 675451 564501
rect 667381 564496 675451 564498
rect 667381 564440 667386 564496
rect 667442 564440 675390 564496
rect 675446 564440 675451 564496
rect 667381 564438 675451 564440
rect 667381 564435 667447 564438
rect 675385 564435 675451 564438
rect 651649 564090 651715 564093
rect 650164 564088 651715 564090
rect 650164 564032 651654 564088
rect 651710 564032 651715 564088
rect 650164 564030 651715 564032
rect 651649 564027 651715 564030
rect 675477 562732 675543 562733
rect 675477 562728 675524 562732
rect 675588 562730 675594 562732
rect 675477 562672 675482 562728
rect 675477 562668 675524 562672
rect 675588 562670 675634 562730
rect 675588 562668 675594 562670
rect 675477 562667 675543 562668
rect 675477 561236 675543 561237
rect 675477 561232 675524 561236
rect 675588 561234 675594 561236
rect 675477 561176 675482 561232
rect 675477 561172 675524 561176
rect 675588 561174 675634 561234
rect 675588 561172 675594 561174
rect 675477 561171 675543 561172
rect 673177 560146 673243 560149
rect 675385 560146 675451 560149
rect 673177 560144 675451 560146
rect 673177 560088 673182 560144
rect 673238 560088 675390 560144
rect 675446 560088 675451 560144
rect 673177 560086 675451 560088
rect 673177 560083 673243 560086
rect 675385 560083 675451 560086
rect 674833 559602 674899 559605
rect 675477 559602 675543 559605
rect 674833 559600 675543 559602
rect 674833 559544 674838 559600
rect 674894 559544 675482 559600
rect 675538 559544 675543 559600
rect 674833 559542 675543 559544
rect 674833 559539 674899 559542
rect 675477 559539 675543 559542
rect 62113 558786 62179 558789
rect 62113 558784 64492 558786
rect 62113 558728 62118 558784
rect 62174 558728 64492 558784
rect 62113 558726 64492 558728
rect 62113 558723 62179 558726
rect 42057 558514 42123 558517
rect 41492 558512 42123 558514
rect 41492 558456 42062 558512
rect 42118 558456 42123 558512
rect 41492 558454 42123 558456
rect 42057 558451 42123 558454
rect 35801 558106 35867 558109
rect 35788 558104 35867 558106
rect 35788 558048 35806 558104
rect 35862 558048 35867 558104
rect 35788 558046 35867 558048
rect 35801 558043 35867 558046
rect 674005 558106 674071 558109
rect 675385 558106 675451 558109
rect 674005 558104 675451 558106
rect 674005 558048 674010 558104
rect 674066 558048 675390 558104
rect 675446 558048 675451 558104
rect 674005 558046 675451 558048
rect 674005 558043 674071 558046
rect 675385 558043 675451 558046
rect 673821 557970 673887 557973
rect 673821 557968 673930 557970
rect 673821 557912 673826 557968
rect 673882 557912 673930 557968
rect 673821 557907 673930 557912
rect 48957 557834 49023 557837
rect 41830 557832 49023 557834
rect 41830 557776 48962 557832
rect 49018 557776 49023 557832
rect 41830 557774 49023 557776
rect 673870 557834 673930 557907
rect 675385 557834 675451 557837
rect 673870 557832 675451 557834
rect 673870 557776 675390 557832
rect 675446 557776 675451 557832
rect 673870 557774 675451 557776
rect 41830 557698 41890 557774
rect 48957 557771 49023 557774
rect 675385 557771 675451 557774
rect 41492 557638 41890 557698
rect 42057 557562 42123 557565
rect 50337 557562 50403 557565
rect 42057 557560 50403 557562
rect 42057 557504 42062 557560
rect 42118 557504 50342 557560
rect 50398 557504 50403 557560
rect 42057 557502 50403 557504
rect 42057 557499 42123 557502
rect 50337 557499 50403 557502
rect 669037 557562 669103 557565
rect 675017 557562 675083 557565
rect 669037 557560 675083 557562
rect 669037 557504 669042 557560
rect 669098 557504 675022 557560
rect 675078 557504 675083 557560
rect 669037 557502 675083 557504
rect 669037 557499 669103 557502
rect 675017 557499 675083 557502
rect 675477 557562 675543 557565
rect 676806 557562 676812 557564
rect 675477 557560 676812 557562
rect 675477 557504 675482 557560
rect 675538 557504 676812 557560
rect 675477 557502 676812 557504
rect 675477 557499 675543 557502
rect 676806 557500 676812 557502
rect 676876 557500 676882 557564
rect 44633 557290 44699 557293
rect 41492 557288 44699 557290
rect 41492 557232 44638 557288
rect 44694 557232 44699 557288
rect 41492 557230 44699 557232
rect 44633 557227 44699 557230
rect 45645 556882 45711 556885
rect 41492 556880 45711 556882
rect 41492 556824 45650 556880
rect 45706 556824 45711 556880
rect 41492 556822 45711 556824
rect 45645 556819 45711 556822
rect 44817 556474 44883 556477
rect 41492 556472 44883 556474
rect 41492 556416 44822 556472
rect 44878 556416 44883 556472
rect 41492 556414 44883 556416
rect 44817 556411 44883 556414
rect 46013 556066 46079 556069
rect 41492 556064 46079 556066
rect 41492 556008 46018 556064
rect 46074 556008 46079 556064
rect 41492 556006 46079 556008
rect 46013 556003 46079 556006
rect 675017 555794 675083 555797
rect 675477 555794 675543 555797
rect 675017 555792 675543 555794
rect 675017 555736 675022 555792
rect 675078 555736 675482 555792
rect 675538 555736 675543 555792
rect 675017 555734 675543 555736
rect 675017 555731 675083 555734
rect 675477 555731 675543 555734
rect 45001 555658 45067 555661
rect 41492 555656 45067 555658
rect 41492 555600 45006 555656
rect 45062 555600 45067 555656
rect 41492 555598 45067 555600
rect 45001 555595 45067 555598
rect 44633 555250 44699 555253
rect 41492 555248 44699 555250
rect 41492 555192 44638 555248
rect 44694 555192 44699 555248
rect 41492 555190 44699 555192
rect 44633 555187 44699 555190
rect 35801 554842 35867 554845
rect 35788 554840 35867 554842
rect 35788 554784 35806 554840
rect 35862 554784 35867 554840
rect 35788 554782 35867 554784
rect 35801 554779 35867 554782
rect 44265 554434 44331 554437
rect 41492 554432 44331 554434
rect 41492 554376 44270 554432
rect 44326 554376 44331 554432
rect 41492 554374 44331 554376
rect 44265 554371 44331 554374
rect 674373 554434 674439 554437
rect 675385 554434 675451 554437
rect 674373 554432 675451 554434
rect 674373 554376 674378 554432
rect 674434 554376 675390 554432
rect 675446 554376 675451 554432
rect 674373 554374 675451 554376
rect 674373 554371 674439 554374
rect 675385 554371 675451 554374
rect 42190 554026 42196 554028
rect 41492 553966 42196 554026
rect 42190 553964 42196 553966
rect 42260 553964 42266 554028
rect 658917 554026 658983 554029
rect 675201 554026 675267 554029
rect 658917 554024 675267 554026
rect 658917 553968 658922 554024
rect 658978 553968 675206 554024
rect 675262 553968 675267 554024
rect 658917 553966 675267 553968
rect 658917 553963 658983 553966
rect 675201 553963 675267 553966
rect 35801 553618 35867 553621
rect 35788 553616 35867 553618
rect 35788 553560 35806 553616
rect 35862 553560 35867 553616
rect 35788 553558 35867 553560
rect 35801 553555 35867 553558
rect 670417 553482 670483 553485
rect 675385 553482 675451 553485
rect 670417 553480 675451 553482
rect 670417 553424 670422 553480
rect 670478 553424 675390 553480
rect 675446 553424 675451 553480
rect 670417 553422 675451 553424
rect 670417 553419 670483 553422
rect 675385 553419 675451 553422
rect 42006 553210 42012 553212
rect 41492 553150 42012 553210
rect 42006 553148 42012 553150
rect 42076 553148 42082 553212
rect 41321 552802 41387 552805
rect 41308 552800 41387 552802
rect 41308 552744 41326 552800
rect 41382 552744 41387 552800
rect 41308 552742 41387 552744
rect 41321 552739 41387 552742
rect 669221 552666 669287 552669
rect 675477 552666 675543 552669
rect 669221 552664 675543 552666
rect 669221 552608 669226 552664
rect 669282 552608 675482 552664
rect 675538 552608 675543 552664
rect 669221 552606 675543 552608
rect 669221 552603 669287 552606
rect 675477 552603 675543 552606
rect 44449 552394 44515 552397
rect 41492 552392 44515 552394
rect 41492 552336 44454 552392
rect 44510 552336 44515 552392
rect 41492 552334 44515 552336
rect 44449 552331 44515 552334
rect 33777 551986 33843 551989
rect 33764 551984 33843 551986
rect 33764 551928 33782 551984
rect 33838 551928 33843 551984
rect 33764 551926 33843 551928
rect 33777 551923 33843 551926
rect 41689 551850 41755 551853
rect 42374 551850 42380 551852
rect 41689 551848 42380 551850
rect 41689 551792 41694 551848
rect 41750 551792 42380 551848
rect 41689 551790 42380 551792
rect 41689 551787 41755 551790
rect 42374 551788 42380 551790
rect 42444 551788 42450 551852
rect 43069 551578 43135 551581
rect 41492 551576 43135 551578
rect 41492 551520 43074 551576
rect 43130 551520 43135 551576
rect 41492 551518 43135 551520
rect 43069 551515 43135 551518
rect 44909 551170 44975 551173
rect 41492 551168 44975 551170
rect 41492 551112 44914 551168
rect 44970 551112 44975 551168
rect 41492 551110 44975 551112
rect 44909 551107 44975 551110
rect 651465 550898 651531 550901
rect 650164 550896 651531 550898
rect 650164 550840 651470 550896
rect 651526 550840 651531 550896
rect 650164 550838 651531 550840
rect 651465 550835 651531 550838
rect 41781 550762 41847 550765
rect 41492 550760 41847 550762
rect 41492 550704 41786 550760
rect 41842 550704 41847 550760
rect 41492 550702 41847 550704
rect 41781 550699 41847 550702
rect 41965 550354 42031 550357
rect 41492 550352 42031 550354
rect 41492 550296 41970 550352
rect 42026 550296 42031 550352
rect 41492 550294 42031 550296
rect 41965 550291 42031 550294
rect 675753 550354 675819 550357
rect 676990 550354 676996 550356
rect 675753 550352 676996 550354
rect 675753 550296 675758 550352
rect 675814 550296 676996 550352
rect 675753 550294 676996 550296
rect 675753 550291 675819 550294
rect 676990 550292 676996 550294
rect 677060 550292 677066 550356
rect 675109 550220 675175 550221
rect 675109 550218 675156 550220
rect 675064 550216 675156 550218
rect 675064 550160 675114 550216
rect 675064 550158 675156 550160
rect 675109 550156 675156 550158
rect 675220 550156 675226 550220
rect 675109 550155 675175 550156
rect 40493 549946 40559 549949
rect 40493 549944 40572 549946
rect 40493 549888 40498 549944
rect 40554 549888 40572 549944
rect 40493 549886 40572 549888
rect 40493 549883 40559 549886
rect 45093 549538 45159 549541
rect 41492 549536 45159 549538
rect 41492 549480 45098 549536
rect 45154 549480 45159 549536
rect 41492 549478 45159 549480
rect 45093 549475 45159 549478
rect 45277 549130 45343 549133
rect 41492 549128 45343 549130
rect 41492 549072 45282 549128
rect 45338 549072 45343 549128
rect 41492 549070 45343 549072
rect 45277 549067 45343 549070
rect 44817 548722 44883 548725
rect 41492 548720 44883 548722
rect 41492 548664 44822 548720
rect 44878 548664 44883 548720
rect 41492 548662 44883 548664
rect 44817 548659 44883 548662
rect 41781 548450 41847 548453
rect 42885 548450 42951 548453
rect 41781 548448 42951 548450
rect 41781 548392 41786 548448
rect 41842 548392 42890 548448
rect 42946 548392 42951 548448
rect 41781 548390 42951 548392
rect 41781 548387 41847 548390
rect 42885 548387 42951 548390
rect 671153 548450 671219 548453
rect 675477 548450 675543 548453
rect 671153 548448 675543 548450
rect 671153 548392 671158 548448
rect 671214 548392 675482 548448
rect 675538 548392 675543 548448
rect 671153 548390 675543 548392
rect 671153 548387 671219 548390
rect 675477 548387 675543 548390
rect 41278 548147 41338 548284
rect 31753 548144 31819 548147
rect 31710 548142 31819 548144
rect 31710 548086 31758 548142
rect 31814 548086 31819 548142
rect 31710 548081 31819 548086
rect 41229 548142 41338 548147
rect 41229 548086 41234 548142
rect 41290 548086 41338 548142
rect 41689 548178 41755 548181
rect 43805 548178 43871 548181
rect 41689 548176 43871 548178
rect 41689 548120 41694 548176
rect 41750 548120 43810 548176
rect 43866 548120 43871 548176
rect 41689 548118 43871 548120
rect 41689 548115 41755 548118
rect 43805 548115 43871 548118
rect 41229 548084 41338 548086
rect 41229 548081 41295 548084
rect 28766 547498 28826 547890
rect 31710 547498 31770 548081
rect 675150 547572 675156 547636
rect 675220 547634 675226 547636
rect 675845 547634 675911 547637
rect 675220 547632 675911 547634
rect 675220 547576 675850 547632
rect 675906 547576 675911 547632
rect 675220 547574 675911 547576
rect 675220 547572 675226 547574
rect 675845 547571 675911 547574
rect 676070 547572 676076 547636
rect 676140 547634 676146 547636
rect 678237 547634 678303 547637
rect 676140 547632 678303 547634
rect 676140 547576 678242 547632
rect 678298 547576 678303 547632
rect 676140 547574 678303 547576
rect 676140 547572 676146 547574
rect 678237 547571 678303 547574
rect 28766 547468 31770 547498
rect 28796 547438 31770 547468
rect 674230 547300 674236 547364
rect 674300 547362 674306 547364
rect 683573 547362 683639 547365
rect 674300 547360 683639 547362
rect 674300 547304 683578 547360
rect 683634 547304 683639 547360
rect 674300 547302 683639 547304
rect 674300 547300 674306 547302
rect 683573 547299 683639 547302
rect 43989 547090 44055 547093
rect 41492 547088 44055 547090
rect 41492 547032 43994 547088
rect 44050 547032 44055 547088
rect 41492 547030 44055 547032
rect 43989 547027 44055 547030
rect 674189 547090 674255 547093
rect 683849 547090 683915 547093
rect 674189 547088 683915 547090
rect 674189 547032 674194 547088
rect 674250 547032 683854 547088
rect 683910 547032 683915 547088
rect 674189 547030 683915 547032
rect 674189 547027 674255 547030
rect 683849 547027 683915 547030
rect 674833 546410 674899 546413
rect 675661 546410 675727 546413
rect 674833 546408 675727 546410
rect 674833 546352 674838 546408
rect 674894 546352 675666 546408
rect 675722 546352 675727 546408
rect 674833 546350 675727 546352
rect 674833 546347 674899 546350
rect 675661 546347 675727 546350
rect 675293 546138 675359 546141
rect 675518 546138 675524 546140
rect 675293 546136 675524 546138
rect 675293 546080 675298 546136
rect 675354 546080 675524 546136
rect 675293 546078 675524 546080
rect 675293 546075 675359 546078
rect 675518 546076 675524 546078
rect 675588 546076 675594 546140
rect 62113 545866 62179 545869
rect 673637 545866 673703 545869
rect 62113 545864 64492 545866
rect 62113 545808 62118 545864
rect 62174 545808 64492 545864
rect 62113 545806 64492 545808
rect 673637 545864 676230 545866
rect 673637 545808 673642 545864
rect 673698 545808 676230 545864
rect 673637 545806 676230 545808
rect 62113 545803 62179 545806
rect 673637 545803 673703 545806
rect 40718 545668 40724 545732
rect 40788 545730 40794 545732
rect 41965 545730 42031 545733
rect 40788 545728 42031 545730
rect 40788 545672 41970 545728
rect 42026 545672 42031 545728
rect 40788 545670 42031 545672
rect 676170 545730 676230 545806
rect 683297 545730 683363 545733
rect 676170 545728 683363 545730
rect 676170 545672 683302 545728
rect 683358 545672 683363 545728
rect 676170 545670 683363 545672
rect 40788 545668 40794 545670
rect 41965 545667 42031 545670
rect 683297 545667 683363 545670
rect 674833 545594 674899 545597
rect 675334 545594 675340 545596
rect 674833 545592 675340 545594
rect 674833 545536 674838 545592
rect 674894 545536 675340 545592
rect 674833 545534 675340 545536
rect 674833 545531 674899 545534
rect 675334 545532 675340 545534
rect 675404 545532 675410 545596
rect 40493 545460 40559 545461
rect 40493 545456 40540 545460
rect 40604 545458 40610 545460
rect 40493 545400 40498 545456
rect 40493 545396 40540 545400
rect 40604 545398 40650 545458
rect 40604 545396 40610 545398
rect 40493 545395 40559 545396
rect 41781 541106 41847 541109
rect 41781 541104 41890 541106
rect 41781 541048 41786 541104
rect 41842 541048 41890 541104
rect 41781 541043 41890 541048
rect 41830 540701 41890 541043
rect 41781 540696 41890 540701
rect 41781 540640 41786 540696
rect 41842 540640 41890 540696
rect 41781 540638 41890 540640
rect 41781 540635 41847 540638
rect 42609 540290 42675 540293
rect 56041 540290 56107 540293
rect 42609 540288 56107 540290
rect 42609 540232 42614 540288
rect 42670 540232 56046 540288
rect 56102 540232 56107 540288
rect 42609 540230 56107 540232
rect 42609 540227 42675 540230
rect 56041 540227 56107 540230
rect 40718 538188 40724 538252
rect 40788 538250 40794 538252
rect 42241 538250 42307 538253
rect 40788 538248 42307 538250
rect 40788 538192 42246 538248
rect 42302 538192 42307 538248
rect 40788 538190 42307 538192
rect 40788 538188 40794 538190
rect 42241 538187 42307 538190
rect 42057 537978 42123 537981
rect 42609 537978 42675 537981
rect 42057 537976 42675 537978
rect 42057 537920 42062 537976
rect 42118 537920 42614 537976
rect 42670 537920 42675 537976
rect 42057 537918 42675 537920
rect 42057 537915 42123 537918
rect 42609 537915 42675 537918
rect 651465 537570 651531 537573
rect 650164 537568 651531 537570
rect 650164 537512 651470 537568
rect 651526 537512 651531 537568
rect 650164 537510 651531 537512
rect 651465 537507 651531 537510
rect 42609 537434 42675 537437
rect 45369 537434 45435 537437
rect 42609 537432 45435 537434
rect 42609 537376 42614 537432
rect 42670 537376 45374 537432
rect 45430 537376 45435 537432
rect 42609 537374 45435 537376
rect 42609 537371 42675 537374
rect 45369 537371 45435 537374
rect 44817 536890 44883 536893
rect 42198 536888 44883 536890
rect 42198 536832 44822 536888
rect 44878 536832 44883 536888
rect 42198 536830 44883 536832
rect 42198 536349 42258 536830
rect 44817 536827 44883 536830
rect 42198 536344 42307 536349
rect 42198 536288 42246 536344
rect 42302 536288 42307 536344
rect 42198 536286 42307 536288
rect 42241 536283 42307 536286
rect 668577 535938 668643 535941
rect 676262 535938 676322 536112
rect 668577 535936 676322 535938
rect 668577 535880 668582 535936
rect 668638 535880 676322 535936
rect 668577 535878 676322 535880
rect 668577 535875 668643 535878
rect 663057 535530 663123 535533
rect 676262 535530 676322 535704
rect 663057 535528 676322 535530
rect 663057 535472 663062 535528
rect 663118 535472 676322 535528
rect 663057 535470 676322 535472
rect 663057 535467 663123 535470
rect 40534 535196 40540 535260
rect 40604 535258 40610 535260
rect 41781 535258 41847 535261
rect 40604 535256 41847 535258
rect 40604 535200 41786 535256
rect 41842 535200 41847 535256
rect 40604 535198 41847 535200
rect 40604 535196 40610 535198
rect 41781 535195 41847 535198
rect 667197 535258 667263 535261
rect 676262 535258 676322 535296
rect 667197 535256 676322 535258
rect 667197 535200 667202 535256
rect 667258 535200 676322 535256
rect 667197 535198 676322 535200
rect 667197 535195 667263 535198
rect 670233 534986 670299 534989
rect 670233 534984 676322 534986
rect 670233 534928 670238 534984
rect 670294 534928 676322 534984
rect 670233 534926 676322 534928
rect 670233 534923 670299 534926
rect 676262 534888 676322 534926
rect 669957 534714 670023 534717
rect 675753 534714 675819 534717
rect 669957 534712 675819 534714
rect 669957 534656 669962 534712
rect 670018 534656 675758 534712
rect 675814 534656 675819 534712
rect 669957 534654 675819 534656
rect 669957 534651 670023 534654
rect 675753 534651 675819 534654
rect 42517 534306 42583 534309
rect 44449 534306 44515 534309
rect 42517 534304 44515 534306
rect 42517 534248 42522 534304
rect 42578 534248 44454 534304
rect 44510 534248 44515 534304
rect 42517 534246 44515 534248
rect 42517 534243 42583 534246
rect 44449 534243 44515 534246
rect 671797 534306 671863 534309
rect 676262 534306 676322 534480
rect 671797 534304 676322 534306
rect 671797 534248 671802 534304
rect 671858 534248 676322 534304
rect 671797 534246 676322 534248
rect 671797 534243 671863 534246
rect 675753 534102 675819 534105
rect 675753 534100 676292 534102
rect 675753 534044 675758 534100
rect 675814 534044 676292 534100
rect 675753 534042 676292 534044
rect 675753 534039 675819 534042
rect 672625 533490 672691 533493
rect 676262 533490 676322 533664
rect 672625 533488 676322 533490
rect 672625 533432 672630 533488
rect 672686 533432 676322 533488
rect 672625 533430 676322 533432
rect 672625 533427 672691 533430
rect 42425 533354 42491 533357
rect 45277 533354 45343 533357
rect 42425 533352 45343 533354
rect 42425 533296 42430 533352
rect 42486 533296 45282 533352
rect 45338 533296 45343 533352
rect 42425 533294 45343 533296
rect 42425 533291 42491 533294
rect 45277 533291 45343 533294
rect 669589 533082 669655 533085
rect 676262 533082 676322 533256
rect 669589 533080 676322 533082
rect 669589 533024 669594 533080
rect 669650 533024 676322 533080
rect 669589 533022 676322 533024
rect 669589 533019 669655 533022
rect 62113 532810 62179 532813
rect 670969 532810 671035 532813
rect 676262 532810 676322 532848
rect 62113 532808 64492 532810
rect 62113 532752 62118 532808
rect 62174 532752 64492 532808
rect 62113 532750 64492 532752
rect 670969 532808 676322 532810
rect 670969 532752 670974 532808
rect 671030 532752 676322 532808
rect 670969 532750 676322 532752
rect 62113 532747 62179 532750
rect 670969 532747 671035 532750
rect 42701 532674 42767 532677
rect 45001 532674 45067 532677
rect 42701 532672 45067 532674
rect 42701 532616 42706 532672
rect 42762 532616 45006 532672
rect 45062 532616 45067 532672
rect 42701 532614 45067 532616
rect 42701 532611 42767 532614
rect 45001 532611 45067 532614
rect 672257 532538 672323 532541
rect 675753 532538 675819 532541
rect 672257 532536 675819 532538
rect 672257 532480 672262 532536
rect 672318 532480 675758 532536
rect 675814 532480 675819 532536
rect 672257 532478 675819 532480
rect 672257 532475 672323 532478
rect 675753 532475 675819 532478
rect 676262 532266 676322 532440
rect 674606 532206 676322 532266
rect 671613 531858 671679 531861
rect 674606 531858 674666 532206
rect 676262 531858 676322 532032
rect 671613 531856 674666 531858
rect 671613 531800 671618 531856
rect 671674 531800 674666 531856
rect 671613 531798 674666 531800
rect 674790 531798 676322 531858
rect 671613 531795 671679 531798
rect 671613 531450 671679 531453
rect 674790 531450 674850 531798
rect 675753 531654 675819 531657
rect 675753 531652 676292 531654
rect 675753 531596 675758 531652
rect 675814 531596 676292 531652
rect 675753 531594 676292 531596
rect 675753 531591 675819 531594
rect 671613 531448 674850 531450
rect 671613 531392 671618 531448
rect 671674 531392 674850 531448
rect 671613 531390 674850 531392
rect 680997 531450 681063 531453
rect 680997 531448 681106 531450
rect 680997 531392 681002 531448
rect 681058 531392 681106 531448
rect 671613 531387 671679 531390
rect 680997 531387 681106 531392
rect 681046 531216 681106 531387
rect 678237 531042 678303 531045
rect 678237 531040 678346 531042
rect 678237 530984 678242 531040
rect 678298 530984 678346 531040
rect 678237 530979 678346 530984
rect 678286 530808 678346 530979
rect 672993 530634 673059 530637
rect 676029 530634 676095 530637
rect 672993 530632 676095 530634
rect 672993 530576 672998 530632
rect 673054 530576 676034 530632
rect 676090 530576 676095 530632
rect 672993 530574 676095 530576
rect 672993 530571 673059 530574
rect 676029 530571 676095 530574
rect 41638 530164 41644 530228
rect 41708 530226 41714 530228
rect 42425 530226 42491 530229
rect 41708 530224 42491 530226
rect 41708 530168 42430 530224
rect 42486 530168 42491 530224
rect 41708 530166 42491 530168
rect 41708 530164 41714 530166
rect 42425 530163 42491 530166
rect 672809 530226 672875 530229
rect 676262 530226 676322 530400
rect 672809 530224 676322 530226
rect 672809 530168 672814 530224
rect 672870 530168 676322 530224
rect 672809 530166 676322 530168
rect 672809 530163 672875 530166
rect 42057 529954 42123 529957
rect 42701 529954 42767 529957
rect 42057 529952 42767 529954
rect 42057 529896 42062 529952
rect 42118 529896 42706 529952
rect 42762 529896 42767 529952
rect 42057 529894 42767 529896
rect 42057 529891 42123 529894
rect 42701 529891 42767 529894
rect 667657 529954 667723 529957
rect 676262 529954 676322 529992
rect 667657 529952 676322 529954
rect 667657 529896 667662 529952
rect 667718 529896 676322 529952
rect 667657 529894 676322 529896
rect 667657 529891 667723 529894
rect 41454 529620 41460 529684
rect 41524 529682 41530 529684
rect 42701 529682 42767 529685
rect 41524 529680 42767 529682
rect 41524 529624 42706 529680
rect 42762 529624 42767 529680
rect 41524 529622 42767 529624
rect 41524 529620 41530 529622
rect 42701 529619 42767 529622
rect 41873 529412 41939 529413
rect 41822 529410 41828 529412
rect 41782 529350 41828 529410
rect 41892 529408 41939 529412
rect 41934 529352 41939 529408
rect 41822 529348 41828 529350
rect 41892 529348 41939 529352
rect 41873 529347 41939 529348
rect 674189 529410 674255 529413
rect 676262 529410 676322 529584
rect 674189 529408 676322 529410
rect 674189 529352 674194 529408
rect 674250 529352 676322 529408
rect 674189 529350 676322 529352
rect 674189 529347 674255 529350
rect 672441 529002 672507 529005
rect 676262 529002 676322 529176
rect 672441 529000 676322 529002
rect 672441 528944 672446 529000
rect 672502 528944 676322 529000
rect 672441 528942 676322 528944
rect 672441 528939 672507 528942
rect 676029 528798 676095 528801
rect 676029 528796 676292 528798
rect 676029 528740 676034 528796
rect 676090 528740 676292 528796
rect 676029 528738 676292 528740
rect 676029 528735 676095 528738
rect 667013 528594 667079 528597
rect 674189 528594 674255 528597
rect 667013 528592 674255 528594
rect 667013 528536 667018 528592
rect 667074 528536 674194 528592
rect 674250 528536 674255 528592
rect 667013 528534 674255 528536
rect 667013 528531 667079 528534
rect 674189 528531 674255 528534
rect 673637 528322 673703 528325
rect 676262 528322 676322 528360
rect 673637 528320 676322 528322
rect 673637 528264 673642 528320
rect 673698 528264 676322 528320
rect 673637 528262 676322 528264
rect 673637 528259 673703 528262
rect 683849 528186 683915 528189
rect 683806 528184 683915 528186
rect 683806 528128 683854 528184
rect 683910 528128 683915 528184
rect 683806 528123 683915 528128
rect 683806 527952 683866 528123
rect 668393 527370 668459 527373
rect 676262 527370 676322 527544
rect 668393 527368 676322 527370
rect 668393 527312 668398 527368
rect 668454 527312 676322 527368
rect 668393 527310 676322 527312
rect 683573 527370 683639 527373
rect 683573 527368 683682 527370
rect 683573 527312 683578 527368
rect 683634 527312 683682 527368
rect 668393 527307 668459 527310
rect 683573 527307 683682 527312
rect 683622 527136 683682 527307
rect 674649 526962 674715 526965
rect 674649 526960 676322 526962
rect 674649 526904 674654 526960
rect 674710 526904 676322 526960
rect 674649 526902 676322 526904
rect 674649 526899 674715 526902
rect 676262 526728 676322 526902
rect 683297 526554 683363 526557
rect 683254 526552 683363 526554
rect 683254 526496 683302 526552
rect 683358 526496 683363 526552
rect 683254 526491 683363 526496
rect 683254 526320 683314 526491
rect 682886 525738 682946 525912
rect 683113 525738 683179 525741
rect 682886 525736 683179 525738
rect 682886 525680 683118 525736
rect 683174 525680 683179 525736
rect 682886 525678 683179 525680
rect 683113 525675 683179 525678
rect 671337 524922 671403 524925
rect 676262 524922 676322 525504
rect 671337 524920 676322 524922
rect 671337 524864 671342 524920
rect 671398 524864 676322 524920
rect 671337 524862 676322 524864
rect 671337 524859 671403 524862
rect 677918 524517 677978 524688
rect 677869 524512 677978 524517
rect 677869 524456 677874 524512
rect 677930 524456 677978 524512
rect 677869 524454 677978 524456
rect 677869 524451 677935 524454
rect 651833 524242 651899 524245
rect 650164 524240 651899 524242
rect 650164 524184 651838 524240
rect 651894 524184 651899 524240
rect 650164 524182 651899 524184
rect 651833 524179 651899 524182
rect 62113 519754 62179 519757
rect 62113 519752 64492 519754
rect 62113 519696 62118 519752
rect 62174 519696 64492 519752
rect 62113 519694 64492 519696
rect 62113 519691 62179 519694
rect 651465 511050 651531 511053
rect 650164 511048 651531 511050
rect 650164 510992 651470 511048
rect 651526 510992 651531 511048
rect 650164 510990 651531 510992
rect 651465 510987 651531 510990
rect 62113 506698 62179 506701
rect 62113 506696 64492 506698
rect 62113 506640 62118 506696
rect 62174 506640 64492 506696
rect 62113 506638 64492 506640
rect 62113 506635 62179 506638
rect 676990 503644 676996 503708
rect 677060 503706 677066 503708
rect 683113 503706 683179 503709
rect 677060 503704 683179 503706
rect 677060 503648 683118 503704
rect 683174 503648 683179 503704
rect 677060 503646 683179 503648
rect 677060 503644 677066 503646
rect 683113 503643 683179 503646
rect 674833 502618 674899 502621
rect 676029 502618 676095 502621
rect 674833 502616 676095 502618
rect 674833 502560 674838 502616
rect 674894 502560 676034 502616
rect 676090 502560 676095 502616
rect 674833 502558 676095 502560
rect 674833 502555 674899 502558
rect 676029 502555 676095 502558
rect 674925 502210 674991 502213
rect 675845 502210 675911 502213
rect 674925 502208 675911 502210
rect 674925 502152 674930 502208
rect 674986 502152 675850 502208
rect 675906 502152 675911 502208
rect 674925 502150 675911 502152
rect 674925 502147 674991 502150
rect 675845 502147 675911 502150
rect 670785 500986 670851 500989
rect 676397 500986 676463 500989
rect 670785 500984 676463 500986
rect 670785 500928 670790 500984
rect 670846 500928 676402 500984
rect 676458 500928 676463 500984
rect 670785 500926 676463 500928
rect 670785 500923 670851 500926
rect 676397 500923 676463 500926
rect 652569 497722 652635 497725
rect 650164 497720 652635 497722
rect 650164 497664 652574 497720
rect 652630 497664 652635 497720
rect 650164 497662 652635 497664
rect 652569 497659 652635 497662
rect 664437 494730 664503 494733
rect 683297 494730 683363 494733
rect 664437 494728 683363 494730
rect 664437 494672 664442 494728
rect 664498 494672 683302 494728
rect 683358 494672 683363 494728
rect 664437 494670 683363 494672
rect 664437 494667 664503 494670
rect 683297 494667 683363 494670
rect 62113 493642 62179 493645
rect 62113 493640 64492 493642
rect 62113 493584 62118 493640
rect 62174 493584 64492 493640
rect 62113 493582 64492 493584
rect 62113 493579 62179 493582
rect 676806 492764 676812 492828
rect 676876 492826 676882 492828
rect 677501 492826 677567 492829
rect 676876 492824 677567 492826
rect 676876 492768 677506 492824
rect 677562 492768 677567 492824
rect 676876 492766 677567 492768
rect 676876 492764 676882 492766
rect 677501 492763 677567 492766
rect 665817 492146 665883 492149
rect 665817 492144 676292 492146
rect 665817 492088 665822 492144
rect 665878 492088 676292 492144
rect 665817 492086 676292 492088
rect 665817 492083 665883 492086
rect 663750 491678 676292 491738
rect 661677 491602 661743 491605
rect 663750 491602 663810 491678
rect 661677 491600 663810 491602
rect 661677 491544 661682 491600
rect 661738 491544 663810 491600
rect 661677 491542 663810 491544
rect 661677 491539 661743 491542
rect 683297 491330 683363 491333
rect 683284 491328 683363 491330
rect 683284 491272 683302 491328
rect 683358 491272 683363 491328
rect 683284 491270 683363 491272
rect 683297 491267 683363 491270
rect 671797 490922 671863 490925
rect 671797 490920 676292 490922
rect 671797 490864 671802 490920
rect 671858 490864 676292 490920
rect 671797 490862 676292 490864
rect 671797 490859 671863 490862
rect 671429 490514 671495 490517
rect 671429 490512 676292 490514
rect 671429 490456 671434 490512
rect 671490 490456 676292 490512
rect 671429 490454 676292 490456
rect 671429 490451 671495 490454
rect 672625 490106 672691 490109
rect 672625 490104 676292 490106
rect 672625 490048 672630 490104
rect 672686 490048 676292 490104
rect 672625 490046 676292 490048
rect 672625 490043 672691 490046
rect 671797 489698 671863 489701
rect 671797 489696 676292 489698
rect 671797 489640 671802 489696
rect 671858 489640 676292 489696
rect 671797 489638 676292 489640
rect 671797 489635 671863 489638
rect 670969 489290 671035 489293
rect 670969 489288 676292 489290
rect 670969 489232 670974 489288
rect 671030 489232 676292 489288
rect 670969 489230 676292 489232
rect 670969 489227 671035 489230
rect 675886 488820 675892 488884
rect 675956 488882 675962 488884
rect 675956 488822 676292 488882
rect 675956 488820 675962 488822
rect 671613 488474 671679 488477
rect 671613 488472 676292 488474
rect 671613 488416 671618 488472
rect 671674 488416 676292 488472
rect 671613 488414 676292 488416
rect 671613 488411 671679 488414
rect 676029 488066 676095 488069
rect 676029 488064 676292 488066
rect 676029 488008 676034 488064
rect 676090 488008 676292 488064
rect 676029 488006 676292 488008
rect 676029 488003 676095 488006
rect 675109 487658 675175 487661
rect 675109 487656 676292 487658
rect 675109 487600 675114 487656
rect 675170 487600 676292 487656
rect 675109 487598 676292 487600
rect 675109 487595 675175 487598
rect 674005 487250 674071 487253
rect 675845 487250 675911 487253
rect 683113 487250 683179 487253
rect 674005 487248 675911 487250
rect 674005 487192 674010 487248
rect 674066 487192 675850 487248
rect 675906 487192 675911 487248
rect 674005 487190 675911 487192
rect 683100 487248 683179 487250
rect 683100 487192 683118 487248
rect 683174 487192 683179 487248
rect 683100 487190 683179 487192
rect 674005 487187 674071 487190
rect 675845 487187 675911 487190
rect 683113 487187 683179 487190
rect 678237 486842 678303 486845
rect 678237 486840 678316 486842
rect 678237 486784 678242 486840
rect 678298 486784 678316 486840
rect 678237 486782 678316 486784
rect 678237 486779 678303 486782
rect 675293 486434 675359 486437
rect 675293 486432 676292 486434
rect 675293 486376 675298 486432
rect 675354 486376 676292 486432
rect 675293 486374 676292 486376
rect 675293 486371 675359 486374
rect 673821 486162 673887 486165
rect 675661 486162 675727 486165
rect 673821 486160 675727 486162
rect 673821 486104 673826 486160
rect 673882 486104 675666 486160
rect 675722 486104 675727 486160
rect 673821 486102 675727 486104
rect 673821 486099 673887 486102
rect 675661 486099 675727 486102
rect 675894 485966 676292 486026
rect 669037 485890 669103 485893
rect 675894 485890 675954 485966
rect 669037 485888 675954 485890
rect 669037 485832 669042 485888
rect 669098 485832 675954 485888
rect 669037 485830 675954 485832
rect 669037 485827 669103 485830
rect 671153 485618 671219 485621
rect 671153 485616 676292 485618
rect 671153 485560 671158 485616
rect 671214 485560 676292 485616
rect 671153 485558 676292 485560
rect 671153 485555 671219 485558
rect 667381 485210 667447 485213
rect 667381 485208 676292 485210
rect 667381 485152 667386 485208
rect 667442 485152 676292 485208
rect 667381 485150 676292 485152
rect 667381 485147 667447 485150
rect 673177 484802 673243 484805
rect 673177 484800 676292 484802
rect 673177 484744 673182 484800
rect 673238 484744 676292 484800
rect 673177 484742 676292 484744
rect 673177 484739 673243 484742
rect 651465 484530 651531 484533
rect 650164 484528 651531 484530
rect 650164 484472 651470 484528
rect 651526 484472 651531 484528
rect 650164 484470 651531 484472
rect 651465 484467 651531 484470
rect 675845 484394 675911 484397
rect 675845 484392 676292 484394
rect 675845 484336 675850 484392
rect 675906 484336 676292 484392
rect 675845 484334 676292 484336
rect 675845 484331 675911 484334
rect 669221 483986 669287 483989
rect 669221 483984 676292 483986
rect 669221 483928 669226 483984
rect 669282 483928 676292 483984
rect 669221 483926 676292 483928
rect 669221 483923 669287 483926
rect 674373 483578 674439 483581
rect 674373 483576 676292 483578
rect 674373 483520 674378 483576
rect 674434 483520 676292 483576
rect 674373 483518 676292 483520
rect 674373 483515 674439 483518
rect 675661 483170 675727 483173
rect 675661 483168 676292 483170
rect 675661 483112 675666 483168
rect 675722 483112 676292 483168
rect 675661 483110 676292 483112
rect 675661 483107 675727 483110
rect 683297 482762 683363 482765
rect 683284 482760 683363 482762
rect 683284 482704 683302 482760
rect 683358 482704 683363 482760
rect 683284 482702 683363 482704
rect 683297 482699 683363 482702
rect 670417 482354 670483 482357
rect 670417 482352 676292 482354
rect 670417 482296 670422 482352
rect 670478 482296 676292 482352
rect 670417 482294 676292 482296
rect 670417 482291 670483 482294
rect 675661 481946 675727 481949
rect 675661 481944 676292 481946
rect 675661 481888 675666 481944
rect 675722 481888 676292 481944
rect 675661 481886 676292 481888
rect 675661 481883 675727 481886
rect 683113 481538 683179 481541
rect 677212 481536 683179 481538
rect 677212 481508 683118 481536
rect 677182 481480 683118 481508
rect 683174 481480 683179 481536
rect 677182 481478 683179 481480
rect 677182 481100 677242 481478
rect 683113 481475 683179 481478
rect 675845 480722 675911 480725
rect 675845 480720 676292 480722
rect 675845 480664 675850 480720
rect 675906 480664 676292 480720
rect 675845 480662 676292 480664
rect 675845 480659 675911 480662
rect 62113 480586 62179 480589
rect 62113 480584 64492 480586
rect 62113 480528 62118 480584
rect 62174 480528 64492 480584
rect 62113 480526 64492 480528
rect 62113 480523 62179 480526
rect 674598 475356 674604 475420
rect 674668 475418 674674 475420
rect 676213 475418 676279 475421
rect 674668 475416 676279 475418
rect 674668 475360 676218 475416
rect 676274 475360 676279 475416
rect 674668 475358 676279 475360
rect 674668 475356 674674 475358
rect 676213 475355 676279 475358
rect 651465 471202 651531 471205
rect 650164 471200 651531 471202
rect 650164 471144 651470 471200
rect 651526 471144 651531 471200
rect 650164 471142 651531 471144
rect 651465 471139 651531 471142
rect 62113 467530 62179 467533
rect 62113 467528 64492 467530
rect 62113 467472 62118 467528
rect 62174 467472 64492 467528
rect 62113 467470 64492 467472
rect 62113 467467 62179 467470
rect 652385 457874 652451 457877
rect 650164 457872 652451 457874
rect 650164 457816 652390 457872
rect 652446 457816 652451 457872
rect 650164 457814 652451 457816
rect 652385 457811 652451 457814
rect 672901 456514 672967 456517
rect 676949 456514 677015 456517
rect 672901 456512 677015 456514
rect 672901 456456 672906 456512
rect 672962 456456 676954 456512
rect 677010 456456 677015 456512
rect 672901 456454 677015 456456
rect 672901 456451 672967 456454
rect 676949 456451 677015 456454
rect 667841 456242 667907 456245
rect 673941 456242 674007 456245
rect 667841 456240 674007 456242
rect 667841 456184 667846 456240
rect 667902 456184 673946 456240
rect 674002 456184 674007 456240
rect 667841 456182 674007 456184
rect 667841 456179 667907 456182
rect 673941 456179 674007 456182
rect 673821 455970 673887 455973
rect 676213 455970 676279 455973
rect 673821 455968 676279 455970
rect 673821 455912 673826 455968
rect 673882 455912 676218 455968
rect 676274 455912 676279 455968
rect 673821 455910 676279 455912
rect 673821 455907 673887 455910
rect 676213 455907 676279 455910
rect 671981 455698 672047 455701
rect 673591 455698 673657 455701
rect 671981 455696 673657 455698
rect 671981 455640 671986 455696
rect 672042 455640 673596 455696
rect 673652 455640 673657 455696
rect 671981 455638 673657 455640
rect 671981 455635 672047 455638
rect 673591 455635 673657 455638
rect 670601 455426 670667 455429
rect 673269 455426 673335 455429
rect 670601 455424 673335 455426
rect 670601 455368 670606 455424
rect 670662 455368 673274 455424
rect 673330 455368 673335 455424
rect 670601 455366 673335 455368
rect 670601 455363 670667 455366
rect 673269 455363 673335 455366
rect 673381 455290 673447 455293
rect 673862 455290 673868 455292
rect 673381 455288 673868 455290
rect 673381 455232 673386 455288
rect 673442 455232 673868 455288
rect 673381 455230 673868 455232
rect 673381 455227 673447 455230
rect 673862 455228 673868 455230
rect 673932 455228 673938 455292
rect 669773 455154 669839 455157
rect 672073 455154 672139 455157
rect 669773 455152 672139 455154
rect 669773 455096 669778 455152
rect 669834 455096 672078 455152
rect 672134 455096 672139 455152
rect 669773 455094 672139 455096
rect 669773 455091 669839 455094
rect 672073 455091 672139 455094
rect 673039 454882 673105 454885
rect 675477 454882 675543 454885
rect 673039 454880 675543 454882
rect 673039 454824 673044 454880
rect 673100 454824 675482 454880
rect 675538 454824 675543 454880
rect 673039 454822 675543 454824
rect 673039 454819 673105 454822
rect 675477 454819 675543 454822
rect 62113 454610 62179 454613
rect 673157 454610 673223 454613
rect 676765 454610 676831 454613
rect 62113 454608 64492 454610
rect 62113 454552 62118 454608
rect 62174 454552 64492 454608
rect 62113 454550 64492 454552
rect 673157 454608 676831 454610
rect 673157 454552 673162 454608
rect 673218 454552 676770 454608
rect 676826 454552 676831 454608
rect 673157 454550 676831 454552
rect 62113 454547 62179 454550
rect 673157 454547 673223 454550
rect 676765 454547 676831 454550
rect 672809 454202 672875 454205
rect 675845 454202 675911 454205
rect 672809 454200 675911 454202
rect 672809 454144 672814 454200
rect 672870 454144 675850 454200
rect 675906 454144 675911 454200
rect 672809 454142 675911 454144
rect 672809 454139 672875 454142
rect 675845 454139 675911 454142
rect 672717 453930 672783 453933
rect 675201 453930 675267 453933
rect 672717 453928 675267 453930
rect 672717 453872 672722 453928
rect 672778 453872 675206 453928
rect 675262 453872 675267 453928
rect 672717 453870 675267 453872
rect 672717 453867 672783 453870
rect 675201 453867 675267 453870
rect 675334 453732 675340 453796
rect 675404 453794 675410 453796
rect 676029 453794 676095 453797
rect 675404 453792 676095 453794
rect 675404 453736 676034 453792
rect 676090 453736 676095 453792
rect 675404 453734 676095 453736
rect 675404 453732 675410 453734
rect 676029 453731 676095 453734
rect 651465 444546 651531 444549
rect 650164 444544 651531 444546
rect 650164 444488 651470 444544
rect 651526 444488 651531 444544
rect 650164 444486 651531 444488
rect 651465 444483 651531 444486
rect 62113 441554 62179 441557
rect 62113 441552 64492 441554
rect 62113 441496 62118 441552
rect 62174 441496 64492 441552
rect 62113 441494 64492 441496
rect 62113 441491 62179 441494
rect 651465 431354 651531 431357
rect 650164 431352 651531 431354
rect 650164 431296 651470 431352
rect 651526 431296 651531 431352
rect 650164 431294 651531 431296
rect 651465 431291 651531 431294
rect 50337 430946 50403 430949
rect 41492 430944 50403 430946
rect 41492 430888 50342 430944
rect 50398 430888 50403 430944
rect 41492 430886 50403 430888
rect 50337 430883 50403 430886
rect 54477 430538 54543 430541
rect 41492 430536 54543 430538
rect 41492 430480 54482 430536
rect 54538 430480 54543 430536
rect 41492 430478 54543 430480
rect 54477 430475 54543 430478
rect 47577 430130 47643 430133
rect 41492 430128 47643 430130
rect 41492 430072 47582 430128
rect 47638 430072 47643 430128
rect 41492 430070 47643 430072
rect 47577 430067 47643 430070
rect 45645 429722 45711 429725
rect 41492 429720 45711 429722
rect 41492 429664 45650 429720
rect 45706 429664 45711 429720
rect 41492 429662 45711 429664
rect 45645 429659 45711 429662
rect 45829 429314 45895 429317
rect 41492 429312 45895 429314
rect 41492 429256 45834 429312
rect 45890 429256 45895 429312
rect 41492 429254 45895 429256
rect 45829 429251 45895 429254
rect 46013 428906 46079 428909
rect 41492 428904 46079 428906
rect 41492 428848 46018 428904
rect 46074 428848 46079 428904
rect 41492 428846 46079 428848
rect 46013 428843 46079 428846
rect 45645 428498 45711 428501
rect 41492 428496 45711 428498
rect 41492 428440 45650 428496
rect 45706 428440 45711 428496
rect 41492 428438 45711 428440
rect 45645 428435 45711 428438
rect 62113 428498 62179 428501
rect 62113 428496 64492 428498
rect 62113 428440 62118 428496
rect 62174 428440 64492 428496
rect 62113 428438 64492 428440
rect 62113 428435 62179 428438
rect 44633 428090 44699 428093
rect 41492 428088 44699 428090
rect 41492 428032 44638 428088
rect 44694 428032 44699 428088
rect 41492 428030 44699 428032
rect 44633 428027 44699 428030
rect 44725 427682 44791 427685
rect 41492 427680 44791 427682
rect 41492 427624 44730 427680
rect 44786 427624 44791 427680
rect 41492 427622 44791 427624
rect 44725 427619 44791 427622
rect 44265 427274 44331 427277
rect 41492 427272 44331 427274
rect 41492 427216 44270 427272
rect 44326 427216 44331 427272
rect 41492 427214 44331 427216
rect 44265 427211 44331 427214
rect 44265 426866 44331 426869
rect 41492 426864 44331 426866
rect 41492 426808 44270 426864
rect 44326 426808 44331 426864
rect 41492 426806 44331 426808
rect 44265 426803 44331 426806
rect 46933 426458 46999 426461
rect 41492 426456 46999 426458
rect 41492 426400 46938 426456
rect 46994 426400 46999 426456
rect 41492 426398 46999 426400
rect 46933 426395 46999 426398
rect 41321 426050 41387 426053
rect 41308 426048 41387 426050
rect 41308 425992 41326 426048
rect 41382 425992 41387 426048
rect 41308 425990 41387 425992
rect 41321 425987 41387 425990
rect 40953 425642 41019 425645
rect 40940 425640 41019 425642
rect 40940 425584 40958 425640
rect 41014 425584 41019 425640
rect 40940 425582 41019 425584
rect 40953 425579 41019 425582
rect 41822 425234 41828 425236
rect 41492 425174 41828 425234
rect 41822 425172 41828 425174
rect 41892 425172 41898 425236
rect 42006 424826 42012 424828
rect 41492 424766 42012 424826
rect 42006 424764 42012 424766
rect 42076 424764 42082 424828
rect 33777 424418 33843 424421
rect 33764 424416 33843 424418
rect 33764 424360 33782 424416
rect 33838 424360 33843 424416
rect 33764 424358 33843 424360
rect 33777 424355 33843 424358
rect 42793 424010 42859 424013
rect 41492 424008 42859 424010
rect 41492 423952 42798 424008
rect 42854 423952 42859 424008
rect 41492 423950 42859 423952
rect 42793 423947 42859 423950
rect 45093 423602 45159 423605
rect 41492 423600 45159 423602
rect 41492 423544 45098 423600
rect 45154 423544 45159 423600
rect 41492 423542 45159 423544
rect 45093 423539 45159 423542
rect 44449 423194 44515 423197
rect 41492 423192 44515 423194
rect 41492 423136 44454 423192
rect 44510 423136 44515 423192
rect 41492 423134 44515 423136
rect 44449 423131 44515 423134
rect 41781 422786 41847 422789
rect 41492 422784 41847 422786
rect 41492 422728 41786 422784
rect 41842 422728 41847 422784
rect 41492 422726 41847 422728
rect 41781 422723 41847 422726
rect 44909 422378 44975 422381
rect 41492 422376 44975 422378
rect 41492 422320 44914 422376
rect 44970 422320 44975 422376
rect 41492 422318 44975 422320
rect 44909 422315 44975 422318
rect 42006 421970 42012 421972
rect 41492 421910 42012 421970
rect 42006 421908 42012 421910
rect 42076 421908 42082 421972
rect 45461 421562 45527 421565
rect 41492 421560 45527 421562
rect 41492 421504 45466 421560
rect 45522 421504 45527 421560
rect 41492 421502 45527 421504
rect 45461 421499 45527 421502
rect 45277 421154 45343 421157
rect 41492 421152 45343 421154
rect 41492 421096 45282 421152
rect 45338 421096 45343 421152
rect 41492 421094 45343 421096
rect 45277 421091 45343 421094
rect 43253 420746 43319 420749
rect 41492 420744 43319 420746
rect 41492 420688 43258 420744
rect 43314 420688 43319 420744
rect 41492 420686 43319 420688
rect 43253 420683 43319 420686
rect 41462 419930 41522 420308
rect 42517 419930 42583 419933
rect 41462 419928 42583 419930
rect 41462 419900 42522 419928
rect 41492 419872 42522 419900
rect 42578 419872 42583 419928
rect 41492 419870 42583 419872
rect 42517 419867 42583 419870
rect 41492 419462 41844 419522
rect 41784 419250 41844 419462
rect 43069 419250 43135 419253
rect 41784 419248 43135 419250
rect 41784 419192 43074 419248
rect 43130 419192 43135 419248
rect 41784 419190 43135 419192
rect 43069 419187 43135 419190
rect 41137 418842 41203 418845
rect 41454 418842 41460 418844
rect 41137 418840 41460 418842
rect 41137 418784 41142 418840
rect 41198 418784 41460 418840
rect 41137 418782 41460 418784
rect 41137 418779 41203 418782
rect 41454 418780 41460 418782
rect 41524 418780 41530 418844
rect 40718 418508 40724 418572
rect 40788 418570 40794 418572
rect 41781 418570 41847 418573
rect 40788 418568 41847 418570
rect 40788 418512 41786 418568
rect 41842 418512 41847 418568
rect 40788 418510 41847 418512
rect 40788 418508 40794 418510
rect 41781 418507 41847 418510
rect 40534 418236 40540 418300
rect 40604 418298 40610 418300
rect 42006 418298 42012 418300
rect 40604 418238 42012 418298
rect 40604 418236 40610 418238
rect 42006 418236 42012 418238
rect 42076 418236 42082 418300
rect 651833 418026 651899 418029
rect 650164 418024 651899 418026
rect 650164 417968 651838 418024
rect 651894 417968 651899 418024
rect 650164 417966 651899 417968
rect 651833 417963 651899 417966
rect 62757 415442 62823 415445
rect 62757 415440 64492 415442
rect 62757 415384 62762 415440
rect 62818 415384 64492 415440
rect 62757 415382 64492 415384
rect 62757 415379 62823 415382
rect 42057 411906 42123 411909
rect 42609 411906 42675 411909
rect 42057 411904 42675 411906
rect 42057 411848 42062 411904
rect 42118 411848 42614 411904
rect 42670 411848 42675 411904
rect 42057 411846 42675 411848
rect 42057 411843 42123 411846
rect 42609 411843 42675 411846
rect 660297 411906 660363 411909
rect 683297 411906 683363 411909
rect 660297 411904 683363 411906
rect 660297 411848 660302 411904
rect 660358 411848 683302 411904
rect 683358 411848 683363 411904
rect 660297 411846 683363 411848
rect 660297 411843 660363 411846
rect 683297 411843 683363 411846
rect 675334 410484 675340 410548
rect 675404 410546 675410 410548
rect 676029 410546 676095 410549
rect 675404 410544 676095 410546
rect 675404 410488 676034 410544
rect 676090 410488 676095 410544
rect 675404 410486 676095 410488
rect 675404 410484 675410 410486
rect 676029 410483 676095 410486
rect 40718 409396 40724 409460
rect 40788 409458 40794 409460
rect 41781 409458 41847 409461
rect 40788 409456 41847 409458
rect 40788 409400 41786 409456
rect 41842 409400 41847 409456
rect 40788 409398 41847 409400
rect 40788 409396 40794 409398
rect 41781 409395 41847 409398
rect 42425 408506 42491 408509
rect 55857 408506 55923 408509
rect 42425 408504 55923 408506
rect 42425 408448 42430 408504
rect 42486 408448 55862 408504
rect 55918 408448 55923 408504
rect 42425 408446 55923 408448
rect 42425 408443 42491 408446
rect 55857 408443 55923 408446
rect 42425 407826 42491 407829
rect 45277 407826 45343 407829
rect 42425 407824 45343 407826
rect 42425 407768 42430 407824
rect 42486 407768 45282 407824
rect 45338 407768 45343 407824
rect 42425 407766 45343 407768
rect 42425 407763 42491 407766
rect 45277 407763 45343 407766
rect 42057 406738 42123 406741
rect 45461 406738 45527 406741
rect 42057 406736 45527 406738
rect 42057 406680 42062 406736
rect 42118 406680 45466 406736
rect 45522 406680 45527 406736
rect 42057 406678 45527 406680
rect 42057 406675 42123 406678
rect 45461 406675 45527 406678
rect 41781 406332 41847 406333
rect 41781 406328 41828 406332
rect 41892 406330 41898 406332
rect 661861 406330 661927 406333
rect 683113 406330 683179 406333
rect 41781 406272 41786 406328
rect 41781 406268 41828 406272
rect 41892 406270 41938 406330
rect 661861 406328 683179 406330
rect 661861 406272 661866 406328
rect 661922 406272 683118 406328
rect 683174 406272 683179 406328
rect 661861 406270 683179 406272
rect 41892 406268 41898 406270
rect 41781 406267 41847 406268
rect 661861 406267 661927 406270
rect 683113 406267 683179 406270
rect 42425 405650 42491 405653
rect 44909 405650 44975 405653
rect 42425 405648 44975 405650
rect 42425 405592 42430 405648
rect 42486 405592 44914 405648
rect 44970 405592 44975 405648
rect 42425 405590 44975 405592
rect 42425 405587 42491 405590
rect 44909 405587 44975 405590
rect 651465 404698 651531 404701
rect 650164 404696 651531 404698
rect 650164 404640 651470 404696
rect 651526 404640 651531 404696
rect 650164 404638 651531 404640
rect 651465 404635 651531 404638
rect 40534 403820 40540 403884
rect 40604 403882 40610 403884
rect 41781 403882 41847 403885
rect 40604 403880 41847 403882
rect 40604 403824 41786 403880
rect 41842 403824 41847 403880
rect 40604 403822 41847 403824
rect 40604 403820 40610 403822
rect 41781 403819 41847 403822
rect 669405 403746 669471 403749
rect 676262 403746 676322 403852
rect 683297 403746 683363 403749
rect 669405 403744 676322 403746
rect 669405 403688 669410 403744
rect 669466 403688 676322 403744
rect 669405 403686 676322 403688
rect 683254 403744 683363 403746
rect 683254 403688 683302 403744
rect 683358 403688 683363 403744
rect 669405 403683 669471 403686
rect 683254 403683 683363 403688
rect 683254 403444 683314 403683
rect 683113 403338 683179 403341
rect 682886 403336 683179 403338
rect 682886 403280 683118 403336
rect 683174 403280 683179 403336
rect 682886 403278 683179 403280
rect 682886 403036 682946 403278
rect 683113 403275 683179 403278
rect 42333 402930 42399 402933
rect 44449 402930 44515 402933
rect 42333 402928 44515 402930
rect 42333 402872 42338 402928
rect 42394 402872 44454 402928
rect 44510 402872 44515 402928
rect 42333 402870 44515 402872
rect 42333 402867 42399 402870
rect 44449 402867 44515 402870
rect 42425 402522 42491 402525
rect 45093 402522 45159 402525
rect 42425 402520 45159 402522
rect 42425 402464 42430 402520
rect 42486 402464 45098 402520
rect 45154 402464 45159 402520
rect 42425 402462 45159 402464
rect 42425 402459 42491 402462
rect 45093 402459 45159 402462
rect 671429 402522 671495 402525
rect 676262 402522 676322 402628
rect 671429 402520 676322 402522
rect 671429 402464 671434 402520
rect 671490 402464 676322 402520
rect 671429 402462 676322 402464
rect 671429 402459 671495 402462
rect 62113 402386 62179 402389
rect 62113 402384 64492 402386
rect 62113 402328 62118 402384
rect 62174 402328 64492 402384
rect 62113 402326 64492 402328
rect 62113 402323 62179 402326
rect 674189 402250 674255 402253
rect 674189 402248 676292 402250
rect 674189 402192 674194 402248
rect 674250 402192 676292 402248
rect 674189 402190 676292 402192
rect 674189 402187 674255 402190
rect 41781 401980 41847 401981
rect 41781 401976 41828 401980
rect 41892 401978 41898 401980
rect 41781 401920 41786 401976
rect 41781 401916 41828 401920
rect 41892 401918 41938 401978
rect 41892 401916 41898 401918
rect 41781 401915 41847 401916
rect 671797 401706 671863 401709
rect 676262 401706 676322 401812
rect 671797 401704 676322 401706
rect 671797 401648 671802 401704
rect 671858 401648 676322 401704
rect 671797 401646 676322 401648
rect 671797 401643 671863 401646
rect 674649 401434 674715 401437
rect 674649 401432 676292 401434
rect 674649 401376 674654 401432
rect 674710 401376 676292 401432
rect 674649 401374 676292 401376
rect 674649 401371 674715 401374
rect 676806 401236 676812 401300
rect 676876 401236 676882 401300
rect 676814 400996 676874 401236
rect 672809 400482 672875 400485
rect 676262 400482 676322 400588
rect 672809 400480 676322 400482
rect 672809 400424 672814 400480
rect 672870 400424 676322 400480
rect 672809 400422 676322 400424
rect 672809 400419 672875 400422
rect 676029 400210 676095 400213
rect 676029 400208 676292 400210
rect 676029 400152 676034 400208
rect 676090 400152 676292 400208
rect 676029 400150 676292 400152
rect 676029 400147 676095 400150
rect 42425 399802 42491 399805
rect 46933 399802 46999 399805
rect 42425 399800 46999 399802
rect 42425 399744 42430 399800
rect 42486 399744 46938 399800
rect 46994 399744 46999 399800
rect 42425 399742 46999 399744
rect 42425 399739 42491 399742
rect 46933 399739 46999 399742
rect 673177 399666 673243 399669
rect 676262 399666 676322 399772
rect 673177 399664 676322 399666
rect 673177 399608 673182 399664
rect 673238 399608 676322 399664
rect 673177 399606 676322 399608
rect 673177 399603 673243 399606
rect 676029 399394 676095 399397
rect 676029 399392 676292 399394
rect 676029 399336 676034 399392
rect 676090 399336 676292 399392
rect 676029 399334 676292 399336
rect 676029 399331 676095 399334
rect 41454 398788 41460 398852
rect 41524 398850 41530 398852
rect 41781 398850 41847 398853
rect 41524 398848 41847 398850
rect 41524 398792 41786 398848
rect 41842 398792 41847 398848
rect 41524 398790 41847 398792
rect 41524 398788 41530 398790
rect 41781 398787 41847 398790
rect 676070 398788 676076 398852
rect 676140 398850 676146 398852
rect 676262 398850 676322 398956
rect 676140 398790 676322 398850
rect 676140 398788 676146 398790
rect 676262 398445 676322 398548
rect 676213 398440 676322 398445
rect 676213 398384 676218 398440
rect 676274 398384 676322 398440
rect 676213 398382 676322 398384
rect 676213 398379 676279 398382
rect 676446 398037 676506 398140
rect 676397 398032 676506 398037
rect 676397 397976 676402 398032
rect 676458 397976 676506 398032
rect 676397 397974 676506 397976
rect 676397 397971 676463 397974
rect 681046 397629 681106 397732
rect 680997 397624 681106 397629
rect 680997 397568 681002 397624
rect 681058 397568 681106 397624
rect 680997 397566 681106 397568
rect 680997 397563 681063 397566
rect 672993 397218 673059 397221
rect 676262 397218 676322 397324
rect 672993 397216 676322 397218
rect 672993 397160 672998 397216
rect 673054 397160 676322 397216
rect 672993 397158 676322 397160
rect 672993 397155 673059 397158
rect 676630 396812 676690 396916
rect 676622 396748 676628 396812
rect 676692 396748 676698 396812
rect 673361 396402 673427 396405
rect 676262 396402 676322 396508
rect 673361 396400 676322 396402
rect 673361 396344 673366 396400
rect 673422 396344 676322 396400
rect 673361 396342 676322 396344
rect 673361 396339 673427 396342
rect 673821 396130 673887 396133
rect 673821 396128 676292 396130
rect 673821 396072 673826 396128
rect 673882 396072 676292 396128
rect 673821 396070 676292 396072
rect 673821 396067 673887 396070
rect 674005 395722 674071 395725
rect 674005 395720 676292 395722
rect 674005 395664 674010 395720
rect 674066 395664 676292 395720
rect 674005 395662 676292 395664
rect 674005 395659 674071 395662
rect 676262 395180 676322 395284
rect 676254 395116 676260 395180
rect 676324 395116 676330 395180
rect 676446 394772 676506 394876
rect 676438 394708 676444 394772
rect 676508 394708 676514 394772
rect 674465 394498 674531 394501
rect 674465 394496 676292 394498
rect 674465 394440 674470 394496
rect 674526 394440 676292 394496
rect 674465 394438 676292 394440
rect 674465 394435 674531 394438
rect 672625 393954 672691 393957
rect 676262 393954 676322 394060
rect 672625 393952 676322 393954
rect 672625 393896 672630 393952
rect 672686 393896 676322 393952
rect 672625 393894 676322 393896
rect 672625 393891 672691 393894
rect 671981 393546 672047 393549
rect 676262 393546 676322 393652
rect 671981 393544 676322 393546
rect 671981 393488 671986 393544
rect 672042 393488 676322 393544
rect 671981 393486 676322 393488
rect 671981 393483 672047 393486
rect 683070 392733 683130 393244
rect 683021 392728 683130 392733
rect 683021 392672 683026 392728
rect 683082 392672 683130 392728
rect 683021 392670 683130 392672
rect 683021 392667 683087 392670
rect 672349 392322 672415 392325
rect 676262 392322 676322 392428
rect 672349 392320 676322 392322
rect 672349 392264 672354 392320
rect 672410 392264 676322 392320
rect 672349 392262 676322 392264
rect 672349 392259 672415 392262
rect 652569 391506 652635 391509
rect 650164 391504 652635 391506
rect 650164 391448 652574 391504
rect 652630 391448 652635 391504
rect 650164 391446 652635 391448
rect 652569 391443 652635 391446
rect 62113 389330 62179 389333
rect 62113 389328 64492 389330
rect 62113 389272 62118 389328
rect 62174 389272 64492 389328
rect 62113 389270 64492 389272
rect 62113 389267 62179 389270
rect 675886 388996 675892 389060
rect 675956 389058 675962 389060
rect 683021 389058 683087 389061
rect 675956 389056 683087 389058
rect 675956 389000 683026 389056
rect 683082 389000 683087 389056
rect 675956 388998 683087 389000
rect 675956 388996 675962 388998
rect 683021 388995 683087 388998
rect 42057 387698 42123 387701
rect 41492 387696 42123 387698
rect 41492 387640 42062 387696
rect 42118 387640 42123 387696
rect 41492 387638 42123 387640
rect 42057 387635 42123 387638
rect 675702 387636 675708 387700
rect 675772 387698 675778 387700
rect 680997 387698 681063 387701
rect 675772 387696 681063 387698
rect 675772 387640 681002 387696
rect 681058 387640 681063 387696
rect 675772 387638 681063 387640
rect 675772 387636 675778 387638
rect 680997 387635 681063 387638
rect 41873 387290 41939 387293
rect 45829 387290 45895 387293
rect 41873 387288 45895 387290
rect 41094 387157 41154 387260
rect 41873 387232 41878 387288
rect 41934 387232 45834 387288
rect 45890 387232 45895 387288
rect 41873 387230 45895 387232
rect 41873 387227 41939 387230
rect 45829 387227 45895 387230
rect 41094 387152 41203 387157
rect 41094 387096 41142 387152
rect 41198 387096 41203 387152
rect 41094 387094 41203 387096
rect 41137 387091 41203 387094
rect 48957 387018 49023 387021
rect 41830 387016 49023 387018
rect 41830 386960 48962 387016
rect 49018 386960 49023 387016
rect 41830 386958 49023 386960
rect 41830 386882 41890 386958
rect 48957 386955 49023 386958
rect 41492 386822 41890 386882
rect 42057 386746 42123 386749
rect 51717 386746 51783 386749
rect 42057 386744 51783 386746
rect 42057 386688 42062 386744
rect 42118 386688 51722 386744
rect 51778 386688 51783 386744
rect 42057 386686 51783 386688
rect 42057 386683 42123 386686
rect 51717 386683 51783 386686
rect 41873 386474 41939 386477
rect 41492 386472 41939 386474
rect 41492 386416 41878 386472
rect 41934 386416 41939 386472
rect 41492 386414 41939 386416
rect 41873 386411 41939 386414
rect 42057 386474 42123 386477
rect 51901 386474 51967 386477
rect 42057 386472 51967 386474
rect 42057 386416 42062 386472
rect 42118 386416 51906 386472
rect 51962 386416 51967 386472
rect 42057 386414 51967 386416
rect 42057 386411 42123 386414
rect 51901 386411 51967 386414
rect 45277 386066 45343 386069
rect 41492 386064 45343 386066
rect 41492 386008 45282 386064
rect 45338 386008 45343 386064
rect 41492 386006 45343 386008
rect 45277 386003 45343 386006
rect 45645 385658 45711 385661
rect 41492 385656 45711 385658
rect 41492 385600 45650 385656
rect 45706 385600 45711 385656
rect 41492 385598 45711 385600
rect 45645 385595 45711 385598
rect 45093 385250 45159 385253
rect 41492 385248 45159 385250
rect 41492 385192 45098 385248
rect 45154 385192 45159 385248
rect 41492 385190 45159 385192
rect 45093 385187 45159 385190
rect 675753 384978 675819 384981
rect 676622 384978 676628 384980
rect 675753 384976 676628 384978
rect 675753 384920 675758 384976
rect 675814 384920 676628 384976
rect 675753 384918 676628 384920
rect 675753 384915 675819 384918
rect 676622 384916 676628 384918
rect 676692 384916 676698 384980
rect 44725 384842 44791 384845
rect 41492 384840 44791 384842
rect 41492 384784 44730 384840
rect 44786 384784 44791 384840
rect 41492 384782 44791 384784
rect 44725 384779 44791 384782
rect 45829 384434 45895 384437
rect 41492 384432 45895 384434
rect 41492 384376 45834 384432
rect 45890 384376 45895 384432
rect 41492 384374 45895 384376
rect 45829 384371 45895 384374
rect 44265 384026 44331 384029
rect 41492 384024 44331 384026
rect 41492 383968 44270 384024
rect 44326 383968 44331 384024
rect 41492 383966 44331 383968
rect 44265 383963 44331 383966
rect 45645 383618 45711 383621
rect 41492 383616 45711 383618
rect 41492 383560 45650 383616
rect 45706 383560 45711 383616
rect 41492 383558 45711 383560
rect 45645 383555 45711 383558
rect 35390 383077 35450 383180
rect 35390 383072 35499 383077
rect 35390 383016 35438 383072
rect 35494 383016 35499 383072
rect 35390 383014 35499 383016
rect 35433 383011 35499 383014
rect 35574 382669 35634 382772
rect 35574 382664 35683 382669
rect 35574 382608 35622 382664
rect 35678 382608 35683 382664
rect 35574 382606 35683 382608
rect 35617 382603 35683 382606
rect 35758 382261 35818 382364
rect 35758 382256 35867 382261
rect 35758 382200 35806 382256
rect 35862 382200 35867 382256
rect 35758 382198 35867 382200
rect 35801 382195 35867 382198
rect 41505 382258 41571 382261
rect 42793 382258 42859 382261
rect 41505 382256 42859 382258
rect 41505 382200 41510 382256
rect 41566 382200 42798 382256
rect 42854 382200 42859 382256
rect 41505 382198 42859 382200
rect 41505 382195 41571 382198
rect 42793 382195 42859 382198
rect 673361 382258 673427 382261
rect 675385 382258 675451 382261
rect 673361 382256 675451 382258
rect 673361 382200 673366 382256
rect 673422 382200 675390 382256
rect 675446 382200 675451 382256
rect 673361 382198 675451 382200
rect 673361 382195 673427 382198
rect 675385 382195 675451 382198
rect 41462 381852 41522 381956
rect 41454 381788 41460 381852
rect 41524 381788 41530 381852
rect 35574 381445 35634 381548
rect 35525 381440 35634 381445
rect 35801 381442 35867 381445
rect 35525 381384 35530 381440
rect 35586 381384 35634 381440
rect 35525 381382 35634 381384
rect 35758 381440 35867 381442
rect 35758 381384 35806 381440
rect 35862 381384 35867 381440
rect 35525 381379 35591 381382
rect 35758 381379 35867 381384
rect 673821 381442 673887 381445
rect 675109 381442 675175 381445
rect 673821 381440 675175 381442
rect 673821 381384 673826 381440
rect 673882 381384 675114 381440
rect 675170 381384 675175 381440
rect 673821 381382 675175 381384
rect 673821 381379 673887 381382
rect 675109 381379 675175 381382
rect 35758 381140 35818 381379
rect 46933 380762 46999 380765
rect 41492 380760 46999 380762
rect 41492 380704 46938 380760
rect 46994 380704 46999 380760
rect 41492 380702 46999 380704
rect 46933 380699 46999 380702
rect 675753 380626 675819 380629
rect 676438 380626 676444 380628
rect 675753 380624 676444 380626
rect 675753 380568 675758 380624
rect 675814 380568 676444 380624
rect 675753 380566 676444 380568
rect 675753 380563 675819 380566
rect 676438 380564 676444 380566
rect 676508 380564 676514 380628
rect 47117 380354 47183 380357
rect 41492 380352 47183 380354
rect 41492 380296 47122 380352
rect 47178 380296 47183 380352
rect 41492 380294 47183 380296
rect 47117 380291 47183 380294
rect 44541 379946 44607 379949
rect 41492 379944 44607 379946
rect 41492 379888 44546 379944
rect 44602 379888 44607 379944
rect 41492 379886 44607 379888
rect 44541 379883 44607 379886
rect 44909 379538 44975 379541
rect 41492 379536 44975 379538
rect 41492 379480 44914 379536
rect 44970 379480 44975 379536
rect 41492 379478 44975 379480
rect 44909 379475 44975 379478
rect 44725 379130 44791 379133
rect 41492 379128 44791 379130
rect 41492 379072 44730 379128
rect 44786 379072 44791 379128
rect 41492 379070 44791 379072
rect 44725 379067 44791 379070
rect 675753 378724 675819 378725
rect 675702 378722 675708 378724
rect 40542 378588 40602 378692
rect 675662 378662 675708 378722
rect 675772 378720 675819 378724
rect 675814 378664 675819 378720
rect 675702 378660 675708 378662
rect 675772 378660 675819 378664
rect 675753 378659 675819 378660
rect 40534 378524 40540 378588
rect 40604 378524 40610 378588
rect 41321 378586 41387 378589
rect 42333 378586 42399 378589
rect 41321 378584 42399 378586
rect 41321 378528 41326 378584
rect 41382 378528 42338 378584
rect 42394 378528 42399 378584
rect 41321 378526 42399 378528
rect 41321 378523 41387 378526
rect 42333 378523 42399 378526
rect 40726 378180 40786 378284
rect 40718 378116 40724 378180
rect 40788 378116 40794 378180
rect 652385 378178 652451 378181
rect 650164 378176 652451 378178
rect 650164 378120 652390 378176
rect 652446 378120 652451 378176
rect 650164 378118 652451 378120
rect 652385 378115 652451 378118
rect 672993 378042 673059 378045
rect 674782 378042 674788 378044
rect 672993 378040 674788 378042
rect 672993 377984 672998 378040
rect 673054 377984 674788 378040
rect 672993 377982 674788 377984
rect 672993 377979 673059 377982
rect 674782 377980 674788 377982
rect 674852 377980 674858 378044
rect 40910 377772 40970 377876
rect 40902 377708 40908 377772
rect 40972 377708 40978 377772
rect 674465 377770 674531 377773
rect 675109 377770 675175 377773
rect 674465 377768 675175 377770
rect 674465 377712 674470 377768
rect 674526 377712 675114 377768
rect 675170 377712 675175 377768
rect 674465 377710 675175 377712
rect 674465 377707 674531 377710
rect 675109 377707 675175 377710
rect 44173 377498 44239 377501
rect 41492 377496 44239 377498
rect 41492 377440 44178 377496
rect 44234 377440 44239 377496
rect 41492 377438 44239 377440
rect 44173 377435 44239 377438
rect 675753 377362 675819 377365
rect 676254 377362 676260 377364
rect 675753 377360 676260 377362
rect 675753 377304 675758 377360
rect 675814 377304 676260 377360
rect 675753 377302 676260 377304
rect 675753 377299 675819 377302
rect 676254 377300 676260 377302
rect 676324 377300 676330 377364
rect 35758 376549 35818 377060
rect 40033 376954 40099 376957
rect 41638 376954 41644 376956
rect 40033 376952 41644 376954
rect 40033 376896 40038 376952
rect 40094 376896 41644 376952
rect 40033 376894 41644 376896
rect 40033 376891 40099 376894
rect 41638 376892 41644 376894
rect 41708 376892 41714 376956
rect 675201 376954 675267 376957
rect 676070 376954 676076 376956
rect 675201 376952 676076 376954
rect 675201 376896 675206 376952
rect 675262 376896 676076 376952
rect 675201 376894 676076 376896
rect 675201 376891 675267 376894
rect 676070 376892 676076 376894
rect 676140 376892 676146 376956
rect 35758 376544 35867 376549
rect 35758 376488 35806 376544
rect 35862 376488 35867 376544
rect 35758 376486 35867 376488
rect 35801 376483 35867 376486
rect 44357 376274 44423 376277
rect 41492 376272 44423 376274
rect 41492 376216 44362 376272
rect 44418 376216 44423 376272
rect 41492 376214 44423 376216
rect 44357 376211 44423 376214
rect 62113 376274 62179 376277
rect 672625 376274 672691 376277
rect 675385 376274 675451 376277
rect 62113 376272 64492 376274
rect 62113 376216 62118 376272
rect 62174 376216 64492 376272
rect 62113 376214 64492 376216
rect 672625 376272 675451 376274
rect 672625 376216 672630 376272
rect 672686 376216 675390 376272
rect 675446 376216 675451 376272
rect 672625 376214 675451 376216
rect 62113 376211 62179 376214
rect 672625 376211 672691 376214
rect 675385 376211 675451 376214
rect 39573 375730 39639 375733
rect 40350 375730 40356 375732
rect 39573 375728 40356 375730
rect 39573 375672 39578 375728
rect 39634 375672 40356 375728
rect 39573 375670 40356 375672
rect 39573 375667 39639 375670
rect 40350 375668 40356 375670
rect 40420 375668 40426 375732
rect 674005 375458 674071 375461
rect 675385 375458 675451 375461
rect 674005 375456 675451 375458
rect 674005 375400 674010 375456
rect 674066 375400 675390 375456
rect 675446 375400 675451 375456
rect 674005 375398 675451 375400
rect 674005 375395 674071 375398
rect 675385 375395 675451 375398
rect 675661 373010 675727 373013
rect 675886 373010 675892 373012
rect 675661 373008 675892 373010
rect 675661 372952 675666 373008
rect 675722 372952 675892 373008
rect 675661 372950 675892 372952
rect 675661 372947 675727 372950
rect 675886 372948 675892 372950
rect 675956 372948 675962 373012
rect 674782 372540 674788 372604
rect 674852 372602 674858 372604
rect 675109 372602 675175 372605
rect 674852 372600 675175 372602
rect 674852 372544 675114 372600
rect 675170 372544 675175 372600
rect 674852 372542 675175 372544
rect 674852 372540 674858 372542
rect 675109 372539 675175 372542
rect 37917 371378 37983 371381
rect 41822 371378 41828 371380
rect 37917 371376 41828 371378
rect 37917 371320 37922 371376
rect 37978 371320 41828 371376
rect 37917 371318 41828 371320
rect 37917 371315 37983 371318
rect 41822 371316 41828 371318
rect 41892 371316 41898 371380
rect 40350 368596 40356 368660
rect 40420 368658 40426 368660
rect 41781 368658 41847 368661
rect 40420 368656 41847 368658
rect 40420 368600 41786 368656
rect 41842 368600 41847 368656
rect 40420 368598 41847 368600
rect 40420 368596 40426 368598
rect 41781 368595 41847 368598
rect 42425 367026 42491 367029
rect 46197 367026 46263 367029
rect 42425 367024 46263 367026
rect 42425 366968 42430 367024
rect 42486 366968 46202 367024
rect 46258 366968 46263 367024
rect 42425 366966 46263 366968
rect 42425 366963 42491 366966
rect 46197 366963 46263 366966
rect 42425 365802 42491 365805
rect 44817 365802 44883 365805
rect 42425 365800 44883 365802
rect 42425 365744 42430 365800
rect 42486 365744 44822 365800
rect 44878 365744 44883 365800
rect 42425 365742 44883 365744
rect 42425 365739 42491 365742
rect 44817 365739 44883 365742
rect 651833 364850 651899 364853
rect 650164 364848 651899 364850
rect 650164 364792 651838 364848
rect 651894 364792 651899 364848
rect 650164 364790 651899 364792
rect 651833 364787 651899 364790
rect 40902 364244 40908 364308
rect 40972 364306 40978 364308
rect 41781 364306 41847 364309
rect 40972 364304 41847 364306
rect 40972 364248 41786 364304
rect 41842 364248 41847 364304
rect 40972 364246 41847 364248
rect 40972 364244 40978 364246
rect 41781 364243 41847 364246
rect 42425 364306 42491 364309
rect 44817 364306 44883 364309
rect 42425 364304 44883 364306
rect 42425 364248 42430 364304
rect 42486 364248 44822 364304
rect 44878 364248 44883 364304
rect 42425 364246 44883 364248
rect 42425 364243 42491 364246
rect 44817 364243 44883 364246
rect 40718 363700 40724 363764
rect 40788 363762 40794 363764
rect 41781 363762 41847 363765
rect 40788 363760 41847 363762
rect 40788 363704 41786 363760
rect 41842 363704 41847 363760
rect 40788 363702 41847 363704
rect 40788 363700 40794 363702
rect 41781 363699 41847 363702
rect 62113 363354 62179 363357
rect 62113 363352 64492 363354
rect 62113 363296 62118 363352
rect 62174 363296 64492 363352
rect 62113 363294 64492 363296
rect 62113 363291 62179 363294
rect 41781 362948 41847 362949
rect 41781 362944 41828 362948
rect 41892 362946 41898 362948
rect 41781 362888 41786 362944
rect 41781 362884 41828 362888
rect 41892 362886 41938 362946
rect 41892 362884 41898 362886
rect 41781 362883 41847 362884
rect 667197 360906 667263 360909
rect 675845 360906 675911 360909
rect 667197 360904 675911 360906
rect 667197 360848 667202 360904
rect 667258 360848 675850 360904
rect 675906 360848 675911 360904
rect 667197 360846 675911 360848
rect 667197 360843 667263 360846
rect 675845 360843 675911 360846
rect 40534 360028 40540 360092
rect 40604 360090 40610 360092
rect 41781 360090 41847 360093
rect 40604 360088 41847 360090
rect 40604 360032 41786 360088
rect 41842 360032 41847 360088
rect 40604 360030 41847 360032
rect 40604 360028 40610 360030
rect 41781 360027 41847 360030
rect 659101 360090 659167 360093
rect 676029 360090 676095 360093
rect 659101 360088 676095 360090
rect 659101 360032 659106 360088
rect 659162 360032 676034 360088
rect 676090 360032 676095 360088
rect 659101 360030 676095 360032
rect 659101 360027 659167 360030
rect 676029 360027 676095 360030
rect 42149 359954 42215 359957
rect 44633 359954 44699 359957
rect 42149 359952 44699 359954
rect 42149 359896 42154 359952
rect 42210 359896 44638 359952
rect 44694 359896 44699 359952
rect 42149 359894 44699 359896
rect 42149 359891 42215 359894
rect 44633 359891 44699 359894
rect 41454 358668 41460 358732
rect 41524 358730 41530 358732
rect 41781 358730 41847 358733
rect 41524 358728 41847 358730
rect 41524 358672 41786 358728
rect 41842 358672 41847 358728
rect 41524 358670 41847 358672
rect 41524 358668 41530 358670
rect 41781 358667 41847 358670
rect 663750 358670 676292 358730
rect 663241 358594 663307 358597
rect 663750 358594 663810 358670
rect 663241 358592 663810 358594
rect 663241 358536 663246 358592
rect 663302 358536 663810 358592
rect 663241 358534 663810 358536
rect 663241 358531 663307 358534
rect 676029 358322 676095 358325
rect 676029 358320 676292 358322
rect 676029 358264 676034 358320
rect 676090 358264 676292 358320
rect 676029 358262 676292 358264
rect 676029 358259 676095 358262
rect 675845 357914 675911 357917
rect 675845 357912 676292 357914
rect 675845 357856 675850 357912
rect 675906 357856 676292 357912
rect 675845 357854 676292 357856
rect 675845 357851 675911 357854
rect 674189 357506 674255 357509
rect 674189 357504 676292 357506
rect 674189 357448 674194 357504
rect 674250 357448 676292 357504
rect 674189 357446 676292 357448
rect 674189 357443 674255 357446
rect 42425 357370 42491 357373
rect 47117 357370 47183 357373
rect 42425 357368 47183 357370
rect 42425 357312 42430 357368
rect 42486 357312 47122 357368
rect 47178 357312 47183 357368
rect 42425 357310 47183 357312
rect 42425 357307 42491 357310
rect 47117 357307 47183 357310
rect 672165 357098 672231 357101
rect 672165 357096 676292 357098
rect 672165 357040 672170 357096
rect 672226 357040 676292 357096
rect 672165 357038 676292 357040
rect 672165 357035 672231 357038
rect 44173 356690 44239 356693
rect 45185 356690 45251 356693
rect 44173 356688 45251 356690
rect 44173 356632 44178 356688
rect 44234 356632 45190 356688
rect 45246 356632 45251 356688
rect 44173 356630 45251 356632
rect 44173 356627 44239 356630
rect 45185 356627 45251 356630
rect 674649 356690 674715 356693
rect 674649 356688 676292 356690
rect 674649 356632 674654 356688
rect 674710 356632 676292 356688
rect 674649 356630 676292 356632
rect 674649 356627 674715 356630
rect 44449 356282 44515 356285
rect 45185 356282 45251 356285
rect 44449 356280 45251 356282
rect 44449 356224 44454 356280
rect 44510 356224 45190 356280
rect 45246 356224 45251 356280
rect 44449 356222 45251 356224
rect 44449 356219 44515 356222
rect 45185 356219 45251 356222
rect 672625 356282 672691 356285
rect 672625 356280 676292 356282
rect 672625 356224 672630 356280
rect 672686 356224 676292 356280
rect 672625 356222 676292 356224
rect 672625 356219 672691 356222
rect 42333 356010 42399 356013
rect 46933 356010 46999 356013
rect 42333 356008 46999 356010
rect 42333 355952 42338 356008
rect 42394 355952 46938 356008
rect 46994 355952 46999 356008
rect 42333 355950 46999 355952
rect 42333 355947 42399 355950
rect 46933 355947 46999 355950
rect 672809 355874 672875 355877
rect 672809 355872 676292 355874
rect 672809 355816 672814 355872
rect 672870 355816 676292 355872
rect 672809 355814 676292 355816
rect 672809 355811 672875 355814
rect 41873 355740 41939 355741
rect 41822 355738 41828 355740
rect 41782 355678 41828 355738
rect 41892 355736 41939 355740
rect 41934 355680 41939 355736
rect 41822 355676 41828 355678
rect 41892 355676 41939 355680
rect 41873 355675 41939 355676
rect 43069 355602 43135 355605
rect 44633 355602 44699 355605
rect 43069 355600 44699 355602
rect 43069 355544 43074 355600
rect 43130 355544 44638 355600
rect 44694 355544 44699 355600
rect 43069 355542 44699 355544
rect 43069 355539 43135 355542
rect 44633 355539 44699 355542
rect 673177 355466 673243 355469
rect 673177 355464 676292 355466
rect 673177 355408 673182 355464
rect 673238 355408 676292 355464
rect 673177 355406 676292 355408
rect 673177 355403 673243 355406
rect 43805 355330 43871 355333
rect 44817 355330 44883 355333
rect 43805 355328 44883 355330
rect 43805 355272 43810 355328
rect 43866 355272 44822 355328
rect 44878 355272 44883 355328
rect 43805 355270 44883 355272
rect 43805 355267 43871 355270
rect 44817 355267 44883 355270
rect 673361 355058 673427 355061
rect 673361 355056 676292 355058
rect 673361 355000 673366 355056
rect 673422 355000 676292 355056
rect 673361 354998 676292 355000
rect 673361 354995 673427 354998
rect 674649 354650 674715 354653
rect 674649 354648 676292 354650
rect 674649 354592 674654 354648
rect 674710 354592 676292 354648
rect 674649 354590 676292 354592
rect 674649 354587 674715 354590
rect 675334 354180 675340 354244
rect 675404 354242 675410 354244
rect 675404 354182 676292 354242
rect 675404 354180 675410 354182
rect 675702 353772 675708 353836
rect 675772 353834 675778 353836
rect 675772 353774 676292 353834
rect 675772 353772 675778 353774
rect 43253 353698 43319 353701
rect 45139 353698 45205 353701
rect 43253 353696 45205 353698
rect 43253 353640 43258 353696
rect 43314 353640 45144 353696
rect 45200 353640 45205 353696
rect 43253 353638 45205 353640
rect 43253 353635 43319 353638
rect 45139 353635 45205 353638
rect 673361 353426 673427 353429
rect 673361 353424 676292 353426
rect 673361 353368 673366 353424
rect 673422 353368 676292 353424
rect 673361 353366 676292 353368
rect 673361 353363 673427 353366
rect 676029 353018 676095 353021
rect 676029 353016 676292 353018
rect 676029 352960 676034 353016
rect 676090 352960 676292 353016
rect 676029 352958 676292 352960
rect 676029 352955 676095 352958
rect 674465 352610 674531 352613
rect 674465 352608 676292 352610
rect 674465 352552 674470 352608
rect 674526 352552 676292 352608
rect 674465 352550 676292 352552
rect 674465 352547 674531 352550
rect 674281 352202 674347 352205
rect 674281 352200 676292 352202
rect 674281 352144 674286 352200
rect 674342 352144 676292 352200
rect 674281 352142 676292 352144
rect 674281 352139 674347 352142
rect 675886 351868 675892 351932
rect 675956 351930 675962 351932
rect 675956 351870 676230 351930
rect 675956 351868 675962 351870
rect 676170 351794 676230 351870
rect 676170 351734 676292 351794
rect 652385 351658 652451 351661
rect 650164 351656 652451 351658
rect 650164 351600 652390 351656
rect 652446 351600 652451 351656
rect 650164 351598 652451 351600
rect 652385 351595 652451 351598
rect 672809 351386 672875 351389
rect 672809 351384 676292 351386
rect 672809 351328 672814 351384
rect 672870 351328 676292 351384
rect 672809 351326 676292 351328
rect 672809 351323 672875 351326
rect 28533 351250 28599 351253
rect 50521 351250 50587 351253
rect 28533 351248 50587 351250
rect 28533 351192 28538 351248
rect 28594 351192 50526 351248
rect 50582 351192 50587 351248
rect 28533 351190 50587 351192
rect 28533 351187 28599 351190
rect 50521 351187 50587 351190
rect 675886 350916 675892 350980
rect 675956 350978 675962 350980
rect 675956 350918 676292 350978
rect 675956 350916 675962 350918
rect 673729 350570 673795 350573
rect 673729 350568 676292 350570
rect 673729 350512 673734 350568
rect 673790 350512 676292 350568
rect 673729 350510 676292 350512
rect 673729 350507 673795 350510
rect 62113 350298 62179 350301
rect 62113 350296 64492 350298
rect 62113 350240 62118 350296
rect 62174 350240 64492 350296
rect 62113 350238 64492 350240
rect 62113 350235 62179 350238
rect 675886 350100 675892 350164
rect 675956 350162 675962 350164
rect 675956 350102 676292 350162
rect 675956 350100 675962 350102
rect 674097 349754 674163 349757
rect 674097 349752 676292 349754
rect 674097 349696 674102 349752
rect 674158 349696 676292 349752
rect 674097 349694 676292 349696
rect 674097 349691 674163 349694
rect 673545 349482 673611 349485
rect 673545 349480 676230 349482
rect 673545 349424 673550 349480
rect 673606 349424 676230 349480
rect 673545 349422 676230 349424
rect 673545 349419 673611 349422
rect 676170 349346 676230 349422
rect 676170 349286 676292 349346
rect 675150 349148 675156 349212
rect 675220 349210 675226 349212
rect 675937 349210 676003 349213
rect 675220 349208 676003 349210
rect 675220 349152 675942 349208
rect 675998 349152 676003 349208
rect 675220 349150 676003 349152
rect 675220 349148 675226 349150
rect 675937 349147 676003 349150
rect 672993 348938 673059 348941
rect 672993 348936 676292 348938
rect 672993 348880 672998 348936
rect 673054 348880 676292 348936
rect 672993 348878 676292 348880
rect 672993 348875 673059 348878
rect 673913 348530 673979 348533
rect 673913 348528 676292 348530
rect 673913 348472 673918 348528
rect 673974 348472 676292 348528
rect 673913 348470 676292 348472
rect 673913 348467 673979 348470
rect 671797 347714 671863 347717
rect 683070 347714 683130 348092
rect 671797 347712 683130 347714
rect 671797 347656 671802 347712
rect 671858 347684 683130 347712
rect 671858 347656 683100 347684
rect 671797 347654 683100 347656
rect 671797 347651 671863 347654
rect 670601 347306 670667 347309
rect 670601 347304 676292 347306
rect 670601 347248 670606 347304
rect 670662 347248 676292 347304
rect 670601 347246 676292 347248
rect 670601 347243 670667 347246
rect 62757 345674 62823 345677
rect 45510 345672 62823 345674
rect 45510 345616 62762 345672
rect 62818 345616 62823 345672
rect 45510 345614 62823 345616
rect 40217 345538 40283 345541
rect 45510 345538 45570 345614
rect 62757 345611 62823 345614
rect 40217 345536 45570 345538
rect 40217 345480 40222 345536
rect 40278 345480 45570 345536
rect 40217 345478 45570 345480
rect 40217 345475 40283 345478
rect 41462 344314 41522 344556
rect 54477 344314 54543 344317
rect 41462 344312 54543 344314
rect 41462 344256 54482 344312
rect 54538 344256 54543 344312
rect 41462 344254 54543 344256
rect 54477 344251 54543 344254
rect 35758 343909 35818 344148
rect 28533 343906 28599 343909
rect 28533 343904 28642 343906
rect 28533 343848 28538 343904
rect 28594 343848 28642 343904
rect 28533 343843 28642 343848
rect 35758 343904 35867 343909
rect 35758 343848 35806 343904
rect 35862 343848 35867 343904
rect 35758 343846 35867 343848
rect 35801 343843 35867 343846
rect 28582 343740 28642 343843
rect 45461 343362 45527 343365
rect 41492 343360 45527 343362
rect 41492 343304 45466 343360
rect 45522 343304 45527 343360
rect 41492 343302 45527 343304
rect 45461 343299 45527 343302
rect 44214 342954 44220 342956
rect 41492 342894 44220 342954
rect 44214 342892 44220 342894
rect 44284 342892 44290 342956
rect 44817 342546 44883 342549
rect 41492 342544 44883 342546
rect 41492 342488 44822 342544
rect 44878 342488 44883 342544
rect 41492 342486 44883 342488
rect 44817 342483 44883 342486
rect 44398 342138 44404 342140
rect 41492 342078 44404 342138
rect 44398 342076 44404 342078
rect 44468 342076 44474 342140
rect 45829 341730 45895 341733
rect 41492 341728 45895 341730
rect 41492 341672 45834 341728
rect 45890 341672 45895 341728
rect 41492 341670 45895 341672
rect 45829 341667 45895 341670
rect 45461 341322 45527 341325
rect 41492 341320 45527 341322
rect 41492 341264 45466 341320
rect 45522 341264 45527 341320
rect 41492 341262 45527 341264
rect 45461 341259 45527 341262
rect 45645 340914 45711 340917
rect 41492 340912 45711 340914
rect 41492 340856 45650 340912
rect 45706 340856 45711 340912
rect 41492 340854 45711 340856
rect 45645 340851 45711 340854
rect 673361 340778 673427 340781
rect 675109 340778 675175 340781
rect 673361 340776 675175 340778
rect 673361 340720 673366 340776
rect 673422 340720 675114 340776
rect 675170 340720 675175 340776
rect 673361 340718 675175 340720
rect 673361 340715 673427 340718
rect 675109 340715 675175 340718
rect 43662 340506 43668 340508
rect 41492 340446 43668 340506
rect 43662 340444 43668 340446
rect 43732 340444 43738 340508
rect 675753 340234 675819 340237
rect 676622 340234 676628 340236
rect 675753 340232 676628 340234
rect 675753 340176 675758 340232
rect 675814 340176 676628 340232
rect 675753 340174 676628 340176
rect 675753 340171 675819 340174
rect 676622 340172 676628 340174
rect 676692 340172 676698 340236
rect 45737 340098 45803 340101
rect 41492 340096 45803 340098
rect 41492 340040 45742 340096
rect 45798 340040 45803 340096
rect 41492 340038 45803 340040
rect 45737 340035 45803 340038
rect 35801 339826 35867 339829
rect 35758 339824 35867 339826
rect 35758 339768 35806 339824
rect 35862 339768 35867 339824
rect 35758 339763 35867 339768
rect 35758 339660 35818 339763
rect 675661 339418 675727 339421
rect 675886 339418 675892 339420
rect 675661 339416 675892 339418
rect 675661 339360 675666 339416
rect 675722 339360 675892 339416
rect 675661 339358 675892 339360
rect 675661 339355 675727 339358
rect 675886 339356 675892 339358
rect 675956 339356 675962 339420
rect 35206 339013 35266 339252
rect 35157 339008 35266 339013
rect 35157 338952 35162 339008
rect 35218 338952 35266 339008
rect 35157 338950 35266 338952
rect 35157 338947 35223 338950
rect 40726 338604 40786 338844
rect 40718 338540 40724 338604
rect 40788 338540 40794 338604
rect 33734 338197 33794 338436
rect 652017 338330 652083 338333
rect 650164 338328 652083 338330
rect 650164 338272 652022 338328
rect 652078 338272 652083 338328
rect 650164 338270 652083 338272
rect 652017 338267 652083 338270
rect 33734 338192 33843 338197
rect 33734 338136 33782 338192
rect 33838 338136 33843 338192
rect 33734 338134 33843 338136
rect 33777 338131 33843 338134
rect 45921 338058 45987 338061
rect 41492 338056 45987 338058
rect 41492 338000 45926 338056
rect 45982 338000 45987 338056
rect 41492 337998 45987 338000
rect 45921 337995 45987 337998
rect 675569 337788 675635 337789
rect 675518 337786 675524 337788
rect 675478 337726 675524 337786
rect 675588 337784 675635 337788
rect 675630 337728 675635 337784
rect 675518 337724 675524 337726
rect 675588 337724 675635 337728
rect 675569 337723 675635 337724
rect 42926 337650 42932 337652
rect 41492 337590 42932 337650
rect 42926 337588 42932 337590
rect 42996 337588 43002 337652
rect 43294 337242 43300 337244
rect 41492 337182 43300 337242
rect 43294 337180 43300 337182
rect 43364 337180 43370 337244
rect 62113 337242 62179 337245
rect 672809 337242 672875 337245
rect 675109 337242 675175 337245
rect 62113 337240 64492 337242
rect 62113 337184 62118 337240
rect 62174 337184 64492 337240
rect 62113 337182 64492 337184
rect 672809 337240 675175 337242
rect 672809 337184 672814 337240
rect 672870 337184 675114 337240
rect 675170 337184 675175 337240
rect 672809 337182 675175 337184
rect 62113 337179 62179 337182
rect 672809 337179 672875 337182
rect 675109 337179 675175 337182
rect 40534 336908 40540 336972
rect 40604 336908 40610 336972
rect 40542 336804 40602 336908
rect 674281 336698 674347 336701
rect 674782 336698 674788 336700
rect 674281 336696 674788 336698
rect 674281 336640 674286 336696
rect 674342 336640 674788 336696
rect 674281 336638 674788 336640
rect 674281 336635 674347 336638
rect 674782 336636 674788 336638
rect 674852 336636 674858 336700
rect 37549 336562 37615 336565
rect 41822 336562 41828 336564
rect 37549 336560 41828 336562
rect 37549 336504 37554 336560
rect 37610 336504 41828 336560
rect 37549 336502 41828 336504
rect 37549 336499 37615 336502
rect 41822 336500 41828 336502
rect 41892 336500 41898 336564
rect 41462 336154 41522 336396
rect 43110 336154 43116 336156
rect 41462 336094 43116 336154
rect 43110 336092 43116 336094
rect 43180 336092 43186 336156
rect 41278 335746 41338 335988
rect 674097 335882 674163 335885
rect 675477 335882 675543 335885
rect 674097 335880 675543 335882
rect 674097 335824 674102 335880
rect 674158 335824 675482 335880
rect 675538 335824 675543 335880
rect 674097 335822 675543 335824
rect 674097 335819 674163 335822
rect 675477 335819 675543 335822
rect 43846 335746 43852 335748
rect 41278 335686 43852 335746
rect 43846 335684 43852 335686
rect 43916 335684 43922 335748
rect 41462 335474 41522 335580
rect 42742 335474 42748 335476
rect 41462 335414 42748 335474
rect 42742 335412 42748 335414
rect 42812 335412 42818 335476
rect 675293 335338 675359 335341
rect 676438 335338 676444 335340
rect 675293 335336 676444 335338
rect 675293 335280 675298 335336
rect 675354 335280 676444 335336
rect 675293 335278 676444 335280
rect 675293 335275 675359 335278
rect 676438 335276 676444 335278
rect 676508 335276 676514 335340
rect 41462 334930 41522 335172
rect 41462 334870 44466 334930
rect 41462 334658 41522 334764
rect 44406 334661 44466 334870
rect 42793 334660 42859 334661
rect 43161 334660 43227 334661
rect 42742 334658 42748 334660
rect 41462 334598 42258 334658
rect 42702 334598 42748 334658
rect 42812 334656 42859 334660
rect 43110 334658 43116 334660
rect 42854 334600 42859 334656
rect 42198 334386 42258 334598
rect 42742 334596 42748 334598
rect 42812 334596 42859 334600
rect 43070 334598 43116 334658
rect 43180 334656 43227 334660
rect 43222 334600 43227 334656
rect 43110 334596 43116 334598
rect 43180 334596 43227 334600
rect 43846 334596 43852 334660
rect 43916 334658 43922 334660
rect 44173 334658 44239 334661
rect 43916 334656 44239 334658
rect 43916 334600 44178 334656
rect 44234 334600 44239 334656
rect 43916 334598 44239 334600
rect 43916 334596 43922 334598
rect 42793 334595 42859 334596
rect 43161 334595 43227 334596
rect 44173 334595 44239 334598
rect 44357 334656 44466 334661
rect 44357 334600 44362 334656
rect 44418 334600 44466 334656
rect 44357 334598 44466 334600
rect 44357 334595 44423 334598
rect 42977 334386 43043 334389
rect 42198 334384 43043 334386
rect 41462 334114 41522 334356
rect 42198 334328 42982 334384
rect 43038 334328 43043 334384
rect 42198 334326 43043 334328
rect 42977 334323 43043 334326
rect 48957 334114 49023 334117
rect 41462 334112 49023 334114
rect 41462 334056 48962 334112
rect 49018 334056 49023 334112
rect 41462 334054 49023 334056
rect 48957 334051 49023 334054
rect 674465 333978 674531 333981
rect 675109 333978 675175 333981
rect 674465 333976 675175 333978
rect 27662 333540 27722 333948
rect 40910 333708 40970 333948
rect 674465 333920 674470 333976
rect 674526 333920 675114 333976
rect 675170 333920 675175 333976
rect 674465 333918 675175 333920
rect 674465 333915 674531 333918
rect 675109 333915 675175 333918
rect 40902 333644 40908 333708
rect 40972 333644 40978 333708
rect 47577 333162 47643 333165
rect 41492 333160 47643 333162
rect 41492 333104 47582 333160
rect 47638 333104 47643 333160
rect 41492 333102 47643 333104
rect 47577 333099 47643 333102
rect 673545 332754 673611 332757
rect 675109 332754 675175 332757
rect 673545 332752 675175 332754
rect 673545 332696 673550 332752
rect 673606 332696 675114 332752
rect 675170 332696 675175 332752
rect 673545 332694 675175 332696
rect 673545 332691 673611 332694
rect 675109 332691 675175 332694
rect 675753 332346 675819 332349
rect 676254 332346 676260 332348
rect 675753 332344 676260 332346
rect 675753 332288 675758 332344
rect 675814 332288 676260 332344
rect 675753 332286 676260 332288
rect 675753 332283 675819 332286
rect 676254 332284 676260 332286
rect 676324 332284 676330 332348
rect 672993 331530 673059 331533
rect 675109 331530 675175 331533
rect 672993 331528 675175 331530
rect 672993 331472 672998 331528
rect 673054 331472 675114 331528
rect 675170 331472 675175 331528
rect 672993 331470 675175 331472
rect 672993 331467 673059 331470
rect 675109 331467 675175 331470
rect 673729 331122 673795 331125
rect 675109 331122 675175 331125
rect 673729 331120 675175 331122
rect 673729 331064 673734 331120
rect 673790 331064 675114 331120
rect 675170 331064 675175 331120
rect 673729 331062 675175 331064
rect 673729 331059 673795 331062
rect 675109 331059 675175 331062
rect 35157 329082 35223 329085
rect 42006 329082 42012 329084
rect 35157 329080 42012 329082
rect 35157 329024 35162 329080
rect 35218 329024 42012 329080
rect 35157 329022 42012 329024
rect 35157 329019 35223 329022
rect 42006 329020 42012 329022
rect 42076 329020 42082 329084
rect 675753 328402 675819 328405
rect 676070 328402 676076 328404
rect 675753 328400 676076 328402
rect 675753 328344 675758 328400
rect 675814 328344 676076 328400
rect 675753 328342 676076 328344
rect 675753 328339 675819 328342
rect 676070 328340 676076 328342
rect 676140 328340 676146 328404
rect 33777 327722 33843 327725
rect 41638 327722 41644 327724
rect 33777 327720 41644 327722
rect 33777 327664 33782 327720
rect 33838 327664 41644 327720
rect 33777 327662 41644 327664
rect 33777 327659 33843 327662
rect 41638 327660 41644 327662
rect 41708 327660 41714 327724
rect 674782 326844 674788 326908
rect 674852 326906 674858 326908
rect 675385 326906 675451 326909
rect 674852 326904 675451 326906
rect 674852 326848 675390 326904
rect 675446 326848 675451 326904
rect 674852 326846 675451 326848
rect 674852 326844 674858 326846
rect 675385 326843 675451 326846
rect 671797 325682 671863 325685
rect 675109 325682 675175 325685
rect 671797 325680 675175 325682
rect 671797 325624 671802 325680
rect 671858 325624 675114 325680
rect 675170 325624 675175 325680
rect 671797 325622 675175 325624
rect 671797 325619 671863 325622
rect 675109 325619 675175 325622
rect 40902 325348 40908 325412
rect 40972 325410 40978 325412
rect 41781 325410 41847 325413
rect 40972 325408 41847 325410
rect 40972 325352 41786 325408
rect 41842 325352 41847 325408
rect 40972 325350 41847 325352
rect 40972 325348 40978 325350
rect 41781 325347 41847 325350
rect 651465 325002 651531 325005
rect 650164 325000 651531 325002
rect 650164 324944 651470 325000
rect 651526 324944 651531 325000
rect 650164 324942 651531 324944
rect 651465 324939 651531 324942
rect 41873 324732 41939 324733
rect 41822 324730 41828 324732
rect 41782 324670 41828 324730
rect 41892 324728 41939 324732
rect 41934 324672 41939 324728
rect 41822 324668 41828 324670
rect 41892 324668 41939 324672
rect 41873 324667 41939 324668
rect 42241 324322 42307 324325
rect 45921 324322 45987 324325
rect 42241 324320 45987 324322
rect 42241 324264 42246 324320
rect 42302 324264 45926 324320
rect 45982 324264 45987 324320
rect 42241 324262 45987 324264
rect 42241 324259 42307 324262
rect 45921 324259 45987 324262
rect 42241 323642 42307 323645
rect 42977 323642 43043 323645
rect 42241 323640 43043 323642
rect 42241 323584 42246 323640
rect 42302 323584 42982 323640
rect 43038 323584 43043 323640
rect 42241 323582 43043 323584
rect 42241 323579 42307 323582
rect 42977 323579 43043 323582
rect 43621 322962 43687 322965
rect 64462 322962 64522 324156
rect 43621 322960 64522 322962
rect 43621 322904 43626 322960
rect 43682 322904 64522 322960
rect 43621 322902 64522 322904
rect 43621 322899 43687 322902
rect 42057 322826 42123 322829
rect 43161 322826 43227 322829
rect 42057 322824 43227 322826
rect 42057 322768 42062 322824
rect 42118 322768 43166 322824
rect 43222 322768 43227 322824
rect 42057 322766 43227 322768
rect 42057 322763 42123 322766
rect 43161 322763 43227 322766
rect 42425 321466 42491 321469
rect 53097 321466 53163 321469
rect 42425 321464 53163 321466
rect 42425 321408 42430 321464
rect 42486 321408 53102 321464
rect 53158 321408 53163 321464
rect 42425 321406 53163 321408
rect 42425 321403 42491 321406
rect 53097 321403 53163 321406
rect 42425 321194 42491 321197
rect 44173 321194 44239 321197
rect 42425 321192 44239 321194
rect 42425 321136 42430 321192
rect 42486 321136 44178 321192
rect 44234 321136 44239 321192
rect 42425 321134 44239 321136
rect 42425 321131 42491 321134
rect 44173 321131 44239 321134
rect 42425 320106 42491 320109
rect 44357 320106 44423 320109
rect 42425 320104 44423 320106
rect 42425 320048 42430 320104
rect 42486 320048 44362 320104
rect 44418 320048 44423 320104
rect 42425 320046 44423 320048
rect 42425 320043 42491 320046
rect 44357 320043 44423 320046
rect 41781 319972 41847 319973
rect 41781 319968 41828 319972
rect 41892 319970 41898 319972
rect 41781 319912 41786 319968
rect 41781 319908 41828 319912
rect 41892 319910 41938 319970
rect 41892 319908 41898 319910
rect 41781 319907 41847 319908
rect 40534 316780 40540 316844
rect 40604 316842 40610 316844
rect 41781 316842 41847 316845
rect 40604 316840 41847 316842
rect 40604 316784 41786 316840
rect 41842 316784 41847 316840
rect 40604 316782 41847 316784
rect 40604 316780 40610 316782
rect 41781 316779 41847 316782
rect 42149 316026 42215 316029
rect 43110 316026 43116 316028
rect 42149 316024 43116 316026
rect 42149 315968 42154 316024
rect 42210 315968 43116 316024
rect 42149 315966 43116 315968
rect 42149 315963 42215 315966
rect 43110 315964 43116 315966
rect 43180 315964 43186 316028
rect 41454 315556 41460 315620
rect 41524 315618 41530 315620
rect 41781 315618 41847 315621
rect 41524 315616 41847 315618
rect 41524 315560 41786 315616
rect 41842 315560 41847 315616
rect 41524 315558 41847 315560
rect 41524 315556 41530 315558
rect 41781 315555 41847 315558
rect 665817 315482 665883 315485
rect 676029 315482 676095 315485
rect 665817 315480 676095 315482
rect 665817 315424 665822 315480
rect 665878 315424 676034 315480
rect 676090 315424 676095 315480
rect 665817 315422 676095 315424
rect 665817 315419 665883 315422
rect 676029 315419 676095 315422
rect 42149 313714 42215 313717
rect 45737 313714 45803 313717
rect 42149 313712 45803 313714
rect 42149 313656 42154 313712
rect 42210 313656 45742 313712
rect 45798 313656 45803 313712
rect 42149 313654 45803 313656
rect 42149 313651 42215 313654
rect 45737 313651 45803 313654
rect 663750 313654 676292 313714
rect 661677 313578 661743 313581
rect 663750 313578 663810 313654
rect 661677 313576 663810 313578
rect 661677 313520 661682 313576
rect 661738 313520 663810 313576
rect 661677 313518 663810 313520
rect 661677 313515 661743 313518
rect 676029 313306 676095 313309
rect 676029 313304 676292 313306
rect 676029 313248 676034 313304
rect 676090 313248 676292 313304
rect 676029 313246 676292 313248
rect 676029 313243 676095 313246
rect 674649 313034 674715 313037
rect 674649 313032 675034 313034
rect 674649 312976 674654 313032
rect 674710 312976 675034 313032
rect 674649 312974 675034 312976
rect 674649 312971 674715 312974
rect 674974 312898 675034 312974
rect 674974 312838 676292 312898
rect 42425 312762 42491 312765
rect 42926 312762 42932 312764
rect 42425 312760 42932 312762
rect 42425 312704 42430 312760
rect 42486 312704 42932 312760
rect 42425 312702 42932 312704
rect 42425 312699 42491 312702
rect 42926 312700 42932 312702
rect 42996 312700 43002 312764
rect 672809 312762 672875 312765
rect 674833 312762 674899 312765
rect 672809 312760 674899 312762
rect 672809 312704 672814 312760
rect 672870 312704 674838 312760
rect 674894 312704 674899 312760
rect 672809 312702 674899 312704
rect 672809 312699 672875 312702
rect 674833 312699 674899 312702
rect 41965 312628 42031 312629
rect 41965 312624 42012 312628
rect 42076 312626 42082 312628
rect 41965 312568 41970 312624
rect 41965 312564 42012 312568
rect 42076 312566 42122 312626
rect 42076 312564 42082 312566
rect 41965 312563 42031 312564
rect 672165 312490 672231 312493
rect 672165 312488 676292 312490
rect 672165 312432 672170 312488
rect 672226 312432 676292 312488
rect 672165 312430 676292 312432
rect 672165 312427 672231 312430
rect 674833 312082 674899 312085
rect 674833 312080 676292 312082
rect 674833 312024 674838 312080
rect 674894 312024 676292 312080
rect 674833 312022 676292 312024
rect 674833 312019 674899 312022
rect 668577 311946 668643 311949
rect 674649 311946 674715 311949
rect 668577 311944 674715 311946
rect 668577 311888 668582 311944
rect 668638 311888 674654 311944
rect 674710 311888 674715 311944
rect 668577 311886 674715 311888
rect 668577 311883 668643 311886
rect 674649 311883 674715 311886
rect 651465 311810 651531 311813
rect 650164 311808 651531 311810
rect 650164 311752 651470 311808
rect 651526 311752 651531 311808
rect 650164 311750 651531 311752
rect 651465 311747 651531 311750
rect 672625 311674 672691 311677
rect 672625 311672 676292 311674
rect 672625 311616 672630 311672
rect 672686 311616 676292 311672
rect 672625 311614 676292 311616
rect 672625 311611 672691 311614
rect 44541 311404 44607 311405
rect 44541 311400 44588 311404
rect 44652 311402 44658 311404
rect 44541 311344 44546 311400
rect 44541 311340 44588 311344
rect 44652 311342 44698 311402
rect 44652 311340 44658 311342
rect 44541 311339 44607 311340
rect 673085 311266 673151 311269
rect 673085 311264 676292 311266
rect 673085 311208 673090 311264
rect 673146 311208 676292 311264
rect 673085 311206 676292 311208
rect 673085 311203 673151 311206
rect 44357 311132 44423 311133
rect 44357 311128 44404 311132
rect 44468 311130 44474 311132
rect 62113 311130 62179 311133
rect 44357 311072 44362 311128
rect 44357 311068 44404 311072
rect 44468 311070 44514 311130
rect 62113 311128 64492 311130
rect 62113 311072 62118 311128
rect 62174 311072 64492 311128
rect 62113 311070 64492 311072
rect 44468 311068 44474 311070
rect 44357 311067 44423 311068
rect 62113 311067 62179 311070
rect 673269 310858 673335 310861
rect 673269 310856 676292 310858
rect 673269 310800 673274 310856
rect 673330 310800 676292 310856
rect 673269 310798 676292 310800
rect 673269 310795 673335 310798
rect 674649 310450 674715 310453
rect 674649 310448 676292 310450
rect 674649 310392 674654 310448
rect 674710 310392 676292 310448
rect 674649 310390 676292 310392
rect 674649 310387 674715 310390
rect 674465 310042 674531 310045
rect 674465 310040 676292 310042
rect 674465 309984 674470 310040
rect 674526 309984 676292 310040
rect 674465 309982 676292 309984
rect 674465 309979 674531 309982
rect 674189 309634 674255 309637
rect 674189 309632 676292 309634
rect 674189 309576 674194 309632
rect 674250 309576 676292 309632
rect 674189 309574 676292 309576
rect 674189 309571 674255 309574
rect 675109 309226 675175 309229
rect 675109 309224 676292 309226
rect 675109 309168 675114 309224
rect 675170 309168 676292 309224
rect 675109 309166 676292 309168
rect 675109 309163 675175 309166
rect 675702 308756 675708 308820
rect 675772 308818 675778 308820
rect 675772 308758 676292 308818
rect 675772 308756 675778 308758
rect 676029 308410 676095 308413
rect 676029 308408 676292 308410
rect 676029 308352 676034 308408
rect 676090 308352 676292 308408
rect 676029 308350 676292 308352
rect 676029 308347 676095 308350
rect 675385 308002 675451 308005
rect 675385 308000 676292 308002
rect 675385 307944 675390 308000
rect 675446 307944 676292 308000
rect 675385 307942 676292 307944
rect 675385 307939 675451 307942
rect 680997 307594 681063 307597
rect 680997 307592 681076 307594
rect 680997 307536 681002 307592
rect 681058 307536 681076 307592
rect 680997 307534 681076 307536
rect 680997 307531 681063 307534
rect 678237 307186 678303 307189
rect 678237 307184 678316 307186
rect 678237 307128 678242 307184
rect 678298 307128 678316 307184
rect 678237 307126 678316 307128
rect 678237 307123 678303 307126
rect 675886 306716 675892 306780
rect 675956 306778 675962 306780
rect 675956 306718 676292 306778
rect 675956 306716 675962 306718
rect 678973 306370 679039 306373
rect 678973 306368 679052 306370
rect 678973 306312 678978 306368
rect 679034 306312 679052 306368
rect 678973 306310 679052 306312
rect 678973 306307 679039 306310
rect 675886 305900 675892 305964
rect 675956 305962 675962 305964
rect 675956 305902 676292 305962
rect 675956 305900 675962 305902
rect 673729 305554 673795 305557
rect 673729 305552 676292 305554
rect 673729 305496 673734 305552
rect 673790 305496 676292 305552
rect 673729 305494 676292 305496
rect 673729 305491 673795 305494
rect 676024 305084 676030 305148
rect 676094 305146 676100 305148
rect 676094 305086 676292 305146
rect 676094 305084 676100 305086
rect 673545 304738 673611 304741
rect 673545 304736 676292 304738
rect 673545 304680 673550 304736
rect 673606 304680 676292 304736
rect 673545 304678 676292 304680
rect 673545 304675 673611 304678
rect 672625 304330 672691 304333
rect 672625 304328 676292 304330
rect 672625 304272 672630 304328
rect 672686 304272 676292 304328
rect 672625 304270 676292 304272
rect 672625 304267 672691 304270
rect 674373 303922 674439 303925
rect 674373 303920 676292 303922
rect 674373 303864 674378 303920
rect 674434 303864 676292 303920
rect 674373 303862 676292 303864
rect 674373 303859 674439 303862
rect 673269 303514 673335 303517
rect 673269 303512 676292 303514
rect 673269 303456 673274 303512
rect 673330 303456 676292 303512
rect 673269 303454 676292 303456
rect 673269 303451 673335 303454
rect 41781 303106 41847 303109
rect 50337 303106 50403 303109
rect 41781 303104 50403 303106
rect 41781 303048 41786 303104
rect 41842 303048 50342 303104
rect 50398 303048 50403 303104
rect 41781 303046 50403 303048
rect 41781 303043 41847 303046
rect 50337 303043 50403 303046
rect 683070 302701 683130 303076
rect 683021 302696 683130 302701
rect 683021 302640 683026 302696
rect 683082 302668 683130 302696
rect 683082 302640 683100 302668
rect 683021 302638 683100 302640
rect 683021 302635 683087 302638
rect 669221 302290 669287 302293
rect 669221 302288 676292 302290
rect 669221 302232 669226 302288
rect 669282 302232 676292 302288
rect 669221 302230 676292 302232
rect 669221 302227 669287 302230
rect 51901 301338 51967 301341
rect 41492 301336 51967 301338
rect 41492 301280 51906 301336
rect 51962 301280 51967 301336
rect 41492 301278 51967 301280
rect 51901 301275 51967 301278
rect 41781 300930 41847 300933
rect 41492 300928 41847 300930
rect 41492 300872 41786 300928
rect 41842 300872 41847 300928
rect 41492 300870 41847 300872
rect 41781 300867 41847 300870
rect 47761 300522 47827 300525
rect 41492 300520 47827 300522
rect 41492 300464 47766 300520
rect 47822 300464 47827 300520
rect 41492 300462 47827 300464
rect 47761 300459 47827 300462
rect 44357 300114 44423 300117
rect 41492 300112 44423 300114
rect 41492 300056 44362 300112
rect 44418 300056 44423 300112
rect 41492 300054 44423 300056
rect 44357 300051 44423 300054
rect 44173 299706 44239 299709
rect 41492 299704 44239 299706
rect 41492 299648 44178 299704
rect 44234 299648 44239 299704
rect 41492 299646 44239 299648
rect 44173 299643 44239 299646
rect 675702 299372 675708 299436
rect 675772 299434 675778 299436
rect 683021 299434 683087 299437
rect 675772 299432 683087 299434
rect 675772 299376 683026 299432
rect 683082 299376 683087 299432
rect 675772 299374 683087 299376
rect 675772 299372 675778 299374
rect 683021 299371 683087 299374
rect 44541 299298 44607 299301
rect 41492 299296 44607 299298
rect 41492 299240 44546 299296
rect 44602 299240 44607 299296
rect 41492 299238 44607 299240
rect 44541 299235 44607 299238
rect 45185 298890 45251 298893
rect 41492 298888 45251 298890
rect 41492 298832 45190 298888
rect 45246 298832 45251 298888
rect 41492 298830 45251 298832
rect 45185 298827 45251 298830
rect 45461 298482 45527 298485
rect 652201 298482 652267 298485
rect 41492 298480 45527 298482
rect 41492 298424 45466 298480
rect 45522 298424 45527 298480
rect 41492 298422 45527 298424
rect 650164 298480 652267 298482
rect 650164 298424 652206 298480
rect 652262 298424 652267 298480
rect 650164 298422 652267 298424
rect 45461 298419 45527 298422
rect 652201 298419 652267 298422
rect 62113 298210 62179 298213
rect 62113 298208 64492 298210
rect 62113 298152 62118 298208
rect 62174 298152 64492 298208
rect 62113 298150 64492 298152
rect 62113 298147 62179 298150
rect 44357 298074 44423 298077
rect 41492 298072 44423 298074
rect 41492 298016 44362 298072
rect 44418 298016 44423 298072
rect 41492 298014 44423 298016
rect 44357 298011 44423 298014
rect 43662 297666 43668 297668
rect 41492 297606 43668 297666
rect 43662 297604 43668 297606
rect 43732 297604 43738 297668
rect 675518 297604 675524 297668
rect 675588 297666 675594 297668
rect 675937 297666 676003 297669
rect 675588 297664 676003 297666
rect 675588 297608 675942 297664
rect 675998 297608 676003 297664
rect 675588 297606 676003 297608
rect 675588 297604 675594 297606
rect 675937 297603 676003 297606
rect 675886 297332 675892 297396
rect 675956 297394 675962 297396
rect 678237 297394 678303 297397
rect 675956 297392 678303 297394
rect 675956 297336 678242 297392
rect 678298 297336 678303 297392
rect 675956 297334 678303 297336
rect 675956 297332 675962 297334
rect 678237 297331 678303 297334
rect 42793 297258 42859 297261
rect 41492 297256 42859 297258
rect 41492 297200 42798 297256
rect 42854 297200 42859 297256
rect 41492 297198 42859 297200
rect 42793 297195 42859 297198
rect 674833 297122 674899 297125
rect 676213 297122 676279 297125
rect 674833 297120 676279 297122
rect 674833 297064 674838 297120
rect 674894 297064 676218 297120
rect 676274 297064 676279 297120
rect 674833 297062 676279 297064
rect 674833 297059 674899 297062
rect 676213 297059 676279 297062
rect 41781 296850 41847 296853
rect 41492 296848 41847 296850
rect 41492 296792 41786 296848
rect 41842 296792 41847 296848
rect 41492 296790 41847 296792
rect 41781 296787 41847 296790
rect 675385 296716 675451 296717
rect 675334 296652 675340 296716
rect 675404 296714 675451 296716
rect 675404 296712 675496 296714
rect 675446 296656 675496 296712
rect 675404 296654 675496 296656
rect 675404 296652 675451 296654
rect 675385 296651 675451 296652
rect 42006 296442 42012 296444
rect 41492 296382 42012 296442
rect 42006 296380 42012 296382
rect 42076 296380 42082 296444
rect 675753 296304 675819 296309
rect 675753 296248 675758 296304
rect 675814 296248 675819 296304
rect 675753 296243 675819 296248
rect 41321 296034 41387 296037
rect 41308 296032 41387 296034
rect 41308 295976 41326 296032
rect 41382 295976 41387 296032
rect 41308 295974 41387 295976
rect 41321 295971 41387 295974
rect 675756 295901 675816 296243
rect 675753 295896 675819 295901
rect 675753 295840 675758 295896
rect 675814 295840 675819 295896
rect 675753 295835 675819 295840
rect 41822 295626 41828 295628
rect 41492 295566 41828 295626
rect 41822 295564 41828 295566
rect 41892 295564 41898 295628
rect 42977 295218 43043 295221
rect 41492 295216 43043 295218
rect 41492 295160 42982 295216
rect 43038 295160 43043 295216
rect 41492 295158 43043 295160
rect 42977 295155 43043 295158
rect 675753 295218 675819 295221
rect 676806 295218 676812 295220
rect 675753 295216 676812 295218
rect 675753 295160 675758 295216
rect 675814 295160 676812 295216
rect 675753 295158 676812 295160
rect 675753 295155 675819 295158
rect 676806 295156 676812 295158
rect 676876 295156 676882 295220
rect 39297 294810 39363 294813
rect 39284 294808 39363 294810
rect 39284 294752 39302 294808
rect 39358 294752 39363 294808
rect 39284 294750 39363 294752
rect 39297 294747 39363 294750
rect 44817 294674 44883 294677
rect 45461 294674 45527 294677
rect 44817 294672 45527 294674
rect 44817 294616 44822 294672
rect 44878 294616 45466 294672
rect 45522 294616 45527 294672
rect 44817 294614 45527 294616
rect 44817 294611 44883 294614
rect 45461 294611 45527 294614
rect 45553 294402 45619 294405
rect 41492 294400 45619 294402
rect 41492 294344 45558 294400
rect 45614 294344 45619 294400
rect 41492 294342 45619 294344
rect 45553 294339 45619 294342
rect 44633 293994 44699 293997
rect 41492 293992 44699 293994
rect 41492 293936 44638 293992
rect 44694 293936 44699 293992
rect 41492 293934 44699 293936
rect 44633 293931 44699 293934
rect 43989 293586 44055 293589
rect 41492 293584 44055 293586
rect 41492 293528 43994 293584
rect 44050 293528 44055 293584
rect 41492 293526 44055 293528
rect 43989 293523 44055 293526
rect 43161 293178 43227 293181
rect 41492 293176 43227 293178
rect 41492 293120 43166 293176
rect 43222 293120 43227 293176
rect 41492 293118 43227 293120
rect 43161 293115 43227 293118
rect 41781 292908 41847 292909
rect 675385 292908 675451 292909
rect 41781 292904 41828 292908
rect 41892 292906 41898 292908
rect 675334 292906 675340 292908
rect 41781 292848 41786 292904
rect 41781 292844 41828 292848
rect 41892 292846 41938 292906
rect 675294 292846 675340 292906
rect 675404 292904 675451 292908
rect 675446 292848 675451 292904
rect 41892 292844 41898 292846
rect 675334 292844 675340 292846
rect 675404 292844 675451 292848
rect 41781 292843 41847 292844
rect 675385 292843 675451 292844
rect 40910 292592 40970 292740
rect 40534 292528 40540 292592
rect 40604 292528 40610 292592
rect 40902 292528 40908 292592
rect 40972 292528 40978 292592
rect 40542 292332 40602 292528
rect 41781 292228 41847 292229
rect 41781 292224 41828 292228
rect 41892 292226 41898 292228
rect 41781 292168 41786 292224
rect 41781 292164 41828 292168
rect 41892 292166 41938 292226
rect 41892 292164 41898 292166
rect 41781 292163 41847 292164
rect 675569 292092 675635 292093
rect 675518 292028 675524 292092
rect 675588 292090 675635 292092
rect 675588 292088 675680 292090
rect 675630 292032 675680 292088
rect 675588 292030 675680 292032
rect 675588 292028 675635 292030
rect 675569 292027 675635 292028
rect 41492 291894 41890 291954
rect 41830 291818 41890 291894
rect 45001 291818 45067 291821
rect 41830 291816 45067 291818
rect 41830 291760 45006 291816
rect 45062 291760 45067 291816
rect 41830 291758 45067 291760
rect 45001 291755 45067 291758
rect 43805 291546 43871 291549
rect 41492 291544 43871 291546
rect 41492 291488 43810 291544
rect 43866 291488 43871 291544
rect 41492 291486 43871 291488
rect 43805 291483 43871 291486
rect 675753 291546 675819 291549
rect 676438 291546 676444 291548
rect 675753 291544 676444 291546
rect 675753 291488 675758 291544
rect 675814 291488 676444 291544
rect 675753 291486 676444 291488
rect 675753 291483 675819 291486
rect 676438 291484 676444 291486
rect 676508 291484 676514 291548
rect 43437 291138 43503 291141
rect 41492 291136 43503 291138
rect 41492 291080 43442 291136
rect 43498 291080 43503 291136
rect 41492 291078 43503 291080
rect 43437 291075 43503 291078
rect 50337 290730 50403 290733
rect 41492 290728 50403 290730
rect 41492 290672 50342 290728
rect 50398 290672 50403 290728
rect 41492 290670 50403 290672
rect 50337 290667 50403 290670
rect 673545 290594 673611 290597
rect 675109 290594 675175 290597
rect 673545 290592 675175 290594
rect 673545 290536 673550 290592
rect 673606 290536 675114 290592
rect 675170 290536 675175 290592
rect 673545 290534 675175 290536
rect 673545 290531 673611 290534
rect 675109 290531 675175 290534
rect 41321 290322 41387 290325
rect 41308 290320 41387 290322
rect 41308 290264 41326 290320
rect 41382 290264 41387 290320
rect 41308 290262 41387 290264
rect 41321 290259 41387 290262
rect 49141 289914 49207 289917
rect 41492 289912 49207 289914
rect 41492 289856 49146 289912
rect 49202 289856 49207 289912
rect 41492 289854 49207 289856
rect 49141 289851 49207 289854
rect 672625 287874 672691 287877
rect 675109 287874 675175 287877
rect 672625 287872 675175 287874
rect 672625 287816 672630 287872
rect 672686 287816 675114 287872
rect 675170 287816 675175 287872
rect 672625 287814 675175 287816
rect 672625 287811 672691 287814
rect 675109 287811 675175 287814
rect 675753 287058 675819 287061
rect 676254 287058 676260 287060
rect 675753 287056 676260 287058
rect 675753 287000 675758 287056
rect 675814 287000 676260 287056
rect 675753 286998 676260 287000
rect 675753 286995 675819 286998
rect 676254 286996 676260 286998
rect 676324 286996 676330 287060
rect 674373 286650 674439 286653
rect 675385 286650 675451 286653
rect 674373 286648 675451 286650
rect 674373 286592 674378 286648
rect 674434 286592 675390 286648
rect 675446 286592 675451 286648
rect 674373 286590 675451 286592
rect 674373 286587 674439 286590
rect 675385 286587 675451 286590
rect 673729 285562 673795 285565
rect 675109 285562 675175 285565
rect 673729 285560 675175 285562
rect 673729 285504 673734 285560
rect 673790 285504 675114 285560
rect 675170 285504 675175 285560
rect 673729 285502 675175 285504
rect 673729 285499 673795 285502
rect 675109 285499 675175 285502
rect 651465 285290 651531 285293
rect 650164 285288 651531 285290
rect 650164 285232 651470 285288
rect 651526 285232 651531 285288
rect 650164 285230 651531 285232
rect 651465 285227 651531 285230
rect 62757 285154 62823 285157
rect 62757 285152 64492 285154
rect 62757 285096 62762 285152
rect 62818 285096 64492 285152
rect 62757 285094 64492 285096
rect 62757 285091 62823 285094
rect 675753 283658 675819 283661
rect 676070 283658 676076 283660
rect 675753 283656 676076 283658
rect 675753 283600 675758 283656
rect 675814 283600 676076 283656
rect 675753 283598 676076 283600
rect 675753 283595 675819 283598
rect 676070 283596 676076 283598
rect 676140 283596 676146 283660
rect 675661 282844 675727 282845
rect 675661 282840 675708 282844
rect 675772 282842 675778 282844
rect 675661 282784 675666 282840
rect 675661 282780 675708 282784
rect 675772 282782 675818 282842
rect 675772 282780 675778 282782
rect 675661 282779 675727 282780
rect 41965 281484 42031 281485
rect 41965 281480 42012 281484
rect 42076 281482 42082 281484
rect 41965 281424 41970 281480
rect 41965 281420 42012 281424
rect 42076 281422 42122 281482
rect 42076 281420 42082 281422
rect 41965 281419 42031 281420
rect 675661 281210 675727 281213
rect 675886 281210 675892 281212
rect 675661 281208 675892 281210
rect 675661 281152 675666 281208
rect 675722 281152 675892 281208
rect 675661 281150 675892 281152
rect 675661 281147 675727 281150
rect 675886 281148 675892 281150
rect 675956 281148 675962 281212
rect 42149 279850 42215 279853
rect 43161 279850 43227 279853
rect 42149 279848 43227 279850
rect 42149 279792 42154 279848
rect 42210 279792 43166 279848
rect 43222 279792 43227 279848
rect 42149 279790 43227 279792
rect 42149 279787 42215 279790
rect 43161 279787 43227 279790
rect 42425 278762 42491 278765
rect 55857 278762 55923 278765
rect 42425 278760 55923 278762
rect 42425 278704 42430 278760
rect 42486 278704 55862 278760
rect 55918 278704 55923 278760
rect 42425 278702 55923 278704
rect 42425 278699 42491 278702
rect 55857 278699 55923 278702
rect 42425 278218 42491 278221
rect 43805 278218 43871 278221
rect 42425 278216 43871 278218
rect 42425 278160 42430 278216
rect 42486 278160 43810 278216
rect 43866 278160 43871 278216
rect 42425 278158 43871 278160
rect 42425 278155 42491 278158
rect 43805 278155 43871 278158
rect 40902 277884 40908 277948
rect 40972 277946 40978 277948
rect 41781 277946 41847 277949
rect 40972 277944 41847 277946
rect 40972 277888 41786 277944
rect 41842 277888 41847 277944
rect 40972 277886 41847 277888
rect 40972 277884 40978 277886
rect 41781 277883 41847 277886
rect 40718 277612 40724 277676
rect 40788 277674 40794 277676
rect 42241 277674 42307 277677
rect 40788 277672 42307 277674
rect 40788 277616 42246 277672
rect 42302 277616 42307 277672
rect 40788 277614 42307 277616
rect 40788 277612 40794 277614
rect 42241 277611 42307 277614
rect 42057 277130 42123 277133
rect 45001 277130 45067 277133
rect 42057 277128 45067 277130
rect 42057 277072 42062 277128
rect 42118 277072 45006 277128
rect 45062 277072 45067 277128
rect 42057 277070 45067 277072
rect 42057 277067 42123 277070
rect 45001 277067 45067 277070
rect 42057 276722 42123 276725
rect 42977 276722 43043 276725
rect 42057 276720 43043 276722
rect 42057 276664 42062 276720
rect 42118 276664 42982 276720
rect 43038 276664 43043 276720
rect 42057 276662 43043 276664
rect 42057 276659 42123 276662
rect 42977 276659 43043 276662
rect 525149 275634 525215 275637
rect 525977 275634 526043 275637
rect 525149 275632 526043 275634
rect 525149 275576 525154 275632
rect 525210 275576 525982 275632
rect 526038 275576 526043 275632
rect 525149 275574 526043 275576
rect 525149 275571 525215 275574
rect 525977 275571 526043 275574
rect 669957 275362 670023 275365
rect 683297 275362 683363 275365
rect 669957 275360 683363 275362
rect 669957 275304 669962 275360
rect 670018 275304 683302 275360
rect 683358 275304 683363 275360
rect 669957 275302 683363 275304
rect 669957 275299 670023 275302
rect 683297 275299 683363 275302
rect 529565 275226 529631 275229
rect 626165 275226 626231 275229
rect 529565 275224 626231 275226
rect 529565 275168 529570 275224
rect 529626 275168 626170 275224
rect 626226 275168 626231 275224
rect 529565 275166 626231 275168
rect 529565 275163 529631 275166
rect 626165 275163 626231 275166
rect 40534 274212 40540 274276
rect 40604 274274 40610 274276
rect 41781 274274 41847 274277
rect 40604 274272 41847 274274
rect 40604 274216 41786 274272
rect 41842 274216 41847 274272
rect 40604 274214 41847 274216
rect 40604 274212 40610 274214
rect 41781 274211 41847 274214
rect 522389 274138 522455 274141
rect 595437 274138 595503 274141
rect 522389 274136 595503 274138
rect 522389 274080 522394 274136
rect 522450 274080 595442 274136
rect 595498 274080 595503 274136
rect 522389 274078 595503 274080
rect 522389 274075 522455 274078
rect 595437 274075 595503 274078
rect 513189 273866 513255 273869
rect 602521 273866 602587 273869
rect 513189 273864 602587 273866
rect 513189 273808 513194 273864
rect 513250 273808 602526 273864
rect 602582 273808 602587 273864
rect 513189 273806 602587 273808
rect 513189 273803 513255 273806
rect 602521 273803 602587 273806
rect 42057 273050 42123 273053
rect 43989 273050 44055 273053
rect 42057 273048 44055 273050
rect 42057 272992 42062 273048
rect 42118 272992 43994 273048
rect 44050 272992 44055 273048
rect 42057 272990 44055 272992
rect 42057 272987 42123 272990
rect 43989 272987 44055 272990
rect 42057 272778 42123 272781
rect 44541 272778 44607 272781
rect 42057 272776 44607 272778
rect 42057 272720 42062 272776
rect 42118 272720 44546 272776
rect 44602 272720 44607 272776
rect 42057 272718 44607 272720
rect 42057 272715 42123 272718
rect 44541 272715 44607 272718
rect 521561 272778 521627 272781
rect 614389 272778 614455 272781
rect 521561 272776 614455 272778
rect 521561 272720 521566 272776
rect 521622 272720 614394 272776
rect 614450 272720 614455 272776
rect 521561 272718 614455 272720
rect 521561 272715 521627 272718
rect 614389 272715 614455 272718
rect 533889 272506 533955 272509
rect 632145 272506 632211 272509
rect 533889 272504 632211 272506
rect 533889 272448 533894 272504
rect 533950 272448 632150 272504
rect 632206 272448 632211 272504
rect 533889 272446 632211 272448
rect 533889 272443 533955 272446
rect 632145 272443 632211 272446
rect 478597 271418 478663 271421
rect 551737 271418 551803 271421
rect 478597 271416 551803 271418
rect 478597 271360 478602 271416
rect 478658 271360 551742 271416
rect 551798 271360 551803 271416
rect 478597 271358 551803 271360
rect 478597 271355 478663 271358
rect 551737 271355 551803 271358
rect 507669 271146 507735 271149
rect 593137 271146 593203 271149
rect 507669 271144 593203 271146
rect 507669 271088 507674 271144
rect 507730 271088 593142 271144
rect 593198 271088 593203 271144
rect 507669 271086 593203 271088
rect 507669 271083 507735 271086
rect 593137 271083 593203 271086
rect 664437 271146 664503 271149
rect 683113 271146 683179 271149
rect 664437 271144 683179 271146
rect 664437 271088 664442 271144
rect 664498 271088 683118 271144
rect 683174 271088 683179 271144
rect 664437 271086 683179 271088
rect 664437 271083 664503 271086
rect 683113 271083 683179 271086
rect 41454 270404 41460 270468
rect 41524 270466 41530 270468
rect 41781 270466 41847 270469
rect 41524 270464 41847 270466
rect 41524 270408 41786 270464
rect 41842 270408 41847 270464
rect 41524 270406 41847 270408
rect 41524 270404 41530 270406
rect 41781 270403 41847 270406
rect 530945 270330 531011 270333
rect 626533 270330 626599 270333
rect 530945 270328 626599 270330
rect 530945 270272 530950 270328
rect 531006 270272 626538 270328
rect 626594 270272 626599 270328
rect 530945 270270 626599 270272
rect 530945 270267 531011 270270
rect 626533 270267 626599 270270
rect 538029 270058 538095 270061
rect 637573 270058 637639 270061
rect 538029 270056 637639 270058
rect 538029 270000 538034 270056
rect 538090 270000 637578 270056
rect 637634 270000 637639 270056
rect 538029 269998 637639 270000
rect 538029 269995 538095 269998
rect 637573 269995 637639 269998
rect 102041 269786 102107 269789
rect 161289 269786 161355 269789
rect 102041 269784 161355 269786
rect 102041 269728 102046 269784
rect 102102 269728 161294 269784
rect 161350 269728 161355 269784
rect 102041 269726 161355 269728
rect 102041 269723 102107 269726
rect 161289 269723 161355 269726
rect 468753 269786 468819 269789
rect 537661 269786 537727 269789
rect 468753 269784 537727 269786
rect 468753 269728 468758 269784
rect 468814 269728 537666 269784
rect 537722 269728 537727 269784
rect 468753 269726 537727 269728
rect 468753 269723 468819 269726
rect 537661 269723 537727 269726
rect 540513 269786 540579 269789
rect 640701 269786 640767 269789
rect 540513 269784 640767 269786
rect 540513 269728 540518 269784
rect 540574 269728 640706 269784
rect 640762 269728 640767 269784
rect 540513 269726 640767 269728
rect 540513 269723 540579 269726
rect 640701 269723 640767 269726
rect 497273 269514 497339 269517
rect 568573 269514 568639 269517
rect 497273 269512 568639 269514
rect 497273 269456 497278 269512
rect 497334 269456 568578 269512
rect 568634 269456 568639 269512
rect 497273 269454 568639 269456
rect 497273 269451 497339 269454
rect 568573 269451 568639 269454
rect 470961 269242 471027 269245
rect 539501 269242 539567 269245
rect 470961 269240 539567 269242
rect 470961 269184 470966 269240
rect 471022 269184 539506 269240
rect 539562 269184 539567 269240
rect 470961 269182 539567 269184
rect 470961 269179 471027 269182
rect 539501 269179 539567 269182
rect 41781 269108 41847 269109
rect 41781 269104 41828 269108
rect 41892 269106 41898 269108
rect 41781 269048 41786 269104
rect 41781 269044 41828 269048
rect 41892 269046 41938 269106
rect 41892 269044 41898 269046
rect 41781 269043 41847 269044
rect 676262 268562 676322 268668
rect 683297 268562 683363 268565
rect 663750 268502 676322 268562
rect 683254 268560 683363 268562
rect 683254 268504 683302 268560
rect 683358 268504 683363 268560
rect 506105 268426 506171 268429
rect 591021 268426 591087 268429
rect 506105 268424 591087 268426
rect 506105 268368 506110 268424
rect 506166 268368 591026 268424
rect 591082 268368 591087 268424
rect 506105 268366 591087 268368
rect 506105 268363 506171 268366
rect 591021 268363 591087 268366
rect 663057 268154 663123 268157
rect 663750 268154 663810 268502
rect 683254 268499 683363 268504
rect 683254 268260 683314 268499
rect 683113 268154 683179 268157
rect 663057 268152 663810 268154
rect 663057 268096 663062 268152
rect 663118 268096 663810 268152
rect 663057 268094 663810 268096
rect 683070 268152 683179 268154
rect 683070 268096 683118 268152
rect 683174 268096 683179 268152
rect 663057 268091 663123 268094
rect 683070 268091 683179 268096
rect 683070 267852 683130 268091
rect 42425 267746 42491 267749
rect 45553 267746 45619 267749
rect 42425 267744 45619 267746
rect 42425 267688 42430 267744
rect 42486 267688 45558 267744
rect 45614 267688 45619 267744
rect 42425 267686 45619 267688
rect 42425 267683 42491 267686
rect 45553 267683 45619 267686
rect 519813 267610 519879 267613
rect 563697 267610 563763 267613
rect 519813 267608 563763 267610
rect 519813 267552 519818 267608
rect 519874 267552 563702 267608
rect 563758 267552 563763 267608
rect 519813 267550 563763 267552
rect 519813 267547 519879 267550
rect 563697 267547 563763 267550
rect 673085 267610 673151 267613
rect 675017 267610 675083 267613
rect 673085 267608 675083 267610
rect 673085 267552 673090 267608
rect 673146 267552 675022 267608
rect 675078 267552 675083 267608
rect 673085 267550 675083 267552
rect 673085 267547 673151 267550
rect 675017 267547 675083 267550
rect 517145 267338 517211 267341
rect 585777 267338 585843 267341
rect 676262 267338 676322 267444
rect 517145 267336 585843 267338
rect 517145 267280 517150 267336
rect 517206 267280 585782 267336
rect 585838 267280 585843 267336
rect 517145 267278 585843 267280
rect 517145 267275 517211 267278
rect 585777 267275 585843 267278
rect 674606 267278 676322 267338
rect 75913 267066 75979 267069
rect 138105 267066 138171 267069
rect 75913 267064 138171 267066
rect 75913 267008 75918 267064
rect 75974 267008 138110 267064
rect 138166 267008 138171 267064
rect 75913 267006 138171 267008
rect 75913 267003 75979 267006
rect 138105 267003 138171 267006
rect 467557 267066 467623 267069
rect 509693 267066 509759 267069
rect 467557 267064 509759 267066
rect 467557 267008 467562 267064
rect 467618 267008 509698 267064
rect 509754 267008 509759 267064
rect 467557 267006 509759 267008
rect 467557 267003 467623 267006
rect 509693 267003 509759 267006
rect 539685 267066 539751 267069
rect 625797 267066 625863 267069
rect 539685 267064 625863 267066
rect 539685 267008 539690 267064
rect 539746 267008 625802 267064
rect 625858 267008 625863 267064
rect 539685 267006 625863 267008
rect 539685 267003 539751 267006
rect 625797 267003 625863 267006
rect 672809 266930 672875 266933
rect 674606 266930 674666 267278
rect 676262 266930 676322 267036
rect 672809 266928 674666 266930
rect 672809 266872 672814 266928
rect 672870 266872 674666 266928
rect 672809 266870 674666 266872
rect 674790 266870 676322 266930
rect 672809 266867 672875 266870
rect 672809 266522 672875 266525
rect 674790 266522 674850 266870
rect 675017 266658 675083 266661
rect 675017 266656 676292 266658
rect 675017 266600 675022 266656
rect 675078 266600 676292 266656
rect 675017 266598 676292 266600
rect 675017 266595 675083 266598
rect 672809 266520 674850 266522
rect 672809 266464 672814 266520
rect 672870 266464 674850 266520
rect 672809 266462 674850 266464
rect 672809 266459 672875 266462
rect 673085 266114 673151 266117
rect 676262 266114 676322 266220
rect 673085 266112 676322 266114
rect 673085 266056 673090 266112
rect 673146 266056 676322 266112
rect 673085 266054 676322 266056
rect 673085 266051 673151 266054
rect 674557 265842 674623 265845
rect 674557 265840 676292 265842
rect 674557 265784 674562 265840
rect 674618 265784 676292 265840
rect 674557 265782 676292 265784
rect 674557 265779 674623 265782
rect 674557 265434 674623 265437
rect 674557 265432 676292 265434
rect 674557 265376 674562 265432
rect 674618 265376 676292 265432
rect 674557 265374 676292 265376
rect 674557 265371 674623 265374
rect 674189 265026 674255 265029
rect 674189 265024 676292 265026
rect 674189 264968 674194 265024
rect 674250 264968 676292 265024
rect 674189 264966 676292 264968
rect 674189 264963 674255 264966
rect 674373 264618 674439 264621
rect 674373 264616 676292 264618
rect 674373 264560 674378 264616
rect 674434 264560 676292 264616
rect 674373 264558 676292 264560
rect 674373 264555 674439 264558
rect 675017 264210 675083 264213
rect 675017 264208 676292 264210
rect 675017 264152 675022 264208
rect 675078 264152 676292 264208
rect 675017 264150 676292 264152
rect 675017 264147 675083 264150
rect 676070 263604 676076 263668
rect 676140 263666 676146 263668
rect 676262 263666 676322 263772
rect 676140 263606 676322 263666
rect 676140 263604 676146 263606
rect 678286 263261 678346 263364
rect 678237 263256 678346 263261
rect 678237 263200 678242 263256
rect 678298 263200 678346 263256
rect 678237 263198 678346 263200
rect 678237 263195 678303 263198
rect 676446 262853 676506 262956
rect 676397 262848 676506 262853
rect 676397 262792 676402 262848
rect 676458 262792 676506 262848
rect 676397 262790 676506 262792
rect 676397 262787 676463 262790
rect 676262 262445 676322 262548
rect 676213 262440 676322 262445
rect 676213 262384 676218 262440
rect 676274 262384 676322 262440
rect 676213 262382 676322 262384
rect 676213 262379 676279 262382
rect 554405 262170 554471 262173
rect 552460 262168 554471 262170
rect 552460 262112 554410 262168
rect 554466 262112 554471 262168
rect 552460 262110 554471 262112
rect 554405 262107 554471 262110
rect 674833 262034 674899 262037
rect 676262 262034 676322 262140
rect 674833 262032 676322 262034
rect 674833 261976 674838 262032
rect 674894 261976 676322 262032
rect 674833 261974 676322 261976
rect 674833 261971 674899 261974
rect 670417 261626 670483 261629
rect 676998 261628 677058 261732
rect 670417 261624 676506 261626
rect 670417 261568 670422 261624
rect 670478 261568 676506 261624
rect 670417 261566 676506 261568
rect 670417 261563 670483 261566
rect 676446 261324 676506 261566
rect 676990 261564 676996 261628
rect 677060 261564 677066 261628
rect 671705 261218 671771 261221
rect 674833 261218 674899 261221
rect 671705 261216 674899 261218
rect 671705 261160 671710 261216
rect 671766 261160 674838 261216
rect 674894 261160 674899 261216
rect 671705 261158 674899 261160
rect 671705 261155 671771 261158
rect 674833 261155 674899 261158
rect 675886 261156 675892 261220
rect 675956 261218 675962 261220
rect 676213 261218 676279 261221
rect 675956 261216 676279 261218
rect 675956 261160 676218 261216
rect 676274 261160 676279 261216
rect 675956 261158 676279 261160
rect 675956 261156 675962 261158
rect 676213 261155 676279 261158
rect 671521 260946 671587 260949
rect 671521 260944 676292 260946
rect 671521 260888 671526 260944
rect 671582 260888 676292 260944
rect 671521 260886 676292 260888
rect 671521 260883 671587 260886
rect 670233 260402 670299 260405
rect 676262 260402 676322 260508
rect 670233 260400 676322 260402
rect 670233 260344 670238 260400
rect 670294 260344 676322 260400
rect 670233 260342 676322 260344
rect 670233 260339 670299 260342
rect 35801 259994 35867 259997
rect 54477 259994 54543 259997
rect 554313 259994 554379 259997
rect 676814 259996 676874 260100
rect 35801 259992 54543 259994
rect 35801 259936 35806 259992
rect 35862 259936 54482 259992
rect 54538 259936 54543 259992
rect 35801 259934 54543 259936
rect 552460 259992 554379 259994
rect 552460 259936 554318 259992
rect 554374 259936 554379 259992
rect 552460 259934 554379 259936
rect 35801 259931 35867 259934
rect 54477 259931 54543 259934
rect 554313 259931 554379 259934
rect 676806 259932 676812 259996
rect 676876 259932 676882 259996
rect 673637 259722 673703 259725
rect 673637 259720 676292 259722
rect 673637 259664 673642 259720
rect 673698 259664 676292 259720
rect 673637 259662 676292 259664
rect 673637 259659 673703 259662
rect 675661 259178 675727 259181
rect 676262 259178 676322 259284
rect 675661 259176 676322 259178
rect 675661 259120 675666 259176
rect 675722 259120 676322 259176
rect 675661 259118 676322 259120
rect 675661 259115 675727 259118
rect 674097 258906 674163 258909
rect 674097 258904 676292 258906
rect 674097 258848 674102 258904
rect 674158 258848 676292 258904
rect 674097 258846 676292 258848
rect 674097 258843 674163 258846
rect 673637 258498 673703 258501
rect 673637 258496 676292 258498
rect 673637 258440 673642 258496
rect 673698 258440 676292 258496
rect 673637 258438 676292 258440
rect 673637 258435 673703 258438
rect 35801 258362 35867 258365
rect 35758 258360 35867 258362
rect 35758 258304 35806 258360
rect 35862 258304 35867 258360
rect 35758 258299 35867 258304
rect 35758 258060 35818 258299
rect 675661 258226 675727 258229
rect 675661 258224 675954 258226
rect 675661 258168 675666 258224
rect 675722 258168 675954 258224
rect 675661 258166 675954 258168
rect 675661 258163 675727 258166
rect 672625 257954 672691 257957
rect 675894 257954 675954 258166
rect 672625 257952 675954 257954
rect 672625 257896 672630 257952
rect 672686 257896 675954 257952
rect 672625 257894 675954 257896
rect 672625 257891 672691 257894
rect 553945 257818 554011 257821
rect 552460 257816 554011 257818
rect 552460 257760 553950 257816
rect 554006 257760 554011 257816
rect 552460 257758 554011 257760
rect 553945 257755 554011 257758
rect 43621 257682 43687 257685
rect 41492 257680 43687 257682
rect 41492 257624 43626 257680
rect 43682 257624 43687 257680
rect 41492 257622 43687 257624
rect 43621 257619 43687 257622
rect 675293 257546 675359 257549
rect 676262 257546 676322 258060
rect 675293 257544 676322 257546
rect 675293 257488 675298 257544
rect 675354 257488 676322 257544
rect 675293 257486 676322 257488
rect 675293 257483 675359 257486
rect 46197 257274 46263 257277
rect 41492 257272 46263 257274
rect 41492 257216 46202 257272
rect 46258 257216 46263 257272
rect 41492 257214 46263 257216
rect 46197 257211 46263 257214
rect 672625 257138 672691 257141
rect 676262 257138 676322 257244
rect 672625 257136 676322 257138
rect 672625 257080 672630 257136
rect 672686 257080 676322 257136
rect 672625 257078 676322 257080
rect 672625 257075 672691 257078
rect 44173 256866 44239 256869
rect 41492 256864 44239 256866
rect 41492 256808 44178 256864
rect 44234 256808 44239 256864
rect 41492 256806 44239 256808
rect 44173 256803 44239 256806
rect 671337 256730 671403 256733
rect 675293 256730 675359 256733
rect 671337 256728 675359 256730
rect 671337 256672 671342 256728
rect 671398 256672 675298 256728
rect 675354 256672 675359 256728
rect 671337 256670 675359 256672
rect 671337 256667 671403 256670
rect 675293 256667 675359 256670
rect 43253 256458 43319 256461
rect 41492 256456 43319 256458
rect 41492 256400 43258 256456
rect 43314 256400 43319 256456
rect 41492 256398 43319 256400
rect 43253 256395 43319 256398
rect 45093 256050 45159 256053
rect 41492 256048 45159 256050
rect 41492 255992 45098 256048
rect 45154 255992 45159 256048
rect 41492 255990 45159 255992
rect 45093 255987 45159 255990
rect 43161 255642 43227 255645
rect 553485 255642 553551 255645
rect 41492 255640 43227 255642
rect 41492 255584 43166 255640
rect 43222 255584 43227 255640
rect 41492 255582 43227 255584
rect 552460 255640 553551 255642
rect 552460 255584 553490 255640
rect 553546 255584 553551 255640
rect 552460 255582 553551 255584
rect 43161 255579 43227 255582
rect 553485 255579 553551 255582
rect 44357 255234 44423 255237
rect 41492 255232 44423 255234
rect 41492 255176 44362 255232
rect 44418 255176 44423 255232
rect 41492 255174 44423 255176
rect 44357 255171 44423 255174
rect 42793 254826 42859 254829
rect 41492 254824 42859 254826
rect 41492 254768 42798 254824
rect 42854 254768 42859 254824
rect 41492 254766 42859 254768
rect 42793 254763 42859 254766
rect 42977 254418 43043 254421
rect 41492 254416 43043 254418
rect 41492 254360 42982 254416
rect 43038 254360 43043 254416
rect 41492 254358 43043 254360
rect 42977 254355 43043 254358
rect 44173 254010 44239 254013
rect 41492 254008 44239 254010
rect 41492 253952 44178 254008
rect 44234 253952 44239 254008
rect 41492 253950 44239 253952
rect 44173 253947 44239 253950
rect 35574 253469 35634 253572
rect 35574 253464 35683 253469
rect 554405 253466 554471 253469
rect 35574 253408 35622 253464
rect 35678 253408 35683 253464
rect 35574 253406 35683 253408
rect 552460 253464 554471 253466
rect 552460 253408 554410 253464
rect 554466 253408 554471 253464
rect 552460 253406 554471 253408
rect 35617 253403 35683 253406
rect 554405 253403 554471 253406
rect 35758 253061 35818 253164
rect 35758 253056 35867 253061
rect 35758 253000 35806 253056
rect 35862 253000 35867 253056
rect 35758 252998 35867 253000
rect 35801 252995 35867 252998
rect 45553 252786 45619 252789
rect 41492 252784 45619 252786
rect 41492 252728 45558 252784
rect 45614 252728 45619 252784
rect 41492 252726 45619 252728
rect 45553 252723 45619 252726
rect 35758 252245 35818 252348
rect 35758 252240 35867 252245
rect 35758 252184 35806 252240
rect 35862 252184 35867 252240
rect 35758 252182 35867 252184
rect 35801 252179 35867 252182
rect 47025 251970 47091 251973
rect 41492 251968 47091 251970
rect 41492 251912 47030 251968
rect 47086 251912 47091 251968
rect 41492 251910 47091 251912
rect 47025 251907 47091 251910
rect 40542 251428 40602 251532
rect 40534 251364 40540 251428
rect 40604 251364 40610 251428
rect 554129 251290 554195 251293
rect 552460 251288 554195 251290
rect 552460 251232 554134 251288
rect 554190 251232 554195 251288
rect 552460 251230 554195 251232
rect 554129 251227 554195 251230
rect 45829 251154 45895 251157
rect 41492 251152 45895 251154
rect 41492 251096 45834 251152
rect 45890 251096 45895 251152
rect 41492 251094 45895 251096
rect 45829 251091 45895 251094
rect 47209 250746 47275 250749
rect 41492 250744 47275 250746
rect 41492 250688 47214 250744
rect 47270 250688 47275 250744
rect 41492 250686 47275 250688
rect 47209 250683 47275 250686
rect 44357 250338 44423 250341
rect 41492 250336 44423 250338
rect 41492 250280 44362 250336
rect 44418 250280 44423 250336
rect 41492 250278 44423 250280
rect 44357 250275 44423 250278
rect 675753 250338 675819 250341
rect 676990 250338 676996 250340
rect 675753 250336 676996 250338
rect 675753 250280 675758 250336
rect 675814 250280 676996 250336
rect 675753 250278 676996 250280
rect 675753 250275 675819 250278
rect 676990 250276 676996 250278
rect 677060 250276 677066 250340
rect 40726 249796 40786 249900
rect 40718 249732 40724 249796
rect 40788 249732 40794 249796
rect 675886 249658 675892 249660
rect 674790 249598 675892 249658
rect 46013 249522 46079 249525
rect 41492 249520 46079 249522
rect 41492 249464 46018 249520
rect 46074 249464 46079 249520
rect 41492 249462 46079 249464
rect 46013 249459 46079 249462
rect 674790 249389 674850 249598
rect 675886 249596 675892 249598
rect 675956 249596 675962 249660
rect 676070 249596 676076 249660
rect 676140 249596 676146 249660
rect 674790 249384 674899 249389
rect 674790 249328 674838 249384
rect 674894 249328 674899 249384
rect 674790 249326 674899 249328
rect 674833 249323 674899 249326
rect 675017 249386 675083 249389
rect 675385 249386 675451 249389
rect 675017 249384 675451 249386
rect 675017 249328 675022 249384
rect 675078 249328 675390 249384
rect 675446 249328 675451 249384
rect 675017 249326 675451 249328
rect 675017 249323 675083 249326
rect 675385 249323 675451 249326
rect 43621 249114 43687 249117
rect 553853 249114 553919 249117
rect 41492 249112 43687 249114
rect 41492 249056 43626 249112
rect 43682 249056 43687 249112
rect 41492 249054 43687 249056
rect 552460 249112 553919 249114
rect 552460 249056 553858 249112
rect 553914 249056 553919 249112
rect 552460 249054 553919 249056
rect 43621 249051 43687 249054
rect 553853 249051 553919 249054
rect 44541 248706 44607 248709
rect 41492 248704 44607 248706
rect 41492 248648 44546 248704
rect 44602 248648 44607 248704
rect 41492 248646 44607 248648
rect 44541 248643 44607 248646
rect 675017 248434 675083 248437
rect 676078 248434 676138 249596
rect 675017 248432 676138 248434
rect 675017 248376 675022 248432
rect 675078 248376 676138 248432
rect 675017 248374 676138 248376
rect 675017 248371 675083 248374
rect 45001 248298 45067 248301
rect 41492 248296 45067 248298
rect 41492 248240 45006 248296
rect 45062 248240 45067 248296
rect 41492 248238 45067 248240
rect 45001 248235 45067 248238
rect 46197 247890 46263 247893
rect 41492 247888 46263 247890
rect 41492 247832 46202 247888
rect 46258 247832 46263 247888
rect 41492 247830 46263 247832
rect 46197 247827 46263 247830
rect 47761 247482 47827 247485
rect 41492 247480 47827 247482
rect 41492 247424 47766 247480
rect 47822 247424 47827 247480
rect 41492 247422 47827 247424
rect 47761 247419 47827 247422
rect 670417 247074 670483 247077
rect 675293 247074 675359 247077
rect 670417 247072 675359 247074
rect 34470 246941 34530 247044
rect 670417 247016 670422 247072
rect 670478 247016 675298 247072
rect 675354 247016 675359 247072
rect 670417 247014 675359 247016
rect 670417 247011 670483 247014
rect 675293 247011 675359 247014
rect 34421 246936 34530 246941
rect 554405 246938 554471 246941
rect 34421 246880 34426 246936
rect 34482 246880 34530 246936
rect 34421 246878 34530 246880
rect 552460 246936 554471 246938
rect 552460 246880 554410 246936
rect 554466 246880 554471 246936
rect 552460 246878 554471 246880
rect 34421 246875 34487 246878
rect 554405 246875 554471 246878
rect 671521 246666 671587 246669
rect 675293 246666 675359 246669
rect 671521 246664 675359 246666
rect 41462 246530 41522 246636
rect 671521 246608 671526 246664
rect 671582 246608 675298 246664
rect 675354 246608 675359 246664
rect 671521 246606 675359 246608
rect 671521 246603 671587 246606
rect 675293 246603 675359 246606
rect 50521 246530 50587 246533
rect 41462 246528 50587 246530
rect 41462 246472 50526 246528
rect 50582 246472 50587 246528
rect 41462 246470 50587 246472
rect 50521 246467 50587 246470
rect 673453 245850 673519 245853
rect 675293 245850 675359 245853
rect 673453 245848 675359 245850
rect 673453 245792 673458 245848
rect 673514 245792 675298 245848
rect 675354 245792 675359 245848
rect 673453 245790 675359 245792
rect 673453 245787 673519 245790
rect 675293 245787 675359 245790
rect 675017 245578 675083 245581
rect 675334 245578 675340 245580
rect 675017 245576 675340 245578
rect 675017 245520 675022 245576
rect 675078 245520 675340 245576
rect 675017 245518 675340 245520
rect 675017 245515 675083 245518
rect 675334 245516 675340 245518
rect 675404 245516 675410 245580
rect 671705 245306 671771 245309
rect 674741 245306 674807 245309
rect 671705 245304 674807 245306
rect 671705 245248 671710 245304
rect 671766 245248 674746 245304
rect 674802 245248 674807 245304
rect 671705 245246 674807 245248
rect 671705 245243 671771 245246
rect 674741 245243 674807 245246
rect 674925 245306 674991 245309
rect 676806 245306 676812 245308
rect 674925 245304 676812 245306
rect 674925 245248 674930 245304
rect 674986 245248 676812 245304
rect 674925 245246 676812 245248
rect 674925 245243 674991 245246
rect 676806 245244 676812 245246
rect 676876 245244 676882 245308
rect 553393 244762 553459 244765
rect 552460 244760 553459 244762
rect 552460 244704 553398 244760
rect 553454 244704 553459 244760
rect 552460 244702 553459 244704
rect 553393 244699 553459 244702
rect 41689 242858 41755 242861
rect 42425 242858 42491 242861
rect 41689 242856 42491 242858
rect 41689 242800 41694 242856
rect 41750 242800 42430 242856
rect 42486 242800 42491 242856
rect 41689 242798 42491 242800
rect 41689 242795 41755 242798
rect 42425 242795 42491 242798
rect 672533 242858 672599 242861
rect 675109 242858 675175 242861
rect 672533 242856 675175 242858
rect 672533 242800 672538 242856
rect 672594 242800 675114 242856
rect 675170 242800 675175 242856
rect 672533 242798 675175 242800
rect 672533 242795 672599 242798
rect 675109 242795 675175 242798
rect 553945 242586 554011 242589
rect 552460 242584 554011 242586
rect 552460 242528 553950 242584
rect 554006 242528 554011 242584
rect 552460 242526 554011 242528
rect 553945 242523 554011 242526
rect 40677 241498 40743 241501
rect 43805 241498 43871 241501
rect 40677 241496 43871 241498
rect 40677 241440 40682 241496
rect 40738 241440 43810 241496
rect 43866 241440 43871 241496
rect 40677 241438 43871 241440
rect 40677 241435 40743 241438
rect 43805 241435 43871 241438
rect 674097 241498 674163 241501
rect 675109 241498 675175 241501
rect 674097 241496 675175 241498
rect 674097 241440 674102 241496
rect 674158 241440 675114 241496
rect 675170 241440 675175 241496
rect 674097 241438 675175 241440
rect 674097 241435 674163 241438
rect 675109 241435 675175 241438
rect 554037 240410 554103 240413
rect 552460 240408 554103 240410
rect 552460 240352 554042 240408
rect 554098 240352 554103 240408
rect 552460 240350 554103 240352
rect 554037 240347 554103 240350
rect 670233 240274 670299 240277
rect 675109 240274 675175 240277
rect 670233 240272 675175 240274
rect 670233 240216 670238 240272
rect 670294 240216 675114 240272
rect 675170 240216 675175 240272
rect 670233 240214 675175 240216
rect 670233 240211 670299 240214
rect 675109 240211 675175 240214
rect 40534 240076 40540 240140
rect 40604 240138 40610 240140
rect 41781 240138 41847 240141
rect 40604 240136 41847 240138
rect 40604 240080 41786 240136
rect 41842 240080 41847 240136
rect 40604 240078 41847 240080
rect 40604 240076 40610 240078
rect 41781 240075 41847 240078
rect 675385 238644 675451 238645
rect 675334 238642 675340 238644
rect 675294 238582 675340 238642
rect 675404 238640 675451 238644
rect 675446 238584 675451 238640
rect 675334 238580 675340 238582
rect 675404 238580 675451 238584
rect 675385 238579 675451 238580
rect 554313 238234 554379 238237
rect 552460 238232 554379 238234
rect 552460 238176 554318 238232
rect 554374 238176 554379 238232
rect 552460 238174 554379 238176
rect 554313 238171 554379 238174
rect 42006 238036 42012 238100
rect 42076 238098 42082 238100
rect 42425 238098 42491 238101
rect 42076 238096 42491 238098
rect 42076 238040 42430 238096
rect 42486 238040 42491 238096
rect 42076 238038 42491 238040
rect 42076 238036 42082 238038
rect 42425 238035 42491 238038
rect 671337 237826 671403 237829
rect 675385 237826 675451 237829
rect 671337 237824 675451 237826
rect 671337 237768 671342 237824
rect 671398 237768 675390 237824
rect 675446 237768 675451 237824
rect 671337 237766 675451 237768
rect 671337 237763 671403 237766
rect 675385 237763 675451 237766
rect 669957 237146 670023 237149
rect 673521 237146 673587 237149
rect 669957 237144 673587 237146
rect 669957 237088 669962 237144
rect 670018 237088 673526 237144
rect 673582 237088 673587 237144
rect 669957 237086 673587 237088
rect 669957 237083 670023 237086
rect 673521 237083 673587 237086
rect 670233 236874 670299 236877
rect 673407 236874 673473 236877
rect 670233 236872 673473 236874
rect 670233 236816 670238 236872
rect 670294 236816 673412 236872
rect 673468 236816 673473 236872
rect 670233 236814 673473 236816
rect 670233 236811 670299 236814
rect 673407 236811 673473 236814
rect 673453 236330 673519 236333
rect 676806 236330 676812 236332
rect 673453 236328 676812 236330
rect 673453 236272 673458 236328
rect 673514 236272 676812 236328
rect 673453 236270 676812 236272
rect 673453 236267 673519 236270
rect 676806 236268 676812 236270
rect 676876 236268 676882 236332
rect 554497 236058 554563 236061
rect 552460 236056 554563 236058
rect 552460 236000 554502 236056
rect 554558 236000 554563 236056
rect 552460 235998 554563 236000
rect 554497 235995 554563 235998
rect 673494 235996 673500 236060
rect 673564 236058 673570 236060
rect 673745 236058 673811 236061
rect 673564 236056 673811 236058
rect 673564 236000 673750 236056
rect 673806 236000 673811 236056
rect 673564 235998 673811 236000
rect 673564 235996 673570 235998
rect 673745 235995 673811 235998
rect 40718 235860 40724 235924
rect 40788 235922 40794 235924
rect 41781 235922 41847 235925
rect 40788 235920 41847 235922
rect 40788 235864 41786 235920
rect 41842 235864 41847 235920
rect 40788 235862 41847 235864
rect 40788 235860 40794 235862
rect 41781 235859 41847 235862
rect 42425 235922 42491 235925
rect 45001 235922 45067 235925
rect 42425 235920 45067 235922
rect 42425 235864 42430 235920
rect 42486 235864 45006 235920
rect 45062 235864 45067 235920
rect 42425 235862 45067 235864
rect 42425 235859 42491 235862
rect 45001 235859 45067 235862
rect 669405 234970 669471 234973
rect 674529 234970 674595 234973
rect 669405 234968 674595 234970
rect 669405 234912 669410 234968
rect 669466 234912 674534 234968
rect 674590 234912 674595 234968
rect 669405 234910 674595 234912
rect 669405 234907 669471 234910
rect 674529 234907 674595 234910
rect 668485 234562 668551 234565
rect 671061 234562 671127 234565
rect 668485 234560 671127 234562
rect 668485 234504 668490 234560
rect 668546 234504 671066 234560
rect 671122 234504 671127 234560
rect 668485 234502 671127 234504
rect 668485 234499 668551 234502
rect 671061 234499 671127 234502
rect 671286 234500 671292 234564
rect 671356 234562 671362 234564
rect 671705 234562 671771 234565
rect 671356 234560 671771 234562
rect 671356 234504 671710 234560
rect 671766 234504 671771 234560
rect 671356 234502 671771 234504
rect 671356 234500 671362 234502
rect 671705 234499 671771 234502
rect 674741 234426 674807 234429
rect 675845 234426 675911 234429
rect 674741 234424 675911 234426
rect 674741 234368 674746 234424
rect 674802 234368 675850 234424
rect 675906 234368 675911 234424
rect 674741 234366 675911 234368
rect 674741 234363 674807 234366
rect 675845 234363 675911 234366
rect 42241 234154 42307 234157
rect 44541 234154 44607 234157
rect 42241 234152 44607 234154
rect 42241 234096 42246 234152
rect 42302 234096 44546 234152
rect 44602 234096 44607 234152
rect 42241 234094 44607 234096
rect 42241 234091 42307 234094
rect 44541 234091 44607 234094
rect 660297 234154 660363 234157
rect 683297 234154 683363 234157
rect 660297 234152 683363 234154
rect 660297 234096 660302 234152
rect 660358 234096 683302 234152
rect 683358 234096 683363 234152
rect 660297 234094 683363 234096
rect 660297 234091 660363 234094
rect 683297 234091 683363 234094
rect 554405 233882 554471 233885
rect 552460 233880 554471 233882
rect 552460 233824 554410 233880
rect 554466 233824 554471 233880
rect 552460 233822 554471 233824
rect 554405 233819 554471 233822
rect 658917 233882 658983 233885
rect 683665 233882 683731 233885
rect 658917 233880 683731 233882
rect 658917 233824 658922 233880
rect 658978 233824 683670 233880
rect 683726 233824 683731 233880
rect 658917 233822 683731 233824
rect 658917 233819 658983 233822
rect 683665 233819 683731 233822
rect 674557 233474 674623 233477
rect 675845 233474 675911 233477
rect 674557 233472 675911 233474
rect 674557 233416 674562 233472
rect 674618 233416 675850 233472
rect 675906 233416 675911 233472
rect 674557 233414 675911 233416
rect 674557 233411 674623 233414
rect 675845 233411 675911 233414
rect 670141 232794 670207 232797
rect 673494 232794 673500 232796
rect 670141 232792 673500 232794
rect 670141 232736 670146 232792
rect 670202 232736 673500 232792
rect 670141 232734 673500 232736
rect 670141 232731 670207 232734
rect 673494 232732 673500 232734
rect 673564 232732 673570 232796
rect 42609 232522 42675 232525
rect 46013 232522 46079 232525
rect 42609 232520 46079 232522
rect 42609 232464 42614 232520
rect 42670 232464 46018 232520
rect 46074 232464 46079 232520
rect 42609 232462 46079 232464
rect 42609 232459 42675 232462
rect 46013 232459 46079 232462
rect 670601 232522 670667 232525
rect 673361 232522 673427 232525
rect 670601 232520 673427 232522
rect 670601 232464 670606 232520
rect 670662 232464 673366 232520
rect 673422 232464 673427 232520
rect 670601 232462 673427 232464
rect 670601 232459 670667 232462
rect 673361 232459 673427 232462
rect 42425 232250 42491 232253
rect 47025 232250 47091 232253
rect 42425 232248 47091 232250
rect 42425 232192 42430 232248
rect 42486 232192 47030 232248
rect 47086 232192 47091 232248
rect 42425 232190 47091 232192
rect 42425 232187 42491 232190
rect 47025 232187 47091 232190
rect 42425 231842 42491 231845
rect 43621 231842 43687 231845
rect 42425 231840 43687 231842
rect 42425 231784 42430 231840
rect 42486 231784 43626 231840
rect 43682 231784 43687 231840
rect 42425 231782 43687 231784
rect 42425 231779 42491 231782
rect 43621 231779 43687 231782
rect 663793 231842 663859 231845
rect 668945 231842 669011 231845
rect 663793 231840 669011 231842
rect 663793 231784 663798 231840
rect 663854 231784 668950 231840
rect 669006 231784 669011 231840
rect 663793 231782 669011 231784
rect 663793 231779 663859 231782
rect 668945 231779 669011 231782
rect 672901 231842 672967 231845
rect 673126 231842 673132 231844
rect 672901 231840 673132 231842
rect 672901 231784 672906 231840
rect 672962 231784 673132 231840
rect 672901 231782 673132 231784
rect 672901 231779 672967 231782
rect 673126 231780 673132 231782
rect 673196 231780 673202 231844
rect 673310 231780 673316 231844
rect 673380 231842 673386 231844
rect 673637 231842 673703 231845
rect 673380 231840 673703 231842
rect 673380 231784 673642 231840
rect 673698 231784 673703 231840
rect 673380 231782 673703 231784
rect 673380 231780 673386 231782
rect 673637 231779 673703 231782
rect 674230 231780 674236 231844
rect 674300 231842 674306 231844
rect 674465 231842 674531 231845
rect 674300 231840 674531 231842
rect 674300 231784 674470 231840
rect 674526 231784 674531 231840
rect 674300 231782 674531 231784
rect 674300 231780 674306 231782
rect 674465 231779 674531 231782
rect 668301 231570 668367 231573
rect 675173 231570 675239 231573
rect 668301 231568 675239 231570
rect 668301 231512 668306 231568
rect 668362 231512 675178 231568
rect 675234 231512 675239 231568
rect 668301 231510 675239 231512
rect 668301 231507 668367 231510
rect 675173 231507 675239 231510
rect 668945 231298 669011 231301
rect 675063 231298 675129 231301
rect 668945 231296 675129 231298
rect 668945 231240 668950 231296
rect 669006 231240 675068 231296
rect 675124 231240 675129 231296
rect 668945 231238 675129 231240
rect 668945 231235 669011 231238
rect 675063 231235 675129 231238
rect 662045 231162 662111 231165
rect 667933 231162 667999 231165
rect 662045 231160 667999 231162
rect 662045 231104 662050 231160
rect 662106 231104 667938 231160
rect 667994 231104 667999 231160
rect 662045 231102 667999 231104
rect 662045 231099 662111 231102
rect 667933 231099 667999 231102
rect 675017 231026 675083 231029
rect 676029 231026 676095 231029
rect 675017 231024 676095 231026
rect 675017 230968 675022 231024
rect 675078 230968 676034 231024
rect 676090 230968 676095 231024
rect 675017 230966 676095 230968
rect 675017 230963 675083 230966
rect 676029 230963 676095 230966
rect 664437 230890 664503 230893
rect 674725 230890 674791 230893
rect 664437 230888 674791 230890
rect 664437 230832 664442 230888
rect 664498 230832 674730 230888
rect 674786 230832 674791 230888
rect 664437 230830 674791 230832
rect 664437 230827 664503 230830
rect 674725 230827 674791 230830
rect 663057 230618 663123 230621
rect 668301 230618 668367 230621
rect 663057 230616 668367 230618
rect 663057 230560 663062 230616
rect 663118 230560 668306 230616
rect 668362 230560 668367 230616
rect 663057 230558 668367 230560
rect 663057 230555 663123 230558
rect 668301 230555 668367 230558
rect 42149 230482 42215 230485
rect 44357 230482 44423 230485
rect 42149 230480 44423 230482
rect 42149 230424 42154 230480
rect 42210 230424 44362 230480
rect 44418 230424 44423 230480
rect 42149 230422 44423 230424
rect 42149 230419 42215 230422
rect 44357 230419 44423 230422
rect 106917 230346 106983 230349
rect 166257 230346 166323 230349
rect 106917 230344 166323 230346
rect 106917 230288 106922 230344
rect 106978 230288 166262 230344
rect 166318 230288 166323 230344
rect 106917 230286 166323 230288
rect 106917 230283 106983 230286
rect 166257 230283 166323 230286
rect 665265 230346 665331 230349
rect 674389 230346 674455 230349
rect 665265 230344 674455 230346
rect 665265 230288 665270 230344
rect 665326 230288 674394 230344
rect 674450 230288 674455 230344
rect 665265 230286 674455 230288
rect 665265 230283 665331 230286
rect 674389 230283 674455 230286
rect 674649 230346 674715 230349
rect 676857 230346 676923 230349
rect 674649 230344 676923 230346
rect 674649 230288 674654 230344
rect 674710 230288 676862 230344
rect 676918 230288 676923 230344
rect 674649 230286 676923 230288
rect 674649 230283 674715 230286
rect 676857 230283 676923 230286
rect 71037 230074 71103 230077
rect 150801 230074 150867 230077
rect 71037 230072 150867 230074
rect 71037 230016 71042 230072
rect 71098 230016 150806 230072
rect 150862 230016 150867 230072
rect 71037 230014 150867 230016
rect 71037 230011 71103 230014
rect 150801 230011 150867 230014
rect 639597 230074 639663 230077
rect 673453 230074 673519 230077
rect 639597 230072 673519 230074
rect 639597 230016 639602 230072
rect 639658 230016 673458 230072
rect 673514 230016 673519 230072
rect 639597 230014 673519 230016
rect 639597 230011 639663 230014
rect 673453 230011 673519 230014
rect 673821 230074 673887 230077
rect 675109 230074 675175 230077
rect 673821 230072 675175 230074
rect 673821 230016 673826 230072
rect 673882 230016 675114 230072
rect 675170 230016 675175 230072
rect 673821 230014 675175 230016
rect 673821 230011 673887 230014
rect 675109 230011 675175 230014
rect 65517 229802 65583 229805
rect 148225 229802 148291 229805
rect 65517 229800 148291 229802
rect 65517 229744 65522 229800
rect 65578 229744 148230 229800
rect 148286 229744 148291 229800
rect 65517 229742 148291 229744
rect 65517 229739 65583 229742
rect 148225 229739 148291 229742
rect 660941 229802 661007 229805
rect 674833 229802 674899 229805
rect 660941 229800 674899 229802
rect 660941 229744 660946 229800
rect 661002 229744 674838 229800
rect 674894 229744 674899 229800
rect 660941 229742 674899 229744
rect 660941 229739 661007 229742
rect 674833 229739 674899 229742
rect 673269 229530 673335 229533
rect 675109 229530 675175 229533
rect 673269 229528 675175 229530
rect 673269 229472 673274 229528
rect 673330 229472 675114 229528
rect 675170 229472 675175 229528
rect 673269 229470 675175 229472
rect 673269 229467 673335 229470
rect 675109 229467 675175 229470
rect 671470 229332 671476 229396
rect 671540 229394 671546 229396
rect 671705 229394 671771 229397
rect 671540 229392 671771 229394
rect 671540 229336 671710 229392
rect 671766 229336 671771 229392
rect 671540 229334 671771 229336
rect 671540 229332 671546 229334
rect 671705 229331 671771 229334
rect 653397 229122 653463 229125
rect 673453 229122 673519 229125
rect 653397 229120 673519 229122
rect 653397 229064 653402 229120
rect 653458 229064 673458 229120
rect 673514 229064 673519 229120
rect 653397 229062 673519 229064
rect 653397 229059 653463 229062
rect 673453 229059 673519 229062
rect 41965 228988 42031 228989
rect 41965 228984 42012 228988
rect 42076 228986 42082 228988
rect 41965 228928 41970 228984
rect 41965 228924 42012 228928
rect 42076 228926 42122 228986
rect 42076 228924 42082 228926
rect 41965 228923 42031 228924
rect 113081 228850 113147 228853
rect 184933 228850 184999 228853
rect 113081 228848 184999 228850
rect 113081 228792 113086 228848
rect 113142 228792 184938 228848
rect 184994 228792 184999 228848
rect 113081 228790 184999 228792
rect 113081 228787 113147 228790
rect 184933 228787 184999 228790
rect 673361 228850 673427 228853
rect 675109 228850 675175 228853
rect 673361 228848 675175 228850
rect 673361 228792 673366 228848
rect 673422 228792 675114 228848
rect 675170 228792 675175 228848
rect 673361 228790 675175 228792
rect 673361 228787 673427 228790
rect 675109 228787 675175 228790
rect 64137 228578 64203 228581
rect 143073 228578 143139 228581
rect 64137 228576 143139 228578
rect 64137 228520 64142 228576
rect 64198 228520 143078 228576
rect 143134 228520 143139 228576
rect 64137 228518 143139 228520
rect 64137 228515 64203 228518
rect 143073 228515 143139 228518
rect 672257 228578 672323 228581
rect 672942 228578 672948 228580
rect 672257 228576 672948 228578
rect 672257 228520 672262 228576
rect 672318 228520 672948 228576
rect 672257 228518 672948 228520
rect 672257 228515 672323 228518
rect 672942 228516 672948 228518
rect 673012 228516 673018 228580
rect 673381 228578 673447 228581
rect 674966 228578 674972 228580
rect 673381 228576 674972 228578
rect 673381 228520 673386 228576
rect 673442 228520 674972 228576
rect 673381 228518 674972 228520
rect 673381 228515 673447 228518
rect 674966 228516 674972 228518
rect 675036 228516 675042 228580
rect 73797 228306 73863 228309
rect 155309 228306 155375 228309
rect 73797 228304 155375 228306
rect 73797 228248 73802 228304
rect 73858 228248 155314 228304
rect 155370 228248 155375 228304
rect 73797 228246 155375 228248
rect 73797 228243 73863 228246
rect 155309 228243 155375 228246
rect 169017 228306 169083 228309
rect 223573 228306 223639 228309
rect 169017 228304 223639 228306
rect 169017 228248 169022 228304
rect 169078 228248 223578 228304
rect 223634 228248 223639 228304
rect 169017 228246 223639 228248
rect 169017 228243 169083 228246
rect 223573 228243 223639 228246
rect 42425 227626 42491 227629
rect 43805 227626 43871 227629
rect 42425 227624 43871 227626
rect 42425 227568 42430 227624
rect 42486 227568 43810 227624
rect 43866 227568 43871 227624
rect 42425 227566 43871 227568
rect 42425 227563 42491 227566
rect 43805 227563 43871 227566
rect 136357 227490 136423 227493
rect 202965 227490 203031 227493
rect 136357 227488 203031 227490
rect 136357 227432 136362 227488
rect 136418 227432 202970 227488
rect 203026 227432 203031 227488
rect 136357 227430 203031 227432
rect 136357 227427 136423 227430
rect 202965 227427 203031 227430
rect 42241 227354 42307 227357
rect 47209 227354 47275 227357
rect 42241 227352 47275 227354
rect 42241 227296 42246 227352
rect 42302 227296 47214 227352
rect 47270 227296 47275 227352
rect 42241 227294 47275 227296
rect 42241 227291 42307 227294
rect 47209 227291 47275 227294
rect 89621 227218 89687 227221
rect 166901 227218 166967 227221
rect 89621 227216 166967 227218
rect 89621 227160 89626 227216
rect 89682 227160 166906 227216
rect 166962 227160 166967 227216
rect 89621 227158 166967 227160
rect 89621 227155 89687 227158
rect 166901 227155 166967 227158
rect 671797 227084 671863 227085
rect 671797 227080 671844 227084
rect 671908 227082 671914 227084
rect 672257 227082 672323 227085
rect 672993 227082 673059 227085
rect 671797 227024 671802 227080
rect 671797 227020 671844 227024
rect 671908 227022 671954 227082
rect 672257 227080 673059 227082
rect 672257 227024 672262 227080
rect 672318 227024 672998 227080
rect 673054 227024 673059 227080
rect 672257 227022 673059 227024
rect 671908 227020 671914 227022
rect 671797 227019 671863 227020
rect 672257 227019 672323 227022
rect 672993 227019 673059 227022
rect 673729 227082 673795 227085
rect 676213 227082 676279 227085
rect 673729 227080 676279 227082
rect 673729 227024 673734 227080
rect 673790 227024 676218 227080
rect 676274 227024 676279 227080
rect 673729 227022 676279 227024
rect 673729 227019 673795 227022
rect 676213 227019 676279 227022
rect 79961 226946 80027 226949
rect 160461 226946 160527 226949
rect 671613 226948 671679 226949
rect 671613 226946 671660 226948
rect 79961 226944 160527 226946
rect 79961 226888 79966 226944
rect 80022 226888 160466 226944
rect 160522 226888 160527 226944
rect 79961 226886 160527 226888
rect 671568 226944 671660 226946
rect 671568 226888 671618 226944
rect 671568 226886 671660 226888
rect 79961 226883 80027 226886
rect 160461 226883 160527 226886
rect 671613 226884 671660 226886
rect 671724 226884 671730 226948
rect 671613 226883 671679 226884
rect 673157 226810 673223 226813
rect 675293 226810 675359 226813
rect 673157 226808 675359 226810
rect 673157 226752 673162 226808
rect 673218 226752 675298 226808
rect 675354 226752 675359 226808
rect 673157 226750 675359 226752
rect 673157 226747 673223 226750
rect 675293 226747 675359 226750
rect 654777 226674 654843 226677
rect 671797 226674 671863 226677
rect 654777 226672 671863 226674
rect 654777 226616 654782 226672
rect 654838 226616 671802 226672
rect 671858 226616 671863 226672
rect 654777 226614 671863 226616
rect 654777 226611 654843 226614
rect 671797 226611 671863 226614
rect 672257 226538 672323 226541
rect 674741 226538 674807 226541
rect 672257 226536 674807 226538
rect 672257 226480 672262 226536
rect 672318 226480 674746 226536
rect 674802 226480 674807 226536
rect 672257 226478 674807 226480
rect 672257 226475 672323 226478
rect 674741 226475 674807 226478
rect 658917 226402 658983 226405
rect 658917 226400 666570 226402
rect 658917 226344 658922 226400
rect 658978 226344 666570 226400
rect 658917 226342 666570 226344
rect 658917 226339 658983 226342
rect 666510 226266 666570 226342
rect 670693 226266 670759 226269
rect 673729 226266 673795 226269
rect 666510 226264 670759 226266
rect 666510 226208 670698 226264
rect 670754 226208 670759 226264
rect 666510 226206 670759 226208
rect 670693 226203 670759 226206
rect 672030 226264 673795 226266
rect 672030 226208 673734 226264
rect 673790 226208 673795 226264
rect 672030 226206 673795 226208
rect 42425 226130 42491 226133
rect 45553 226130 45619 226133
rect 42425 226128 45619 226130
rect 42425 226072 42430 226128
rect 42486 226072 45558 226128
rect 45614 226072 45619 226128
rect 42425 226070 45619 226072
rect 42425 226067 42491 226070
rect 45553 226067 45619 226070
rect 125501 226130 125567 226133
rect 196525 226130 196591 226133
rect 125501 226128 196591 226130
rect 125501 226072 125506 226128
rect 125562 226072 196530 226128
rect 196586 226072 196591 226128
rect 125501 226070 196591 226072
rect 125501 226067 125567 226070
rect 196525 226067 196591 226070
rect 671797 226130 671863 226133
rect 672030 226130 672090 226206
rect 673729 226203 673795 226206
rect 671797 226128 672090 226130
rect 671797 226072 671802 226128
rect 671858 226072 672090 226128
rect 671797 226070 672090 226072
rect 671797 226067 671863 226070
rect 672165 225994 672231 225997
rect 674949 225994 675015 225997
rect 672165 225992 675015 225994
rect 672165 225936 672170 225992
rect 672226 225936 674954 225992
rect 675010 225936 675015 225992
rect 672165 225934 675015 225936
rect 672165 225931 672231 225934
rect 674949 225931 675015 225934
rect 89161 225858 89227 225861
rect 168189 225858 168255 225861
rect 89161 225856 168255 225858
rect 89161 225800 89166 225856
rect 89222 225800 168194 225856
rect 168250 225800 168255 225856
rect 89161 225798 168255 225800
rect 89161 225795 89227 225798
rect 168189 225795 168255 225798
rect 671153 225722 671219 225725
rect 663750 225720 671219 225722
rect 663750 225664 671158 225720
rect 671214 225664 671219 225720
rect 663750 225662 671219 225664
rect 42241 225586 42307 225589
rect 62757 225586 62823 225589
rect 42241 225584 62823 225586
rect 42241 225528 42246 225584
rect 42302 225528 62762 225584
rect 62818 225528 62823 225584
rect 42241 225526 62823 225528
rect 42241 225523 42307 225526
rect 62757 225523 62823 225526
rect 82537 225586 82603 225589
rect 163037 225586 163103 225589
rect 82537 225584 163103 225586
rect 82537 225528 82542 225584
rect 82598 225528 163042 225584
rect 163098 225528 163103 225584
rect 82537 225526 163103 225528
rect 82537 225523 82603 225526
rect 163037 225523 163103 225526
rect 650637 225586 650703 225589
rect 663750 225586 663810 225662
rect 671153 225659 671219 225662
rect 671813 225722 671879 225725
rect 672758 225722 672764 225724
rect 671813 225720 672764 225722
rect 671813 225664 671818 225720
rect 671874 225664 672764 225720
rect 671813 225662 672764 225664
rect 671813 225659 671879 225662
rect 672758 225660 672764 225662
rect 672828 225660 672834 225724
rect 673729 225722 673795 225725
rect 674373 225722 674439 225725
rect 673729 225720 674439 225722
rect 673729 225664 673734 225720
rect 673790 225664 674378 225720
rect 674434 225664 674439 225720
rect 673729 225662 674439 225664
rect 673729 225659 673795 225662
rect 674373 225659 674439 225662
rect 650637 225584 663810 225586
rect 650637 225528 650642 225584
rect 650698 225528 663810 225584
rect 650637 225526 663810 225528
rect 650637 225523 650703 225526
rect 665817 225450 665883 225453
rect 670693 225450 670759 225453
rect 665817 225448 670759 225450
rect 665817 225392 665822 225448
rect 665878 225392 670698 225448
rect 670754 225392 670759 225448
rect 665817 225390 670759 225392
rect 665817 225387 665883 225390
rect 670693 225387 670759 225390
rect 671153 225450 671219 225453
rect 673729 225450 673795 225453
rect 671153 225448 673795 225450
rect 671153 225392 671158 225448
rect 671214 225392 673734 225448
rect 673790 225392 673795 225448
rect 671153 225390 673795 225392
rect 671153 225387 671219 225390
rect 673729 225387 673795 225390
rect 671797 225178 671863 225181
rect 674557 225178 674623 225181
rect 671797 225176 674623 225178
rect 671797 225120 671802 225176
rect 671858 225120 674562 225176
rect 674618 225120 674623 225176
rect 671797 225118 674623 225120
rect 671797 225115 671863 225118
rect 674557 225115 674623 225118
rect 656709 225042 656775 225045
rect 670693 225042 670759 225045
rect 656709 225040 670759 225042
rect 656709 224984 656714 225040
rect 656770 224984 670698 225040
rect 670754 224984 670759 225040
rect 656709 224982 670759 224984
rect 656709 224979 656775 224982
rect 670693 224979 670759 224982
rect 42609 224906 42675 224909
rect 45829 224906 45895 224909
rect 42609 224904 45895 224906
rect 42609 224848 42614 224904
rect 42670 224848 45834 224904
rect 45890 224848 45895 224904
rect 42609 224846 45895 224848
rect 42609 224843 42675 224846
rect 45829 224843 45895 224846
rect 671470 224844 671476 224908
rect 671540 224906 671546 224908
rect 671705 224906 671771 224909
rect 671540 224904 671771 224906
rect 671540 224848 671710 224904
rect 671766 224848 671771 224904
rect 671540 224846 671771 224848
rect 671540 224844 671546 224846
rect 671705 224843 671771 224846
rect 72417 224770 72483 224773
rect 152733 224770 152799 224773
rect 72417 224768 152799 224770
rect 72417 224712 72422 224768
rect 72478 224712 152738 224768
rect 152794 224712 152799 224768
rect 72417 224710 152799 224712
rect 72417 224707 72483 224710
rect 152733 224707 152799 224710
rect 670877 224634 670943 224637
rect 672165 224634 672231 224637
rect 670877 224632 672231 224634
rect 670877 224576 670882 224632
rect 670938 224576 672170 224632
rect 672226 224576 672231 224632
rect 670877 224574 672231 224576
rect 670877 224571 670943 224574
rect 672165 224571 672231 224574
rect 66897 224498 66963 224501
rect 149789 224498 149855 224501
rect 66897 224496 149855 224498
rect 66897 224440 66902 224496
rect 66958 224440 149794 224496
rect 149850 224440 149855 224496
rect 66897 224438 149855 224440
rect 66897 224435 66963 224438
rect 149789 224435 149855 224438
rect 519537 224498 519603 224501
rect 606753 224498 606819 224501
rect 519537 224496 528570 224498
rect 519537 224440 519542 224496
rect 519598 224440 528570 224496
rect 519537 224438 528570 224440
rect 519537 224435 519603 224438
rect 59261 224226 59327 224229
rect 145005 224226 145071 224229
rect 59261 224224 145071 224226
rect 59261 224168 59266 224224
rect 59322 224168 145010 224224
rect 145066 224168 145071 224224
rect 59261 224166 145071 224168
rect 59261 224163 59327 224166
rect 145005 224163 145071 224166
rect 167545 224226 167611 224229
rect 199745 224226 199811 224229
rect 167545 224224 199811 224226
rect 167545 224168 167550 224224
rect 167606 224168 199750 224224
rect 199806 224168 199811 224224
rect 167545 224166 199811 224168
rect 167545 224163 167611 224166
rect 199745 224163 199811 224166
rect 512269 224226 512335 224229
rect 528510 224226 528570 224438
rect 601650 224496 606819 224498
rect 601650 224440 606758 224496
rect 606814 224440 606819 224496
rect 601650 224438 606819 224440
rect 601650 224226 601710 224438
rect 606753 224435 606819 224438
rect 656157 224498 656223 224501
rect 656157 224496 659670 224498
rect 656157 224440 656162 224496
rect 656218 224440 659670 224496
rect 656157 224438 659670 224440
rect 656157 224435 656223 224438
rect 659610 224362 659670 224438
rect 669037 224362 669103 224365
rect 659610 224360 669103 224362
rect 659610 224304 669042 224360
rect 669098 224304 669103 224360
rect 659610 224302 669103 224304
rect 669037 224299 669103 224302
rect 671654 224300 671660 224364
rect 671724 224362 671730 224364
rect 675569 224362 675635 224365
rect 671724 224360 675635 224362
rect 671724 224304 675574 224360
rect 675630 224304 675635 224360
rect 671724 224302 675635 224304
rect 671724 224300 671730 224302
rect 675569 224299 675635 224302
rect 617149 224226 617215 224229
rect 512269 224224 524430 224226
rect 512269 224168 512274 224224
rect 512330 224168 524430 224224
rect 512269 224166 524430 224168
rect 528510 224166 601710 224226
rect 606526 224224 617215 224226
rect 606526 224168 617154 224224
rect 617210 224168 617215 224224
rect 606526 224166 617215 224168
rect 512269 224163 512335 224166
rect 146845 223954 146911 223957
rect 176285 223954 176351 223957
rect 146845 223952 176351 223954
rect 146845 223896 146850 223952
rect 146906 223896 176290 223952
rect 176346 223896 176351 223952
rect 146845 223894 176351 223896
rect 146845 223891 146911 223894
rect 176285 223891 176351 223894
rect 496813 223954 496879 223957
rect 497825 223954 497891 223957
rect 519537 223954 519603 223957
rect 496813 223952 519603 223954
rect 496813 223896 496818 223952
rect 496874 223896 497830 223952
rect 497886 223896 519542 223952
rect 519598 223896 519603 223952
rect 496813 223894 519603 223896
rect 524370 223954 524430 224166
rect 606526 223954 606586 224166
rect 617149 224163 617215 224166
rect 524370 223894 606586 223954
rect 606753 223954 606819 223957
rect 630949 223954 631015 223957
rect 606753 223952 631015 223954
rect 606753 223896 606758 223952
rect 606814 223896 630954 223952
rect 631010 223896 631015 223952
rect 606753 223894 631015 223896
rect 496813 223891 496879 223894
rect 497825 223891 497891 223894
rect 519537 223891 519603 223894
rect 606753 223891 606819 223894
rect 630949 223891 631015 223894
rect 658181 223954 658247 223957
rect 670923 223954 670989 223957
rect 658181 223952 670989 223954
rect 658181 223896 658186 223952
rect 658242 223896 670928 223952
rect 670984 223896 670989 223952
rect 658181 223894 670989 223896
rect 658181 223891 658247 223894
rect 670923 223891 670989 223894
rect 672758 223892 672764 223956
rect 672828 223954 672834 223956
rect 673177 223954 673243 223957
rect 672828 223952 673243 223954
rect 672828 223896 673182 223952
rect 673238 223896 673243 223952
rect 672828 223894 673243 223896
rect 672828 223892 672834 223894
rect 673177 223891 673243 223894
rect 485865 223682 485931 223685
rect 486601 223682 486667 223685
rect 611629 223682 611695 223685
rect 485865 223680 611695 223682
rect 485865 223624 485870 223680
rect 485926 223624 486606 223680
rect 486662 223624 611634 223680
rect 611690 223624 611695 223680
rect 485865 223622 611695 223624
rect 485865 223619 485931 223622
rect 486601 223619 486667 223622
rect 611629 223619 611695 223622
rect 656893 223682 656959 223685
rect 670509 223682 670575 223685
rect 656893 223680 670575 223682
rect 656893 223624 656898 223680
rect 656954 223624 670514 223680
rect 670570 223624 670575 223680
rect 656893 223622 670575 223624
rect 656893 223619 656959 223622
rect 670509 223619 670575 223622
rect 683297 223546 683363 223549
rect 683284 223544 683363 223546
rect 683284 223488 683302 223544
rect 683358 223488 683363 223544
rect 683284 223486 683363 223488
rect 683297 223483 683363 223486
rect 92381 223410 92447 223413
rect 170765 223410 170831 223413
rect 92381 223408 170831 223410
rect 92381 223352 92386 223408
rect 92442 223352 170770 223408
rect 170826 223352 170831 223408
rect 92381 223350 170831 223352
rect 92381 223347 92447 223350
rect 170765 223347 170831 223350
rect 660205 223410 660271 223413
rect 675109 223410 675175 223413
rect 660205 223408 675175 223410
rect 660205 223352 660210 223408
rect 660266 223352 675114 223408
rect 675170 223352 675175 223408
rect 660205 223350 675175 223352
rect 660205 223347 660271 223350
rect 675109 223347 675175 223350
rect 71681 223138 71747 223141
rect 152089 223138 152155 223141
rect 71681 223136 152155 223138
rect 71681 223080 71686 223136
rect 71742 223080 152094 223136
rect 152150 223080 152155 223136
rect 71681 223078 152155 223080
rect 71681 223075 71747 223078
rect 152089 223075 152155 223078
rect 657537 223138 657603 223141
rect 667933 223138 667999 223141
rect 683665 223138 683731 223141
rect 657537 223136 667999 223138
rect 657537 223080 657542 223136
rect 657598 223080 667938 223136
rect 667994 223080 667999 223136
rect 657537 223078 667999 223080
rect 683652 223136 683731 223138
rect 683652 223080 683670 223136
rect 683726 223080 683731 223136
rect 683652 223078 683731 223080
rect 657537 223075 657603 223078
rect 667933 223075 667999 223078
rect 683665 223075 683731 223078
rect 28533 222866 28599 222869
rect 51717 222866 51783 222869
rect 28533 222864 51783 222866
rect 28533 222808 28538 222864
rect 28594 222808 51722 222864
rect 51778 222808 51783 222864
rect 28533 222806 51783 222808
rect 28533 222803 28599 222806
rect 51717 222803 51783 222806
rect 64781 222866 64847 222869
rect 146661 222866 146727 222869
rect 64781 222864 146727 222866
rect 64781 222808 64786 222864
rect 64842 222808 146666 222864
rect 146722 222808 146727 222864
rect 64781 222806 146727 222808
rect 64781 222803 64847 222806
rect 146661 222803 146727 222806
rect 151261 222866 151327 222869
rect 213913 222866 213979 222869
rect 151261 222864 213979 222866
rect 151261 222808 151266 222864
rect 151322 222808 213918 222864
rect 213974 222808 213979 222864
rect 151261 222806 213979 222808
rect 151261 222803 151327 222806
rect 213913 222803 213979 222806
rect 652385 222866 652451 222869
rect 673913 222866 673979 222869
rect 652385 222864 673979 222866
rect 652385 222808 652390 222864
rect 652446 222808 673918 222864
rect 673974 222808 673979 222864
rect 652385 222806 673979 222808
rect 652385 222803 652451 222806
rect 673913 222803 673979 222806
rect 683481 222730 683547 222733
rect 683468 222728 683547 222730
rect 683468 222672 683486 222728
rect 683542 222672 683547 222728
rect 683468 222670 683547 222672
rect 683481 222667 683547 222670
rect 482737 222322 482803 222325
rect 593965 222322 594031 222325
rect 482737 222320 594031 222322
rect 482737 222264 482742 222320
rect 482798 222264 593970 222320
rect 594026 222264 594031 222320
rect 482737 222262 594031 222264
rect 482737 222259 482803 222262
rect 593965 222259 594031 222262
rect 673126 222260 673132 222324
rect 673196 222322 673202 222324
rect 673196 222262 676292 222322
rect 673196 222260 673202 222262
rect 108941 222050 109007 222053
rect 183645 222050 183711 222053
rect 108941 222048 183711 222050
rect 108941 221992 108946 222048
rect 109002 221992 183650 222048
rect 183706 221992 183711 222048
rect 108941 221990 183711 221992
rect 108941 221987 109007 221990
rect 183645 221987 183711 221990
rect 523033 222050 523099 222053
rect 523401 222050 523467 222053
rect 532693 222050 532759 222053
rect 523033 222048 532759 222050
rect 523033 221992 523038 222048
rect 523094 221992 523406 222048
rect 523462 221992 532698 222048
rect 532754 221992 532759 222048
rect 523033 221990 532759 221992
rect 523033 221987 523099 221990
rect 523401 221987 523467 221990
rect 532693 221987 532759 221990
rect 532877 222050 532943 222053
rect 600681 222050 600747 222053
rect 532877 222048 600747 222050
rect 532877 221992 532882 222048
rect 532938 221992 600686 222048
rect 600742 221992 600747 222048
rect 532877 221990 600747 221992
rect 532877 221987 532943 221990
rect 600681 221987 600747 221990
rect 670785 222050 670851 222053
rect 673729 222050 673795 222053
rect 670785 222048 673795 222050
rect 670785 221992 670790 222048
rect 670846 221992 673734 222048
rect 673790 221992 673795 222048
rect 670785 221990 673795 221992
rect 670785 221987 670851 221990
rect 673729 221987 673795 221990
rect 669037 221914 669103 221917
rect 669037 221912 669882 221914
rect 669037 221856 669042 221912
rect 669098 221856 669882 221912
rect 669037 221854 669882 221856
rect 669037 221851 669103 221854
rect 97717 221778 97783 221781
rect 172697 221778 172763 221781
rect 97717 221776 172763 221778
rect 97717 221720 97722 221776
rect 97778 221720 172702 221776
rect 172758 221720 172763 221776
rect 97717 221718 172763 221720
rect 97717 221715 97783 221718
rect 172697 221715 172763 221718
rect 513465 221778 513531 221781
rect 599025 221778 599091 221781
rect 513465 221776 599091 221778
rect 513465 221720 513470 221776
rect 513526 221720 599030 221776
rect 599086 221720 599091 221776
rect 513465 221718 599091 221720
rect 669822 221778 669882 221854
rect 676170 221854 676292 221914
rect 676170 221778 676230 221854
rect 669822 221718 676230 221778
rect 513465 221715 513531 221718
rect 599025 221715 599091 221718
rect 659610 221582 666570 221642
rect 95693 221506 95759 221509
rect 172973 221506 173039 221509
rect 95693 221504 173039 221506
rect 95693 221448 95698 221504
rect 95754 221448 172978 221504
rect 173034 221448 173039 221504
rect 95693 221446 173039 221448
rect 95693 221443 95759 221446
rect 172973 221443 173039 221446
rect 518433 221506 518499 221509
rect 532877 221506 532943 221509
rect 518433 221504 532943 221506
rect 518433 221448 518438 221504
rect 518494 221448 532882 221504
rect 532938 221448 532943 221504
rect 518433 221446 532943 221448
rect 518433 221443 518499 221446
rect 532877 221443 532943 221446
rect 533061 221506 533127 221509
rect 601969 221506 602035 221509
rect 533061 221504 602035 221506
rect 533061 221448 533066 221504
rect 533122 221448 601974 221504
rect 602030 221448 602035 221504
rect 533061 221446 602035 221448
rect 533061 221443 533127 221446
rect 601969 221443 602035 221446
rect 649717 221506 649783 221509
rect 659610 221506 659670 221582
rect 649717 221504 659670 221506
rect 649717 221448 649722 221504
rect 649778 221448 659670 221504
rect 649717 221446 659670 221448
rect 666510 221506 666570 221582
rect 673361 221506 673427 221509
rect 683113 221506 683179 221509
rect 666510 221504 673427 221506
rect 666510 221448 673366 221504
rect 673422 221448 673427 221504
rect 666510 221446 673427 221448
rect 683100 221504 683179 221506
rect 683100 221448 683118 221504
rect 683174 221448 683179 221504
rect 683100 221446 683179 221448
rect 649717 221443 649783 221446
rect 673361 221443 673427 221446
rect 683113 221443 683179 221446
rect 170581 221234 170647 221237
rect 229553 221234 229619 221237
rect 170581 221232 229619 221234
rect 170581 221176 170586 221232
rect 170642 221176 229558 221232
rect 229614 221176 229619 221232
rect 170581 221174 229619 221176
rect 170581 221171 170647 221174
rect 229553 221171 229619 221174
rect 515765 221234 515831 221237
rect 600865 221234 600931 221237
rect 515765 221232 600931 221234
rect 515765 221176 515770 221232
rect 515826 221176 600870 221232
rect 600926 221176 600931 221232
rect 515765 221174 600931 221176
rect 515765 221171 515831 221174
rect 600865 221171 600931 221174
rect 652937 221234 653003 221237
rect 667933 221234 667999 221237
rect 673545 221234 673611 221237
rect 652937 221232 667999 221234
rect 652937 221176 652942 221232
rect 652998 221176 667938 221232
rect 667994 221176 667999 221232
rect 652937 221174 667999 221176
rect 652937 221171 653003 221174
rect 667933 221171 667999 221174
rect 669638 221232 673611 221234
rect 669638 221176 673550 221232
rect 673606 221176 673611 221232
rect 669638 221174 673611 221176
rect 510705 220962 510771 220965
rect 599209 220962 599275 220965
rect 510705 220960 599275 220962
rect 510705 220904 510710 220960
rect 510766 220904 599214 220960
rect 599270 220904 599275 220960
rect 510705 220902 599275 220904
rect 510705 220899 510771 220902
rect 599209 220899 599275 220902
rect 665449 220962 665515 220965
rect 669638 220962 669698 221174
rect 673545 221171 673611 221174
rect 676170 221038 676292 221098
rect 665449 220960 669698 220962
rect 665449 220904 665454 220960
rect 665510 220904 669698 220960
rect 665449 220902 669698 220904
rect 665449 220899 665515 220902
rect 669814 220900 669820 220964
rect 669884 220962 669890 220964
rect 670601 220962 670667 220965
rect 676170 220962 676230 221038
rect 669884 220960 670667 220962
rect 669884 220904 670606 220960
rect 670662 220904 670667 220960
rect 669884 220902 670667 220904
rect 669884 220900 669890 220902
rect 670601 220899 670667 220902
rect 670926 220902 676230 220962
rect 147581 220690 147647 220693
rect 211337 220690 211403 220693
rect 147581 220688 211403 220690
rect 147581 220632 147586 220688
rect 147642 220632 211342 220688
rect 211398 220632 211403 220688
rect 147581 220630 211403 220632
rect 147581 220627 147647 220630
rect 211337 220627 211403 220630
rect 653121 220690 653187 220693
rect 670366 220690 670372 220692
rect 653121 220688 670372 220690
rect 653121 220632 653126 220688
rect 653182 220632 670372 220688
rect 653121 220630 670372 220632
rect 653121 220627 653187 220630
rect 670366 220628 670372 220630
rect 670436 220628 670442 220692
rect 670601 220690 670667 220693
rect 670926 220690 670986 220902
rect 670601 220688 670986 220690
rect 670601 220632 670606 220688
rect 670662 220632 670986 220688
rect 670601 220630 670986 220632
rect 670601 220627 670667 220630
rect 671102 220628 671108 220692
rect 671172 220690 671178 220692
rect 674373 220690 674439 220693
rect 671172 220688 674439 220690
rect 671172 220632 674378 220688
rect 674434 220632 674439 220688
rect 671172 220630 674439 220632
rect 671172 220628 671178 220630
rect 674373 220627 674439 220630
rect 680997 220690 681063 220693
rect 680997 220688 681076 220690
rect 680997 220632 681002 220688
rect 681058 220632 681076 220688
rect 680997 220630 681076 220632
rect 680997 220627 681063 220630
rect 518801 220554 518867 220557
rect 617701 220554 617767 220557
rect 518801 220552 617767 220554
rect 518801 220496 518806 220552
rect 518862 220496 617706 220552
rect 617762 220496 617767 220552
rect 518801 220494 617767 220496
rect 518801 220491 518867 220494
rect 617701 220491 617767 220494
rect 124673 220418 124739 220421
rect 193305 220418 193371 220421
rect 124673 220416 193371 220418
rect 124673 220360 124678 220416
rect 124734 220360 193310 220416
rect 193366 220360 193371 220416
rect 124673 220358 193371 220360
rect 124673 220355 124739 220358
rect 193305 220355 193371 220358
rect 644749 220418 644815 220421
rect 671838 220418 671844 220420
rect 644749 220416 671844 220418
rect 644749 220360 644754 220416
rect 644810 220360 671844 220416
rect 644749 220358 671844 220360
rect 644749 220355 644815 220358
rect 671838 220356 671844 220358
rect 671908 220356 671914 220420
rect 673453 220418 673519 220421
rect 674373 220418 674439 220421
rect 673453 220416 674439 220418
rect 673453 220360 673458 220416
rect 673514 220360 674378 220416
rect 674434 220360 674439 220416
rect 673453 220358 674439 220360
rect 673453 220355 673519 220358
rect 674373 220355 674439 220358
rect 507761 220282 507827 220285
rect 528553 220282 528619 220285
rect 507761 220280 528619 220282
rect 507761 220224 507766 220280
rect 507822 220224 528558 220280
rect 528614 220224 528619 220280
rect 507761 220222 528619 220224
rect 507761 220219 507827 220222
rect 528553 220219 528619 220222
rect 528737 220282 528803 220285
rect 534073 220282 534139 220285
rect 528737 220280 534139 220282
rect 528737 220224 528742 220280
rect 528798 220224 534078 220280
rect 534134 220224 534139 220280
rect 528737 220222 534139 220224
rect 528737 220219 528803 220222
rect 534073 220219 534139 220222
rect 534257 220282 534323 220285
rect 543733 220282 543799 220285
rect 534257 220280 543799 220282
rect 534257 220224 534262 220280
rect 534318 220224 543738 220280
rect 543794 220224 543799 220280
rect 534257 220222 543799 220224
rect 534257 220219 534323 220222
rect 543733 220219 543799 220222
rect 543917 220282 543983 220285
rect 553117 220282 553183 220285
rect 543917 220280 553183 220282
rect 543917 220224 543922 220280
rect 543978 220224 553122 220280
rect 553178 220224 553183 220280
rect 543917 220222 553183 220224
rect 543917 220219 543983 220222
rect 553117 220219 553183 220222
rect 553301 220282 553367 220285
rect 604637 220282 604703 220285
rect 615677 220282 615743 220285
rect 553301 220280 604703 220282
rect 553301 220224 553306 220280
rect 553362 220224 604642 220280
rect 604698 220224 604703 220280
rect 553301 220222 604703 220224
rect 553301 220219 553367 220222
rect 604637 220219 604703 220222
rect 611310 220280 615743 220282
rect 611310 220224 615682 220280
rect 615738 220224 615743 220280
rect 611310 220222 615743 220224
rect 118049 220146 118115 220149
rect 187877 220146 187943 220149
rect 118049 220144 187943 220146
rect 118049 220088 118054 220144
rect 118110 220088 187882 220144
rect 187938 220088 187943 220144
rect 118049 220086 187943 220088
rect 118049 220083 118115 220086
rect 187877 220083 187943 220086
rect 505921 220010 505987 220013
rect 582373 220010 582439 220013
rect 505921 220008 582439 220010
rect 505921 219952 505926 220008
rect 505982 219952 582378 220008
rect 582434 219952 582439 220008
rect 505921 219950 582439 219952
rect 505921 219947 505987 219950
rect 582373 219947 582439 219950
rect 582557 220010 582623 220013
rect 611310 220010 611370 220222
rect 615677 220219 615743 220222
rect 676170 220222 676292 220282
rect 670785 220146 670851 220149
rect 676170 220146 676230 220222
rect 670785 220144 676230 220146
rect 670785 220088 670790 220144
rect 670846 220088 676230 220144
rect 670785 220086 676230 220088
rect 670785 220083 670851 220086
rect 582557 220008 611370 220010
rect 582557 219952 582562 220008
rect 582618 219952 611370 220008
rect 582557 219950 611370 219952
rect 582557 219947 582623 219950
rect 648613 219874 648679 219877
rect 673453 219874 673519 219877
rect 648613 219872 673519 219874
rect 648613 219816 648618 219872
rect 648674 219816 673458 219872
rect 673514 219816 673519 219872
rect 648613 219814 673519 219816
rect 648613 219811 648679 219814
rect 673453 219811 673519 219814
rect 684493 219874 684559 219877
rect 684493 219872 684572 219874
rect 684493 219816 684498 219872
rect 684554 219816 684572 219872
rect 684493 219814 684572 219816
rect 684493 219811 684559 219814
rect 501321 219738 501387 219741
rect 582373 219738 582439 219741
rect 594793 219738 594859 219741
rect 501321 219736 582439 219738
rect 501321 219680 501326 219736
rect 501382 219680 582378 219736
rect 582434 219680 582439 219736
rect 501321 219678 582439 219680
rect 501321 219675 501387 219678
rect 582373 219675 582439 219678
rect 582790 219736 594859 219738
rect 582790 219680 594798 219736
rect 594854 219680 594859 219736
rect 582790 219678 594859 219680
rect 582790 219602 582850 219678
rect 594793 219675 594859 219678
rect 582606 219542 582850 219602
rect 488993 219466 489059 219469
rect 582606 219466 582666 219542
rect 488993 219464 582666 219466
rect 488993 219408 488998 219464
rect 489054 219408 582666 219464
rect 488993 219406 582666 219408
rect 583109 219466 583175 219469
rect 618805 219466 618871 219469
rect 583109 219464 618871 219466
rect 583109 219408 583114 219464
rect 583170 219408 618810 219464
rect 618866 219408 618871 219464
rect 583109 219406 618871 219408
rect 488993 219403 489059 219406
rect 583109 219403 583175 219406
rect 618805 219403 618871 219406
rect 667841 219466 667907 219469
rect 667841 219464 676292 219466
rect 667841 219408 667846 219464
rect 667902 219408 676292 219464
rect 667841 219406 676292 219408
rect 667841 219403 667907 219406
rect 490741 219194 490807 219197
rect 494789 219194 494855 219197
rect 500217 219194 500283 219197
rect 490741 219192 494530 219194
rect 490741 219136 490746 219192
rect 490802 219136 494530 219192
rect 490741 219134 494530 219136
rect 490741 219131 490807 219134
rect 77201 218922 77267 218925
rect 157517 218922 157583 218925
rect 77201 218920 157583 218922
rect 77201 218864 77206 218920
rect 77262 218864 157522 218920
rect 157578 218864 157583 218920
rect 77201 218862 157583 218864
rect 77201 218859 77267 218862
rect 157517 218859 157583 218862
rect 490557 218922 490623 218925
rect 491201 218922 491267 218925
rect 494470 218922 494530 219134
rect 494789 219192 500283 219194
rect 494789 219136 494794 219192
rect 494850 219136 500222 219192
rect 500278 219136 500283 219192
rect 494789 219134 500283 219136
rect 494789 219131 494855 219134
rect 500217 219131 500283 219134
rect 500401 219194 500467 219197
rect 504541 219194 504607 219197
rect 500401 219192 504607 219194
rect 500401 219136 500406 219192
rect 500462 219136 504546 219192
rect 504602 219136 504607 219192
rect 500401 219134 504607 219136
rect 500401 219131 500467 219134
rect 504541 219131 504607 219134
rect 504725 219194 504791 219197
rect 506289 219194 506355 219197
rect 524045 219194 524111 219197
rect 504725 219192 505018 219194
rect 504725 219136 504730 219192
rect 504786 219136 505018 219192
rect 504725 219134 505018 219136
rect 504725 219131 504791 219134
rect 504725 218922 504791 218925
rect 490557 218920 494346 218922
rect 490557 218864 490562 218920
rect 490618 218864 491206 218920
rect 491262 218864 494346 218920
rect 490557 218862 494346 218864
rect 494470 218920 504791 218922
rect 494470 218864 504730 218920
rect 504786 218864 504791 218920
rect 494470 218862 504791 218864
rect 504958 218922 505018 219134
rect 506289 219192 524111 219194
rect 506289 219136 506294 219192
rect 506350 219136 524050 219192
rect 524106 219136 524111 219192
rect 506289 219134 524111 219136
rect 506289 219131 506355 219134
rect 524045 219131 524111 219134
rect 524229 219194 524295 219197
rect 528277 219194 528343 219197
rect 524229 219192 528343 219194
rect 524229 219136 524234 219192
rect 524290 219136 528282 219192
rect 528338 219136 528343 219192
rect 524229 219134 528343 219136
rect 524229 219131 524295 219134
rect 528277 219131 528343 219134
rect 528461 219194 528527 219197
rect 534257 219194 534323 219197
rect 528461 219192 534323 219194
rect 528461 219136 528466 219192
rect 528522 219136 534262 219192
rect 534318 219136 534323 219192
rect 528461 219134 534323 219136
rect 528461 219131 528527 219134
rect 534257 219131 534323 219134
rect 534441 219194 534507 219197
rect 543457 219194 543523 219197
rect 534441 219192 543523 219194
rect 534441 219136 534446 219192
rect 534502 219136 543462 219192
rect 543518 219136 543523 219192
rect 534441 219134 543523 219136
rect 534441 219131 534507 219134
rect 543457 219131 543523 219134
rect 543641 219194 543707 219197
rect 543917 219194 543983 219197
rect 543641 219192 543983 219194
rect 543641 219136 543646 219192
rect 543702 219136 543922 219192
rect 543978 219136 543983 219192
rect 543641 219134 543983 219136
rect 543641 219131 543707 219134
rect 543917 219131 543983 219134
rect 544101 219194 544167 219197
rect 552565 219194 552631 219197
rect 544101 219192 552631 219194
rect 544101 219136 544106 219192
rect 544162 219136 552570 219192
rect 552626 219136 552631 219192
rect 544101 219134 552631 219136
rect 544101 219131 544167 219134
rect 552565 219131 552631 219134
rect 552933 219194 552999 219197
rect 623773 219194 623839 219197
rect 552933 219192 623839 219194
rect 552933 219136 552938 219192
rect 552994 219136 623778 219192
rect 623834 219136 623839 219192
rect 552933 219134 623839 219136
rect 552933 219131 552999 219134
rect 623773 219131 623839 219134
rect 651281 219194 651347 219197
rect 673177 219194 673243 219197
rect 651281 219192 673243 219194
rect 651281 219136 651286 219192
rect 651342 219136 673182 219192
rect 673238 219136 673243 219192
rect 651281 219134 673243 219136
rect 651281 219131 651347 219134
rect 673177 219131 673243 219134
rect 679617 219058 679683 219061
rect 679604 219056 679683 219058
rect 679604 219000 679622 219056
rect 679678 219000 679683 219056
rect 679604 218998 679683 219000
rect 679617 218995 679683 218998
rect 553485 218922 553551 218925
rect 504958 218920 553551 218922
rect 504958 218864 553490 218920
rect 553546 218864 553551 218920
rect 504958 218862 553551 218864
rect 490557 218859 490623 218862
rect 491201 218859 491267 218862
rect 70853 218650 70919 218653
rect 153469 218650 153535 218653
rect 70853 218648 153535 218650
rect 70853 218592 70858 218648
rect 70914 218592 153474 218648
rect 153530 218592 153535 218648
rect 70853 218590 153535 218592
rect 70853 218587 70919 218590
rect 153469 218587 153535 218590
rect 166901 218650 166967 218653
rect 206277 218650 206343 218653
rect 166901 218648 206343 218650
rect 166901 218592 166906 218648
rect 166962 218592 206282 218648
rect 206338 218592 206343 218648
rect 166901 218590 206343 218592
rect 166901 218587 166967 218590
rect 206277 218587 206343 218590
rect 491937 218650 492003 218653
rect 494286 218650 494346 218862
rect 504725 218859 504791 218862
rect 553485 218859 553551 218862
rect 553853 218922 553919 218925
rect 562777 218922 562843 218925
rect 553853 218920 562843 218922
rect 553853 218864 553858 218920
rect 553914 218864 562782 218920
rect 562838 218864 562843 218920
rect 553853 218862 562843 218864
rect 553853 218859 553919 218862
rect 562777 218859 562843 218862
rect 563053 218922 563119 218925
rect 595897 218922 595963 218925
rect 563053 218920 595963 218922
rect 563053 218864 563058 218920
rect 563114 218864 595902 218920
rect 595958 218864 595963 218920
rect 563053 218862 595963 218864
rect 563053 218859 563119 218862
rect 595897 218859 595963 218862
rect 596081 218922 596147 218925
rect 630673 218922 630739 218925
rect 596081 218920 630739 218922
rect 596081 218864 596086 218920
rect 596142 218864 630678 218920
rect 630734 218864 630739 218920
rect 596081 218862 630739 218864
rect 596081 218859 596147 218862
rect 630673 218859 630739 218862
rect 643829 218922 643895 218925
rect 675569 218922 675635 218925
rect 643829 218920 675635 218922
rect 643829 218864 643834 218920
rect 643890 218864 675574 218920
rect 675630 218864 675635 218920
rect 643829 218862 675635 218864
rect 643829 218859 643895 218862
rect 675569 218859 675635 218862
rect 500033 218650 500099 218653
rect 491937 218648 494162 218650
rect 491937 218592 491942 218648
rect 491998 218592 494162 218648
rect 491937 218590 494162 218592
rect 494286 218648 500099 218650
rect 494286 218592 500038 218648
rect 500094 218592 500099 218648
rect 494286 218590 500099 218592
rect 491937 218587 492003 218590
rect 492673 218378 492739 218381
rect 493910 218378 493916 218380
rect 492673 218376 493916 218378
rect 492673 218320 492678 218376
rect 492734 218320 493916 218376
rect 492673 218318 493916 218320
rect 492673 218315 492739 218318
rect 493910 218316 493916 218318
rect 493980 218316 493986 218380
rect 494102 218378 494162 218590
rect 500033 218587 500099 218590
rect 500217 218650 500283 218653
rect 514753 218650 514819 218653
rect 500217 218648 514819 218650
rect 500217 218592 500222 218648
rect 500278 218592 514758 218648
rect 514814 218592 514819 218648
rect 500217 218590 514819 218592
rect 500217 218587 500283 218590
rect 514753 218587 514819 218590
rect 514937 218650 515003 218653
rect 523769 218650 523835 218653
rect 514937 218648 523835 218650
rect 514937 218592 514942 218648
rect 514998 218592 523774 218648
rect 523830 218592 523835 218648
rect 514937 218590 523835 218592
rect 514937 218587 515003 218590
rect 523769 218587 523835 218590
rect 524229 218650 524295 218653
rect 528277 218650 528343 218653
rect 524229 218648 528343 218650
rect 524229 218592 524234 218648
rect 524290 218592 528282 218648
rect 528338 218592 528343 218648
rect 524229 218590 528343 218592
rect 524229 218587 524295 218590
rect 528277 218587 528343 218590
rect 528461 218650 528527 218653
rect 528645 218650 528711 218653
rect 528461 218648 528711 218650
rect 528461 218592 528466 218648
rect 528522 218592 528650 218648
rect 528706 218592 528711 218648
rect 528461 218590 528711 218592
rect 528461 218587 528527 218590
rect 528645 218587 528711 218590
rect 529013 218650 529079 218653
rect 534073 218650 534139 218653
rect 529013 218648 534139 218650
rect 529013 218592 529018 218648
rect 529074 218592 534078 218648
rect 534134 218592 534139 218648
rect 529013 218590 534139 218592
rect 529013 218587 529079 218590
rect 534073 218587 534139 218590
rect 534257 218650 534323 218653
rect 543457 218650 543523 218653
rect 534257 218648 543523 218650
rect 534257 218592 534262 218648
rect 534318 218592 543462 218648
rect 543518 218592 543523 218648
rect 534257 218590 543523 218592
rect 534257 218587 534323 218590
rect 543457 218587 543523 218590
rect 543917 218650 543983 218653
rect 553117 218650 553183 218653
rect 543917 218648 553183 218650
rect 543917 218592 543922 218648
rect 543978 218592 553122 218648
rect 553178 218592 553183 218648
rect 543917 218590 553183 218592
rect 543917 218587 543983 218590
rect 553117 218587 553183 218590
rect 553301 218650 553367 218653
rect 553526 218650 553532 218652
rect 553301 218648 553532 218650
rect 553301 218592 553306 218648
rect 553362 218592 553532 218648
rect 553301 218590 553532 218592
rect 553301 218587 553367 218590
rect 553526 218588 553532 218590
rect 553596 218588 553602 218652
rect 553853 218650 553919 218653
rect 605097 218650 605163 218653
rect 622945 218650 623011 218653
rect 553853 218648 605163 218650
rect 553853 218592 553858 218648
rect 553914 218592 605102 218648
rect 605158 218592 605163 218648
rect 553853 218590 605163 218592
rect 553853 218587 553919 218590
rect 605097 218587 605163 218590
rect 611310 218648 623011 218650
rect 611310 218592 622950 218648
rect 623006 218592 623011 218648
rect 611310 218590 623011 218592
rect 505042 218378 505048 218380
rect 494102 218318 505048 218378
rect 505042 218316 505048 218318
rect 505112 218316 505118 218380
rect 505277 218378 505343 218381
rect 563053 218378 563119 218381
rect 505277 218376 563119 218378
rect 505277 218320 505282 218376
rect 505338 218320 563058 218376
rect 563114 218320 563119 218376
rect 505277 218318 563119 218320
rect 505277 218315 505343 218318
rect 563053 218315 563119 218318
rect 563237 218378 563303 218381
rect 572437 218378 572503 218381
rect 563237 218376 572503 218378
rect 563237 218320 563242 218376
rect 563298 218320 572442 218376
rect 572498 218320 572503 218376
rect 563237 218318 572503 218320
rect 563237 218315 563303 218318
rect 572437 218315 572503 218318
rect 572662 218316 572668 218380
rect 572732 218378 572738 218380
rect 576577 218378 576643 218381
rect 572732 218376 576643 218378
rect 572732 218320 576582 218376
rect 576638 218320 576643 218376
rect 572732 218318 576643 218320
rect 572732 218316 572738 218318
rect 576577 218315 576643 218318
rect 576761 218378 576827 218381
rect 611310 218378 611370 218590
rect 622945 218587 623011 218590
rect 640609 218650 640675 218653
rect 640609 218648 659670 218650
rect 640609 218592 640614 218648
rect 640670 218592 659670 218648
rect 640609 218590 659670 218592
rect 640609 218587 640675 218590
rect 576761 218376 611370 218378
rect 576761 218320 576766 218376
rect 576822 218320 611370 218376
rect 576761 218318 611370 218320
rect 659610 218378 659670 218590
rect 675518 218588 675524 218652
rect 675588 218650 675594 218652
rect 675588 218590 676292 218650
rect 675588 218588 675594 218590
rect 676029 218378 676095 218381
rect 659610 218376 676095 218378
rect 659610 218320 676034 218376
rect 676090 218320 676095 218376
rect 659610 218318 676095 218320
rect 576761 218315 576827 218318
rect 676029 218315 676095 218318
rect 676170 218182 676292 218242
rect 487797 218106 487863 218109
rect 629385 218106 629451 218109
rect 487797 218104 629451 218106
rect 487797 218048 487802 218104
rect 487858 218048 629390 218104
rect 629446 218048 629451 218104
rect 487797 218046 629451 218048
rect 487797 218043 487863 218046
rect 629385 218043 629451 218046
rect 667013 218106 667079 218109
rect 674649 218106 674715 218109
rect 667013 218104 674715 218106
rect 667013 218048 667018 218104
rect 667074 218048 674654 218104
rect 674710 218048 674715 218104
rect 667013 218046 674715 218048
rect 667013 218043 667079 218046
rect 674649 218043 674715 218046
rect 675702 218044 675708 218108
rect 675772 218106 675778 218108
rect 676170 218106 676230 218182
rect 675772 218046 676230 218106
rect 675772 218044 675778 218046
rect 508865 217834 508931 217837
rect 553485 217834 553551 217837
rect 508865 217832 553551 217834
rect 508865 217776 508870 217832
rect 508926 217776 553490 217832
rect 553546 217776 553551 217832
rect 508865 217774 553551 217776
rect 508865 217771 508931 217774
rect 553485 217771 553551 217774
rect 553710 217772 553716 217836
rect 553780 217834 553786 217836
rect 562542 217834 562548 217836
rect 553780 217774 562548 217834
rect 553780 217772 553786 217774
rect 562542 217772 562548 217774
rect 562612 217772 562618 217836
rect 562869 217834 562935 217837
rect 608961 217834 609027 217837
rect 562869 217832 609027 217834
rect 562869 217776 562874 217832
rect 562930 217776 608966 217832
rect 609022 217776 609027 217832
rect 562869 217774 609027 217776
rect 562869 217771 562935 217774
rect 608961 217771 609027 217774
rect 639965 217834 640031 217837
rect 674966 217834 674972 217836
rect 639965 217832 674972 217834
rect 639965 217776 639970 217832
rect 640026 217776 674972 217832
rect 639965 217774 674972 217776
rect 639965 217771 640031 217774
rect 674966 217772 674972 217774
rect 675036 217772 675042 217836
rect 676029 217834 676095 217837
rect 676029 217832 676292 217834
rect 676029 217776 676034 217832
rect 676090 217776 676292 217832
rect 676029 217774 676292 217776
rect 676029 217771 676095 217774
rect 493869 217700 493935 217701
rect 493869 217698 493916 217700
rect 493824 217696 493916 217698
rect 493824 217640 493874 217696
rect 493824 217638 493916 217640
rect 493869 217636 493916 217638
rect 493980 217636 493986 217700
rect 493869 217635 493935 217636
rect 500217 217562 500283 217565
rect 553209 217562 553275 217565
rect 500217 217560 553275 217562
rect 500217 217504 500222 217560
rect 500278 217504 553214 217560
rect 553270 217504 553275 217560
rect 500217 217502 553275 217504
rect 500217 217499 500283 217502
rect 553209 217499 553275 217502
rect 554221 217562 554287 217565
rect 576577 217562 576643 217565
rect 554221 217560 576643 217562
rect 554221 217504 554226 217560
rect 554282 217504 576582 217560
rect 576638 217504 576643 217560
rect 554221 217502 576643 217504
rect 554221 217499 554287 217502
rect 576577 217499 576643 217502
rect 576761 217562 576827 217565
rect 610065 217562 610131 217565
rect 576761 217560 610131 217562
rect 576761 217504 576766 217560
rect 576822 217504 610070 217560
rect 610126 217504 610131 217560
rect 576761 217502 610131 217504
rect 576761 217499 576827 217502
rect 610065 217499 610131 217502
rect 644565 217562 644631 217565
rect 674833 217562 674899 217565
rect 644565 217560 674899 217562
rect 644565 217504 644570 217560
rect 644626 217504 674838 217560
rect 674894 217504 674899 217560
rect 644565 217502 674899 217504
rect 644565 217499 644631 217502
rect 674833 217499 674899 217502
rect 553350 217366 553778 217426
rect 498837 217290 498903 217293
rect 553350 217290 553410 217366
rect 498837 217288 553410 217290
rect 498837 217232 498842 217288
rect 498898 217232 553410 217288
rect 498837 217230 553410 217232
rect 553718 217290 553778 217366
rect 676170 217366 676292 217426
rect 563053 217290 563119 217293
rect 553718 217288 563119 217290
rect 553718 217232 563058 217288
rect 563114 217232 563119 217288
rect 553718 217230 563119 217232
rect 498837 217227 498903 217230
rect 563053 217227 563119 217230
rect 563237 217290 563303 217293
rect 572345 217290 572411 217293
rect 563237 217288 572411 217290
rect 563237 217232 563242 217288
rect 563298 217232 572350 217288
rect 572406 217232 572411 217288
rect 563237 217230 572411 217232
rect 563237 217227 563303 217230
rect 572345 217227 572411 217230
rect 572529 217290 572595 217293
rect 575381 217290 575447 217293
rect 572529 217288 575447 217290
rect 572529 217232 572534 217288
rect 572590 217232 575386 217288
rect 575442 217232 575447 217288
rect 572529 217230 575447 217232
rect 572529 217227 572595 217230
rect 575381 217227 575447 217230
rect 576802 217228 576808 217292
rect 576872 217290 576878 217292
rect 591757 217290 591823 217293
rect 576872 217288 591823 217290
rect 576872 217232 591762 217288
rect 591818 217232 591823 217288
rect 576872 217230 591823 217232
rect 576872 217228 576878 217230
rect 591757 217227 591823 217230
rect 591941 217290 592007 217293
rect 591941 217288 596190 217290
rect 591941 217232 591946 217288
rect 592002 217232 596190 217288
rect 591941 217230 596190 217232
rect 591941 217227 592007 217230
rect 596130 217154 596190 217230
rect 666318 217228 666324 217292
rect 666388 217290 666394 217292
rect 676170 217290 676230 217366
rect 666388 217230 676230 217290
rect 666388 217228 666394 217230
rect 597553 217154 597619 217157
rect 596130 217152 597619 217154
rect 596130 217096 597558 217152
rect 597614 217096 597619 217152
rect 596130 217094 597619 217096
rect 597553 217091 597619 217094
rect 503713 217018 503779 217021
rect 508865 217018 508931 217021
rect 503713 217016 508931 217018
rect 503713 216960 503718 217016
rect 503774 216960 508870 217016
rect 508926 216960 508931 217016
rect 503713 216958 508931 216960
rect 503713 216955 503779 216958
rect 508865 216955 508931 216958
rect 553485 217018 553551 217021
rect 571701 217018 571767 217021
rect 553485 217016 571767 217018
rect 553485 216960 553490 217016
rect 553546 216960 571706 217016
rect 571762 216960 571767 217016
rect 553485 216958 571767 216960
rect 553485 216955 553551 216958
rect 571701 216955 571767 216958
rect 576945 217018 577011 217021
rect 591573 217018 591639 217021
rect 576945 217016 591639 217018
rect 576945 216960 576950 217016
rect 577006 216960 591578 217016
rect 591634 216960 591639 217016
rect 576945 216958 591639 216960
rect 576945 216955 577011 216958
rect 591573 216955 591639 216958
rect 591941 217018 592007 217021
rect 656525 217018 656591 217021
rect 672165 217018 672231 217021
rect 591941 217016 596098 217018
rect 591941 216960 591946 217016
rect 592002 216960 596098 217016
rect 591941 216958 596098 216960
rect 591941 216955 592007 216958
rect 596038 216882 596098 216958
rect 656525 217016 672231 217018
rect 656525 216960 656530 217016
rect 656586 216960 672170 217016
rect 672226 216960 672231 217016
rect 656525 216958 672231 216960
rect 656525 216955 656591 216958
rect 672165 216955 672231 216958
rect 675702 216956 675708 217020
rect 675772 217018 675778 217020
rect 675772 216958 676292 217018
rect 675772 216956 675778 216958
rect 627821 216882 627887 216885
rect 596038 216880 627887 216882
rect 596038 216824 627826 216880
rect 627882 216824 627887 216880
rect 596038 216822 627887 216824
rect 627821 216819 627887 216822
rect 577129 216746 577195 216749
rect 582373 216746 582439 216749
rect 577129 216744 582439 216746
rect 577129 216688 577134 216744
rect 577190 216688 582378 216744
rect 582434 216688 582439 216744
rect 577129 216686 582439 216688
rect 577129 216683 577195 216686
rect 582373 216683 582439 216686
rect 582557 216746 582623 216749
rect 582557 216744 595914 216746
rect 582557 216688 582562 216744
rect 582618 216688 595914 216744
rect 582557 216686 595914 216688
rect 582557 216683 582623 216686
rect 595854 216610 595914 216686
rect 596265 216610 596331 216613
rect 595854 216608 596331 216610
rect 595854 216552 596270 216608
rect 596326 216552 596331 216608
rect 595854 216550 596331 216552
rect 596265 216547 596331 216550
rect 674557 216610 674623 216613
rect 674557 216608 676292 216610
rect 674557 216552 674562 216608
rect 674618 216552 676292 216608
rect 674557 216550 676292 216552
rect 674557 216547 674623 216550
rect 575381 216474 575447 216477
rect 591757 216474 591823 216477
rect 575381 216472 591823 216474
rect 575381 216416 575386 216472
rect 575442 216416 591762 216472
rect 591818 216416 591823 216472
rect 575381 216414 591823 216416
rect 575381 216411 575447 216414
rect 591757 216411 591823 216414
rect 597921 216338 597987 216341
rect 591990 216336 597987 216338
rect 591990 216280 597926 216336
rect 597982 216280 597987 216336
rect 591990 216278 597987 216280
rect 582925 216202 582991 216205
rect 591990 216202 592050 216278
rect 597921 216275 597987 216278
rect 582925 216200 592050 216202
rect 582925 216144 582930 216200
rect 582986 216144 592050 216200
rect 582925 216142 592050 216144
rect 646589 216202 646655 216205
rect 672993 216202 673059 216205
rect 646589 216200 673059 216202
rect 646589 216144 646594 216200
rect 646650 216144 672998 216200
rect 673054 216144 673059 216200
rect 646589 216142 673059 216144
rect 582925 216139 582991 216142
rect 646589 216139 646655 216142
rect 672993 216139 673059 216142
rect 675569 216202 675635 216205
rect 675569 216200 676292 216202
rect 675569 216144 675574 216200
rect 675630 216144 676292 216200
rect 675569 216142 676292 216144
rect 675569 216139 675635 216142
rect 675109 216066 675175 216069
rect 673134 216064 675175 216066
rect 673134 216008 675114 216064
rect 675170 216008 675175 216064
rect 673134 216006 675175 216008
rect 643001 215930 643067 215933
rect 673134 215930 673194 216006
rect 675109 216003 675175 216006
rect 643001 215928 673194 215930
rect 643001 215872 643006 215928
rect 643062 215872 673194 215928
rect 643001 215870 673194 215872
rect 643001 215867 643067 215870
rect 673361 215794 673427 215797
rect 673361 215792 676292 215794
rect 673361 215736 673366 215792
rect 673422 215736 676292 215792
rect 673361 215734 676292 215736
rect 673361 215731 673427 215734
rect 673637 215386 673703 215389
rect 673637 215384 676292 215386
rect 673637 215328 673642 215384
rect 673698 215328 676292 215384
rect 673637 215326 676292 215328
rect 673637 215323 673703 215326
rect 666277 215114 666343 215117
rect 675845 215114 675911 215117
rect 666277 215112 675911 215114
rect 666277 215056 666282 215112
rect 666338 215056 675850 215112
rect 675906 215056 675911 215112
rect 676254 215086 676260 215150
rect 676324 215086 676330 215150
rect 666277 215054 675911 215056
rect 666277 215051 666343 215054
rect 675845 215051 675911 215054
rect 44817 214978 44883 214981
rect 41492 214976 44883 214978
rect 41492 214920 44822 214976
rect 44878 214920 44883 214976
rect 676262 214948 676322 215086
rect 41492 214918 44883 214920
rect 44817 214915 44883 214918
rect 674833 214706 674899 214709
rect 675753 214706 675819 214709
rect 674833 214704 675819 214706
rect 674833 214648 674838 214704
rect 674894 214648 675758 214704
rect 675814 214648 675819 214704
rect 674833 214646 675819 214648
rect 674833 214643 674899 214646
rect 675753 214643 675819 214646
rect 659377 214570 659443 214573
rect 676029 214570 676095 214573
rect 659377 214568 663810 214570
rect 41278 214301 41338 214540
rect 659377 214512 659382 214568
rect 659438 214512 663810 214568
rect 659377 214510 663810 214512
rect 659377 214507 659443 214510
rect 663750 214434 663810 214510
rect 676029 214568 676292 214570
rect 676029 214512 676034 214568
rect 676090 214512 676292 214568
rect 676029 214510 676292 214512
rect 676029 214507 676095 214510
rect 675845 214434 675911 214437
rect 663750 214432 675911 214434
rect 28533 214298 28599 214301
rect 28533 214296 28642 214298
rect 28533 214240 28538 214296
rect 28594 214240 28642 214296
rect 28533 214235 28642 214240
rect 41278 214296 41387 214301
rect 41278 214240 41326 214296
rect 41382 214240 41387 214296
rect 41278 214238 41387 214240
rect 41321 214235 41387 214238
rect 28582 214132 28642 214235
rect 575982 214026 576042 214404
rect 663750 214376 675850 214432
rect 675906 214376 675911 214432
rect 663750 214374 675911 214376
rect 675845 214371 675911 214374
rect 673177 214162 673243 214165
rect 673177 214160 676292 214162
rect 673177 214104 673182 214160
rect 673238 214104 676292 214160
rect 673177 214102 676292 214104
rect 673177 214099 673243 214102
rect 578877 214026 578943 214029
rect 575982 214024 578943 214026
rect 575982 213968 578882 214024
rect 578938 213968 578943 214024
rect 575982 213966 578943 213968
rect 578877 213963 578943 213966
rect 43253 213754 43319 213757
rect 41492 213752 43319 213754
rect 41492 213696 43258 213752
rect 43314 213696 43319 213752
rect 41492 213694 43319 213696
rect 43253 213691 43319 213694
rect 674649 213754 674715 213757
rect 674649 213752 676292 213754
rect 674649 213696 674654 213752
rect 674710 213696 676292 213752
rect 674649 213694 676292 213696
rect 674649 213691 674715 213694
rect 664805 213482 664871 213485
rect 675845 213482 675911 213485
rect 664805 213480 675911 213482
rect 664805 213424 664810 213480
rect 664866 213424 675850 213480
rect 675906 213424 675911 213480
rect 664805 213422 675911 213424
rect 664805 213419 664871 213422
rect 675845 213419 675911 213422
rect 47945 213346 48011 213349
rect 683297 213346 683363 213349
rect 41492 213344 48011 213346
rect 41492 213288 47950 213344
rect 48006 213288 48011 213344
rect 41492 213286 48011 213288
rect 683284 213344 683363 213346
rect 683284 213288 683302 213344
rect 683358 213288 683363 213344
rect 683284 213286 683363 213288
rect 47945 213283 48011 213286
rect 683297 213283 683363 213286
rect 578182 213148 578188 213212
rect 578252 213210 578258 213212
rect 612825 213210 612891 213213
rect 578252 213208 612891 213210
rect 578252 213152 612830 213208
rect 612886 213152 612891 213208
rect 578252 213150 612891 213152
rect 578252 213148 578258 213150
rect 612825 213147 612891 213150
rect 647141 213210 647207 213213
rect 667013 213210 667079 213213
rect 647141 213208 667079 213210
rect 647141 213152 647146 213208
rect 647202 213152 667018 213208
rect 667074 213152 667079 213208
rect 647141 213150 667079 213152
rect 647141 213147 647207 213150
rect 667013 213147 667079 213150
rect 42977 212938 43043 212941
rect 41492 212936 43043 212938
rect 41492 212880 42982 212936
rect 43038 212880 43043 212936
rect 41492 212878 43043 212880
rect 42977 212875 43043 212878
rect 683070 212533 683130 212908
rect 683070 212528 683179 212533
rect 683070 212500 683118 212528
rect 41094 212261 41154 212500
rect 683100 212472 683118 212500
rect 683174 212472 683179 212528
rect 683100 212470 683179 212472
rect 683113 212467 683179 212470
rect 41094 212256 41203 212261
rect 41094 212200 41142 212256
rect 41198 212200 41203 212256
rect 41094 212198 41203 212200
rect 41137 212195 41203 212198
rect 42793 212122 42859 212125
rect 41492 212120 42859 212122
rect 41492 212064 42798 212120
rect 42854 212064 42859 212120
rect 41492 212062 42859 212064
rect 42793 212059 42859 212062
rect 41321 211850 41387 211853
rect 41278 211848 41387 211850
rect 41278 211792 41326 211848
rect 41382 211792 41387 211848
rect 41278 211787 41387 211792
rect 41278 211684 41338 211787
rect 575982 211714 576042 212228
rect 674046 212060 674052 212124
rect 674116 212122 674122 212124
rect 674116 212062 676292 212122
rect 674116 212060 674122 212062
rect 578509 211714 578575 211717
rect 575982 211712 578575 211714
rect 575982 211656 578514 211712
rect 578570 211656 578575 211712
rect 575982 211654 578575 211656
rect 578509 211651 578575 211654
rect 672165 211442 672231 211445
rect 676765 211444 676831 211445
rect 677041 211444 677107 211445
rect 676765 211442 676812 211444
rect 672165 211440 676506 211442
rect 672165 211384 672170 211440
rect 672226 211384 676506 211440
rect 672165 211382 676506 211384
rect 676720 211440 676812 211442
rect 676720 211384 676770 211440
rect 676720 211382 676812 211384
rect 672165 211379 672231 211382
rect 44173 211306 44239 211309
rect 41492 211304 44239 211306
rect 41492 211248 44178 211304
rect 44234 211248 44239 211304
rect 41492 211246 44239 211248
rect 676446 211306 676506 211382
rect 676765 211380 676812 211382
rect 676876 211380 676882 211444
rect 676990 211380 676996 211444
rect 677060 211442 677107 211444
rect 677060 211440 677152 211442
rect 677102 211384 677152 211440
rect 677060 211382 677152 211384
rect 677060 211380 677107 211382
rect 676765 211379 676831 211380
rect 677041 211379 677107 211380
rect 676446 211246 676690 211306
rect 44173 211243 44239 211246
rect 670734 211108 670740 211172
rect 670804 211170 670810 211172
rect 671981 211170 672047 211173
rect 670804 211168 672047 211170
rect 670804 211112 671986 211168
rect 672042 211112 672047 211168
rect 670804 211110 672047 211112
rect 670804 211108 670810 211110
rect 671981 211107 672047 211110
rect 673821 211170 673887 211173
rect 676305 211170 676371 211173
rect 673821 211168 676371 211170
rect 673821 211112 673826 211168
rect 673882 211112 676310 211168
rect 676366 211112 676371 211168
rect 673821 211110 676371 211112
rect 676630 211170 676690 211246
rect 683113 211170 683179 211173
rect 676630 211168 683179 211170
rect 676630 211112 683118 211168
rect 683174 211112 683179 211168
rect 676630 211110 683179 211112
rect 673821 211107 673887 211110
rect 676305 211107 676371 211110
rect 683113 211107 683179 211110
rect 48129 210898 48195 210901
rect 41492 210896 48195 210898
rect 41492 210840 48134 210896
rect 48190 210840 48195 210896
rect 41492 210838 48195 210840
rect 48129 210835 48195 210838
rect 41278 210221 41338 210460
rect 683297 210354 683363 210357
rect 678930 210352 683363 210354
rect 678930 210296 683302 210352
rect 683358 210296 683363 210352
rect 678930 210294 683363 210296
rect 41278 210216 41387 210221
rect 41278 210160 41326 210216
rect 41382 210160 41387 210216
rect 41278 210158 41387 210160
rect 41321 210155 41387 210158
rect 672257 210218 672323 210221
rect 678930 210218 678990 210294
rect 683297 210291 683363 210294
rect 672257 210216 678990 210218
rect 672257 210160 672262 210216
rect 672318 210160 678990 210216
rect 672257 210158 678990 210160
rect 672257 210155 672323 210158
rect 41094 209813 41154 210052
rect 41094 209808 41203 209813
rect 41094 209752 41142 209808
rect 41198 209752 41203 209808
rect 41094 209750 41203 209752
rect 575982 209810 576042 210052
rect 578417 209810 578483 209813
rect 575982 209808 578483 209810
rect 575982 209752 578422 209808
rect 578478 209752 578483 209808
rect 575982 209750 578483 209752
rect 41137 209747 41203 209750
rect 578417 209747 578483 209750
rect 46933 209674 46999 209677
rect 41492 209672 46999 209674
rect 41492 209616 46938 209672
rect 46994 209616 46999 209672
rect 41492 209614 46999 209616
rect 46933 209611 46999 209614
rect 672901 209674 672967 209677
rect 673126 209674 673132 209676
rect 672901 209672 673132 209674
rect 672901 209616 672906 209672
rect 672962 209616 673132 209672
rect 672901 209614 673132 209616
rect 672901 209611 672967 209614
rect 673126 209612 673132 209614
rect 673196 209612 673202 209676
rect 674557 209674 674623 209677
rect 675477 209674 675543 209677
rect 674557 209672 675543 209674
rect 674557 209616 674562 209672
rect 674618 209616 675482 209672
rect 675538 209616 675543 209672
rect 674557 209614 675543 209616
rect 674557 209611 674623 209614
rect 675477 209611 675543 209614
rect 41321 209402 41387 209405
rect 41638 209402 41644 209404
rect 41321 209400 41644 209402
rect 41321 209344 41326 209400
rect 41382 209344 41644 209400
rect 41321 209342 41644 209344
rect 41321 209339 41387 209342
rect 41638 209340 41644 209342
rect 41708 209340 41714 209404
rect 672073 209402 672139 209405
rect 677685 209402 677751 209405
rect 672073 209400 677751 209402
rect 672073 209344 672078 209400
rect 672134 209344 677690 209400
rect 677746 209344 677751 209400
rect 672073 209342 677751 209344
rect 672073 209339 672139 209342
rect 677685 209339 677751 209342
rect 41278 208997 41338 209236
rect 41278 208992 41387 208997
rect 41278 208936 41326 208992
rect 41382 208936 41387 208992
rect 41278 208934 41387 208936
rect 41321 208931 41387 208934
rect 47117 208858 47183 208861
rect 41492 208856 47183 208858
rect 41492 208800 47122 208856
rect 47178 208800 47183 208856
rect 41492 208798 47183 208800
rect 47117 208795 47183 208798
rect 41689 208586 41755 208589
rect 49325 208586 49391 208589
rect 41689 208584 49391 208586
rect 41689 208528 41694 208584
rect 41750 208528 49330 208584
rect 49386 208528 49391 208584
rect 41689 208526 49391 208528
rect 41689 208523 41755 208526
rect 49325 208523 49391 208526
rect 40542 208180 40602 208420
rect 674005 208314 674071 208317
rect 676765 208314 676831 208317
rect 674005 208312 676831 208314
rect 674005 208256 674010 208312
rect 674066 208256 676770 208312
rect 676826 208256 676831 208312
rect 674005 208254 676831 208256
rect 674005 208251 674071 208254
rect 676765 208251 676831 208254
rect 40534 208116 40540 208180
rect 40604 208116 40610 208180
rect 44173 208042 44239 208045
rect 41492 208040 44239 208042
rect 41492 207984 44178 208040
rect 44234 207984 44239 208040
rect 41492 207982 44239 207984
rect 44173 207979 44239 207982
rect 589457 208042 589523 208045
rect 589457 208040 592572 208042
rect 589457 207984 589462 208040
rect 589518 207984 592572 208040
rect 589457 207982 592572 207984
rect 589457 207979 589523 207982
rect 42793 207634 42859 207637
rect 41492 207632 42859 207634
rect 41492 207576 42798 207632
rect 42854 207576 42859 207632
rect 41492 207574 42859 207576
rect 42793 207571 42859 207574
rect 575982 207498 576042 207876
rect 579521 207498 579587 207501
rect 575982 207496 579587 207498
rect 575982 207440 579526 207496
rect 579582 207440 579587 207496
rect 575982 207438 579587 207440
rect 579521 207435 579587 207438
rect 41137 207362 41203 207365
rect 41822 207362 41828 207364
rect 41137 207360 41828 207362
rect 41137 207304 41142 207360
rect 41198 207304 41828 207360
rect 41137 207302 41828 207304
rect 41137 207299 41203 207302
rect 41822 207300 41828 207302
rect 41892 207300 41898 207364
rect 675017 207362 675083 207365
rect 666878 207360 675083 207362
rect 666878 207304 675022 207360
rect 675078 207304 675083 207360
rect 666878 207302 675083 207304
rect 666878 207294 666938 207302
rect 675017 207299 675083 207302
rect 666356 207234 666938 207294
rect 40910 206957 40970 207196
rect 675702 207028 675708 207092
rect 675772 207090 675778 207092
rect 679617 207090 679683 207093
rect 675772 207088 679683 207090
rect 675772 207032 679622 207088
rect 679678 207032 679683 207088
rect 675772 207030 679683 207032
rect 675772 207028 675778 207030
rect 679617 207027 679683 207030
rect 40910 206952 41019 206957
rect 40910 206896 40958 206952
rect 41014 206896 41019 206952
rect 40910 206894 41019 206896
rect 40953 206891 41019 206894
rect 44357 206818 44423 206821
rect 41492 206816 44423 206818
rect 41492 206760 44362 206816
rect 44418 206760 44423 206816
rect 41492 206758 44423 206760
rect 44357 206755 44423 206758
rect 667974 206484 667980 206548
rect 668044 206546 668050 206548
rect 669221 206546 669287 206549
rect 668044 206544 669287 206546
rect 668044 206488 669226 206544
rect 669282 206488 669287 206544
rect 668044 206486 669287 206488
rect 668044 206484 668050 206486
rect 669221 206483 669287 206486
rect 42977 206410 43043 206413
rect 41492 206408 43043 206410
rect 41492 206352 42982 206408
rect 43038 206352 43043 206408
rect 41492 206350 43043 206352
rect 42977 206347 43043 206350
rect 589457 206410 589523 206413
rect 677869 206410 677935 206413
rect 589457 206408 592572 206410
rect 589457 206352 589462 206408
rect 589518 206352 592572 206408
rect 589457 206350 592572 206352
rect 669454 206408 677935 206410
rect 669454 206352 677874 206408
rect 677930 206352 677935 206408
rect 669454 206350 677935 206352
rect 589457 206347 589523 206350
rect 669078 206212 669084 206276
rect 669148 206274 669154 206276
rect 669454 206274 669514 206350
rect 677869 206347 677935 206350
rect 669148 206214 669514 206274
rect 669148 206212 669154 206214
rect 44633 206002 44699 206005
rect 41492 206000 44699 206002
rect 41492 205944 44638 206000
rect 44694 205944 44699 206000
rect 41492 205942 44699 205944
rect 44633 205939 44699 205942
rect 579521 205866 579587 205869
rect 575798 205864 579587 205866
rect 575798 205808 579526 205864
rect 579582 205808 579587 205864
rect 575798 205806 579587 205808
rect 575798 205700 575858 205806
rect 579521 205803 579587 205806
rect 43805 205594 43871 205597
rect 41492 205592 43871 205594
rect 41492 205536 43810 205592
rect 43866 205536 43871 205592
rect 41492 205534 43871 205536
rect 43805 205531 43871 205534
rect 675753 205594 675819 205597
rect 676438 205594 676444 205596
rect 675753 205592 676444 205594
rect 675753 205536 675758 205592
rect 675814 205536 676444 205592
rect 675753 205534 676444 205536
rect 675753 205531 675819 205534
rect 676438 205532 676444 205534
rect 676508 205532 676514 205596
rect 43989 205186 44055 205189
rect 41492 205184 44055 205186
rect 41492 205128 43994 205184
rect 44050 205128 44055 205184
rect 41492 205126 44055 205128
rect 43989 205123 44055 205126
rect 44817 204778 44883 204781
rect 41492 204776 44883 204778
rect 41492 204720 44822 204776
rect 44878 204720 44883 204776
rect 41492 204718 44883 204720
rect 44817 204715 44883 204718
rect 589641 204778 589707 204781
rect 589641 204776 592572 204778
rect 589641 204720 589646 204776
rect 589702 204720 592572 204776
rect 589641 204718 592572 204720
rect 589641 204715 589707 204718
rect 41321 204506 41387 204509
rect 41638 204506 41644 204508
rect 41321 204504 41644 204506
rect 41321 204448 41326 204504
rect 41382 204448 41644 204504
rect 41321 204446 41644 204448
rect 41321 204443 41387 204446
rect 41638 204444 41644 204446
rect 41708 204444 41714 204508
rect 35758 204101 35818 204340
rect 675661 204236 675727 204237
rect 675661 204232 675708 204236
rect 675772 204234 675778 204236
rect 675661 204176 675666 204232
rect 675661 204172 675708 204176
rect 675772 204174 675818 204234
rect 675772 204172 675778 204174
rect 675661 204171 675727 204172
rect 35758 204096 35867 204101
rect 35758 204040 35806 204096
rect 35862 204040 35867 204096
rect 35758 204038 35867 204040
rect 35801 204035 35867 204038
rect 666356 203970 666938 204030
rect 44541 203962 44607 203965
rect 41492 203960 44607 203962
rect 41492 203904 44546 203960
rect 44602 203904 44607 203960
rect 41492 203902 44607 203904
rect 666878 203962 666938 203970
rect 673821 203962 673887 203965
rect 666878 203960 673887 203962
rect 666878 203904 673826 203960
rect 673882 203904 673887 203960
rect 666878 203902 673887 203904
rect 44541 203899 44607 203902
rect 673821 203899 673887 203902
rect 46381 203554 46447 203557
rect 41492 203552 46447 203554
rect 41492 203496 46386 203552
rect 46442 203496 46447 203552
rect 41492 203494 46447 203496
rect 46381 203491 46447 203494
rect 40953 203282 41019 203285
rect 43253 203282 43319 203285
rect 40953 203280 43319 203282
rect 40953 203224 40958 203280
rect 41014 203224 43258 203280
rect 43314 203224 43319 203280
rect 40953 203222 43319 203224
rect 575982 203282 576042 203524
rect 578509 203282 578575 203285
rect 575982 203280 578575 203282
rect 575982 203224 578514 203280
rect 578570 203224 578575 203280
rect 575982 203222 578575 203224
rect 40953 203219 41019 203222
rect 43253 203219 43319 203222
rect 578509 203219 578575 203222
rect 589457 203146 589523 203149
rect 589457 203144 592572 203146
rect 589457 203088 589462 203144
rect 589518 203088 592572 203144
rect 589457 203086 592572 203088
rect 589457 203083 589523 203086
rect 674925 202602 674991 202605
rect 675385 202602 675451 202605
rect 674925 202600 675451 202602
rect 674925 202544 674930 202600
rect 674986 202544 675390 202600
rect 675446 202544 675451 202600
rect 674925 202542 675451 202544
rect 674925 202539 674991 202542
rect 675385 202539 675451 202542
rect 669078 202466 669084 202468
rect 666694 202406 669084 202466
rect 666694 202398 666754 202406
rect 669078 202404 669084 202406
rect 669148 202404 669154 202468
rect 666356 202338 666754 202398
rect 35801 202194 35867 202197
rect 43621 202194 43687 202197
rect 35801 202192 43687 202194
rect 35801 202136 35806 202192
rect 35862 202136 43626 202192
rect 43682 202136 43687 202192
rect 35801 202134 43687 202136
rect 35801 202131 35867 202134
rect 43621 202131 43687 202134
rect 589457 201514 589523 201517
rect 589457 201512 592572 201514
rect 589457 201456 589462 201512
rect 589518 201456 592572 201512
rect 589457 201454 592572 201456
rect 589457 201451 589523 201454
rect 673361 201378 673427 201381
rect 675109 201378 675175 201381
rect 673361 201376 675175 201378
rect 575982 200834 576042 201348
rect 673361 201320 673366 201376
rect 673422 201320 675114 201376
rect 675170 201320 675175 201376
rect 673361 201318 675175 201320
rect 673361 201315 673427 201318
rect 675109 201315 675175 201318
rect 578785 200834 578851 200837
rect 575982 200832 578851 200834
rect 575982 200776 578790 200832
rect 578846 200776 578851 200832
rect 575982 200774 578851 200776
rect 578785 200771 578851 200774
rect 672257 200834 672323 200837
rect 672901 200834 672967 200837
rect 672257 200832 672967 200834
rect 672257 200776 672262 200832
rect 672318 200776 672906 200832
rect 672962 200776 672967 200832
rect 672257 200774 672967 200776
rect 672257 200771 672323 200774
rect 672901 200771 672967 200774
rect 673637 200834 673703 200837
rect 674833 200834 674899 200837
rect 673637 200832 674899 200834
rect 673637 200776 673642 200832
rect 673698 200776 674838 200832
rect 674894 200776 674899 200832
rect 673637 200774 674899 200776
rect 673637 200771 673703 200774
rect 674833 200771 674899 200774
rect 675753 200834 675819 200837
rect 676990 200834 676996 200836
rect 675753 200832 676996 200834
rect 675753 200776 675758 200832
rect 675814 200776 676996 200832
rect 675753 200774 676996 200776
rect 675753 200771 675819 200774
rect 676990 200772 676996 200774
rect 677060 200772 677066 200836
rect 41505 200698 41571 200701
rect 49509 200698 49575 200701
rect 41505 200696 49575 200698
rect 41505 200640 41510 200696
rect 41566 200640 49514 200696
rect 49570 200640 49575 200696
rect 41505 200638 49575 200640
rect 41505 200635 41571 200638
rect 49509 200635 49575 200638
rect 589457 199882 589523 199885
rect 589457 199880 592572 199882
rect 589457 199824 589462 199880
rect 589518 199824 592572 199880
rect 589457 199822 592572 199824
rect 589457 199819 589523 199822
rect 670969 199202 671035 199205
rect 666694 199200 671035 199202
rect 575982 198930 576042 199172
rect 666694 199144 670974 199200
rect 671030 199144 671035 199200
rect 666694 199142 671035 199144
rect 666694 199134 666754 199142
rect 670969 199139 671035 199142
rect 666356 199074 666754 199134
rect 579521 198930 579587 198933
rect 575982 198928 579587 198930
rect 575982 198872 579526 198928
rect 579582 198872 579587 198928
rect 575982 198870 579587 198872
rect 579521 198867 579587 198870
rect 666686 198324 666692 198388
rect 666756 198386 666762 198388
rect 675385 198386 675451 198389
rect 666756 198384 675451 198386
rect 666756 198328 675390 198384
rect 675446 198328 675451 198384
rect 666756 198326 675451 198328
rect 666756 198324 666762 198326
rect 675385 198323 675451 198326
rect 590377 198250 590443 198253
rect 590377 198248 592572 198250
rect 590377 198192 590382 198248
rect 590438 198192 592572 198248
rect 590377 198190 592572 198192
rect 590377 198187 590443 198190
rect 673177 197706 673243 197709
rect 675477 197706 675543 197709
rect 673177 197704 675543 197706
rect 673177 197648 673182 197704
rect 673238 197648 675482 197704
rect 675538 197648 675543 197704
rect 673177 197646 675543 197648
rect 673177 197643 673243 197646
rect 675477 197643 675543 197646
rect 672165 197570 672231 197573
rect 666694 197568 672231 197570
rect 666694 197512 672170 197568
rect 672226 197512 672231 197568
rect 666694 197510 672231 197512
rect 666694 197502 666754 197510
rect 672165 197507 672231 197510
rect 666356 197442 666754 197502
rect 40534 197100 40540 197164
rect 40604 197162 40610 197164
rect 41781 197162 41847 197165
rect 40604 197160 41847 197162
rect 40604 197104 41786 197160
rect 41842 197104 41847 197160
rect 40604 197102 41847 197104
rect 40604 197100 40610 197102
rect 41781 197099 41847 197102
rect 675753 197162 675819 197165
rect 676254 197162 676260 197164
rect 675753 197160 676260 197162
rect 675753 197104 675758 197160
rect 675814 197104 676260 197160
rect 675753 197102 676260 197104
rect 675753 197099 675819 197102
rect 676254 197100 676260 197102
rect 676324 197100 676330 197164
rect 49325 196482 49391 196485
rect 575982 196482 576042 196996
rect 589457 196618 589523 196621
rect 589457 196616 592572 196618
rect 589457 196560 589462 196616
rect 589518 196560 592572 196616
rect 589457 196558 592572 196560
rect 589457 196555 589523 196558
rect 578509 196482 578575 196485
rect 49325 196480 52164 196482
rect 49325 196424 49330 196480
rect 49386 196424 52164 196480
rect 49325 196422 52164 196424
rect 575982 196480 578575 196482
rect 575982 196424 578514 196480
rect 578570 196424 578575 196480
rect 575982 196422 578575 196424
rect 49325 196419 49391 196422
rect 578509 196419 578575 196422
rect 674649 196074 674715 196077
rect 675201 196074 675267 196077
rect 674649 196072 675267 196074
rect 674649 196016 674654 196072
rect 674710 196016 675206 196072
rect 675262 196016 675267 196072
rect 674649 196014 675267 196016
rect 674649 196011 674715 196014
rect 675201 196011 675267 196014
rect 42149 195802 42215 195805
rect 44541 195802 44607 195805
rect 42149 195800 44607 195802
rect 42149 195744 42154 195800
rect 42210 195744 44546 195800
rect 44602 195744 44607 195800
rect 42149 195742 44607 195744
rect 42149 195739 42215 195742
rect 44541 195739 44607 195742
rect 41873 195260 41939 195261
rect 41822 195258 41828 195260
rect 41782 195198 41828 195258
rect 41892 195256 41939 195260
rect 41934 195200 41939 195256
rect 41822 195196 41828 195198
rect 41892 195196 41939 195200
rect 41873 195195 41939 195196
rect 579521 194986 579587 194989
rect 575798 194984 579587 194986
rect 575798 194928 579526 194984
rect 579582 194928 579587 194984
rect 575798 194926 579587 194928
rect 575798 194820 575858 194926
rect 579521 194923 579587 194926
rect 589273 194986 589339 194989
rect 589273 194984 592572 194986
rect 589273 194928 589278 194984
rect 589334 194928 592572 194984
rect 589273 194926 592572 194928
rect 589273 194923 589339 194926
rect 48129 194442 48195 194445
rect 48129 194440 52164 194442
rect 48129 194384 48134 194440
rect 48190 194384 52164 194440
rect 48129 194382 52164 194384
rect 48129 194379 48195 194382
rect 671153 194306 671219 194309
rect 666694 194304 671219 194306
rect 666694 194248 671158 194304
rect 671214 194248 671219 194304
rect 666694 194246 671219 194248
rect 666694 194238 666754 194246
rect 671153 194243 671219 194246
rect 666356 194178 666754 194238
rect 589457 193354 589523 193357
rect 589457 193352 592572 193354
rect 589457 193296 589462 193352
rect 589518 193296 592572 193352
rect 589457 193294 592572 193296
rect 589457 193291 589523 193294
rect 42425 193218 42491 193221
rect 44357 193218 44423 193221
rect 42425 193216 44423 193218
rect 42425 193160 42430 193216
rect 42486 193160 44362 193216
rect 44418 193160 44423 193216
rect 42425 193158 44423 193160
rect 42425 193155 42491 193158
rect 44357 193155 44423 193158
rect 675661 193218 675727 193221
rect 675886 193218 675892 193220
rect 675661 193216 675892 193218
rect 675661 193160 675666 193216
rect 675722 193160 675892 193216
rect 675661 193158 675892 193160
rect 675661 193155 675727 193158
rect 675886 193156 675892 193158
rect 675956 193156 675962 193220
rect 668117 192674 668183 192677
rect 666694 192672 668183 192674
rect 49509 192402 49575 192405
rect 49509 192400 52164 192402
rect 49509 192344 49514 192400
rect 49570 192344 52164 192400
rect 49509 192342 52164 192344
rect 49509 192339 49575 192342
rect 575982 192266 576042 192644
rect 666694 192616 668122 192672
rect 668178 192616 668183 192672
rect 666694 192614 668183 192616
rect 666694 192606 666754 192614
rect 668117 192611 668183 192614
rect 666356 192546 666754 192606
rect 671981 192402 672047 192405
rect 675109 192402 675175 192405
rect 671981 192400 675175 192402
rect 671981 192344 671986 192400
rect 672042 192344 675114 192400
rect 675170 192344 675175 192400
rect 671981 192342 675175 192344
rect 671981 192339 672047 192342
rect 675109 192339 675175 192342
rect 579521 192266 579587 192269
rect 575982 192264 579587 192266
rect 575982 192208 579526 192264
rect 579582 192208 579587 192264
rect 575982 192206 579587 192208
rect 579521 192203 579587 192206
rect 42333 191722 42399 191725
rect 43989 191722 44055 191725
rect 42333 191720 44055 191722
rect 42333 191664 42338 191720
rect 42394 191664 43994 191720
rect 44050 191664 44055 191720
rect 42333 191662 44055 191664
rect 42333 191659 42399 191662
rect 43989 191659 44055 191662
rect 589457 191722 589523 191725
rect 589457 191720 592572 191722
rect 589457 191664 589462 191720
rect 589518 191664 592572 191720
rect 589457 191662 592572 191664
rect 589457 191659 589523 191662
rect 675753 191586 675819 191589
rect 676070 191586 676076 191588
rect 675753 191584 676076 191586
rect 675753 191528 675758 191584
rect 675814 191528 676076 191584
rect 675753 191526 676076 191528
rect 675753 191523 675819 191526
rect 676070 191524 676076 191526
rect 676140 191524 676146 191588
rect 42425 191178 42491 191181
rect 42977 191178 43043 191181
rect 42425 191176 43043 191178
rect 42425 191120 42430 191176
rect 42486 191120 42982 191176
rect 43038 191120 43043 191176
rect 42425 191118 43043 191120
rect 42425 191115 42491 191118
rect 42977 191115 43043 191118
rect 579521 190770 579587 190773
rect 575798 190768 579587 190770
rect 575798 190712 579526 190768
rect 579582 190712 579587 190768
rect 575798 190710 579587 190712
rect 42425 190498 42491 190501
rect 43805 190498 43871 190501
rect 42425 190496 43871 190498
rect 42425 190440 42430 190496
rect 42486 190440 43810 190496
rect 43866 190440 43871 190496
rect 42425 190438 43871 190440
rect 42425 190435 42491 190438
rect 43805 190435 43871 190438
rect 47945 190498 48011 190501
rect 47945 190496 52164 190498
rect 47945 190440 47950 190496
rect 48006 190440 52164 190496
rect 575798 190468 575858 190710
rect 579521 190707 579587 190710
rect 47945 190438 52164 190440
rect 47945 190435 48011 190438
rect 590561 190090 590627 190093
rect 590561 190088 592572 190090
rect 590561 190032 590566 190088
rect 590622 190032 592572 190088
rect 590561 190030 592572 190032
rect 590561 190027 590627 190030
rect 42425 189954 42491 189957
rect 47117 189954 47183 189957
rect 42425 189952 47183 189954
rect 42425 189896 42430 189952
rect 42486 189896 47122 189952
rect 47178 189896 47183 189952
rect 42425 189894 47183 189896
rect 42425 189891 42491 189894
rect 47117 189891 47183 189894
rect 671705 189410 671771 189413
rect 666694 189408 671771 189410
rect 666694 189352 671710 189408
rect 671766 189352 671771 189408
rect 666694 189350 671771 189352
rect 666694 189342 666754 189350
rect 671705 189347 671771 189350
rect 666356 189282 666754 189342
rect 589641 188458 589707 188461
rect 669313 188458 669379 188461
rect 672533 188458 672599 188461
rect 589641 188456 592572 188458
rect 589641 188400 589646 188456
rect 589702 188400 592572 188456
rect 589641 188398 592572 188400
rect 669313 188456 672599 188458
rect 669313 188400 669318 188456
rect 669374 188400 672538 188456
rect 672594 188400 672599 188456
rect 669313 188398 672599 188400
rect 589641 188395 589707 188398
rect 669313 188395 669379 188398
rect 672533 188395 672599 188398
rect 575982 188050 576042 188292
rect 579521 188050 579587 188053
rect 575982 188048 579587 188050
rect 575982 187992 579526 188048
rect 579582 187992 579587 188048
rect 575982 187990 579587 187992
rect 579521 187987 579587 187990
rect 666356 187650 666754 187710
rect 42425 187642 42491 187645
rect 44633 187642 44699 187645
rect 42425 187640 44699 187642
rect 42425 187584 42430 187640
rect 42486 187584 44638 187640
rect 44694 187584 44699 187640
rect 42425 187582 44699 187584
rect 666694 187642 666754 187650
rect 668025 187642 668091 187645
rect 666694 187640 668091 187642
rect 666694 187584 668030 187640
rect 668086 187584 668091 187640
rect 666694 187582 668091 187584
rect 42425 187579 42491 187582
rect 44633 187579 44699 187582
rect 668025 187579 668091 187582
rect 42425 186826 42491 186829
rect 43253 186826 43319 186829
rect 42425 186824 43319 186826
rect 42425 186768 42430 186824
rect 42486 186768 43258 186824
rect 43314 186768 43319 186824
rect 42425 186766 43319 186768
rect 42425 186763 42491 186766
rect 43253 186763 43319 186766
rect 589457 186826 589523 186829
rect 589457 186824 592572 186826
rect 589457 186768 589462 186824
rect 589518 186768 592572 186824
rect 589457 186766 592572 186768
rect 589457 186763 589523 186766
rect 579521 186282 579587 186285
rect 575798 186280 579587 186282
rect 575798 186224 579526 186280
rect 579582 186224 579587 186280
rect 575798 186222 579587 186224
rect 575798 186116 575858 186222
rect 579521 186219 579587 186222
rect 41781 185876 41847 185877
rect 41781 185872 41828 185876
rect 41892 185874 41898 185876
rect 41781 185816 41786 185872
rect 41781 185812 41828 185816
rect 41892 185814 41938 185874
rect 41892 185812 41898 185814
rect 41781 185811 41847 185812
rect 589457 185194 589523 185197
rect 589457 185192 592572 185194
rect 589457 185136 589462 185192
rect 589518 185136 592572 185192
rect 589457 185134 592572 185136
rect 589457 185131 589523 185134
rect 667933 184514 667999 184517
rect 666694 184512 667999 184514
rect 666694 184456 667938 184512
rect 667994 184456 667999 184512
rect 666694 184454 667999 184456
rect 666694 184446 666754 184454
rect 667933 184451 667999 184454
rect 666356 184386 666754 184446
rect 579521 184378 579587 184381
rect 575798 184376 579587 184378
rect 575798 184320 579526 184376
rect 579582 184320 579587 184376
rect 575798 184318 579587 184320
rect 41454 184044 41460 184108
rect 41524 184106 41530 184108
rect 41781 184106 41847 184109
rect 41524 184104 41847 184106
rect 41524 184048 41786 184104
rect 41842 184048 41847 184104
rect 41524 184046 41847 184048
rect 41524 184044 41530 184046
rect 41781 184043 41847 184046
rect 575798 183940 575858 184318
rect 579521 184315 579587 184318
rect 589457 183562 589523 183565
rect 672073 183562 672139 183565
rect 672942 183562 672948 183564
rect 589457 183560 592572 183562
rect 589457 183504 589462 183560
rect 589518 183504 592572 183560
rect 589457 183502 592572 183504
rect 672073 183560 672948 183562
rect 672073 183504 672078 183560
rect 672134 183504 672948 183560
rect 672073 183502 672948 183504
rect 589457 183499 589523 183502
rect 672073 183499 672139 183502
rect 672942 183500 672948 183502
rect 673012 183500 673018 183564
rect 42425 183154 42491 183157
rect 44173 183154 44239 183157
rect 42425 183152 44239 183154
rect 42425 183096 42430 183152
rect 42486 183096 44178 183152
rect 44234 183096 44239 183152
rect 42425 183094 44239 183096
rect 42425 183091 42491 183094
rect 44173 183091 44239 183094
rect 668301 182882 668367 182885
rect 666694 182880 668367 182882
rect 666694 182824 668306 182880
rect 668362 182824 668367 182880
rect 666694 182822 668367 182824
rect 666694 182814 666754 182822
rect 668301 182819 668367 182822
rect 666356 182754 666754 182814
rect 579521 181930 579587 181933
rect 575798 181928 579587 181930
rect 575798 181872 579526 181928
rect 579582 181872 579587 181928
rect 575798 181870 579587 181872
rect 575798 181764 575858 181870
rect 579521 181867 579587 181870
rect 590561 181930 590627 181933
rect 590561 181928 592572 181930
rect 590561 181872 590566 181928
rect 590622 181872 592572 181928
rect 590561 181870 592572 181872
rect 590561 181867 590627 181870
rect 667197 181386 667263 181389
rect 675845 181386 675911 181389
rect 667197 181384 675911 181386
rect 667197 181328 667202 181384
rect 667258 181328 675850 181384
rect 675906 181328 675911 181384
rect 667197 181326 675911 181328
rect 667197 181323 667263 181326
rect 675845 181323 675911 181326
rect 42425 180706 42491 180709
rect 46933 180706 46999 180709
rect 42425 180704 46999 180706
rect 42425 180648 42430 180704
rect 42486 180648 46938 180704
rect 46994 180648 46999 180704
rect 42425 180646 46999 180648
rect 42425 180643 42491 180646
rect 46933 180643 46999 180646
rect 589641 180298 589707 180301
rect 589641 180296 592572 180298
rect 589641 180240 589646 180296
rect 589702 180240 592572 180296
rect 589641 180238 592572 180240
rect 589641 180235 589707 180238
rect 578785 180162 578851 180165
rect 575798 180160 578851 180162
rect 575798 180104 578790 180160
rect 578846 180104 578851 180160
rect 575798 180102 578851 180104
rect 575798 179588 575858 180102
rect 578785 180099 578851 180102
rect 666356 179490 666938 179550
rect 666878 179482 666938 179490
rect 674281 179482 674347 179485
rect 666878 179480 674347 179482
rect 666878 179424 674286 179480
rect 674342 179424 674347 179480
rect 666878 179422 674347 179424
rect 674281 179419 674347 179422
rect 666645 178802 666711 178805
rect 676029 178802 676095 178805
rect 666645 178800 676095 178802
rect 666645 178744 666650 178800
rect 666706 178744 676034 178800
rect 676090 178744 676095 178800
rect 666645 178742 676095 178744
rect 666645 178739 666711 178742
rect 676029 178739 676095 178742
rect 589457 178666 589523 178669
rect 589457 178664 592572 178666
rect 589457 178608 589462 178664
rect 589518 178608 592572 178664
rect 589457 178606 592572 178608
rect 589457 178603 589523 178606
rect 666829 178530 666895 178533
rect 666829 178528 676292 178530
rect 666829 178472 666834 178528
rect 666890 178472 676292 178528
rect 666829 178470 676292 178472
rect 666829 178467 666895 178470
rect 675845 178122 675911 178125
rect 675845 178120 676292 178122
rect 675845 178064 675850 178120
rect 675906 178064 676292 178120
rect 675845 178062 676292 178064
rect 675845 178059 675911 178062
rect 672441 177986 672507 177989
rect 666694 177984 672507 177986
rect 666694 177928 672446 177984
rect 672502 177928 672507 177984
rect 666694 177926 672507 177928
rect 666694 177918 666754 177926
rect 672441 177923 672507 177926
rect 666356 177858 666754 177918
rect 579521 177714 579587 177717
rect 575798 177712 579587 177714
rect 575798 177656 579526 177712
rect 579582 177656 579587 177712
rect 575798 177654 579587 177656
rect 575798 177412 575858 177654
rect 579521 177651 579587 177654
rect 676029 177714 676095 177717
rect 676029 177712 676292 177714
rect 676029 177656 676034 177712
rect 676090 177656 676292 177712
rect 676029 177654 676292 177656
rect 676029 177651 676095 177654
rect 669405 177306 669471 177309
rect 669405 177304 676292 177306
rect 669405 177248 669410 177304
rect 669466 177248 676292 177304
rect 669405 177246 676292 177248
rect 669405 177243 669471 177246
rect 589641 177034 589707 177037
rect 589641 177032 592572 177034
rect 589641 176976 589646 177032
rect 589702 176976 592572 177032
rect 589641 176974 592572 176976
rect 589641 176971 589707 176974
rect 674281 176898 674347 176901
rect 674281 176896 676292 176898
rect 674281 176840 674286 176896
rect 674342 176840 676292 176896
rect 674281 176838 676292 176840
rect 674281 176835 674347 176838
rect 670601 176490 670667 176493
rect 670601 176488 676292 176490
rect 670601 176432 670606 176488
rect 670662 176432 676292 176488
rect 670601 176430 676292 176432
rect 670601 176427 670667 176430
rect 674649 176082 674715 176085
rect 674649 176080 676292 176082
rect 674649 176024 674654 176080
rect 674710 176024 676292 176080
rect 674649 176022 676292 176024
rect 674649 176019 674715 176022
rect 670785 175674 670851 175677
rect 670785 175672 676292 175674
rect 670785 175616 670790 175672
rect 670846 175616 676292 175672
rect 670785 175614 676292 175616
rect 670785 175611 670851 175614
rect 589457 175402 589523 175405
rect 589457 175400 592572 175402
rect 589457 175344 589462 175400
rect 589518 175344 592572 175400
rect 589457 175342 592572 175344
rect 589457 175339 589523 175342
rect 672533 175266 672599 175269
rect 672533 175264 676292 175266
rect 575982 175130 576042 175236
rect 672533 175208 672538 175264
rect 672594 175208 676292 175264
rect 672533 175206 676292 175208
rect 672533 175203 672599 175206
rect 578785 175130 578851 175133
rect 575982 175128 578851 175130
rect 575982 175072 578790 175128
rect 578846 175072 578851 175128
rect 575982 175070 578851 175072
rect 578785 175067 578851 175070
rect 667749 174994 667815 174997
rect 667749 174992 669330 174994
rect 667749 174936 667754 174992
rect 667810 174936 669330 174992
rect 667749 174934 669330 174936
rect 667749 174931 667815 174934
rect 669270 174858 669330 174934
rect 669270 174798 676292 174858
rect 667933 174722 667999 174725
rect 666694 174720 667999 174722
rect 666694 174664 667938 174720
rect 667994 174664 667999 174720
rect 666694 174662 667999 174664
rect 666694 174654 666754 174662
rect 667933 174659 667999 174662
rect 666356 174594 666754 174654
rect 673361 174450 673427 174453
rect 673361 174448 676292 174450
rect 673361 174392 673366 174448
rect 673422 174392 676292 174448
rect 673361 174390 676292 174392
rect 673361 174387 673427 174390
rect 675886 173980 675892 174044
rect 675956 174042 675962 174044
rect 675956 173982 676292 174042
rect 675956 173980 675962 173982
rect 589457 173770 589523 173773
rect 589457 173768 592572 173770
rect 589457 173712 589462 173768
rect 589518 173712 592572 173768
rect 589457 173710 592572 173712
rect 589457 173707 589523 173710
rect 675702 173572 675708 173636
rect 675772 173634 675778 173636
rect 675772 173574 676292 173634
rect 675772 173572 675778 173574
rect 578417 173498 578483 173501
rect 575798 173496 578483 173498
rect 575798 173440 578422 173496
rect 578478 173440 578483 173496
rect 575798 173438 578483 173440
rect 575798 173060 575858 173438
rect 578417 173435 578483 173438
rect 676029 173226 676095 173229
rect 676029 173224 676292 173226
rect 676029 173168 676034 173224
rect 676090 173168 676292 173224
rect 676029 173166 676292 173168
rect 676029 173163 676095 173166
rect 666356 172962 666938 173022
rect 666878 172954 666938 172962
rect 673913 172954 673979 172957
rect 666878 172952 673979 172954
rect 666878 172896 673918 172952
rect 673974 172896 673979 172952
rect 666878 172894 673979 172896
rect 673913 172891 673979 172894
rect 674833 172818 674899 172821
rect 674833 172816 676292 172818
rect 674833 172760 674838 172816
rect 674894 172760 676292 172816
rect 674833 172758 676292 172760
rect 674833 172755 674899 172758
rect 675886 172348 675892 172412
rect 675956 172410 675962 172412
rect 675956 172350 676292 172410
rect 675956 172348 675962 172350
rect 589457 172138 589523 172141
rect 589457 172136 592572 172138
rect 589457 172080 589462 172136
rect 589518 172080 592572 172136
rect 589457 172078 592572 172080
rect 589457 172075 589523 172078
rect 670601 172002 670667 172005
rect 670601 172000 676292 172002
rect 670601 171944 670606 172000
rect 670662 171944 676292 172000
rect 670601 171942 676292 171944
rect 670601 171939 670667 171942
rect 680997 171594 681063 171597
rect 680997 171592 681076 171594
rect 680997 171536 681002 171592
rect 681058 171536 681076 171592
rect 680997 171534 681076 171536
rect 680997 171531 681063 171534
rect 675017 171186 675083 171189
rect 675017 171184 676292 171186
rect 675017 171128 675022 171184
rect 675078 171128 676292 171184
rect 675017 171126 676292 171128
rect 675017 171123 675083 171126
rect 578233 171050 578299 171053
rect 575798 171048 578299 171050
rect 575798 170992 578238 171048
rect 578294 170992 578299 171048
rect 575798 170990 578299 170992
rect 575798 170884 575858 170990
rect 578233 170987 578299 170990
rect 676581 170778 676647 170781
rect 676581 170776 676660 170778
rect 676581 170720 676586 170776
rect 676642 170720 676660 170776
rect 676581 170718 676660 170720
rect 676581 170715 676647 170718
rect 589181 170506 589247 170509
rect 589181 170504 592572 170506
rect 589181 170448 589186 170504
rect 589242 170448 592572 170504
rect 589181 170446 592572 170448
rect 589181 170443 589247 170446
rect 675702 170308 675708 170372
rect 675772 170370 675778 170372
rect 675772 170310 676292 170370
rect 675772 170308 675778 170310
rect 671889 169962 671955 169965
rect 671889 169960 676292 169962
rect 671889 169904 671894 169960
rect 671950 169904 676292 169960
rect 671889 169902 676292 169904
rect 671889 169899 671955 169902
rect 666356 169698 666754 169758
rect 666694 169690 666754 169698
rect 668025 169690 668091 169693
rect 666694 169688 668091 169690
rect 666694 169632 668030 169688
rect 668086 169632 668091 169688
rect 666694 169630 668091 169632
rect 668025 169627 668091 169630
rect 670417 169554 670483 169557
rect 670417 169552 676292 169554
rect 670417 169496 670422 169552
rect 670478 169496 676292 169552
rect 670417 169494 676292 169496
rect 670417 169491 670483 169494
rect 578417 169282 578483 169285
rect 575798 169280 578483 169282
rect 575798 169224 578422 169280
rect 578478 169224 578483 169280
rect 575798 169222 578483 169224
rect 575798 168708 575858 169222
rect 578417 169219 578483 169222
rect 673177 169146 673243 169149
rect 673177 169144 676292 169146
rect 673177 169088 673182 169144
rect 673238 169088 676292 169144
rect 673177 169086 676292 169088
rect 673177 169083 673243 169086
rect 589825 168874 589891 168877
rect 589825 168872 592572 168874
rect 589825 168816 589830 168872
rect 589886 168816 592572 168872
rect 589825 168814 592572 168816
rect 589825 168811 589891 168814
rect 674465 168738 674531 168741
rect 674465 168736 676292 168738
rect 674465 168680 674470 168736
rect 674526 168680 676292 168736
rect 674465 168678 676292 168680
rect 674465 168675 674531 168678
rect 669773 168330 669839 168333
rect 669773 168328 676292 168330
rect 669773 168272 669778 168328
rect 669834 168272 676292 168328
rect 669773 168270 676292 168272
rect 669773 168267 669839 168270
rect 669221 168194 669287 168197
rect 666694 168192 669287 168194
rect 666694 168136 669226 168192
rect 669282 168136 669287 168192
rect 666694 168134 669287 168136
rect 666694 168126 666754 168134
rect 669221 168131 669287 168134
rect 666356 168066 666754 168126
rect 676029 167922 676095 167925
rect 676029 167920 676292 167922
rect 676029 167864 676034 167920
rect 676090 167864 676292 167920
rect 676029 167862 676292 167864
rect 676029 167859 676095 167862
rect 675886 167452 675892 167516
rect 675956 167514 675962 167516
rect 675956 167454 676292 167514
rect 675956 167452 675962 167454
rect 589457 167242 589523 167245
rect 589457 167240 592572 167242
rect 589457 167184 589462 167240
rect 589518 167184 592572 167240
rect 589457 167182 592572 167184
rect 589457 167179 589523 167182
rect 676170 167046 676292 167106
rect 579521 166970 579587 166973
rect 575798 166968 579587 166970
rect 575798 166912 579526 166968
rect 579582 166912 579587 166968
rect 575798 166910 579587 166912
rect 575798 166532 575858 166910
rect 579521 166907 579587 166910
rect 671705 166970 671771 166973
rect 676170 166970 676230 167046
rect 671705 166968 676230 166970
rect 671705 166912 671710 166968
rect 671766 166912 676230 166968
rect 671705 166910 676230 166912
rect 671705 166907 671771 166910
rect 676581 166428 676647 166429
rect 676581 166424 676628 166428
rect 676692 166426 676698 166428
rect 676581 166368 676586 166424
rect 676581 166364 676628 166368
rect 676692 166366 676738 166426
rect 676692 166364 676698 166366
rect 676581 166363 676647 166364
rect 589641 165610 589707 165613
rect 589641 165608 592572 165610
rect 589641 165552 589646 165608
rect 589702 165552 592572 165608
rect 589641 165550 592572 165552
rect 589641 165547 589707 165550
rect 670141 165066 670207 165069
rect 676029 165066 676095 165069
rect 670141 165064 676095 165066
rect 670141 165008 670146 165064
rect 670202 165008 676034 165064
rect 676090 165008 676095 165064
rect 670141 165006 676095 165008
rect 670141 165003 670207 165006
rect 676029 165003 676095 165006
rect 667933 164930 667999 164933
rect 666694 164928 667999 164930
rect 666694 164872 667938 164928
rect 667994 164872 667999 164928
rect 666694 164870 667999 164872
rect 666694 164862 666754 164870
rect 667933 164867 667999 164870
rect 666356 164802 666754 164862
rect 579521 164522 579587 164525
rect 575798 164520 579587 164522
rect 575798 164464 579526 164520
rect 579582 164464 579587 164520
rect 575798 164462 579587 164464
rect 575798 164356 575858 164462
rect 579521 164459 579587 164462
rect 669129 164250 669195 164253
rect 670734 164250 670740 164252
rect 669129 164248 670740 164250
rect 669129 164192 669134 164248
rect 669190 164192 670740 164248
rect 669129 164190 670740 164192
rect 669129 164187 669195 164190
rect 670734 164188 670740 164190
rect 670804 164188 670810 164252
rect 589457 163978 589523 163981
rect 589457 163976 592572 163978
rect 589457 163920 589462 163976
rect 589518 163920 592572 163976
rect 589457 163918 592572 163920
rect 589457 163915 589523 163918
rect 668945 163298 669011 163301
rect 666694 163296 669011 163298
rect 666694 163240 668950 163296
rect 669006 163240 669011 163296
rect 666694 163238 669011 163240
rect 666694 163230 666754 163238
rect 668945 163235 669011 163238
rect 666356 163170 666754 163230
rect 579337 162754 579403 162757
rect 575798 162752 579403 162754
rect 575798 162696 579342 162752
rect 579398 162696 579403 162752
rect 575798 162694 579403 162696
rect 575798 162180 575858 162694
rect 579337 162691 579403 162694
rect 590561 162346 590627 162349
rect 590561 162344 592572 162346
rect 590561 162288 590566 162344
rect 590622 162288 592572 162344
rect 590561 162286 592572 162288
rect 590561 162283 590627 162286
rect 675201 161394 675267 161397
rect 675845 161394 675911 161397
rect 675201 161392 675911 161394
rect 675201 161336 675206 161392
rect 675262 161336 675850 161392
rect 675906 161336 675911 161392
rect 675201 161334 675911 161336
rect 675201 161331 675267 161334
rect 675845 161331 675911 161334
rect 589457 160714 589523 160717
rect 589457 160712 592572 160714
rect 589457 160656 589462 160712
rect 589518 160656 592572 160712
rect 589457 160654 592572 160656
rect 589457 160651 589523 160654
rect 667933 160034 667999 160037
rect 666694 160032 667999 160034
rect 575982 159898 576042 160004
rect 666694 159976 667938 160032
rect 667994 159976 667999 160032
rect 666694 159974 667999 159976
rect 666694 159966 666754 159974
rect 667933 159971 667999 159974
rect 666356 159906 666754 159966
rect 578233 159898 578299 159901
rect 575982 159896 578299 159898
rect 575982 159840 578238 159896
rect 578294 159840 578299 159896
rect 575982 159838 578299 159840
rect 578233 159835 578299 159838
rect 675753 159354 675819 159357
rect 676438 159354 676444 159356
rect 675753 159352 676444 159354
rect 675753 159296 675758 159352
rect 675814 159296 676444 159352
rect 675753 159294 676444 159296
rect 675753 159291 675819 159294
rect 676438 159292 676444 159294
rect 676508 159292 676514 159356
rect 588537 159082 588603 159085
rect 588537 159080 592572 159082
rect 588537 159024 588542 159080
rect 588598 159024 592572 159080
rect 588537 159022 592572 159024
rect 588537 159019 588603 159022
rect 578417 158402 578483 158405
rect 671521 158402 671587 158405
rect 575798 158400 578483 158402
rect 575798 158344 578422 158400
rect 578478 158344 578483 158400
rect 575798 158342 578483 158344
rect 575798 157828 575858 158342
rect 578417 158339 578483 158342
rect 666694 158400 671587 158402
rect 666694 158344 671526 158400
rect 671582 158344 671587 158400
rect 666694 158342 671587 158344
rect 666694 158334 666754 158342
rect 671521 158339 671587 158342
rect 666356 158274 666754 158334
rect 674833 157586 674899 157589
rect 675477 157586 675543 157589
rect 674833 157584 675543 157586
rect 674833 157528 674838 157584
rect 674894 157528 675482 157584
rect 675538 157528 675543 157584
rect 674833 157526 675543 157528
rect 674833 157523 674899 157526
rect 675477 157523 675543 157526
rect 589273 157450 589339 157453
rect 589273 157448 592572 157450
rect 589273 157392 589278 157448
rect 589334 157392 592572 157448
rect 589273 157390 592572 157392
rect 589273 157387 589339 157390
rect 675753 156362 675819 156365
rect 676622 156362 676628 156364
rect 675753 156360 676628 156362
rect 675753 156304 675758 156360
rect 675814 156304 676628 156360
rect 675753 156302 676628 156304
rect 675753 156299 675819 156302
rect 676622 156300 676628 156302
rect 676692 156300 676698 156364
rect 578509 155954 578575 155957
rect 575798 155952 578575 155954
rect 575798 155896 578514 155952
rect 578570 155896 578575 155952
rect 575798 155894 578575 155896
rect 575798 155652 575858 155894
rect 578509 155891 578575 155894
rect 589457 155818 589523 155821
rect 589457 155816 592572 155818
rect 589457 155760 589462 155816
rect 589518 155760 592572 155816
rect 589457 155758 592572 155760
rect 589457 155755 589523 155758
rect 666356 155010 666938 155070
rect 666878 154594 666938 155010
rect 670417 154866 670483 154869
rect 675109 154866 675175 154869
rect 670417 154864 675175 154866
rect 670417 154808 670422 154864
rect 670478 154808 675114 154864
rect 675170 154808 675175 154864
rect 670417 154806 675175 154808
rect 670417 154803 670483 154806
rect 675109 154803 675175 154806
rect 674097 154594 674163 154597
rect 666878 154592 674163 154594
rect 666878 154536 674102 154592
rect 674158 154536 674163 154592
rect 666878 154534 674163 154536
rect 674097 154531 674163 154534
rect 589457 154186 589523 154189
rect 589457 154184 592572 154186
rect 589457 154128 589462 154184
rect 589518 154128 592572 154184
rect 589457 154126 592572 154128
rect 589457 154123 589523 154126
rect 578693 154050 578759 154053
rect 575798 154048 578759 154050
rect 575798 153992 578698 154048
rect 578754 153992 578759 154048
rect 575798 153990 578759 153992
rect 575798 153476 575858 153990
rect 578693 153987 578759 153990
rect 668761 153506 668827 153509
rect 666694 153504 668827 153506
rect 666694 153448 668766 153504
rect 668822 153448 668827 153504
rect 666694 153446 668827 153448
rect 666694 153438 666754 153446
rect 668761 153443 668827 153446
rect 666356 153378 666754 153438
rect 668761 153098 668827 153101
rect 672717 153098 672783 153101
rect 668761 153096 672783 153098
rect 668761 153040 668766 153096
rect 668822 153040 672722 153096
rect 672778 153040 672783 153096
rect 668761 153038 672783 153040
rect 668761 153035 668827 153038
rect 672717 153035 672783 153038
rect 589457 152554 589523 152557
rect 673177 152554 673243 152557
rect 675477 152554 675543 152557
rect 589457 152552 592572 152554
rect 589457 152496 589462 152552
rect 589518 152496 592572 152552
rect 589457 152494 592572 152496
rect 673177 152552 675543 152554
rect 673177 152496 673182 152552
rect 673238 152496 675482 152552
rect 675538 152496 675543 152552
rect 673177 152494 675543 152496
rect 589457 152491 589523 152494
rect 673177 152491 673243 152494
rect 675477 152491 675543 152494
rect 671889 151874 671955 151877
rect 675477 151874 675543 151877
rect 671889 151872 675543 151874
rect 671889 151816 671894 151872
rect 671950 151816 675482 151872
rect 675538 151816 675543 151872
rect 671889 151814 675543 151816
rect 671889 151811 671955 151814
rect 675477 151811 675543 151814
rect 578233 151738 578299 151741
rect 575798 151736 578299 151738
rect 575798 151680 578238 151736
rect 578294 151680 578299 151736
rect 575798 151678 578299 151680
rect 575798 151300 575858 151678
rect 578233 151675 578299 151678
rect 675293 151602 675359 151605
rect 676254 151602 676260 151604
rect 675293 151600 676260 151602
rect 675293 151544 675298 151600
rect 675354 151544 676260 151600
rect 675293 151542 676260 151544
rect 675293 151539 675359 151542
rect 676254 151540 676260 151542
rect 676324 151540 676330 151604
rect 674465 151058 674531 151061
rect 675109 151058 675175 151061
rect 674465 151056 675175 151058
rect 674465 151000 674470 151056
rect 674526 151000 675114 151056
rect 675170 151000 675175 151056
rect 674465 150998 675175 151000
rect 674465 150995 674531 150998
rect 675109 150995 675175 150998
rect 589917 150922 589983 150925
rect 589917 150920 592572 150922
rect 589917 150864 589922 150920
rect 589978 150864 592572 150920
rect 589917 150862 592572 150864
rect 589917 150859 589983 150862
rect 675661 150380 675727 150381
rect 675661 150376 675708 150380
rect 675772 150378 675778 150380
rect 675661 150320 675666 150376
rect 675661 150316 675708 150320
rect 675772 150318 675818 150378
rect 675772 150316 675778 150318
rect 675661 150315 675727 150316
rect 668301 150242 668367 150245
rect 666694 150240 668367 150242
rect 666694 150184 668306 150240
rect 668362 150184 668367 150240
rect 666694 150182 668367 150184
rect 666694 150174 666754 150182
rect 668301 150179 668367 150182
rect 666356 150114 666754 150174
rect 578325 149698 578391 149701
rect 575798 149696 578391 149698
rect 575798 149640 578330 149696
rect 578386 149640 578391 149696
rect 575798 149638 578391 149640
rect 575798 149124 575858 149638
rect 578325 149635 578391 149638
rect 589181 149290 589247 149293
rect 589181 149288 592572 149290
rect 589181 149232 589186 149288
rect 589242 149232 592572 149288
rect 589181 149230 592572 149232
rect 589181 149227 589247 149230
rect 670601 149018 670667 149021
rect 675293 149018 675359 149021
rect 670601 149016 675359 149018
rect 670601 148960 670606 149016
rect 670662 148960 675298 149016
rect 675354 148960 675359 149016
rect 670601 148958 675359 148960
rect 670601 148955 670667 148958
rect 675293 148955 675359 148958
rect 668485 148610 668551 148613
rect 666694 148608 668551 148610
rect 666694 148552 668490 148608
rect 668546 148552 668551 148608
rect 666694 148550 668551 148552
rect 666694 148542 666754 148550
rect 668485 148547 668551 148550
rect 666356 148482 666754 148542
rect 675753 148474 675819 148477
rect 676070 148474 676076 148476
rect 675753 148472 676076 148474
rect 675753 148416 675758 148472
rect 675814 148416 676076 148472
rect 675753 148414 676076 148416
rect 675753 148411 675819 148414
rect 676070 148412 676076 148414
rect 676140 148412 676146 148476
rect 589457 147658 589523 147661
rect 675661 147658 675727 147661
rect 675886 147658 675892 147660
rect 589457 147656 592572 147658
rect 589457 147600 589462 147656
rect 589518 147600 592572 147656
rect 589457 147598 592572 147600
rect 675661 147656 675892 147658
rect 675661 147600 675666 147656
rect 675722 147600 675892 147656
rect 675661 147598 675892 147600
rect 589457 147595 589523 147598
rect 675661 147595 675727 147598
rect 675886 147596 675892 147598
rect 675956 147596 675962 147660
rect 579521 147522 579587 147525
rect 575798 147520 579587 147522
rect 575798 147464 579526 147520
rect 579582 147464 579587 147520
rect 575798 147462 579587 147464
rect 575798 146948 575858 147462
rect 579521 147459 579587 147462
rect 588721 146026 588787 146029
rect 588721 146024 592572 146026
rect 588721 145968 588726 146024
rect 588782 145968 592572 146024
rect 588721 145966 592572 145968
rect 588721 145963 588787 145966
rect 671286 145346 671292 145348
rect 666694 145286 671292 145346
rect 666694 145278 666754 145286
rect 671286 145284 671292 145286
rect 671356 145284 671362 145348
rect 666356 145218 666754 145278
rect 575982 144666 576042 144772
rect 579429 144666 579495 144669
rect 575982 144664 579495 144666
rect 575982 144608 579434 144664
rect 579490 144608 579495 144664
rect 575982 144606 579495 144608
rect 579429 144603 579495 144606
rect 589457 144394 589523 144397
rect 589457 144392 592572 144394
rect 589457 144336 589462 144392
rect 589518 144336 592572 144392
rect 589457 144334 592572 144336
rect 589457 144331 589523 144334
rect 669129 143714 669195 143717
rect 666694 143712 669195 143714
rect 666694 143656 669134 143712
rect 669190 143656 669195 143712
rect 666694 143654 669195 143656
rect 666694 143646 666754 143654
rect 669129 143651 669195 143654
rect 666356 143586 666754 143646
rect 579521 143034 579587 143037
rect 575798 143032 579587 143034
rect 575798 142976 579526 143032
rect 579582 142976 579587 143032
rect 575798 142974 579587 142976
rect 575798 142596 575858 142974
rect 579521 142971 579587 142974
rect 589641 142762 589707 142765
rect 667381 142762 667447 142765
rect 683297 142762 683363 142765
rect 589641 142760 592572 142762
rect 589641 142704 589646 142760
rect 589702 142704 592572 142760
rect 589641 142702 592572 142704
rect 667381 142760 683363 142762
rect 667381 142704 667386 142760
rect 667442 142704 683302 142760
rect 683358 142704 683363 142760
rect 667381 142702 683363 142704
rect 589641 142699 589707 142702
rect 667381 142699 667447 142702
rect 683297 142699 683363 142702
rect 589457 141130 589523 141133
rect 669221 141130 669287 141133
rect 673678 141130 673684 141132
rect 589457 141128 592572 141130
rect 589457 141072 589462 141128
rect 589518 141072 592572 141128
rect 589457 141070 592572 141072
rect 669221 141128 673684 141130
rect 669221 141072 669226 141128
rect 669282 141072 673684 141128
rect 669221 141070 673684 141072
rect 589457 141067 589523 141070
rect 669221 141067 669287 141070
rect 673678 141068 673684 141070
rect 673748 141068 673754 141132
rect 579521 140586 579587 140589
rect 575798 140584 579587 140586
rect 575798 140528 579526 140584
rect 579582 140528 579587 140584
rect 575798 140526 579587 140528
rect 575798 140420 575858 140526
rect 579521 140523 579587 140526
rect 672073 140450 672139 140453
rect 666694 140448 672139 140450
rect 666694 140392 672078 140448
rect 672134 140392 672139 140448
rect 666694 140390 672139 140392
rect 666694 140382 666754 140390
rect 672073 140387 672139 140390
rect 666356 140322 666754 140382
rect 589457 139498 589523 139501
rect 589457 139496 592572 139498
rect 589457 139440 589462 139496
rect 589518 139440 592572 139496
rect 589457 139438 592572 139440
rect 589457 139435 589523 139438
rect 578601 138818 578667 138821
rect 669221 138818 669287 138821
rect 575798 138816 578667 138818
rect 575798 138760 578606 138816
rect 578662 138760 578667 138816
rect 575798 138758 578667 138760
rect 575798 138244 575858 138758
rect 578601 138755 578667 138758
rect 666694 138816 669287 138818
rect 666694 138760 669226 138816
rect 669282 138760 669287 138816
rect 666694 138758 669287 138760
rect 666694 138750 666754 138758
rect 669221 138755 669287 138758
rect 666356 138690 666754 138750
rect 588537 137866 588603 137869
rect 667933 137866 667999 137869
rect 669262 137866 669268 137868
rect 588537 137864 592572 137866
rect 588537 137808 588542 137864
rect 588598 137808 592572 137864
rect 588537 137806 592572 137808
rect 667933 137864 669268 137866
rect 667933 137808 667938 137864
rect 667994 137808 669268 137864
rect 667933 137806 669268 137808
rect 588537 137803 588603 137806
rect 667933 137803 667999 137806
rect 669262 137804 669268 137806
rect 669332 137804 669338 137868
rect 578877 136642 578943 136645
rect 575798 136640 578943 136642
rect 575798 136584 578882 136640
rect 578938 136584 578943 136640
rect 575798 136582 578943 136584
rect 575798 136068 575858 136582
rect 578877 136579 578943 136582
rect 589457 136234 589523 136237
rect 589457 136232 592572 136234
rect 589457 136176 589462 136232
rect 589518 136176 592572 136232
rect 589457 136174 592572 136176
rect 589457 136171 589523 136174
rect 667565 135962 667631 135965
rect 683113 135962 683179 135965
rect 667565 135960 683179 135962
rect 667565 135904 667570 135960
rect 667626 135904 683118 135960
rect 683174 135904 683179 135960
rect 667565 135902 683179 135904
rect 667565 135899 667631 135902
rect 683113 135899 683179 135902
rect 667933 135554 667999 135557
rect 666694 135552 667999 135554
rect 666694 135496 667938 135552
rect 667994 135496 667999 135552
rect 666694 135494 667999 135496
rect 666694 135486 666754 135494
rect 667933 135491 667999 135494
rect 666356 135426 666754 135486
rect 590285 134602 590351 134605
rect 590285 134600 592572 134602
rect 590285 134544 590290 134600
rect 590346 134544 592572 134600
rect 590285 134542 592572 134544
rect 590285 134539 590351 134542
rect 579521 134466 579587 134469
rect 575798 134464 579587 134466
rect 575798 134408 579526 134464
rect 579582 134408 579587 134464
rect 575798 134406 579587 134408
rect 575798 133892 575858 134406
rect 579521 134403 579587 134406
rect 673126 133922 673132 133924
rect 667982 133862 673132 133922
rect 666356 133794 666938 133854
rect 666878 133650 666938 133794
rect 667982 133650 668042 133862
rect 673126 133860 673132 133862
rect 673196 133860 673202 133924
rect 666878 133590 668042 133650
rect 667013 133106 667079 133109
rect 676262 133106 676322 133348
rect 683297 133106 683363 133109
rect 667013 133104 676322 133106
rect 667013 133048 667018 133104
rect 667074 133048 676322 133104
rect 667013 133046 676322 133048
rect 683254 133104 683363 133106
rect 683254 133048 683302 133104
rect 683358 133048 683363 133104
rect 667013 133043 667079 133046
rect 683254 133043 683363 133048
rect 589917 132970 589983 132973
rect 589917 132968 592572 132970
rect 589917 132912 589922 132968
rect 589978 132912 592572 132968
rect 683254 132940 683314 133043
rect 589917 132910 592572 132912
rect 589917 132907 589983 132910
rect 683113 132698 683179 132701
rect 683070 132696 683179 132698
rect 683070 132640 683118 132696
rect 683174 132640 683179 132696
rect 683070 132635 683179 132640
rect 683070 132532 683130 132635
rect 579061 132290 579127 132293
rect 575798 132288 579127 132290
rect 575798 132232 579066 132288
rect 579122 132232 579127 132288
rect 575798 132230 579127 132232
rect 575798 131716 575858 132230
rect 579061 132227 579127 132230
rect 674281 132154 674347 132157
rect 674281 132152 676292 132154
rect 674281 132096 674286 132152
rect 674342 132096 676292 132152
rect 674281 132094 676292 132096
rect 674281 132091 674347 132094
rect 671337 131746 671403 131749
rect 671337 131744 676292 131746
rect 671337 131688 671342 131744
rect 671398 131688 676292 131744
rect 671337 131686 676292 131688
rect 671337 131683 671403 131686
rect 590101 131338 590167 131341
rect 674649 131338 674715 131341
rect 590101 131336 592572 131338
rect 590101 131280 590106 131336
rect 590162 131280 592572 131336
rect 590101 131278 592572 131280
rect 674649 131336 676292 131338
rect 674649 131280 674654 131336
rect 674710 131280 676292 131336
rect 674649 131278 676292 131280
rect 590101 131275 590167 131278
rect 674649 131275 674715 131278
rect 671521 130930 671587 130933
rect 671521 130928 676292 130930
rect 671521 130872 671526 130928
rect 671582 130872 676292 130928
rect 671521 130870 676292 130872
rect 671521 130867 671587 130870
rect 667974 130658 667980 130660
rect 666694 130598 667980 130658
rect 666694 130590 666754 130598
rect 667974 130596 667980 130598
rect 668044 130596 668050 130660
rect 666356 130530 666754 130590
rect 672533 130522 672599 130525
rect 672533 130520 676292 130522
rect 672533 130464 672538 130520
rect 672594 130464 676292 130520
rect 672533 130462 676292 130464
rect 672533 130459 672599 130462
rect 676213 130250 676279 130253
rect 676213 130248 676322 130250
rect 676213 130192 676218 130248
rect 676274 130192 676322 130248
rect 676213 130187 676322 130192
rect 676262 130084 676322 130187
rect 578693 129706 578759 129709
rect 575798 129704 578759 129706
rect 575798 129648 578698 129704
rect 578754 129648 578759 129704
rect 575798 129646 578759 129648
rect 575798 129540 575858 129646
rect 578693 129643 578759 129646
rect 589273 129706 589339 129709
rect 673361 129706 673427 129709
rect 589273 129704 592572 129706
rect 589273 129648 589278 129704
rect 589334 129648 592572 129704
rect 589273 129646 592572 129648
rect 673361 129704 676292 129706
rect 673361 129648 673366 129704
rect 673422 129648 676292 129704
rect 673361 129646 676292 129648
rect 589273 129643 589339 129646
rect 673361 129643 673427 129646
rect 674097 129298 674163 129301
rect 674097 129296 676292 129298
rect 674097 129240 674102 129296
rect 674158 129240 676292 129296
rect 674097 129238 676292 129240
rect 674097 129235 674163 129238
rect 666356 128898 666938 128958
rect 666878 128890 666938 128898
rect 673494 128890 673500 128892
rect 666878 128830 673500 128890
rect 673494 128828 673500 128830
rect 673564 128828 673570 128892
rect 676262 128620 676322 128860
rect 676254 128556 676260 128620
rect 676324 128556 676330 128620
rect 668945 128346 669011 128349
rect 674046 128346 674052 128348
rect 668945 128344 674052 128346
rect 668945 128288 668950 128344
rect 669006 128288 674052 128344
rect 668945 128286 674052 128288
rect 668945 128283 669011 128286
rect 674046 128284 674052 128286
rect 674116 128284 674122 128348
rect 676814 128213 676874 128452
rect 674281 128210 674347 128213
rect 676213 128210 676279 128213
rect 674281 128208 676279 128210
rect 674281 128152 674286 128208
rect 674342 128152 676218 128208
rect 676274 128152 676279 128208
rect 674281 128150 676279 128152
rect 676814 128208 676923 128213
rect 676814 128152 676862 128208
rect 676918 128152 676923 128208
rect 676814 128150 676923 128152
rect 674281 128147 674347 128150
rect 676213 128147 676279 128150
rect 676857 128147 676923 128150
rect 589457 128074 589523 128077
rect 589457 128072 592572 128074
rect 589457 128016 589462 128072
rect 589518 128016 592572 128072
rect 589457 128014 592572 128016
rect 589457 128011 589523 128014
rect 679574 127805 679634 128044
rect 578509 127802 578575 127805
rect 575798 127800 578575 127802
rect 575798 127744 578514 127800
rect 578570 127744 578575 127800
rect 575798 127742 578575 127744
rect 679574 127800 679683 127805
rect 679574 127744 679622 127800
rect 679678 127744 679683 127800
rect 679574 127742 679683 127744
rect 575798 127364 575858 127742
rect 578509 127739 578575 127742
rect 679617 127739 679683 127742
rect 674833 127666 674899 127669
rect 674833 127664 676292 127666
rect 674833 127608 674838 127664
rect 674894 127608 676292 127664
rect 674833 127606 676292 127608
rect 674833 127603 674899 127606
rect 676070 126924 676076 126988
rect 676140 126986 676146 126988
rect 676262 126986 676322 127228
rect 676140 126926 676322 126986
rect 676140 126924 676146 126926
rect 676630 126580 676690 126820
rect 676622 126516 676628 126580
rect 676692 126516 676698 126580
rect 589457 126442 589523 126445
rect 675017 126442 675083 126445
rect 589457 126440 592572 126442
rect 589457 126384 589462 126440
rect 589518 126384 592572 126440
rect 589457 126382 592572 126384
rect 675017 126440 676292 126442
rect 675017 126384 675022 126440
rect 675078 126384 676292 126440
rect 675017 126382 676292 126384
rect 589457 126379 589523 126382
rect 675017 126379 675083 126382
rect 672349 126034 672415 126037
rect 672349 126032 676292 126034
rect 672349 125976 672354 126032
rect 672410 125976 676292 126032
rect 672349 125974 676292 125976
rect 672349 125971 672415 125974
rect 668761 125762 668827 125765
rect 666694 125760 668827 125762
rect 666694 125704 668766 125760
rect 668822 125704 668827 125760
rect 666694 125702 668827 125704
rect 666694 125694 666754 125702
rect 668761 125699 668827 125702
rect 666356 125634 666754 125694
rect 674649 125626 674715 125629
rect 674649 125624 676292 125626
rect 674649 125568 674654 125624
rect 674710 125568 676292 125624
rect 674649 125566 676292 125568
rect 674649 125563 674715 125566
rect 579521 125354 579587 125357
rect 575798 125352 579587 125354
rect 575798 125296 579526 125352
rect 579582 125296 579587 125352
rect 575798 125294 579587 125296
rect 575798 125188 575858 125294
rect 579521 125291 579587 125294
rect 674465 125218 674531 125221
rect 674465 125216 676292 125218
rect 674465 125160 674470 125216
rect 674526 125160 676292 125216
rect 674465 125158 676292 125160
rect 674465 125155 674531 125158
rect 589733 124810 589799 124813
rect 589733 124808 592572 124810
rect 589733 124752 589738 124808
rect 589794 124752 592572 124808
rect 589733 124750 592572 124752
rect 589733 124747 589799 124750
rect 676446 124540 676506 124780
rect 676438 124476 676444 124540
rect 676508 124476 676514 124540
rect 673177 124402 673243 124405
rect 673177 124400 676292 124402
rect 673177 124344 673182 124400
rect 673238 124344 676292 124400
rect 673177 124342 676292 124344
rect 673177 124339 673243 124342
rect 672901 124130 672967 124133
rect 666694 124128 672967 124130
rect 666694 124072 672906 124128
rect 672962 124072 672967 124128
rect 666694 124070 672967 124072
rect 666694 124062 666754 124070
rect 672901 124067 672967 124070
rect 666356 124002 666754 124062
rect 673134 123934 676292 123994
rect 672901 123858 672967 123861
rect 673134 123858 673194 123934
rect 672901 123856 673194 123858
rect 672901 123800 672906 123856
rect 672962 123800 673194 123856
rect 672901 123798 673194 123800
rect 672901 123795 672967 123798
rect 579245 123586 579311 123589
rect 575798 123584 579311 123586
rect 575798 123528 579250 123584
rect 579306 123528 579311 123584
rect 575798 123526 579311 123528
rect 575798 123012 575858 123526
rect 579245 123523 579311 123526
rect 673361 123586 673427 123589
rect 673361 123584 676292 123586
rect 673361 123528 673366 123584
rect 673422 123528 676292 123584
rect 673361 123526 676292 123528
rect 673361 123523 673427 123526
rect 589457 123178 589523 123181
rect 672717 123178 672783 123181
rect 589457 123176 592572 123178
rect 589457 123120 589462 123176
rect 589518 123120 592572 123176
rect 589457 123118 592572 123120
rect 672717 123176 676292 123178
rect 672717 123120 672722 123176
rect 672778 123120 676292 123176
rect 672717 123118 676292 123120
rect 589457 123115 589523 123118
rect 672717 123115 672783 123118
rect 672533 122770 672599 122773
rect 672533 122768 676292 122770
rect 672533 122712 672538 122768
rect 672594 122712 676292 122768
rect 672533 122710 676292 122712
rect 672533 122707 672599 122710
rect 675886 122300 675892 122364
rect 675956 122362 675962 122364
rect 675956 122302 676292 122362
rect 675956 122300 675962 122302
rect 669221 122226 669287 122229
rect 672717 122226 672783 122229
rect 669221 122224 672783 122226
rect 669221 122168 669226 122224
rect 669282 122168 672722 122224
rect 672778 122168 672783 122224
rect 669221 122166 672783 122168
rect 669221 122163 669287 122166
rect 672717 122163 672783 122166
rect 676262 121682 676322 121924
rect 675894 121622 676322 121682
rect 589273 121546 589339 121549
rect 589273 121544 592572 121546
rect 589273 121488 589278 121544
rect 589334 121488 592572 121544
rect 589273 121486 592572 121488
rect 589273 121483 589339 121486
rect 669957 121410 670023 121413
rect 675894 121410 675954 121622
rect 669957 121408 675954 121410
rect 669957 121352 669962 121408
rect 670018 121352 675954 121408
rect 669957 121350 675954 121352
rect 669957 121347 670023 121350
rect 578509 121138 578575 121141
rect 575798 121136 578575 121138
rect 575798 121080 578514 121136
rect 578570 121080 578575 121136
rect 575798 121078 578575 121080
rect 575798 120836 575858 121078
rect 578509 121075 578575 121078
rect 668945 120866 669011 120869
rect 666694 120864 669011 120866
rect 666694 120808 668950 120864
rect 669006 120808 669011 120864
rect 666694 120806 669011 120808
rect 666694 120798 666754 120806
rect 668945 120803 669011 120806
rect 666356 120738 666754 120798
rect 588721 119914 588787 119917
rect 588721 119912 592572 119914
rect 588721 119856 588726 119912
rect 588782 119856 592572 119912
rect 588721 119854 592572 119856
rect 588721 119851 588787 119854
rect 667933 119234 667999 119237
rect 666694 119232 667999 119234
rect 666694 119176 667938 119232
rect 667994 119176 667999 119232
rect 666694 119174 667999 119176
rect 666694 119166 666754 119174
rect 667933 119171 667999 119174
rect 666356 119106 666754 119166
rect 575982 118418 576042 118660
rect 579521 118418 579587 118421
rect 575982 118416 579587 118418
rect 575982 118360 579526 118416
rect 579582 118360 579587 118416
rect 575982 118358 579587 118360
rect 579521 118355 579587 118358
rect 589457 118282 589523 118285
rect 589457 118280 592572 118282
rect 589457 118224 589462 118280
rect 589518 118224 592572 118280
rect 589457 118222 592572 118224
rect 589457 118219 589523 118222
rect 667933 117602 667999 117605
rect 666694 117600 667999 117602
rect 666694 117544 667938 117600
rect 667994 117544 667999 117600
rect 666694 117542 667999 117544
rect 666694 117534 666754 117542
rect 667933 117539 667999 117542
rect 666356 117474 666754 117534
rect 675702 117268 675708 117332
rect 675772 117330 675778 117332
rect 676857 117330 676923 117333
rect 675772 117328 676923 117330
rect 675772 117272 676862 117328
rect 676918 117272 676923 117328
rect 675772 117270 676923 117272
rect 675772 117268 675778 117270
rect 676857 117267 676923 117270
rect 579337 116922 579403 116925
rect 575798 116920 579403 116922
rect 575798 116864 579342 116920
rect 579398 116864 579403 116920
rect 575798 116862 579403 116864
rect 575798 116484 575858 116862
rect 579337 116859 579403 116862
rect 589457 116650 589523 116653
rect 589457 116648 592572 116650
rect 589457 116592 589462 116648
rect 589518 116592 592572 116648
rect 589457 116590 592572 116592
rect 589457 116587 589523 116590
rect 666356 115842 666754 115902
rect 666694 115834 666754 115842
rect 671705 115834 671771 115837
rect 666694 115832 671771 115834
rect 666694 115776 671710 115832
rect 671766 115776 671771 115832
rect 666694 115774 671771 115776
rect 671705 115771 671771 115774
rect 589549 115018 589615 115021
rect 589549 115016 592572 115018
rect 589549 114960 589554 115016
rect 589610 114960 592572 115016
rect 589549 114958 592572 114960
rect 589549 114955 589615 114958
rect 578509 114474 578575 114477
rect 575798 114472 578575 114474
rect 575798 114416 578514 114472
rect 578570 114416 578575 114472
rect 575798 114414 578575 114416
rect 575798 114308 575858 114414
rect 578509 114411 578575 114414
rect 669221 114338 669287 114341
rect 666694 114336 669287 114338
rect 666694 114280 669226 114336
rect 669282 114280 669287 114336
rect 666694 114278 669287 114280
rect 666694 114270 666754 114278
rect 669221 114275 669287 114278
rect 666356 114210 666754 114270
rect 590285 113386 590351 113389
rect 590285 113384 592572 113386
rect 590285 113328 590290 113384
rect 590346 113328 592572 113384
rect 590285 113326 592572 113328
rect 590285 113323 590351 113326
rect 675293 113114 675359 113117
rect 676254 113114 676260 113116
rect 675293 113112 676260 113114
rect 675293 113056 675298 113112
rect 675354 113056 676260 113112
rect 675293 113054 676260 113056
rect 675293 113051 675359 113054
rect 676254 113052 676260 113054
rect 676324 113052 676330 113116
rect 579521 112706 579587 112709
rect 672533 112706 672599 112709
rect 575798 112704 579587 112706
rect 575798 112648 579526 112704
rect 579582 112648 579587 112704
rect 575798 112646 579587 112648
rect 575798 112132 575858 112646
rect 579521 112643 579587 112646
rect 666694 112704 672599 112706
rect 666694 112648 672538 112704
rect 672594 112648 672599 112704
rect 666694 112646 672599 112648
rect 666694 112638 666754 112646
rect 672533 112643 672599 112646
rect 666356 112578 666754 112638
rect 589365 111754 589431 111757
rect 589365 111752 592572 111754
rect 589365 111696 589370 111752
rect 589426 111696 592572 111752
rect 589365 111694 592572 111696
rect 589365 111691 589431 111694
rect 672349 111482 672415 111485
rect 675109 111482 675175 111485
rect 672349 111480 675175 111482
rect 672349 111424 672354 111480
rect 672410 111424 675114 111480
rect 675170 111424 675175 111480
rect 672349 111422 675175 111424
rect 672349 111419 672415 111422
rect 675109 111419 675175 111422
rect 667933 111074 667999 111077
rect 666694 111072 667999 111074
rect 666694 111016 667938 111072
rect 667994 111016 667999 111072
rect 666694 111014 667999 111016
rect 666694 111006 666754 111014
rect 667933 111011 667999 111014
rect 668577 111074 668643 111077
rect 674097 111074 674163 111077
rect 668577 111072 674163 111074
rect 668577 111016 668582 111072
rect 668638 111016 674102 111072
rect 674158 111016 674163 111072
rect 668577 111014 674163 111016
rect 668577 111011 668643 111014
rect 674097 111011 674163 111014
rect 666356 110946 666754 111006
rect 578877 110394 578943 110397
rect 575798 110392 578943 110394
rect 575798 110336 578882 110392
rect 578938 110336 578943 110392
rect 575798 110334 578943 110336
rect 575798 109956 575858 110334
rect 578877 110331 578943 110334
rect 673177 110394 673243 110397
rect 675109 110394 675175 110397
rect 673177 110392 675175 110394
rect 673177 110336 673182 110392
rect 673238 110336 675114 110392
rect 675170 110336 675175 110392
rect 673177 110334 675175 110336
rect 673177 110331 673243 110334
rect 675109 110331 675175 110334
rect 590101 110122 590167 110125
rect 590101 110120 592572 110122
rect 590101 110064 590106 110120
rect 590162 110064 592572 110120
rect 590101 110062 592572 110064
rect 590101 110059 590167 110062
rect 666356 109314 666754 109374
rect 666694 109306 666754 109314
rect 667933 109306 667999 109309
rect 666694 109304 667999 109306
rect 666694 109248 667938 109304
rect 667994 109248 667999 109304
rect 666694 109246 667999 109248
rect 667933 109243 667999 109246
rect 589457 108490 589523 108493
rect 589457 108488 592572 108490
rect 589457 108432 589462 108488
rect 589518 108432 592572 108488
rect 589457 108430 592572 108432
rect 589457 108427 589523 108430
rect 578325 108354 578391 108357
rect 575798 108352 578391 108354
rect 575798 108296 578330 108352
rect 578386 108296 578391 108352
rect 575798 108294 578391 108296
rect 575798 107780 575858 108294
rect 578325 108291 578391 108294
rect 675753 108218 675819 108221
rect 676070 108218 676076 108220
rect 675753 108216 676076 108218
rect 675753 108160 675758 108216
rect 675814 108160 676076 108216
rect 675753 108158 676076 108160
rect 675753 108155 675819 108158
rect 676070 108156 676076 108158
rect 676140 108156 676146 108220
rect 671521 107810 671587 107813
rect 666694 107808 671587 107810
rect 666694 107752 671526 107808
rect 671582 107752 671587 107808
rect 666694 107750 671587 107752
rect 666694 107742 666754 107750
rect 671521 107747 671587 107750
rect 666356 107682 666754 107742
rect 589457 106858 589523 106861
rect 589457 106856 592572 106858
rect 589457 106800 589462 106856
rect 589518 106800 592572 106856
rect 589457 106798 592572 106800
rect 589457 106795 589523 106798
rect 672809 106314 672875 106317
rect 675109 106314 675175 106317
rect 672809 106312 675175 106314
rect 672809 106256 672814 106312
rect 672870 106256 675114 106312
rect 675170 106256 675175 106312
rect 672809 106254 675175 106256
rect 672809 106251 672875 106254
rect 675109 106251 675175 106254
rect 668117 106178 668183 106181
rect 668393 106178 668459 106181
rect 666694 106176 668459 106178
rect 666694 106120 668122 106176
rect 668178 106120 668398 106176
rect 668454 106120 668459 106176
rect 666694 106118 668459 106120
rect 666694 106110 666754 106118
rect 668117 106115 668183 106118
rect 668393 106115 668459 106118
rect 675753 106178 675819 106181
rect 676438 106178 676444 106180
rect 675753 106176 676444 106178
rect 675753 106120 675758 106176
rect 675814 106120 676444 106176
rect 675753 106118 676444 106120
rect 675753 106115 675819 106118
rect 676438 106116 676444 106118
rect 676508 106116 676514 106180
rect 666356 106050 666754 106110
rect 579061 105906 579127 105909
rect 575798 105904 579127 105906
rect 575798 105848 579066 105904
rect 579122 105848 579127 105904
rect 575798 105846 579127 105848
rect 575798 105604 575858 105846
rect 579061 105843 579127 105846
rect 673361 105634 673427 105637
rect 675109 105634 675175 105637
rect 673361 105632 675175 105634
rect 673361 105576 673366 105632
rect 673422 105576 675114 105632
rect 675170 105576 675175 105632
rect 673361 105574 675175 105576
rect 673361 105571 673427 105574
rect 675109 105571 675175 105574
rect 589825 105226 589891 105229
rect 589825 105224 592572 105226
rect 589825 105168 589830 105224
rect 589886 105168 592572 105224
rect 589825 105166 592572 105168
rect 589825 105163 589891 105166
rect 666356 104418 666754 104478
rect 666694 104410 666754 104418
rect 668577 104410 668643 104413
rect 666694 104408 668643 104410
rect 666694 104352 668582 104408
rect 668638 104352 668643 104408
rect 666694 104350 668643 104352
rect 668577 104347 668643 104350
rect 590285 103594 590351 103597
rect 590285 103592 592572 103594
rect 590285 103536 590290 103592
rect 590346 103536 592572 103592
rect 590285 103534 592572 103536
rect 590285 103531 590351 103534
rect 575982 103322 576042 103428
rect 579245 103322 579311 103325
rect 575982 103320 579311 103322
rect 575982 103264 579250 103320
rect 579306 103264 579311 103320
rect 575982 103262 579311 103264
rect 579245 103259 579311 103262
rect 675661 103188 675727 103189
rect 675661 103184 675708 103188
rect 675772 103186 675778 103188
rect 675661 103128 675666 103184
rect 675661 103124 675708 103128
rect 675772 103126 675818 103186
rect 675772 103124 675778 103126
rect 675661 103123 675727 103124
rect 666645 102846 666711 102849
rect 666356 102844 666711 102846
rect 666356 102788 666650 102844
rect 666706 102788 666711 102844
rect 666356 102786 666711 102788
rect 666645 102783 666711 102786
rect 675661 102506 675727 102509
rect 675886 102506 675892 102508
rect 675661 102504 675892 102506
rect 675661 102448 675666 102504
rect 675722 102448 675892 102504
rect 675661 102446 675892 102448
rect 675661 102443 675727 102446
rect 675886 102444 675892 102446
rect 675956 102444 675962 102508
rect 666645 102370 666711 102373
rect 674281 102370 674347 102373
rect 666645 102368 674347 102370
rect 666645 102312 666650 102368
rect 666706 102312 674286 102368
rect 674342 102312 674347 102368
rect 666645 102310 674347 102312
rect 666645 102307 666711 102310
rect 674281 102307 674347 102310
rect 589917 101962 589983 101965
rect 589917 101960 592572 101962
rect 589917 101904 589922 101960
rect 589978 101904 592572 101960
rect 589917 101902 592572 101904
rect 589917 101899 589983 101902
rect 578325 101690 578391 101693
rect 575798 101688 578391 101690
rect 575798 101632 578330 101688
rect 578386 101632 578391 101688
rect 575798 101630 578391 101632
rect 575798 101252 575858 101630
rect 578325 101627 578391 101630
rect 675753 101418 675819 101421
rect 676622 101418 676628 101420
rect 675753 101416 676628 101418
rect 675753 101360 675758 101416
rect 675814 101360 676628 101416
rect 675753 101358 676628 101360
rect 675753 101355 675819 101358
rect 676622 101356 676628 101358
rect 676692 101356 676698 101420
rect 578601 99378 578667 99381
rect 575798 99376 578667 99378
rect 575798 99320 578606 99376
rect 578662 99320 578667 99376
rect 575798 99318 578667 99320
rect 575798 99076 575858 99318
rect 578601 99315 578667 99318
rect 579245 97474 579311 97477
rect 575798 97472 579311 97474
rect 575798 97416 579250 97472
rect 579306 97416 579311 97472
rect 575798 97414 579311 97416
rect 575798 96900 575858 97414
rect 579245 97411 579311 97414
rect 637021 96930 637087 96933
rect 637246 96930 637252 96932
rect 637021 96928 637252 96930
rect 637021 96872 637026 96928
rect 637082 96872 637252 96928
rect 637021 96870 637252 96872
rect 637021 96867 637087 96870
rect 637246 96868 637252 96870
rect 637316 96868 637322 96932
rect 635549 96386 635615 96389
rect 647417 96386 647483 96389
rect 635549 96384 647483 96386
rect 635549 96328 635554 96384
rect 635610 96328 647422 96384
rect 647478 96328 647483 96384
rect 635549 96326 647483 96328
rect 635549 96323 635615 96326
rect 647417 96323 647483 96326
rect 633934 96052 633940 96116
rect 634004 96114 634010 96116
rect 635733 96114 635799 96117
rect 634004 96112 635799 96114
rect 634004 96056 635738 96112
rect 635794 96056 635799 96112
rect 634004 96054 635799 96056
rect 634004 96052 634010 96054
rect 635733 96051 635799 96054
rect 641989 96114 642055 96117
rect 647182 96114 647188 96116
rect 641989 96112 647188 96114
rect 641989 96056 641994 96112
rect 642050 96056 647188 96112
rect 641989 96054 647188 96056
rect 641989 96051 642055 96054
rect 647182 96052 647188 96054
rect 647252 96052 647258 96116
rect 611997 95842 612063 95845
rect 668301 95842 668367 95845
rect 611997 95840 668367 95842
rect 611997 95784 612002 95840
rect 612058 95784 668306 95840
rect 668362 95784 668367 95840
rect 611997 95782 668367 95784
rect 611997 95779 612063 95782
rect 668301 95779 668367 95782
rect 579245 95026 579311 95029
rect 575798 95024 579311 95026
rect 575798 94968 579250 95024
rect 579306 94968 579311 95024
rect 575798 94966 579311 94968
rect 575798 94724 575858 94966
rect 579245 94963 579311 94966
rect 647141 95026 647207 95029
rect 647141 95024 647434 95026
rect 647141 94968 647146 95024
rect 647202 94968 647434 95024
rect 647141 94966 647434 94968
rect 647141 94963 647207 94966
rect 626441 94482 626507 94485
rect 626441 94480 628268 94482
rect 626441 94424 626446 94480
rect 626502 94424 628268 94480
rect 647374 94452 647434 94966
rect 626441 94422 628268 94424
rect 626441 94419 626507 94422
rect 655053 94210 655119 94213
rect 655053 94208 656788 94210
rect 655053 94152 655058 94208
rect 655114 94152 656788 94208
rect 655053 94150 656788 94152
rect 655053 94147 655119 94150
rect 625981 93666 626047 93669
rect 625981 93664 628268 93666
rect 625981 93608 625986 93664
rect 626042 93608 628268 93664
rect 625981 93606 628268 93608
rect 625981 93603 626047 93606
rect 655421 93394 655487 93397
rect 665357 93394 665423 93397
rect 655421 93392 656788 93394
rect 655421 93336 655426 93392
rect 655482 93336 656788 93392
rect 655421 93334 656788 93336
rect 663596 93392 665423 93394
rect 663596 93336 665362 93392
rect 665418 93336 665423 93392
rect 663596 93334 665423 93336
rect 655421 93331 655487 93334
rect 665357 93331 665423 93334
rect 579337 93122 579403 93125
rect 575798 93120 579403 93122
rect 575798 93064 579342 93120
rect 579398 93064 579403 93120
rect 575798 93062 579403 93064
rect 575798 92548 575858 93062
rect 579337 93059 579403 93062
rect 650310 93060 650316 93124
rect 650380 93122 650386 93124
rect 650380 93062 656818 93122
rect 650380 93060 650386 93062
rect 626441 92850 626507 92853
rect 626441 92848 628268 92850
rect 626441 92792 626446 92848
rect 626502 92792 628268 92848
rect 626441 92790 628268 92792
rect 626441 92787 626507 92790
rect 656758 92548 656818 93062
rect 663701 92850 663767 92853
rect 663382 92848 663767 92850
rect 663382 92792 663706 92848
rect 663762 92792 663767 92848
rect 663382 92790 663767 92792
rect 663382 92548 663442 92790
rect 663701 92787 663767 92790
rect 625797 92034 625863 92037
rect 648613 92034 648679 92037
rect 625797 92032 628268 92034
rect 625797 91976 625802 92032
rect 625858 91976 628268 92032
rect 625797 91974 628268 91976
rect 648140 92032 648679 92034
rect 648140 91976 648618 92032
rect 648674 91976 648679 92032
rect 648140 91974 648679 91976
rect 625797 91971 625863 91974
rect 648613 91971 648679 91974
rect 664529 91762 664595 91765
rect 663596 91760 664595 91762
rect 663596 91704 664534 91760
rect 664590 91704 664595 91760
rect 663596 91702 664595 91704
rect 664529 91699 664595 91702
rect 654685 91490 654751 91493
rect 654685 91488 656788 91490
rect 654685 91432 654690 91488
rect 654746 91432 656788 91488
rect 654685 91430 656788 91432
rect 654685 91427 654751 91430
rect 626441 91218 626507 91221
rect 626441 91216 628268 91218
rect 626441 91160 626446 91216
rect 626502 91160 628268 91216
rect 626441 91158 628268 91160
rect 626441 91155 626507 91158
rect 578233 90946 578299 90949
rect 575798 90944 578299 90946
rect 575798 90888 578238 90944
rect 578294 90888 578299 90944
rect 575798 90886 578299 90888
rect 575798 90372 575858 90886
rect 578233 90883 578299 90886
rect 655421 90674 655487 90677
rect 664161 90674 664227 90677
rect 655421 90672 656788 90674
rect 655421 90616 655426 90672
rect 655482 90616 656788 90672
rect 655421 90614 656788 90616
rect 663596 90672 664227 90674
rect 663596 90616 664166 90672
rect 664222 90616 664227 90672
rect 663596 90614 664227 90616
rect 655421 90611 655487 90614
rect 664161 90611 664227 90614
rect 626441 90402 626507 90405
rect 626441 90400 628268 90402
rect 626441 90344 626446 90400
rect 626502 90344 628268 90400
rect 626441 90342 628268 90344
rect 626441 90339 626507 90342
rect 655789 89858 655855 89861
rect 664345 89858 664411 89861
rect 655789 89856 656788 89858
rect 655789 89800 655794 89856
rect 655850 89800 656788 89856
rect 655789 89798 656788 89800
rect 663596 89856 664411 89858
rect 663596 89800 664350 89856
rect 664406 89800 664411 89856
rect 663596 89798 664411 89800
rect 655789 89795 655855 89798
rect 664345 89795 664411 89798
rect 626441 89586 626507 89589
rect 650177 89586 650243 89589
rect 626441 89584 628268 89586
rect 626441 89528 626446 89584
rect 626502 89528 628268 89584
rect 626441 89526 628268 89528
rect 648140 89584 650243 89586
rect 648140 89528 650182 89584
rect 650238 89528 650243 89584
rect 648140 89526 650243 89528
rect 626441 89523 626507 89526
rect 650177 89523 650243 89526
rect 665173 89042 665239 89045
rect 663596 89040 665239 89042
rect 663596 88984 665178 89040
rect 665234 88984 665239 89040
rect 663596 88982 665239 88984
rect 665173 88979 665239 88982
rect 625429 88770 625495 88773
rect 625429 88768 628268 88770
rect 625429 88712 625434 88768
rect 625490 88712 628268 88768
rect 625429 88710 628268 88712
rect 625429 88707 625495 88710
rect 575982 88090 576042 88196
rect 579337 88090 579403 88093
rect 575982 88088 579403 88090
rect 575982 88032 579342 88088
rect 579398 88032 579403 88088
rect 575982 88030 579403 88032
rect 579337 88027 579403 88030
rect 626257 87954 626323 87957
rect 626257 87952 628268 87954
rect 626257 87896 626262 87952
rect 626318 87896 628268 87952
rect 626257 87894 628268 87896
rect 626257 87891 626323 87894
rect 626441 87138 626507 87141
rect 650545 87138 650611 87141
rect 626441 87136 628268 87138
rect 626441 87080 626446 87136
rect 626502 87080 628268 87136
rect 626441 87078 628268 87080
rect 648140 87136 650611 87138
rect 648140 87080 650550 87136
rect 650606 87080 650611 87136
rect 648140 87078 650611 87080
rect 626441 87075 626507 87078
rect 650545 87075 650611 87078
rect 578785 86458 578851 86461
rect 575798 86456 578851 86458
rect 575798 86400 578790 86456
rect 578846 86400 578851 86456
rect 575798 86398 578851 86400
rect 575798 86020 575858 86398
rect 578785 86395 578851 86398
rect 626441 86322 626507 86325
rect 626441 86320 628268 86322
rect 626441 86264 626446 86320
rect 626502 86264 628268 86320
rect 626441 86262 628268 86264
rect 626441 86259 626507 86262
rect 626441 85506 626507 85509
rect 626441 85504 628268 85506
rect 626441 85448 626446 85504
rect 626502 85448 628268 85504
rect 626441 85446 628268 85448
rect 626441 85443 626507 85446
rect 625245 84690 625311 84693
rect 649993 84690 650059 84693
rect 625245 84688 628268 84690
rect 625245 84632 625250 84688
rect 625306 84632 628268 84688
rect 625245 84630 628268 84632
rect 648140 84688 650059 84690
rect 648140 84632 649998 84688
rect 650054 84632 650059 84688
rect 648140 84630 650059 84632
rect 625245 84627 625311 84630
rect 649993 84627 650059 84630
rect 579337 84010 579403 84013
rect 575798 84008 579403 84010
rect 575798 83952 579342 84008
rect 579398 83952 579403 84008
rect 575798 83950 579403 83952
rect 575798 83844 575858 83950
rect 579337 83947 579403 83950
rect 625797 83874 625863 83877
rect 625797 83872 628268 83874
rect 625797 83816 625802 83872
rect 625858 83816 628268 83872
rect 625797 83814 628268 83816
rect 625797 83811 625863 83814
rect 628741 83330 628807 83333
rect 628741 83328 628850 83330
rect 628741 83272 628746 83328
rect 628802 83272 628850 83328
rect 628741 83267 628850 83272
rect 628790 83028 628850 83267
rect 578693 82242 578759 82245
rect 648889 82242 648955 82245
rect 575798 82240 578759 82242
rect 575798 82184 578698 82240
rect 578754 82184 578759 82240
rect 648140 82240 648955 82242
rect 575798 82182 578759 82184
rect 575798 81668 575858 82182
rect 578693 82179 578759 82182
rect 628790 81698 628850 82212
rect 648140 82184 648894 82240
rect 648950 82184 648955 82240
rect 648140 82182 648955 82184
rect 648889 82179 648955 82182
rect 629201 81698 629267 81701
rect 628790 81696 629267 81698
rect 628790 81640 629206 81696
rect 629262 81640 629267 81696
rect 628790 81638 629267 81640
rect 629201 81635 629267 81638
rect 579521 80066 579587 80069
rect 575798 80064 579587 80066
rect 575798 80008 579526 80064
rect 579582 80008 579587 80064
rect 575798 80006 579587 80008
rect 575798 79492 575858 80006
rect 579521 80003 579587 80006
rect 633893 78572 633959 78573
rect 633893 78570 633940 78572
rect 633848 78568 633940 78570
rect 633848 78512 633898 78568
rect 633848 78510 633940 78512
rect 633893 78508 633940 78510
rect 634004 78508 634010 78572
rect 633893 78507 633959 78508
rect 578601 77890 578667 77893
rect 575798 77888 578667 77890
rect 575798 77832 578606 77888
rect 578662 77832 578667 77888
rect 575798 77830 578667 77832
rect 575798 77316 575858 77830
rect 578601 77827 578667 77830
rect 625797 77754 625863 77757
rect 637062 77754 637068 77756
rect 625797 77752 637068 77754
rect 625797 77696 625802 77752
rect 625858 77696 637068 77752
rect 625797 77694 637068 77696
rect 625797 77691 625863 77694
rect 637062 77692 637068 77694
rect 637132 77754 637138 77756
rect 639597 77754 639663 77757
rect 637132 77752 639663 77754
rect 637132 77696 639602 77752
rect 639658 77696 639663 77752
rect 637132 77694 639663 77696
rect 637132 77692 637138 77694
rect 639597 77691 639663 77694
rect 617517 77346 617583 77349
rect 633893 77346 633959 77349
rect 617517 77344 633959 77346
rect 617517 77288 617522 77344
rect 617578 77288 633898 77344
rect 633954 77288 633959 77344
rect 617517 77286 633959 77288
rect 617517 77283 617583 77286
rect 633893 77283 633959 77286
rect 578877 75714 578943 75717
rect 575798 75712 578943 75714
rect 575798 75656 578882 75712
rect 578938 75656 578943 75712
rect 575798 75654 578943 75656
rect 575798 75140 575858 75654
rect 578877 75651 578943 75654
rect 646497 74218 646563 74221
rect 646454 74216 646563 74218
rect 646454 74160 646502 74216
rect 646558 74160 646563 74216
rect 646454 74155 646563 74160
rect 646454 73848 646514 74155
rect 579521 73130 579587 73133
rect 575798 73128 579587 73130
rect 575798 73072 579526 73128
rect 579582 73072 579587 73128
rect 575798 73070 579587 73072
rect 575798 72964 575858 73070
rect 579521 73067 579587 73070
rect 648981 71770 649047 71773
rect 646638 71768 649047 71770
rect 646638 71712 648986 71768
rect 649042 71712 649047 71768
rect 646638 71710 649047 71712
rect 646638 71400 646698 71710
rect 648981 71707 649047 71710
rect 579245 71226 579311 71229
rect 575798 71224 579311 71226
rect 575798 71168 579250 71224
rect 579306 71168 579311 71224
rect 575798 71166 579311 71168
rect 575798 70788 575858 71166
rect 579245 71163 579311 71166
rect 646865 68982 646931 68985
rect 646668 68980 646931 68982
rect 646668 68924 646870 68980
rect 646926 68924 646931 68980
rect 646668 68922 646931 68924
rect 646865 68919 646931 68922
rect 646129 67146 646195 67149
rect 646086 67144 646195 67146
rect 646086 67088 646134 67144
rect 646190 67088 646195 67144
rect 646086 67083 646195 67088
rect 646086 66504 646146 67083
rect 575982 66330 576042 66436
rect 579521 66330 579587 66333
rect 575982 66328 579587 66330
rect 575982 66272 579526 66328
rect 579582 66272 579587 66328
rect 575982 66270 579587 66272
rect 579521 66267 579587 66270
rect 579061 64834 579127 64837
rect 575798 64832 579127 64834
rect 575798 64776 579066 64832
rect 579122 64776 579127 64832
rect 575798 64774 579127 64776
rect 575798 64260 575858 64774
rect 579061 64771 579127 64774
rect 649165 64426 649231 64429
rect 646638 64424 649231 64426
rect 646638 64368 649170 64424
rect 649226 64368 649231 64424
rect 646638 64366 649231 64368
rect 646638 64056 646698 64366
rect 649165 64363 649231 64366
rect 648613 62114 648679 62117
rect 646638 62112 648679 62114
rect 575982 61842 576042 62084
rect 646638 62056 648618 62112
rect 648674 62056 648679 62112
rect 646638 62054 648679 62056
rect 578509 61842 578575 61845
rect 575982 61840 578575 61842
rect 575982 61784 578514 61840
rect 578570 61784 578575 61840
rect 575982 61782 578575 61784
rect 578509 61779 578575 61782
rect 646638 61608 646698 62054
rect 648613 62051 648679 62054
rect 579521 60346 579587 60349
rect 575798 60344 579587 60346
rect 575798 60288 579526 60344
rect 579582 60288 579587 60344
rect 575798 60286 579587 60288
rect 575798 59908 575858 60286
rect 579521 60283 579587 60286
rect 646313 59394 646379 59397
rect 646270 59392 646379 59394
rect 646270 59336 646318 59392
rect 646374 59336 646379 59392
rect 646270 59331 646379 59336
rect 646270 59160 646330 59331
rect 579521 57898 579587 57901
rect 575798 57896 579587 57898
rect 575798 57840 579526 57896
rect 579582 57840 579587 57896
rect 575798 57838 579587 57840
rect 575798 57732 575858 57838
rect 579521 57835 579587 57838
rect 647233 57354 647299 57357
rect 646638 57352 647299 57354
rect 646638 57296 647238 57352
rect 647294 57296 647299 57352
rect 646638 57294 647299 57296
rect 646638 56712 646698 57294
rect 647233 57291 647299 57294
rect 579521 56130 579587 56133
rect 575798 56128 579587 56130
rect 575798 56072 579526 56128
rect 579582 56072 579587 56128
rect 575798 56070 579587 56072
rect 575798 55556 575858 56070
rect 579521 56067 579587 56070
rect 462589 52322 462655 52325
rect 466637 52322 466703 52325
rect 462589 52320 466703 52322
rect 462589 52264 462594 52320
rect 462650 52264 466642 52320
rect 466698 52264 466703 52320
rect 462589 52262 466703 52264
rect 462589 52259 462655 52262
rect 466637 52259 466703 52262
rect 461761 52050 461827 52053
rect 461761 52048 470610 52050
rect 461761 51992 461766 52048
rect 461822 51992 470610 52048
rect 461761 51990 470610 51992
rect 461761 51987 461827 51990
rect 470550 51914 470610 51990
rect 603073 51914 603139 51917
rect 470550 51912 603139 51914
rect 470550 51856 603078 51912
rect 603134 51856 603139 51912
rect 470550 51854 603139 51856
rect 603073 51851 603139 51854
rect 43437 51778 43503 51781
rect 129181 51778 129247 51781
rect 43437 51776 129247 51778
rect 43437 51720 43442 51776
rect 43498 51720 129186 51776
rect 129242 51720 129247 51776
rect 43437 51718 129247 51720
rect 43437 51715 43503 51718
rect 129181 51715 129247 51718
rect 466637 51642 466703 51645
rect 604453 51642 604519 51645
rect 466637 51640 604519 51642
rect 466637 51584 466642 51640
rect 466698 51584 604458 51640
rect 604514 51584 604519 51640
rect 466637 51582 604519 51584
rect 466637 51579 466703 51582
rect 604453 51579 604519 51582
rect 194358 50220 194364 50284
rect 194428 50282 194434 50284
rect 308029 50282 308095 50285
rect 194428 50280 308095 50282
rect 194428 50224 308034 50280
rect 308090 50224 308095 50280
rect 194428 50222 308095 50224
rect 194428 50220 194434 50222
rect 308029 50219 308095 50222
rect 522798 49404 522804 49468
rect 522868 49466 522874 49468
rect 545665 49466 545731 49469
rect 522868 49464 545731 49466
rect 522868 49408 545670 49464
rect 545726 49408 545731 49464
rect 522868 49406 545731 49408
rect 522868 49404 522874 49406
rect 545665 49403 545731 49406
rect 529790 49132 529796 49196
rect 529860 49194 529866 49196
rect 553669 49194 553735 49197
rect 529860 49192 553735 49194
rect 529860 49136 553674 49192
rect 553730 49136 553735 49192
rect 529860 49134 553735 49136
rect 529860 49132 529866 49134
rect 553669 49131 553735 49134
rect 518750 48860 518756 48924
rect 518820 48922 518826 48924
rect 549989 48922 550055 48925
rect 518820 48920 550055 48922
rect 518820 48864 549994 48920
rect 550050 48864 550055 48920
rect 518820 48862 550055 48864
rect 518820 48860 518826 48862
rect 549989 48859 550055 48862
rect 662413 48514 662479 48517
rect 662094 48512 662479 48514
rect 661480 48456 662418 48512
rect 662474 48456 662479 48512
rect 661480 48454 662479 48456
rect 661480 48452 662154 48454
rect 662413 48451 662479 48454
rect 458081 48242 458147 48245
rect 466453 48242 466519 48245
rect 458081 48240 466519 48242
rect 458081 48184 458086 48240
rect 458142 48184 466458 48240
rect 466514 48184 466519 48240
rect 458081 48182 466519 48184
rect 458081 48179 458147 48182
rect 466453 48179 466519 48182
rect 457897 47970 457963 47973
rect 466637 47970 466703 47973
rect 457897 47968 466703 47970
rect 457897 47912 457902 47968
rect 457958 47912 466642 47968
rect 466698 47912 466703 47968
rect 457897 47910 466703 47912
rect 457897 47907 457963 47910
rect 466637 47907 466703 47910
rect 526478 47772 526484 47836
rect 526548 47834 526554 47836
rect 552013 47834 552079 47837
rect 526548 47832 552079 47834
rect 526548 47776 552018 47832
rect 552074 47776 552079 47832
rect 661585 47791 661651 47794
rect 526548 47774 552079 47776
rect 526548 47772 526554 47774
rect 552013 47771 552079 47774
rect 661388 47789 661651 47791
rect 661388 47733 661590 47789
rect 661646 47733 661651 47789
rect 661388 47731 661651 47733
rect 661585 47728 661651 47731
rect 457713 47698 457779 47701
rect 466821 47698 466887 47701
rect 457713 47696 466887 47698
rect 457713 47640 457718 47696
rect 457774 47640 466826 47696
rect 466882 47640 466887 47696
rect 457713 47638 466887 47640
rect 457713 47635 457779 47638
rect 466821 47635 466887 47638
rect 520958 47500 520964 47564
rect 521028 47562 521034 47564
rect 547873 47562 547939 47565
rect 521028 47560 547939 47562
rect 521028 47504 547878 47560
rect 547934 47504 547939 47560
rect 521028 47502 547939 47504
rect 521028 47500 521034 47502
rect 547873 47499 547939 47502
rect 459001 47426 459067 47429
rect 467005 47426 467071 47429
rect 662597 47426 662663 47429
rect 459001 47424 467071 47426
rect 459001 47368 459006 47424
rect 459062 47368 467010 47424
rect 467066 47368 467071 47424
rect 459001 47366 467071 47368
rect 661388 47424 662663 47426
rect 661388 47368 662602 47424
rect 662658 47368 662663 47424
rect 661388 47366 662663 47368
rect 459001 47363 459067 47366
rect 467005 47363 467071 47366
rect 662597 47363 662663 47366
rect 515438 46956 515444 47020
rect 515508 47018 515514 47020
rect 521101 47018 521167 47021
rect 515508 47016 521167 47018
rect 515508 46960 521106 47016
rect 521162 46960 521167 47016
rect 515508 46958 521167 46960
rect 515508 46956 515514 46958
rect 521101 46955 521167 46958
rect 458265 46882 458331 46885
rect 465073 46882 465139 46885
rect 458265 46880 465139 46882
rect 458265 46824 458270 46880
rect 458326 46824 465078 46880
rect 465134 46824 465139 46880
rect 458265 46822 465139 46824
rect 458265 46819 458331 46822
rect 465073 46819 465139 46822
rect 458449 46610 458515 46613
rect 465257 46610 465323 46613
rect 458449 46608 465323 46610
rect 458449 46552 458454 46608
rect 458510 46552 465262 46608
rect 465318 46552 465323 46608
rect 458449 46550 465323 46552
rect 458449 46547 458515 46550
rect 465257 46547 465323 46550
rect 431217 44842 431283 44845
rect 460105 44842 460171 44845
rect 431217 44840 460171 44842
rect 431217 44784 431222 44840
rect 431278 44784 460110 44840
rect 460166 44784 460171 44840
rect 431217 44782 460171 44784
rect 431217 44779 431283 44782
rect 460105 44779 460171 44782
rect 463693 44436 463759 44437
rect 463693 44432 463740 44436
rect 463804 44434 463810 44436
rect 463693 44376 463698 44432
rect 463693 44372 463740 44376
rect 463804 44374 463850 44434
rect 463804 44372 463810 44374
rect 463693 44371 463759 44372
rect 130469 44298 130535 44301
rect 132585 44298 132651 44301
rect 142613 44298 142679 44301
rect 130469 44296 132651 44298
rect 130469 44240 130474 44296
rect 130530 44240 132590 44296
rect 132646 44240 132651 44296
rect 130469 44238 132651 44240
rect 130469 44235 130535 44238
rect 132585 44235 132651 44238
rect 142110 44296 142679 44298
rect 142110 44240 142618 44296
rect 142674 44240 142679 44296
rect 142110 44238 142679 44240
rect 141734 43964 141740 44028
rect 141804 44026 141810 44028
rect 142110 44026 142170 44238
rect 142613 44235 142679 44238
rect 464102 44236 464108 44300
rect 464172 44298 464178 44300
rect 464705 44298 464771 44301
rect 464172 44296 464771 44298
rect 464172 44240 464710 44296
rect 464766 44240 464771 44296
rect 464172 44238 464771 44240
rect 464172 44236 464178 44238
rect 464705 44235 464771 44238
rect 307293 44162 307359 44165
rect 463877 44162 463943 44165
rect 307293 44160 463943 44162
rect 307293 44104 307298 44160
rect 307354 44104 463882 44160
rect 463938 44104 463943 44160
rect 307293 44102 463943 44104
rect 307293 44099 307359 44102
rect 463877 44099 463943 44102
rect 141804 43966 142170 44026
rect 141804 43964 141810 43966
rect 419717 43890 419783 43893
rect 440182 43890 440188 43892
rect 419717 43888 440188 43890
rect 419717 43832 419722 43888
rect 419778 43832 440188 43888
rect 419717 43830 440188 43832
rect 419717 43827 419783 43830
rect 440182 43828 440188 43830
rect 440252 43828 440258 43892
rect 440918 43828 440924 43892
rect 440988 43890 440994 43892
rect 462865 43890 462931 43893
rect 440988 43888 462931 43890
rect 440988 43832 462870 43888
rect 462926 43832 462931 43888
rect 440988 43830 462931 43832
rect 440988 43828 440994 43830
rect 462865 43827 462931 43830
rect 415393 43618 415459 43621
rect 439589 43618 439655 43621
rect 415393 43616 439655 43618
rect 415393 43560 415398 43616
rect 415454 43560 439594 43616
rect 439650 43560 439655 43616
rect 415393 43558 439655 43560
rect 415393 43555 415459 43558
rect 439589 43555 439655 43558
rect 441613 43618 441679 43621
rect 461577 43618 461643 43621
rect 441613 43616 461643 43618
rect 441613 43560 441618 43616
rect 441674 43560 461582 43616
rect 461638 43560 461643 43616
rect 441613 43558 461643 43560
rect 441613 43555 441679 43558
rect 461577 43555 461643 43558
rect 462681 43618 462747 43621
rect 465809 43618 465875 43621
rect 462681 43616 465875 43618
rect 462681 43560 462686 43616
rect 462742 43560 465814 43616
rect 465870 43560 465875 43616
rect 462681 43558 465875 43560
rect 462681 43555 462747 43558
rect 465809 43555 465875 43558
rect 460749 43346 460815 43349
rect 471053 43346 471119 43349
rect 460749 43344 471119 43346
rect 460749 43288 460754 43344
rect 460810 43288 471058 43344
rect 471114 43288 471119 43344
rect 460749 43286 471119 43288
rect 460749 43283 460815 43286
rect 471053 43283 471119 43286
rect 461393 42938 461459 42941
rect 463693 42938 463759 42941
rect 461393 42936 463759 42938
rect 461393 42880 461398 42936
rect 461454 42880 463698 42936
rect 463754 42880 463759 42936
rect 461393 42878 463759 42880
rect 461393 42875 461459 42878
rect 463693 42875 463759 42878
rect 518801 42804 518867 42805
rect 518750 42802 518756 42804
rect 518710 42742 518756 42802
rect 518820 42800 518867 42804
rect 518862 42744 518867 42800
rect 518750 42740 518756 42742
rect 518820 42740 518867 42744
rect 518801 42739 518867 42740
rect 460933 42394 460999 42397
rect 451230 42392 460999 42394
rect 451230 42336 460938 42392
rect 460994 42336 460999 42392
rect 451230 42334 460999 42336
rect 416681 42258 416747 42261
rect 446397 42258 446463 42261
rect 451230 42258 451290 42334
rect 460933 42331 460999 42334
rect 416681 42256 427830 42258
rect 416681 42200 416686 42256
rect 416742 42200 427830 42256
rect 416681 42198 427830 42200
rect 416681 42195 416747 42198
rect 194317 42124 194383 42125
rect 194317 42122 194364 42124
rect 194272 42120 194364 42122
rect 194272 42064 194322 42120
rect 194272 42062 194364 42064
rect 194317 42060 194364 42062
rect 194428 42060 194434 42124
rect 194317 42059 194383 42060
rect 361941 41852 362007 41853
rect 361941 41848 361988 41852
rect 362052 41850 362058 41852
rect 365161 41850 365227 41853
rect 365478 41850 365484 41852
rect 361941 41792 361946 41848
rect 361941 41788 361988 41792
rect 362052 41790 362098 41850
rect 365161 41848 365484 41850
rect 365161 41792 365166 41848
rect 365222 41792 365484 41848
rect 365161 41790 365484 41792
rect 362052 41788 362058 41790
rect 361941 41787 362007 41788
rect 365161 41787 365227 41790
rect 365478 41788 365484 41790
rect 365548 41788 365554 41852
rect 403014 41788 403020 41852
rect 403084 41850 403090 41852
rect 421966 41850 421972 41852
rect 403084 41790 421972 41850
rect 403084 41788 403090 41790
rect 421966 41788 421972 41790
rect 422036 41788 422042 41852
rect 427770 41578 427830 42198
rect 446397 42256 451290 42258
rect 446397 42200 446402 42256
rect 446458 42200 451290 42256
rect 446397 42198 451290 42200
rect 446397 42195 446463 42198
rect 515397 42124 515463 42125
rect 520917 42124 520983 42125
rect 515397 42122 515444 42124
rect 515352 42120 515444 42122
rect 515352 42064 515402 42120
rect 515352 42062 515444 42064
rect 515397 42060 515444 42062
rect 515508 42060 515514 42124
rect 520917 42122 520964 42124
rect 520872 42120 520964 42122
rect 520872 42064 520922 42120
rect 520872 42062 520964 42064
rect 520917 42060 520964 42062
rect 521028 42060 521034 42124
rect 522113 42122 522179 42125
rect 526437 42124 526503 42125
rect 522798 42122 522804 42124
rect 522113 42120 522804 42122
rect 522113 42064 522118 42120
rect 522174 42064 522804 42120
rect 522113 42062 522804 42064
rect 515397 42059 515463 42060
rect 520917 42059 520983 42060
rect 522113 42059 522179 42062
rect 522798 42060 522804 42062
rect 522868 42060 522874 42124
rect 526437 42122 526484 42124
rect 526392 42120 526484 42122
rect 526392 42064 526442 42120
rect 526392 42062 526484 42064
rect 526437 42060 526484 42062
rect 526548 42060 526554 42124
rect 529565 42122 529631 42125
rect 529790 42122 529796 42124
rect 529565 42120 529796 42122
rect 529565 42064 529570 42120
rect 529626 42064 529796 42120
rect 529565 42062 529796 42064
rect 526437 42059 526503 42060
rect 529565 42059 529631 42062
rect 529790 42060 529796 42062
rect 529860 42060 529866 42124
rect 441838 41788 441844 41852
rect 441908 41850 441914 41852
rect 460790 41850 460796 41852
rect 441908 41790 460796 41850
rect 441908 41788 441914 41790
rect 460790 41788 460796 41790
rect 460860 41788 460866 41852
rect 460974 41788 460980 41852
rect 461044 41850 461050 41852
rect 464102 41850 464108 41852
rect 461044 41790 464108 41850
rect 461044 41788 461050 41790
rect 464102 41788 464108 41790
rect 464172 41788 464178 41852
rect 446397 41578 446463 41581
rect 427770 41576 446463 41578
rect 427770 41520 446402 41576
rect 446458 41520 446463 41576
rect 427770 41518 446463 41520
rect 446397 41515 446463 41518
rect 141693 40492 141759 40493
rect 141693 40488 141740 40492
rect 141804 40490 141810 40492
rect 141693 40432 141698 40488
rect 141693 40428 141740 40432
rect 141804 40430 141850 40490
rect 141804 40428 141810 40430
rect 141693 40427 141759 40428
<< via3 >>
rect 84516 997188 84580 997252
rect 245700 997188 245764 997252
rect 293540 997188 293604 997252
rect 86540 996916 86604 996980
rect 293724 996916 293788 996980
rect 387932 997188 387996 997252
rect 482692 997188 482756 997252
rect 530164 997188 530228 997252
rect 627132 996916 627196 996980
rect 90220 996644 90284 996708
rect 141924 996644 141988 996708
rect 87828 996372 87892 996436
rect 86540 995616 86604 995620
rect 86540 995560 86554 995616
rect 86554 995560 86604 995616
rect 86540 995556 86604 995560
rect 87828 995616 87892 995620
rect 87828 995560 87842 995616
rect 87842 995560 87892 995616
rect 87828 995556 87892 995560
rect 90220 995616 90284 995620
rect 90220 995560 90234 995616
rect 90234 995560 90284 995616
rect 90220 995556 90284 995560
rect 84516 995072 84580 995076
rect 84516 995016 84530 995072
rect 84530 995016 84580 995072
rect 84516 995012 84580 995016
rect 141924 995420 141988 995484
rect 242020 996644 242084 996708
rect 288020 996644 288084 996708
rect 243860 996372 243924 996436
rect 172468 995344 172532 995348
rect 172468 995288 172482 995344
rect 172482 995288 172532 995344
rect 172468 995284 172532 995288
rect 242020 995480 242084 995484
rect 242020 995424 242034 995480
rect 242034 995424 242084 995480
rect 242020 995420 242084 995424
rect 243860 995480 243924 995484
rect 243860 995424 243874 995480
rect 243874 995424 243924 995480
rect 243860 995420 243924 995424
rect 293724 996372 293788 996436
rect 386644 996644 386708 996708
rect 476252 996644 476316 996708
rect 626580 996644 626644 996708
rect 295012 996508 295076 996572
rect 388116 996372 388180 996436
rect 288020 995752 288084 995756
rect 288020 995696 288034 995752
rect 288034 995696 288084 995752
rect 288020 995692 288084 995696
rect 293540 995752 293604 995756
rect 293540 995696 293554 995752
rect 293554 995696 293604 995752
rect 293540 995692 293604 995696
rect 295012 995752 295076 995756
rect 295012 995696 295062 995752
rect 295062 995696 295076 995752
rect 295012 995692 295076 995696
rect 386644 995752 386708 995756
rect 386644 995696 386694 995752
rect 386694 995696 386708 995752
rect 386644 995692 386708 995696
rect 387932 995752 387996 995756
rect 387932 995696 387946 995752
rect 387946 995696 387996 995752
rect 387932 995692 387996 995696
rect 388116 995752 388180 995756
rect 474780 996372 474844 996436
rect 388116 995696 388166 995752
rect 388166 995696 388180 995752
rect 388116 995692 388180 995696
rect 474780 995752 474844 995756
rect 474780 995696 474794 995752
rect 474794 995696 474844 995752
rect 474780 995692 474844 995696
rect 476252 995692 476316 995756
rect 479932 995692 479996 995756
rect 482692 995752 482756 995756
rect 482692 995696 482742 995752
rect 482742 995696 482756 995752
rect 482692 995692 482756 995696
rect 526300 996100 526364 996164
rect 525012 995828 525076 995892
rect 627868 996372 627932 996436
rect 530164 995480 530228 995484
rect 530164 995424 530214 995480
rect 530214 995424 530228 995480
rect 530164 995420 530228 995424
rect 525012 995284 525076 995348
rect 626580 995752 626644 995756
rect 626580 995696 626630 995752
rect 626630 995696 626644 995752
rect 626580 995692 626644 995696
rect 627132 995752 627196 995756
rect 627132 995696 627182 995752
rect 627182 995696 627196 995752
rect 627132 995692 627196 995696
rect 627868 995752 627932 995756
rect 627868 995696 627918 995752
rect 627918 995696 627932 995752
rect 627868 995692 627932 995696
rect 142292 994468 142356 994532
rect 526300 994800 526364 994804
rect 526300 994744 526350 994800
rect 526350 994744 526364 994800
rect 526300 994740 526364 994744
rect 536788 994800 536852 994804
rect 536788 994744 536802 994800
rect 536802 994744 536852 994800
rect 536788 994740 536852 994744
rect 142108 993924 142172 993988
rect 479932 993924 479996 993988
rect 572668 990932 572732 990996
rect 42012 967192 42076 967196
rect 42012 967136 42026 967192
rect 42026 967136 42076 967192
rect 42012 967132 42076 967136
rect 675340 966512 675404 966516
rect 675340 966456 675390 966512
rect 675390 966456 675404 966512
rect 675340 966452 675404 966456
rect 676812 964684 676876 964748
rect 676076 963324 676140 963388
rect 41460 962100 41524 962164
rect 41276 959788 41340 959852
rect 40540 959108 40604 959172
rect 42564 957884 42628 957948
rect 676996 957748 677060 957812
rect 676628 956388 676692 956452
rect 40724 955436 40788 955500
rect 41460 952172 41524 952236
rect 42564 951900 42628 951964
rect 41276 951764 41340 951828
rect 42012 951628 42076 951692
rect 675340 951552 675404 951556
rect 675340 951496 675390 951552
rect 675390 951496 675404 951552
rect 675340 951492 675404 951496
rect 676812 950676 676876 950740
rect 676076 949452 676140 949516
rect 41828 941020 41892 941084
rect 675156 938164 675220 938228
rect 674604 937348 674668 937412
rect 40172 937178 40236 937242
rect 41828 937212 41892 937276
rect 41828 936532 41892 936596
rect 41828 935716 41892 935780
rect 676628 931908 676692 931972
rect 676996 931500 677060 931564
rect 42012 911916 42076 911980
rect 42196 911644 42260 911708
rect 42012 885396 42076 885460
rect 42196 885124 42260 885188
rect 676812 876556 676876 876620
rect 676076 875876 676140 875940
rect 675156 873972 675220 874036
rect 673868 873156 673932 873220
rect 675156 866764 675220 866828
rect 40172 815594 40236 815658
rect 42012 811956 42076 812020
rect 41828 809100 41892 809164
rect 40540 808648 40604 808712
rect 41828 807256 41892 807260
rect 41828 807200 41842 807256
rect 41842 807200 41892 807256
rect 41828 807196 41892 807200
rect 41460 805564 41524 805628
rect 40724 805020 40788 805084
rect 40908 794412 40972 794476
rect 40724 793732 40788 793796
rect 40540 792508 40604 792572
rect 41644 789108 41708 789172
rect 41828 788700 41892 788764
rect 41460 788156 41524 788220
rect 674420 782988 674484 783052
rect 675340 780464 675404 780468
rect 675340 780408 675354 780464
rect 675354 780408 675404 780464
rect 675340 780404 675404 780408
rect 675524 778364 675588 778428
rect 674972 777200 675036 777204
rect 674972 777144 675022 777200
rect 675022 777144 675036 777200
rect 674972 777140 675036 777144
rect 675524 776248 675588 776252
rect 675524 776192 675538 776248
rect 675538 776192 675588 776248
rect 675524 776188 675588 776192
rect 675340 776112 675404 776116
rect 675340 776056 675354 776112
rect 675354 776056 675404 776112
rect 675340 776052 675404 776056
rect 674972 773332 675036 773396
rect 673868 772244 673932 772308
rect 41460 769796 41524 769860
rect 676076 768708 676140 768772
rect 675892 766532 675956 766596
rect 40908 765716 40972 765780
rect 40540 765308 40604 765372
rect 676076 765036 676140 765100
rect 40724 764900 40788 764964
rect 676812 761832 676876 761836
rect 676812 761776 676826 761832
rect 676826 761776 676876 761832
rect 676812 761772 676876 761776
rect 41644 759052 41708 759116
rect 41092 757964 41156 758028
rect 42380 757828 42444 757892
rect 42012 757692 42076 757756
rect 40356 757480 40420 757484
rect 40356 757424 40370 757480
rect 40370 757424 40420 757480
rect 40356 757420 40420 757424
rect 40356 755380 40420 755444
rect 42196 754836 42260 754900
rect 41092 753612 41156 753676
rect 42380 753340 42444 753404
rect 42196 752932 42260 752996
rect 42196 752040 42260 752044
rect 42196 751984 42246 752040
rect 42246 751984 42260 752040
rect 42196 751980 42260 751984
rect 40908 751028 40972 751092
rect 40724 750348 40788 750412
rect 40540 749396 40604 749460
rect 41460 746540 41524 746604
rect 41644 746268 41708 746332
rect 42196 745996 42260 746060
rect 41828 745044 41892 745108
rect 674604 741508 674668 741572
rect 674236 739332 674300 739396
rect 675892 728724 675956 728788
rect 676812 728724 676876 728788
rect 41828 726820 41892 726884
rect 676076 725732 676140 725796
rect 41828 722332 41892 722396
rect 40724 721708 40788 721772
rect 41644 721708 41708 721772
rect 40540 717980 40604 718044
rect 41828 717980 41892 718044
rect 41828 715396 41892 715460
rect 40908 714172 40972 714236
rect 42012 714172 42076 714236
rect 675892 711996 675956 712060
rect 40908 709820 40972 709884
rect 40724 709412 40788 709476
rect 674420 707508 674484 707572
rect 42012 706752 42076 706756
rect 42012 706696 42062 706752
rect 42062 706696 42076 706752
rect 42012 706692 42076 706696
rect 40540 704244 40604 704308
rect 41460 702476 41524 702540
rect 41828 702340 41892 702404
rect 41644 701524 41708 701588
rect 675340 696824 675404 696828
rect 675340 696768 675390 696824
rect 675390 696768 675404 696824
rect 675340 696764 675404 696768
rect 676812 694044 676876 694108
rect 674420 692956 674484 693020
rect 675340 685884 675404 685948
rect 41828 683572 41892 683636
rect 674604 682348 674668 682412
rect 674236 680988 674300 681052
rect 40724 678928 40788 678992
rect 40908 678928 40972 678992
rect 41828 678600 41892 678604
rect 41828 678544 41842 678600
rect 41842 678544 41892 678600
rect 41828 678540 41892 678544
rect 41828 672692 41892 672756
rect 41276 672480 41340 672484
rect 41276 672424 41326 672480
rect 41326 672424 41340 672480
rect 41276 672420 41340 672424
rect 42196 672208 42260 672212
rect 42196 672152 42210 672208
rect 42210 672152 42260 672208
rect 42196 672148 42260 672152
rect 40356 670924 40420 670988
rect 42012 669292 42076 669356
rect 41276 669020 41340 669084
rect 42196 668944 42260 668948
rect 42196 668888 42246 668944
rect 42246 668888 42260 668944
rect 42196 668884 42260 668888
rect 40356 668068 40420 668132
rect 42012 667720 42076 667724
rect 42012 667664 42026 667720
rect 42026 667664 42076 667720
rect 42012 667660 42076 667664
rect 40724 666980 40788 667044
rect 42012 665680 42076 665684
rect 42012 665624 42062 665680
rect 42062 665624 42076 665680
rect 42012 665620 42076 665624
rect 40540 665348 40604 665412
rect 42012 664048 42076 664052
rect 42012 663992 42026 664048
rect 42026 663992 42076 664048
rect 42012 663988 42076 663992
rect 42196 662900 42260 662964
rect 41460 659772 41524 659836
rect 42196 659016 42260 659020
rect 42196 658960 42210 659016
rect 42210 658960 42260 659016
rect 42196 658956 42260 658960
rect 41828 658548 41892 658612
rect 41644 658276 41708 658340
rect 675340 652836 675404 652900
rect 675524 651536 675588 651540
rect 675524 651480 675574 651536
rect 675574 651480 675588 651536
rect 675524 651476 675588 651480
rect 674972 645824 675036 645828
rect 674972 645768 675022 645824
rect 675022 645768 675036 645824
rect 674972 645764 675036 645768
rect 676996 644268 677060 644332
rect 674236 642152 674300 642156
rect 674236 642096 674250 642152
rect 674250 642096 674300 642152
rect 674236 642092 674300 642096
rect 674604 640732 674668 640796
rect 41460 640596 41524 640660
rect 674052 640460 674116 640524
rect 675156 639780 675220 639844
rect 41644 638964 41708 639028
rect 675156 637876 675220 637940
rect 675340 637876 675404 637940
rect 674972 637664 675036 637668
rect 674972 637608 674986 637664
rect 674986 637608 675036 637664
rect 674972 637604 675036 637608
rect 675524 637604 675588 637668
rect 674236 636788 674300 636852
rect 674052 636244 674116 636308
rect 40724 634884 40788 634948
rect 40540 634476 40604 634540
rect 674972 631348 675036 631412
rect 676076 631408 676140 631412
rect 676076 631352 676090 631408
rect 676090 631352 676140 631408
rect 676076 631348 676140 631352
rect 41828 630668 41892 630732
rect 42196 626588 42260 626652
rect 42012 625228 42076 625292
rect 42196 624472 42260 624476
rect 42196 624416 42210 624472
rect 42210 624416 42260 624472
rect 42196 624412 42260 624416
rect 40724 623732 40788 623796
rect 42012 623384 42076 623388
rect 42012 623328 42062 623384
rect 42062 623328 42076 623384
rect 42012 623324 42076 623328
rect 40540 620332 40604 620396
rect 676812 619108 676876 619172
rect 41644 618292 41708 618356
rect 42196 617672 42260 617676
rect 42196 617616 42246 617672
rect 42246 617616 42260 617672
rect 42196 617612 42260 617616
rect 674420 617340 674484 617404
rect 673868 616116 673932 616180
rect 42196 615904 42260 615908
rect 42196 615848 42210 615904
rect 42210 615848 42260 615904
rect 42196 615844 42260 615848
rect 41828 615436 41892 615500
rect 41460 614076 41524 614140
rect 675524 607880 675588 607884
rect 675524 607824 675538 607880
rect 675538 607824 675588 607880
rect 675524 607820 675588 607824
rect 674236 602924 674300 602988
rect 41828 597212 41892 597276
rect 41828 596396 41892 596460
rect 675340 595368 675404 595372
rect 675340 595312 675390 595368
rect 675390 595312 675404 595368
rect 675340 595308 675404 595312
rect 675524 593192 675588 593196
rect 675524 593136 675574 593192
rect 675574 593136 675588 593192
rect 675524 593132 675588 593136
rect 675156 592860 675220 592924
rect 675340 592104 675404 592108
rect 675340 592048 675354 592104
rect 675354 592048 675404 592104
rect 675340 592044 675404 592048
rect 676076 591636 676140 591700
rect 40724 589596 40788 589660
rect 40908 589460 40972 589524
rect 40540 589324 40604 589388
rect 42012 586800 42076 586804
rect 42012 586744 42062 586800
rect 42062 586744 42076 586800
rect 42012 586740 42076 586744
rect 676076 586196 676140 586260
rect 41828 584564 41892 584628
rect 42196 584292 42260 584356
rect 42012 581496 42076 581500
rect 42012 581440 42026 581496
rect 42026 581440 42076 581496
rect 42012 581436 42076 581440
rect 42196 580212 42260 580276
rect 40724 578172 40788 578236
rect 42564 577900 42628 577964
rect 40908 577492 40972 577556
rect 40540 576812 40604 576876
rect 42564 574092 42628 574156
rect 41460 573276 41524 573340
rect 676996 572732 677060 572796
rect 41644 572052 41708 572116
rect 41828 570208 41892 570212
rect 41828 570152 41842 570208
rect 41842 570152 41892 570208
rect 41828 570148 41892 570152
rect 675524 562728 675588 562732
rect 675524 562672 675538 562728
rect 675538 562672 675588 562728
rect 675524 562668 675588 562672
rect 675524 561232 675588 561236
rect 675524 561176 675538 561232
rect 675538 561176 675588 561232
rect 675524 561172 675588 561176
rect 676812 557500 676876 557564
rect 42196 553964 42260 554028
rect 42012 553148 42076 553212
rect 42380 551788 42444 551852
rect 676996 550292 677060 550356
rect 675156 550216 675220 550220
rect 675156 550160 675170 550216
rect 675170 550160 675220 550216
rect 675156 550156 675220 550160
rect 675156 547572 675220 547636
rect 676076 547572 676140 547636
rect 674236 547300 674300 547364
rect 675524 546076 675588 546140
rect 40724 545668 40788 545732
rect 675340 545532 675404 545596
rect 40540 545456 40604 545460
rect 40540 545400 40554 545456
rect 40554 545400 40604 545456
rect 40540 545396 40604 545400
rect 40724 538188 40788 538252
rect 40540 535196 40604 535260
rect 41644 530164 41708 530228
rect 41460 529620 41524 529684
rect 41828 529408 41892 529412
rect 41828 529352 41878 529408
rect 41878 529352 41892 529408
rect 41828 529348 41892 529352
rect 676996 503644 677060 503708
rect 676812 492764 676876 492828
rect 675892 488820 675956 488884
rect 674604 475356 674668 475420
rect 673868 455228 673932 455292
rect 675340 453732 675404 453796
rect 41828 425172 41892 425236
rect 42012 424764 42076 424828
rect 42012 421908 42076 421972
rect 41460 418780 41524 418844
rect 40724 418508 40788 418572
rect 40540 418236 40604 418300
rect 42012 418236 42076 418300
rect 675340 410484 675404 410548
rect 40724 409396 40788 409460
rect 41828 406328 41892 406332
rect 41828 406272 41842 406328
rect 41842 406272 41892 406328
rect 41828 406268 41892 406272
rect 40540 403820 40604 403884
rect 41828 401976 41892 401980
rect 41828 401920 41842 401976
rect 41842 401920 41892 401976
rect 41828 401916 41892 401920
rect 676812 401236 676876 401300
rect 41460 398788 41524 398852
rect 676076 398788 676140 398852
rect 676628 396748 676692 396812
rect 676260 395116 676324 395180
rect 676444 394708 676508 394772
rect 675892 388996 675956 389060
rect 675708 387636 675772 387700
rect 676628 384916 676692 384980
rect 41460 381788 41524 381852
rect 676444 380564 676508 380628
rect 675708 378720 675772 378724
rect 675708 378664 675758 378720
rect 675758 378664 675772 378720
rect 675708 378660 675772 378664
rect 40540 378524 40604 378588
rect 40724 378116 40788 378180
rect 674788 377980 674852 378044
rect 40908 377708 40972 377772
rect 676260 377300 676324 377364
rect 41644 376892 41708 376956
rect 676076 376892 676140 376956
rect 40356 375668 40420 375732
rect 675892 372948 675956 373012
rect 674788 372540 674852 372604
rect 41828 371316 41892 371380
rect 40356 368596 40420 368660
rect 40908 364244 40972 364308
rect 40724 363700 40788 363764
rect 41828 362944 41892 362948
rect 41828 362888 41842 362944
rect 41842 362888 41892 362944
rect 41828 362884 41892 362888
rect 40540 360028 40604 360092
rect 41460 358668 41524 358732
rect 41828 355736 41892 355740
rect 41828 355680 41878 355736
rect 41878 355680 41892 355736
rect 41828 355676 41892 355680
rect 675340 354180 675404 354244
rect 675708 353772 675772 353836
rect 675892 351868 675956 351932
rect 675892 350916 675956 350980
rect 675892 350100 675956 350164
rect 675156 349148 675220 349212
rect 44220 342892 44284 342956
rect 44404 342076 44468 342140
rect 43668 340444 43732 340508
rect 676628 340172 676692 340236
rect 675892 339356 675956 339420
rect 40724 338540 40788 338604
rect 675524 337784 675588 337788
rect 675524 337728 675574 337784
rect 675574 337728 675588 337784
rect 675524 337724 675588 337728
rect 42932 337588 42996 337652
rect 43300 337180 43364 337244
rect 40540 336908 40604 336972
rect 674788 336636 674852 336700
rect 41828 336500 41892 336564
rect 43116 336092 43180 336156
rect 43852 335684 43916 335748
rect 42748 335412 42812 335476
rect 676444 335276 676508 335340
rect 42748 334656 42812 334660
rect 42748 334600 42798 334656
rect 42798 334600 42812 334656
rect 42748 334596 42812 334600
rect 43116 334656 43180 334660
rect 43116 334600 43166 334656
rect 43166 334600 43180 334656
rect 43116 334596 43180 334600
rect 43852 334596 43916 334660
rect 40908 333644 40972 333708
rect 676260 332284 676324 332348
rect 42012 329020 42076 329084
rect 676076 328340 676140 328404
rect 41644 327660 41708 327724
rect 674788 326844 674852 326908
rect 40908 325348 40972 325412
rect 41828 324728 41892 324732
rect 41828 324672 41878 324728
rect 41878 324672 41892 324728
rect 41828 324668 41892 324672
rect 41828 319968 41892 319972
rect 41828 319912 41842 319968
rect 41842 319912 41892 319968
rect 41828 319908 41892 319912
rect 40540 316780 40604 316844
rect 43116 315964 43180 316028
rect 41460 315556 41524 315620
rect 42932 312700 42996 312764
rect 42012 312624 42076 312628
rect 42012 312568 42026 312624
rect 42026 312568 42076 312624
rect 42012 312564 42076 312568
rect 44588 311400 44652 311404
rect 44588 311344 44602 311400
rect 44602 311344 44652 311400
rect 44588 311340 44652 311344
rect 44404 311128 44468 311132
rect 44404 311072 44418 311128
rect 44418 311072 44468 311128
rect 44404 311068 44468 311072
rect 675708 308756 675772 308820
rect 675892 306716 675956 306780
rect 675892 305900 675956 305964
rect 676030 305084 676094 305148
rect 675708 299372 675772 299436
rect 43668 297604 43732 297668
rect 675524 297604 675588 297668
rect 675892 297332 675956 297396
rect 675340 296712 675404 296716
rect 675340 296656 675390 296712
rect 675390 296656 675404 296712
rect 675340 296652 675404 296656
rect 42012 296380 42076 296444
rect 41828 295564 41892 295628
rect 676812 295156 676876 295220
rect 41828 292904 41892 292908
rect 41828 292848 41842 292904
rect 41842 292848 41892 292904
rect 41828 292844 41892 292848
rect 675340 292904 675404 292908
rect 675340 292848 675390 292904
rect 675390 292848 675404 292904
rect 675340 292844 675404 292848
rect 40540 292528 40604 292592
rect 40908 292528 40972 292592
rect 41828 292224 41892 292228
rect 41828 292168 41842 292224
rect 41842 292168 41892 292224
rect 41828 292164 41892 292168
rect 675524 292088 675588 292092
rect 675524 292032 675574 292088
rect 675574 292032 675588 292088
rect 675524 292028 675588 292032
rect 676444 291484 676508 291548
rect 676260 286996 676324 287060
rect 676076 283596 676140 283660
rect 675708 282840 675772 282844
rect 675708 282784 675722 282840
rect 675722 282784 675772 282840
rect 675708 282780 675772 282784
rect 42012 281480 42076 281484
rect 42012 281424 42026 281480
rect 42026 281424 42076 281480
rect 42012 281420 42076 281424
rect 675892 281148 675956 281212
rect 40908 277884 40972 277948
rect 40724 277612 40788 277676
rect 40540 274212 40604 274276
rect 41460 270404 41524 270468
rect 41828 269104 41892 269108
rect 41828 269048 41842 269104
rect 41842 269048 41892 269104
rect 41828 269044 41892 269048
rect 676076 263604 676140 263668
rect 676996 261564 677060 261628
rect 675892 261156 675956 261220
rect 676812 259932 676876 259996
rect 40540 251364 40604 251428
rect 676996 250276 677060 250340
rect 40724 249732 40788 249796
rect 675892 249596 675956 249660
rect 676076 249596 676140 249660
rect 675340 245516 675404 245580
rect 676812 245244 676876 245308
rect 40540 240076 40604 240140
rect 675340 238640 675404 238644
rect 675340 238584 675390 238640
rect 675390 238584 675404 238640
rect 675340 238580 675404 238584
rect 42012 238036 42076 238100
rect 676812 236268 676876 236332
rect 673500 235996 673564 236060
rect 40724 235860 40788 235924
rect 671292 234500 671356 234564
rect 673500 232732 673564 232796
rect 673132 231780 673196 231844
rect 673316 231780 673380 231844
rect 674236 231780 674300 231844
rect 671476 229332 671540 229396
rect 42012 228984 42076 228988
rect 42012 228928 42026 228984
rect 42026 228928 42076 228984
rect 42012 228924 42076 228928
rect 672948 228516 673012 228580
rect 674972 228516 675036 228580
rect 671844 227080 671908 227084
rect 671844 227024 671858 227080
rect 671858 227024 671908 227080
rect 671844 227020 671908 227024
rect 671660 226944 671724 226948
rect 671660 226888 671674 226944
rect 671674 226888 671724 226944
rect 671660 226884 671724 226888
rect 672764 225660 672828 225724
rect 671476 224844 671540 224908
rect 671660 224300 671724 224364
rect 672764 223892 672828 223956
rect 673132 222260 673196 222324
rect 669820 220900 669884 220964
rect 670372 220628 670436 220692
rect 671108 220628 671172 220692
rect 671844 220356 671908 220420
rect 493916 218316 493980 218380
rect 553532 218588 553596 218652
rect 505048 218316 505112 218380
rect 572668 218316 572732 218380
rect 675524 218588 675588 218652
rect 675708 218044 675772 218108
rect 553716 217772 553780 217836
rect 562548 217772 562612 217836
rect 674972 217772 675036 217836
rect 493916 217696 493980 217700
rect 493916 217640 493930 217696
rect 493930 217640 493980 217696
rect 493916 217636 493980 217640
rect 576808 217228 576872 217292
rect 666324 217228 666388 217292
rect 675708 216956 675772 217020
rect 676260 215086 676324 215150
rect 578188 213148 578252 213212
rect 674052 212060 674116 212124
rect 676812 211440 676876 211444
rect 676812 211384 676826 211440
rect 676826 211384 676876 211440
rect 676812 211380 676876 211384
rect 676996 211440 677060 211444
rect 676996 211384 677046 211440
rect 677046 211384 677060 211440
rect 676996 211380 677060 211384
rect 670740 211108 670804 211172
rect 673132 209612 673196 209676
rect 41644 209340 41708 209404
rect 40540 208116 40604 208180
rect 41828 207300 41892 207364
rect 675708 207028 675772 207092
rect 667980 206484 668044 206548
rect 669084 206212 669148 206276
rect 676444 205532 676508 205596
rect 41644 204444 41708 204508
rect 675708 204232 675772 204236
rect 675708 204176 675722 204232
rect 675722 204176 675772 204232
rect 675708 204172 675772 204176
rect 669084 202404 669148 202468
rect 676996 200772 677060 200836
rect 666692 198324 666756 198388
rect 40540 197100 40604 197164
rect 676260 197100 676324 197164
rect 41828 195256 41892 195260
rect 41828 195200 41878 195256
rect 41878 195200 41892 195256
rect 41828 195196 41892 195200
rect 675892 193156 675956 193220
rect 676076 191524 676140 191588
rect 41828 185872 41892 185876
rect 41828 185816 41842 185872
rect 41842 185816 41892 185872
rect 41828 185812 41892 185816
rect 41460 184044 41524 184108
rect 672948 183500 673012 183564
rect 675892 173980 675956 174044
rect 675708 173572 675772 173636
rect 675892 172348 675956 172412
rect 675708 170308 675772 170372
rect 675892 167452 675956 167516
rect 676628 166424 676692 166428
rect 676628 166368 676642 166424
rect 676642 166368 676692 166424
rect 676628 166364 676692 166368
rect 670740 164188 670804 164252
rect 676444 159292 676508 159356
rect 676628 156300 676692 156364
rect 676260 151540 676324 151604
rect 675708 150376 675772 150380
rect 675708 150320 675722 150376
rect 675722 150320 675772 150376
rect 675708 150316 675772 150320
rect 676076 148412 676140 148476
rect 675892 147596 675956 147660
rect 671292 145284 671356 145348
rect 673684 141068 673748 141132
rect 669268 137804 669332 137868
rect 673132 133860 673196 133924
rect 667980 130596 668044 130660
rect 673500 128828 673564 128892
rect 676260 128556 676324 128620
rect 674052 128284 674116 128348
rect 676076 126924 676140 126988
rect 676628 126516 676692 126580
rect 676444 124476 676508 124540
rect 675892 122300 675956 122364
rect 675708 117268 675772 117332
rect 676260 113052 676324 113116
rect 676076 108156 676140 108220
rect 676444 106116 676508 106180
rect 675708 103184 675772 103188
rect 675708 103128 675722 103184
rect 675722 103128 675772 103184
rect 675708 103124 675772 103128
rect 675892 102444 675956 102508
rect 676628 101356 676692 101420
rect 637252 96868 637316 96932
rect 633940 96052 634004 96116
rect 647188 96052 647252 96116
rect 650316 93060 650380 93124
rect 633940 78568 634004 78572
rect 633940 78512 633954 78568
rect 633954 78512 634004 78568
rect 633940 78508 634004 78512
rect 637068 77692 637132 77756
rect 194364 50220 194428 50284
rect 522804 49404 522868 49468
rect 529796 49132 529860 49196
rect 518756 48860 518820 48924
rect 526484 47772 526548 47836
rect 520964 47500 521028 47564
rect 515444 46956 515508 47020
rect 463740 44432 463804 44436
rect 463740 44376 463754 44432
rect 463754 44376 463804 44432
rect 463740 44372 463804 44376
rect 141740 43964 141804 44028
rect 464108 44236 464172 44300
rect 440188 43828 440252 43892
rect 440924 43828 440988 43892
rect 518756 42800 518820 42804
rect 518756 42744 518806 42800
rect 518806 42744 518820 42800
rect 518756 42740 518820 42744
rect 194364 42120 194428 42124
rect 194364 42064 194378 42120
rect 194378 42064 194428 42120
rect 194364 42060 194428 42064
rect 361988 41848 362052 41852
rect 361988 41792 362002 41848
rect 362002 41792 362052 41848
rect 361988 41788 362052 41792
rect 365484 41788 365548 41852
rect 403020 41788 403084 41852
rect 421972 41788 422036 41852
rect 515444 42120 515508 42124
rect 515444 42064 515458 42120
rect 515458 42064 515508 42120
rect 515444 42060 515508 42064
rect 520964 42120 521028 42124
rect 520964 42064 520978 42120
rect 520978 42064 521028 42120
rect 520964 42060 521028 42064
rect 522804 42060 522868 42124
rect 526484 42120 526548 42124
rect 526484 42064 526498 42120
rect 526498 42064 526548 42120
rect 526484 42060 526548 42064
rect 529796 42060 529860 42124
rect 441844 41788 441908 41852
rect 460796 41788 460860 41852
rect 460980 41788 461044 41852
rect 464108 41788 464172 41852
rect 141740 40488 141804 40492
rect 141740 40432 141754 40488
rect 141754 40432 141804 40488
rect 141740 40428 141804 40432
<< metal4 >>
rect 84515 997252 84581 997253
rect 84515 997188 84516 997252
rect 84580 997188 84581 997252
rect 84515 997187 84581 997188
rect 84518 995077 84578 997187
rect 293539 997252 293605 997253
rect 293539 997188 293540 997252
rect 293604 997188 293605 997252
rect 293539 997187 293605 997188
rect 387931 997252 387997 997253
rect 387931 997188 387932 997252
rect 387996 997188 387997 997252
rect 387931 997187 387997 997188
rect 482691 997252 482757 997253
rect 482691 997188 482692 997252
rect 482756 997188 482757 997252
rect 482691 997187 482757 997188
rect 530163 997252 530229 997253
rect 530163 997188 530164 997252
rect 530228 997188 530229 997252
rect 530163 997187 530229 997188
rect 86539 996980 86605 996981
rect 86539 996916 86540 996980
rect 86604 996916 86605 996980
rect 86539 996915 86605 996916
rect 86542 995621 86602 996915
rect 90219 996708 90285 996709
rect 90219 996644 90220 996708
rect 90284 996644 90285 996708
rect 90219 996643 90285 996644
rect 141923 996708 141989 996709
rect 141923 996644 141924 996708
rect 141988 996644 141989 996708
rect 141923 996643 141989 996644
rect 87827 996436 87893 996437
rect 87827 996372 87828 996436
rect 87892 996372 87893 996436
rect 87827 996371 87893 996372
rect 87830 995621 87890 996371
rect 90222 995621 90282 996643
rect 86539 995620 86605 995621
rect 86539 995556 86540 995620
rect 86604 995556 86605 995620
rect 86539 995555 86605 995556
rect 87827 995620 87893 995621
rect 87827 995556 87828 995620
rect 87892 995556 87893 995620
rect 87827 995555 87893 995556
rect 90219 995620 90285 995621
rect 90219 995556 90220 995620
rect 90284 995556 90285 995620
rect 90219 995555 90285 995556
rect 141926 995485 141986 996643
rect 141923 995484 141989 995485
rect 141923 995420 141924 995484
rect 141988 995420 141989 995484
rect 141923 995419 141989 995420
rect 172470 995349 172530 997102
rect 242019 996708 242085 996709
rect 242019 996644 242020 996708
rect 242084 996644 242085 996708
rect 242019 996643 242085 996644
rect 288019 996708 288085 996709
rect 288019 996644 288020 996708
rect 288084 996644 288085 996708
rect 288019 996643 288085 996644
rect 242022 995485 242082 996643
rect 243859 996436 243925 996437
rect 243859 996372 243860 996436
rect 243924 996372 243925 996436
rect 243859 996371 243925 996372
rect 243862 995485 243922 996371
rect 288022 995757 288082 996643
rect 293542 995757 293602 997187
rect 293723 996980 293789 996981
rect 293723 996916 293724 996980
rect 293788 996916 293789 996980
rect 293723 996915 293789 996916
rect 293726 996437 293786 996915
rect 386643 996708 386709 996709
rect 386643 996644 386644 996708
rect 386708 996644 386709 996708
rect 386643 996643 386709 996644
rect 295011 996572 295077 996573
rect 295011 996508 295012 996572
rect 295076 996508 295077 996572
rect 295011 996507 295077 996508
rect 293723 996436 293789 996437
rect 293723 996372 293724 996436
rect 293788 996372 293789 996436
rect 293723 996371 293789 996372
rect 295014 995757 295074 996507
rect 386646 995757 386706 996643
rect 387934 995757 387994 997187
rect 476251 996708 476317 996709
rect 476251 996644 476252 996708
rect 476316 996644 476317 996708
rect 476251 996643 476317 996644
rect 388115 996436 388181 996437
rect 388115 996372 388116 996436
rect 388180 996372 388181 996436
rect 388115 996371 388181 996372
rect 474779 996436 474845 996437
rect 474779 996372 474780 996436
rect 474844 996372 474845 996436
rect 474779 996371 474845 996372
rect 388118 995757 388178 996371
rect 474782 995757 474842 996371
rect 476254 995757 476314 996643
rect 482694 995757 482754 997187
rect 526299 996164 526365 996165
rect 526299 996100 526300 996164
rect 526364 996100 526365 996164
rect 526299 996099 526365 996100
rect 525011 995892 525077 995893
rect 525011 995828 525012 995892
rect 525076 995828 525077 995892
rect 525011 995827 525077 995828
rect 288019 995756 288085 995757
rect 288019 995692 288020 995756
rect 288084 995692 288085 995756
rect 288019 995691 288085 995692
rect 293539 995756 293605 995757
rect 293539 995692 293540 995756
rect 293604 995692 293605 995756
rect 293539 995691 293605 995692
rect 295011 995756 295077 995757
rect 295011 995692 295012 995756
rect 295076 995692 295077 995756
rect 295011 995691 295077 995692
rect 386643 995756 386709 995757
rect 386643 995692 386644 995756
rect 386708 995692 386709 995756
rect 386643 995691 386709 995692
rect 387931 995756 387997 995757
rect 387931 995692 387932 995756
rect 387996 995692 387997 995756
rect 387931 995691 387997 995692
rect 388115 995756 388181 995757
rect 388115 995692 388116 995756
rect 388180 995692 388181 995756
rect 388115 995691 388181 995692
rect 474779 995756 474845 995757
rect 474779 995692 474780 995756
rect 474844 995692 474845 995756
rect 474779 995691 474845 995692
rect 476251 995756 476317 995757
rect 476251 995692 476252 995756
rect 476316 995692 476317 995756
rect 476251 995691 476317 995692
rect 479931 995756 479997 995757
rect 479931 995692 479932 995756
rect 479996 995692 479997 995756
rect 479931 995691 479997 995692
rect 482691 995756 482757 995757
rect 482691 995692 482692 995756
rect 482756 995692 482757 995756
rect 482691 995691 482757 995692
rect 242019 995484 242085 995485
rect 242019 995420 242020 995484
rect 242084 995420 242085 995484
rect 242019 995419 242085 995420
rect 243859 995484 243925 995485
rect 243859 995420 243860 995484
rect 243924 995420 243925 995484
rect 243859 995419 243925 995420
rect 172467 995348 172533 995349
rect 172467 995284 172468 995348
rect 172532 995284 172533 995348
rect 172467 995283 172533 995284
rect 84515 995076 84581 995077
rect 84515 995012 84516 995076
rect 84580 995012 84581 995076
rect 84515 995011 84581 995012
rect 142291 994532 142357 994533
rect 142291 994530 142292 994532
rect 142110 994470 142292 994530
rect 142110 993989 142170 994470
rect 142291 994468 142292 994470
rect 142356 994468 142357 994532
rect 142291 994467 142357 994468
rect 479934 993989 479994 995691
rect 525014 995349 525074 995827
rect 525011 995348 525077 995349
rect 525011 995284 525012 995348
rect 525076 995284 525077 995348
rect 525011 995283 525077 995284
rect 526302 994805 526362 996099
rect 530166 995485 530226 997187
rect 627131 996980 627197 996981
rect 627131 996916 627132 996980
rect 627196 996916 627197 996980
rect 627131 996915 627197 996916
rect 626579 996708 626645 996709
rect 626579 996644 626580 996708
rect 626644 996644 626645 996708
rect 626579 996643 626645 996644
rect 626582 995757 626642 996643
rect 627134 995757 627194 996915
rect 627867 996436 627933 996437
rect 627867 996372 627868 996436
rect 627932 996372 627933 996436
rect 627867 996371 627933 996372
rect 627870 995757 627930 996371
rect 626579 995756 626645 995757
rect 626579 995692 626580 995756
rect 626644 995692 626645 995756
rect 626579 995691 626645 995692
rect 627131 995756 627197 995757
rect 627131 995692 627132 995756
rect 627196 995692 627197 995756
rect 627131 995691 627197 995692
rect 627867 995756 627933 995757
rect 627867 995692 627868 995756
rect 627932 995692 627933 995756
rect 627867 995691 627933 995692
rect 530163 995484 530229 995485
rect 530163 995420 530164 995484
rect 530228 995420 530229 995484
rect 530163 995419 530229 995420
rect 526299 994804 526365 994805
rect 526299 994740 526300 994804
rect 526364 994740 526365 994804
rect 526299 994739 526365 994740
rect 536787 994804 536853 994805
rect 536787 994740 536788 994804
rect 536852 994740 536853 994804
rect 536787 994739 536853 994740
rect 142107 993988 142173 993989
rect 142107 993924 142108 993988
rect 142172 993924 142173 993988
rect 142107 993923 142173 993924
rect 479931 993988 479997 993989
rect 479931 993924 479932 993988
rect 479996 993924 479997 993988
rect 479931 993923 479997 993924
rect 536790 993258 536850 994739
rect 572670 990997 572730 993022
rect 572667 990996 572733 990997
rect 572667 990932 572668 990996
rect 572732 990932 572733 990996
rect 572667 990931 572733 990932
rect 42011 967196 42077 967197
rect 42011 967132 42012 967196
rect 42076 967132 42077 967196
rect 42011 967131 42077 967132
rect 41459 962164 41525 962165
rect 41459 962100 41460 962164
rect 41524 962100 41525 962164
rect 41459 962099 41525 962100
rect 41275 959852 41341 959853
rect 41275 959788 41276 959852
rect 41340 959788 41341 959852
rect 41275 959787 41341 959788
rect 40539 959172 40605 959173
rect 40539 959108 40540 959172
rect 40604 959108 40605 959172
rect 40539 959107 40605 959108
rect 40542 939810 40602 959107
rect 40723 955500 40789 955501
rect 40723 955436 40724 955500
rect 40788 955436 40789 955500
rect 40723 955435 40789 955436
rect 40358 939750 40602 939810
rect 40171 937242 40237 937243
rect 40171 937178 40172 937242
rect 40236 937178 40237 937242
rect 40171 937177 40237 937178
rect 40174 930150 40234 937177
rect 40358 936050 40418 939750
rect 40726 937050 40786 955435
rect 41278 951829 41338 959787
rect 41462 952237 41522 962099
rect 41459 952236 41525 952237
rect 41459 952172 41460 952236
rect 41524 952172 41525 952236
rect 41459 952171 41525 952172
rect 41275 951828 41341 951829
rect 41275 951764 41276 951828
rect 41340 951764 41341 951828
rect 41275 951763 41341 951764
rect 42014 951693 42074 967131
rect 675339 966516 675405 966517
rect 675339 966452 675340 966516
rect 675404 966452 675405 966516
rect 675339 966451 675405 966452
rect 42563 957948 42629 957949
rect 42563 957884 42564 957948
rect 42628 957884 42629 957948
rect 42563 957883 42629 957884
rect 42566 951965 42626 957883
rect 42563 951964 42629 951965
rect 42563 951900 42564 951964
rect 42628 951900 42629 951964
rect 42563 951899 42629 951900
rect 42011 951692 42077 951693
rect 42011 951628 42012 951692
rect 42076 951628 42077 951692
rect 42011 951627 42077 951628
rect 675342 951557 675402 966451
rect 676811 964748 676877 964749
rect 676811 964684 676812 964748
rect 676876 964684 676877 964748
rect 676811 964683 676877 964684
rect 676075 963388 676141 963389
rect 676075 963324 676076 963388
rect 676140 963324 676141 963388
rect 676075 963323 676141 963324
rect 675339 951556 675405 951557
rect 675339 951492 675340 951556
rect 675404 951492 675405 951556
rect 675339 951491 675405 951492
rect 676078 949517 676138 963323
rect 676627 956452 676693 956453
rect 676627 956388 676628 956452
rect 676692 956388 676693 956452
rect 676627 956387 676693 956388
rect 676075 949516 676141 949517
rect 676075 949452 676076 949516
rect 676140 949452 676141 949516
rect 676075 949451 676141 949452
rect 41827 941084 41893 941085
rect 41827 941020 41828 941084
rect 41892 941020 41893 941084
rect 41827 941019 41893 941020
rect 41830 937277 41890 941019
rect 675155 938228 675221 938229
rect 675155 938164 675156 938228
rect 675220 938164 675221 938228
rect 675155 938163 675221 938164
rect 674603 937412 674669 937413
rect 674603 937348 674604 937412
rect 674668 937410 674669 937412
rect 675158 937410 675218 938163
rect 674668 937350 675218 937410
rect 674668 937348 674669 937350
rect 674603 937347 674669 937348
rect 41827 937276 41893 937277
rect 41827 937212 41828 937276
rect 41892 937212 41893 937276
rect 41827 937211 41893 937212
rect 40726 936990 41890 937050
rect 41830 936597 41890 936990
rect 41827 936596 41893 936597
rect 41827 936532 41828 936596
rect 41892 936532 41893 936596
rect 41827 936531 41893 936532
rect 40358 935990 41890 936050
rect 41830 935781 41890 935990
rect 41827 935780 41893 935781
rect 41827 935716 41828 935780
rect 41892 935716 41893 935780
rect 41827 935715 41893 935716
rect 676630 931973 676690 956387
rect 676814 950741 676874 964683
rect 676995 957812 677061 957813
rect 676995 957748 676996 957812
rect 677060 957748 677061 957812
rect 676995 957747 677061 957748
rect 676811 950740 676877 950741
rect 676811 950676 676812 950740
rect 676876 950676 676877 950740
rect 676811 950675 676877 950676
rect 676627 931972 676693 931973
rect 676627 931908 676628 931972
rect 676692 931908 676693 931972
rect 676627 931907 676693 931908
rect 676998 931565 677058 957747
rect 676995 931564 677061 931565
rect 676995 931500 676996 931564
rect 677060 931500 677061 931564
rect 676995 931499 677061 931500
rect 39990 930090 40234 930150
rect 39990 828030 40050 930090
rect 42011 911980 42077 911981
rect 42011 911916 42012 911980
rect 42076 911916 42077 911980
rect 42011 911915 42077 911916
rect 42014 885461 42074 911915
rect 42195 911708 42261 911709
rect 42195 911644 42196 911708
rect 42260 911644 42261 911708
rect 42195 911643 42261 911644
rect 42011 885460 42077 885461
rect 42011 885396 42012 885460
rect 42076 885396 42077 885460
rect 42011 885395 42077 885396
rect 42198 885189 42258 911643
rect 42195 885188 42261 885189
rect 42195 885124 42196 885188
rect 42260 885124 42261 885188
rect 42195 885123 42261 885124
rect 676811 876620 676877 876621
rect 676811 876556 676812 876620
rect 676876 876556 676877 876620
rect 676811 876555 676877 876556
rect 676075 875940 676141 875941
rect 676075 875876 676076 875940
rect 676140 875876 676141 875940
rect 676075 875875 676141 875876
rect 675155 874036 675221 874037
rect 675155 873972 675156 874036
rect 675220 873972 675221 874036
rect 675155 873971 675221 873972
rect 673867 873220 673933 873221
rect 673867 873156 673868 873220
rect 673932 873156 673933 873220
rect 673867 873155 673933 873156
rect 39990 827970 40234 828030
rect 40174 815659 40234 827970
rect 40171 815658 40237 815659
rect 40171 815594 40172 815658
rect 40236 815594 40237 815658
rect 40171 815593 40237 815594
rect 42011 812020 42077 812021
rect 42011 811956 42012 812020
rect 42076 811956 42077 812020
rect 42011 811955 42077 811956
rect 41827 809164 41893 809165
rect 41827 809100 41828 809164
rect 41892 809100 41893 809164
rect 41827 809099 41893 809100
rect 41830 808890 41890 809099
rect 40910 808830 41890 808890
rect 40539 808712 40605 808713
rect 40539 808648 40540 808712
rect 40604 808648 40605 808712
rect 40539 808647 40605 808648
rect 40542 792573 40602 808647
rect 40723 805084 40789 805085
rect 40723 805020 40724 805084
rect 40788 805020 40789 805084
rect 40723 805019 40789 805020
rect 40726 793797 40786 805019
rect 40910 794477 40970 808830
rect 42014 808210 42074 811955
rect 41646 808150 42074 808210
rect 41459 805628 41525 805629
rect 41459 805564 41460 805628
rect 41524 805564 41525 805628
rect 41459 805563 41525 805564
rect 40907 794476 40973 794477
rect 40907 794412 40908 794476
rect 40972 794412 40973 794476
rect 40907 794411 40973 794412
rect 40723 793796 40789 793797
rect 40723 793732 40724 793796
rect 40788 793732 40789 793796
rect 40723 793731 40789 793732
rect 40539 792572 40605 792573
rect 40539 792508 40540 792572
rect 40604 792508 40605 792572
rect 40539 792507 40605 792508
rect 41462 788221 41522 805563
rect 41646 789173 41706 808150
rect 41827 807260 41893 807261
rect 41827 807196 41828 807260
rect 41892 807196 41893 807260
rect 41827 807195 41893 807196
rect 41643 789172 41709 789173
rect 41643 789108 41644 789172
rect 41708 789108 41709 789172
rect 41643 789107 41709 789108
rect 41830 788765 41890 807195
rect 41827 788764 41893 788765
rect 41827 788700 41828 788764
rect 41892 788700 41893 788764
rect 41827 788699 41893 788700
rect 41459 788220 41525 788221
rect 41459 788156 41460 788220
rect 41524 788156 41525 788220
rect 41459 788155 41525 788156
rect 673870 772309 673930 873155
rect 675158 866829 675218 873971
rect 675155 866828 675221 866829
rect 675155 866764 675156 866828
rect 675220 866764 675221 866828
rect 675155 866763 675221 866764
rect 674419 783052 674485 783053
rect 674419 782988 674420 783052
rect 674484 782988 674485 783052
rect 674419 782987 674485 782988
rect 673867 772308 673933 772309
rect 673867 772244 673868 772308
rect 673932 772244 673933 772308
rect 673867 772243 673933 772244
rect 41459 769860 41525 769861
rect 41459 769796 41460 769860
rect 41524 769796 41525 769860
rect 41459 769795 41525 769796
rect 40907 765780 40973 765781
rect 40907 765716 40908 765780
rect 40972 765716 40973 765780
rect 40907 765715 40973 765716
rect 40539 765372 40605 765373
rect 40539 765308 40540 765372
rect 40604 765308 40605 765372
rect 40539 765307 40605 765308
rect 40355 757484 40421 757485
rect 40355 757420 40356 757484
rect 40420 757420 40421 757484
rect 40355 757419 40421 757420
rect 40358 755445 40418 757419
rect 40355 755444 40421 755445
rect 40355 755380 40356 755444
rect 40420 755380 40421 755444
rect 40355 755379 40421 755380
rect 40542 749461 40602 765307
rect 40723 764964 40789 764965
rect 40723 764900 40724 764964
rect 40788 764900 40789 764964
rect 40723 764899 40789 764900
rect 40726 750413 40786 764899
rect 40910 751093 40970 765715
rect 41091 758028 41157 758029
rect 41091 757964 41092 758028
rect 41156 757964 41157 758028
rect 41091 757963 41157 757964
rect 41094 753677 41154 757963
rect 41091 753676 41157 753677
rect 41091 753612 41092 753676
rect 41156 753612 41157 753676
rect 41091 753611 41157 753612
rect 40907 751092 40973 751093
rect 40907 751028 40908 751092
rect 40972 751028 40973 751092
rect 40907 751027 40973 751028
rect 40723 750412 40789 750413
rect 40723 750348 40724 750412
rect 40788 750348 40789 750412
rect 40723 750347 40789 750348
rect 40539 749460 40605 749461
rect 40539 749396 40540 749460
rect 40604 749396 40605 749460
rect 40539 749395 40605 749396
rect 41462 746605 41522 769795
rect 41643 759116 41709 759117
rect 41643 759052 41644 759116
rect 41708 759052 41709 759116
rect 41643 759051 41709 759052
rect 41459 746604 41525 746605
rect 41459 746540 41460 746604
rect 41524 746540 41525 746604
rect 41459 746539 41525 746540
rect 41646 746333 41706 759051
rect 42379 757892 42445 757893
rect 42379 757828 42380 757892
rect 42444 757828 42445 757892
rect 42379 757827 42445 757828
rect 42011 757756 42077 757757
rect 42011 757692 42012 757756
rect 42076 757692 42077 757756
rect 42011 757691 42077 757692
rect 42014 746610 42074 757691
rect 42195 754900 42261 754901
rect 42195 754836 42196 754900
rect 42260 754836 42261 754900
rect 42195 754835 42261 754836
rect 42198 752997 42258 754835
rect 42382 753405 42442 757827
rect 42379 753404 42445 753405
rect 42379 753340 42380 753404
rect 42444 753340 42445 753404
rect 42379 753339 42445 753340
rect 42195 752996 42261 752997
rect 42195 752932 42196 752996
rect 42260 752932 42261 752996
rect 42195 752931 42261 752932
rect 42195 752044 42261 752045
rect 42195 751980 42196 752044
rect 42260 751980 42261 752044
rect 42195 751979 42261 751980
rect 41830 746550 42074 746610
rect 41643 746332 41709 746333
rect 41643 746268 41644 746332
rect 41708 746268 41709 746332
rect 41643 746267 41709 746268
rect 41830 745109 41890 746550
rect 42198 746061 42258 751979
rect 42195 746060 42261 746061
rect 42195 745996 42196 746060
rect 42260 745996 42261 746060
rect 42195 745995 42261 745996
rect 41827 745108 41893 745109
rect 41827 745044 41828 745108
rect 41892 745044 41893 745108
rect 41827 745043 41893 745044
rect 674235 739396 674301 739397
rect 674235 739332 674236 739396
rect 674300 739332 674301 739396
rect 674235 739331 674301 739332
rect 41827 726884 41893 726885
rect 41827 726820 41828 726884
rect 41892 726820 41893 726884
rect 41827 726819 41893 726820
rect 41830 726610 41890 726819
rect 41462 726550 41890 726610
rect 40723 721772 40789 721773
rect 40723 721708 40724 721772
rect 40788 721708 40789 721772
rect 40723 721707 40789 721708
rect 40539 718044 40605 718045
rect 40539 717980 40540 718044
rect 40604 717980 40605 718044
rect 40539 717979 40605 717980
rect 40542 704309 40602 717979
rect 40726 709477 40786 721707
rect 40907 714236 40973 714237
rect 40907 714172 40908 714236
rect 40972 714172 40973 714236
rect 40907 714171 40973 714172
rect 40910 709885 40970 714171
rect 40907 709884 40973 709885
rect 40907 709820 40908 709884
rect 40972 709820 40973 709884
rect 40907 709819 40973 709820
rect 40723 709476 40789 709477
rect 40723 709412 40724 709476
rect 40788 709412 40789 709476
rect 40723 709411 40789 709412
rect 40539 704308 40605 704309
rect 40539 704244 40540 704308
rect 40604 704244 40605 704308
rect 40539 704243 40605 704244
rect 41462 702541 41522 726550
rect 41827 722396 41893 722397
rect 41827 722332 41828 722396
rect 41892 722332 41893 722396
rect 41827 722331 41893 722332
rect 41643 721772 41709 721773
rect 41643 721708 41644 721772
rect 41708 721708 41709 721772
rect 41643 721707 41709 721708
rect 41459 702540 41525 702541
rect 41459 702476 41460 702540
rect 41524 702476 41525 702540
rect 41459 702475 41525 702476
rect 41646 701589 41706 721707
rect 41830 718045 41890 722331
rect 41827 718044 41893 718045
rect 41827 717980 41828 718044
rect 41892 717980 41893 718044
rect 41827 717979 41893 717980
rect 41827 715460 41893 715461
rect 41827 715396 41828 715460
rect 41892 715396 41893 715460
rect 41827 715395 41893 715396
rect 41830 702405 41890 715395
rect 42011 714236 42077 714237
rect 42011 714172 42012 714236
rect 42076 714172 42077 714236
rect 42011 714171 42077 714172
rect 42014 706757 42074 714171
rect 42011 706756 42077 706757
rect 42011 706692 42012 706756
rect 42076 706692 42077 706756
rect 42011 706691 42077 706692
rect 41827 702404 41893 702405
rect 41827 702340 41828 702404
rect 41892 702340 41893 702404
rect 41827 702339 41893 702340
rect 41643 701588 41709 701589
rect 41643 701524 41644 701588
rect 41708 701524 41709 701588
rect 41643 701523 41709 701524
rect 41827 683636 41893 683637
rect 41827 683572 41828 683636
rect 41892 683572 41893 683636
rect 41827 683571 41893 683572
rect 40542 679630 40970 679690
rect 40355 670988 40421 670989
rect 40355 670924 40356 670988
rect 40420 670924 40421 670988
rect 40355 670923 40421 670924
rect 40358 668133 40418 670923
rect 40355 668132 40421 668133
rect 40355 668068 40356 668132
rect 40420 668068 40421 668132
rect 40355 668067 40421 668068
rect 40542 665413 40602 679630
rect 40910 678993 40970 679630
rect 41830 679010 41890 683571
rect 674238 681053 674298 739331
rect 674422 707573 674482 782987
rect 675339 780468 675405 780469
rect 675339 780404 675340 780468
rect 675404 780404 675405 780468
rect 675339 780403 675405 780404
rect 674971 777204 675037 777205
rect 674971 777140 674972 777204
rect 675036 777140 675037 777204
rect 674971 777139 675037 777140
rect 674974 773397 675034 777139
rect 675342 776117 675402 780403
rect 675523 778428 675589 778429
rect 675523 778364 675524 778428
rect 675588 778364 675589 778428
rect 675523 778363 675589 778364
rect 675526 776253 675586 778363
rect 675523 776252 675589 776253
rect 675523 776188 675524 776252
rect 675588 776188 675589 776252
rect 675523 776187 675589 776188
rect 675339 776116 675405 776117
rect 675339 776052 675340 776116
rect 675404 776052 675405 776116
rect 675339 776051 675405 776052
rect 674971 773396 675037 773397
rect 674971 773332 674972 773396
rect 675036 773332 675037 773396
rect 674971 773331 675037 773332
rect 676078 768773 676138 875875
rect 676075 768772 676141 768773
rect 676075 768708 676076 768772
rect 676140 768708 676141 768772
rect 676075 768707 676141 768708
rect 675891 766596 675957 766597
rect 675891 766532 675892 766596
rect 675956 766532 675957 766596
rect 675891 766531 675957 766532
rect 674603 741572 674669 741573
rect 674603 741508 674604 741572
rect 674668 741508 674669 741572
rect 674603 741507 674669 741508
rect 674419 707572 674485 707573
rect 674419 707508 674420 707572
rect 674484 707508 674485 707572
rect 674419 707507 674485 707508
rect 674419 693020 674485 693021
rect 674419 692956 674420 693020
rect 674484 692956 674485 693020
rect 674419 692955 674485 692956
rect 674235 681052 674301 681053
rect 674235 680988 674236 681052
rect 674300 680988 674301 681052
rect 674235 680987 674301 680988
rect 40723 678992 40789 678993
rect 40723 678928 40724 678992
rect 40788 678928 40789 678992
rect 40723 678927 40789 678928
rect 40907 678992 40973 678993
rect 40907 678928 40908 678992
rect 40972 678928 40973 678992
rect 40907 678927 40973 678928
rect 41462 678950 41890 679010
rect 40726 667045 40786 678927
rect 41275 672484 41341 672485
rect 41275 672420 41276 672484
rect 41340 672420 41341 672484
rect 41275 672419 41341 672420
rect 41278 669085 41338 672419
rect 41275 669084 41341 669085
rect 41275 669020 41276 669084
rect 41340 669020 41341 669084
rect 41275 669019 41341 669020
rect 40723 667044 40789 667045
rect 40723 666980 40724 667044
rect 40788 666980 40789 667044
rect 40723 666979 40789 666980
rect 40539 665412 40605 665413
rect 40539 665348 40540 665412
rect 40604 665348 40605 665412
rect 40539 665347 40605 665348
rect 41462 659837 41522 678950
rect 41827 678604 41893 678605
rect 41827 678540 41828 678604
rect 41892 678540 41893 678604
rect 41827 678539 41893 678540
rect 41830 676230 41890 678539
rect 41646 676170 41890 676230
rect 41459 659836 41525 659837
rect 41459 659772 41460 659836
rect 41524 659772 41525 659836
rect 41459 659771 41525 659772
rect 41646 658341 41706 676170
rect 41827 672756 41893 672757
rect 41827 672692 41828 672756
rect 41892 672692 41893 672756
rect 41827 672691 41893 672692
rect 41830 658613 41890 672691
rect 42195 672212 42261 672213
rect 42195 672148 42196 672212
rect 42260 672148 42261 672212
rect 42195 672147 42261 672148
rect 42011 669356 42077 669357
rect 42011 669292 42012 669356
rect 42076 669292 42077 669356
rect 42011 669291 42077 669292
rect 42014 667725 42074 669291
rect 42198 668949 42258 672147
rect 42195 668948 42261 668949
rect 42195 668884 42196 668948
rect 42260 668884 42261 668948
rect 42195 668883 42261 668884
rect 42011 667724 42077 667725
rect 42011 667660 42012 667724
rect 42076 667660 42077 667724
rect 42011 667659 42077 667660
rect 42011 665684 42077 665685
rect 42011 665620 42012 665684
rect 42076 665620 42077 665684
rect 42011 665619 42077 665620
rect 42014 664053 42074 665619
rect 42011 664052 42077 664053
rect 42011 663988 42012 664052
rect 42076 663988 42077 664052
rect 42011 663987 42077 663988
rect 42195 662964 42261 662965
rect 42195 662900 42196 662964
rect 42260 662900 42261 662964
rect 42195 662899 42261 662900
rect 42198 659021 42258 662899
rect 42195 659020 42261 659021
rect 42195 658956 42196 659020
rect 42260 658956 42261 659020
rect 42195 658955 42261 658956
rect 41827 658612 41893 658613
rect 41827 658548 41828 658612
rect 41892 658548 41893 658612
rect 41827 658547 41893 658548
rect 41643 658340 41709 658341
rect 41643 658276 41644 658340
rect 41708 658276 41709 658340
rect 41643 658275 41709 658276
rect 674235 642156 674301 642157
rect 674235 642092 674236 642156
rect 674300 642092 674301 642156
rect 674235 642091 674301 642092
rect 41459 640660 41525 640661
rect 41459 640596 41460 640660
rect 41524 640596 41525 640660
rect 41459 640595 41525 640596
rect 40723 634948 40789 634949
rect 40723 634884 40724 634948
rect 40788 634884 40789 634948
rect 40723 634883 40789 634884
rect 40539 634540 40605 634541
rect 40539 634476 40540 634540
rect 40604 634476 40605 634540
rect 40539 634475 40605 634476
rect 40542 620397 40602 634475
rect 40726 623797 40786 634883
rect 40723 623796 40789 623797
rect 40723 623732 40724 623796
rect 40788 623732 40789 623796
rect 40723 623731 40789 623732
rect 40539 620396 40605 620397
rect 40539 620332 40540 620396
rect 40604 620332 40605 620396
rect 40539 620331 40605 620332
rect 41462 614141 41522 640595
rect 674051 640524 674117 640525
rect 674051 640460 674052 640524
rect 674116 640460 674117 640524
rect 674051 640459 674117 640460
rect 41643 639028 41709 639029
rect 41643 638964 41644 639028
rect 41708 638964 41709 639028
rect 41643 638963 41709 638964
rect 41646 618357 41706 638963
rect 674054 636309 674114 640459
rect 674238 636853 674298 642091
rect 674235 636852 674301 636853
rect 674235 636788 674236 636852
rect 674300 636788 674301 636852
rect 674235 636787 674301 636788
rect 674051 636308 674117 636309
rect 674051 636244 674052 636308
rect 674116 636244 674117 636308
rect 674051 636243 674117 636244
rect 41827 630732 41893 630733
rect 41827 630668 41828 630732
rect 41892 630668 41893 630732
rect 41827 630667 41893 630668
rect 41643 618356 41709 618357
rect 41643 618292 41644 618356
rect 41708 618292 41709 618356
rect 41643 618291 41709 618292
rect 41830 615501 41890 630667
rect 42195 626652 42261 626653
rect 42195 626588 42196 626652
rect 42260 626588 42261 626652
rect 42195 626587 42261 626588
rect 42011 625292 42077 625293
rect 42011 625228 42012 625292
rect 42076 625228 42077 625292
rect 42011 625227 42077 625228
rect 42014 623389 42074 625227
rect 42198 624477 42258 626587
rect 42195 624476 42261 624477
rect 42195 624412 42196 624476
rect 42260 624412 42261 624476
rect 42195 624411 42261 624412
rect 42011 623388 42077 623389
rect 42011 623324 42012 623388
rect 42076 623324 42077 623388
rect 42011 623323 42077 623324
rect 42195 617676 42261 617677
rect 42195 617612 42196 617676
rect 42260 617612 42261 617676
rect 42195 617611 42261 617612
rect 42198 615909 42258 617611
rect 674422 617405 674482 692955
rect 674606 682413 674666 741507
rect 675894 728789 675954 766531
rect 676075 765100 676141 765101
rect 676075 765036 676076 765100
rect 676140 765036 676141 765100
rect 676075 765035 676141 765036
rect 675891 728788 675957 728789
rect 675891 728724 675892 728788
rect 675956 728724 675957 728788
rect 675891 728723 675957 728724
rect 676078 725797 676138 765035
rect 676814 761837 676874 876555
rect 676811 761836 676877 761837
rect 676811 761772 676812 761836
rect 676876 761772 676877 761836
rect 676811 761771 676877 761772
rect 676811 728788 676877 728789
rect 676811 728724 676812 728788
rect 676876 728724 676877 728788
rect 676811 728723 676877 728724
rect 676075 725796 676141 725797
rect 676075 725732 676076 725796
rect 676140 725732 676141 725796
rect 676075 725731 676141 725732
rect 676814 712330 676874 728723
rect 675894 712270 676874 712330
rect 675894 712061 675954 712270
rect 675891 712060 675957 712061
rect 675891 711996 675892 712060
rect 675956 711996 675957 712060
rect 675891 711995 675957 711996
rect 675339 696828 675405 696829
rect 675339 696764 675340 696828
rect 675404 696764 675405 696828
rect 675339 696763 675405 696764
rect 675342 685949 675402 696763
rect 676811 694108 676877 694109
rect 676811 694044 676812 694108
rect 676876 694044 676877 694108
rect 676811 694043 676877 694044
rect 675339 685948 675405 685949
rect 675339 685884 675340 685948
rect 675404 685884 675405 685948
rect 675339 685883 675405 685884
rect 674603 682412 674669 682413
rect 674603 682348 674604 682412
rect 674668 682348 674669 682412
rect 674603 682347 674669 682348
rect 675339 652900 675405 652901
rect 675339 652836 675340 652900
rect 675404 652836 675405 652900
rect 675339 652835 675405 652836
rect 674971 645828 675037 645829
rect 674971 645764 674972 645828
rect 675036 645764 675037 645828
rect 674971 645763 675037 645764
rect 674603 640796 674669 640797
rect 674603 640732 674604 640796
rect 674668 640732 674669 640796
rect 674603 640731 674669 640732
rect 674419 617404 674485 617405
rect 674419 617340 674420 617404
rect 674484 617340 674485 617404
rect 674419 617339 674485 617340
rect 673867 616180 673933 616181
rect 673867 616116 673868 616180
rect 673932 616116 673933 616180
rect 673867 616115 673933 616116
rect 42195 615908 42261 615909
rect 42195 615844 42196 615908
rect 42260 615844 42261 615908
rect 42195 615843 42261 615844
rect 41827 615500 41893 615501
rect 41827 615436 41828 615500
rect 41892 615436 41893 615500
rect 41827 615435 41893 615436
rect 41459 614140 41525 614141
rect 41459 614076 41460 614140
rect 41524 614076 41525 614140
rect 41459 614075 41525 614076
rect 41827 597276 41893 597277
rect 41827 597212 41828 597276
rect 41892 597212 41893 597276
rect 41827 597211 41893 597212
rect 41830 596730 41890 597211
rect 41462 596670 41890 596730
rect 40723 589660 40789 589661
rect 40723 589596 40724 589660
rect 40788 589596 40789 589660
rect 40723 589595 40789 589596
rect 40539 589388 40605 589389
rect 40539 589324 40540 589388
rect 40604 589324 40605 589388
rect 40539 589323 40605 589324
rect 40542 576877 40602 589323
rect 40726 578237 40786 589595
rect 40907 589524 40973 589525
rect 40907 589460 40908 589524
rect 40972 589460 40973 589524
rect 40907 589459 40973 589460
rect 40723 578236 40789 578237
rect 40723 578172 40724 578236
rect 40788 578172 40789 578236
rect 40723 578171 40789 578172
rect 40910 577557 40970 589459
rect 40907 577556 40973 577557
rect 40907 577492 40908 577556
rect 40972 577492 40973 577556
rect 40907 577491 40973 577492
rect 40539 576876 40605 576877
rect 40539 576812 40540 576876
rect 40604 576812 40605 576876
rect 40539 576811 40605 576812
rect 41462 573341 41522 596670
rect 41827 596460 41893 596461
rect 41827 596396 41828 596460
rect 41892 596396 41893 596460
rect 41827 596395 41893 596396
rect 41830 589290 41890 596395
rect 41646 589230 41890 589290
rect 41459 573340 41525 573341
rect 41459 573276 41460 573340
rect 41524 573276 41525 573340
rect 41459 573275 41525 573276
rect 41646 572117 41706 589230
rect 42011 586804 42077 586805
rect 42011 586740 42012 586804
rect 42076 586740 42077 586804
rect 42011 586739 42077 586740
rect 41827 584628 41893 584629
rect 41827 584564 41828 584628
rect 41892 584564 41893 584628
rect 41827 584563 41893 584564
rect 41643 572116 41709 572117
rect 41643 572052 41644 572116
rect 41708 572052 41709 572116
rect 41643 572051 41709 572052
rect 41830 570213 41890 584563
rect 42014 581501 42074 586739
rect 42195 584356 42261 584357
rect 42195 584292 42196 584356
rect 42260 584292 42261 584356
rect 42195 584291 42261 584292
rect 42011 581500 42077 581501
rect 42011 581436 42012 581500
rect 42076 581436 42077 581500
rect 42011 581435 42077 581436
rect 42198 580277 42258 584291
rect 42195 580276 42261 580277
rect 42195 580212 42196 580276
rect 42260 580212 42261 580276
rect 42195 580211 42261 580212
rect 42563 577964 42629 577965
rect 42563 577900 42564 577964
rect 42628 577900 42629 577964
rect 42563 577899 42629 577900
rect 42566 574157 42626 577899
rect 42563 574156 42629 574157
rect 42563 574092 42564 574156
rect 42628 574092 42629 574156
rect 42563 574091 42629 574092
rect 41827 570212 41893 570213
rect 41827 570148 41828 570212
rect 41892 570148 41893 570212
rect 41827 570147 41893 570148
rect 42195 554028 42261 554029
rect 42195 553964 42196 554028
rect 42260 553964 42261 554028
rect 42195 553963 42261 553964
rect 42011 553212 42077 553213
rect 42011 553148 42012 553212
rect 42076 553148 42077 553212
rect 42011 553147 42077 553148
rect 42014 549130 42074 553147
rect 41462 549070 42074 549130
rect 40723 545732 40789 545733
rect 40723 545668 40724 545732
rect 40788 545668 40789 545732
rect 40723 545667 40789 545668
rect 40539 545460 40605 545461
rect 40539 545396 40540 545460
rect 40604 545396 40605 545460
rect 40539 545395 40605 545396
rect 40542 535261 40602 545395
rect 40726 538253 40786 545667
rect 40723 538252 40789 538253
rect 40723 538188 40724 538252
rect 40788 538188 40789 538252
rect 40723 538187 40789 538188
rect 40539 535260 40605 535261
rect 40539 535196 40540 535260
rect 40604 535196 40605 535260
rect 40539 535195 40605 535196
rect 41462 529685 41522 549070
rect 42198 548450 42258 553963
rect 42379 551852 42445 551853
rect 42379 551788 42380 551852
rect 42444 551788 42445 551852
rect 42379 551787 42445 551788
rect 41646 548390 42258 548450
rect 41646 530229 41706 548390
rect 42382 547890 42442 551787
rect 41830 547830 42442 547890
rect 41643 530228 41709 530229
rect 41643 530164 41644 530228
rect 41708 530164 41709 530228
rect 41643 530163 41709 530164
rect 41459 529684 41525 529685
rect 41459 529620 41460 529684
rect 41524 529620 41525 529684
rect 41459 529619 41525 529620
rect 41830 529413 41890 547830
rect 41827 529412 41893 529413
rect 41827 529348 41828 529412
rect 41892 529348 41893 529412
rect 41827 529347 41893 529348
rect 673870 455293 673930 616115
rect 674235 602988 674301 602989
rect 674235 602924 674236 602988
rect 674300 602924 674301 602988
rect 674235 602923 674301 602924
rect 674238 547365 674298 602923
rect 674235 547364 674301 547365
rect 674235 547300 674236 547364
rect 674300 547300 674301 547364
rect 674235 547299 674301 547300
rect 674606 475421 674666 640731
rect 674974 637669 675034 645763
rect 675155 639844 675221 639845
rect 675155 639780 675156 639844
rect 675220 639780 675221 639844
rect 675155 639779 675221 639780
rect 675158 637941 675218 639779
rect 675342 637941 675402 652835
rect 675523 651540 675589 651541
rect 675523 651476 675524 651540
rect 675588 651476 675589 651540
rect 675523 651475 675589 651476
rect 675155 637940 675221 637941
rect 675155 637876 675156 637940
rect 675220 637876 675221 637940
rect 675155 637875 675221 637876
rect 675339 637940 675405 637941
rect 675339 637876 675340 637940
rect 675404 637876 675405 637940
rect 675339 637875 675405 637876
rect 675526 637669 675586 651475
rect 674971 637668 675037 637669
rect 674971 637604 674972 637668
rect 675036 637604 675037 637668
rect 674971 637603 675037 637604
rect 675523 637668 675589 637669
rect 675523 637604 675524 637668
rect 675588 637604 675589 637668
rect 675523 637603 675589 637604
rect 674971 631412 675037 631413
rect 674971 631348 674972 631412
rect 675036 631348 675037 631412
rect 674971 631347 675037 631348
rect 676075 631412 676141 631413
rect 676075 631348 676076 631412
rect 676140 631348 676141 631412
rect 676075 631347 676141 631348
rect 674974 630690 675034 631347
rect 674974 630630 675218 630690
rect 675158 592925 675218 630630
rect 675523 607884 675589 607885
rect 675523 607820 675524 607884
rect 675588 607820 675589 607884
rect 675523 607819 675589 607820
rect 675339 595372 675405 595373
rect 675339 595308 675340 595372
rect 675404 595308 675405 595372
rect 675339 595307 675405 595308
rect 675155 592924 675221 592925
rect 675155 592860 675156 592924
rect 675220 592860 675221 592924
rect 675155 592859 675221 592860
rect 675342 592109 675402 595307
rect 675526 593197 675586 607819
rect 675523 593196 675589 593197
rect 675523 593132 675524 593196
rect 675588 593132 675589 593196
rect 675523 593131 675589 593132
rect 675339 592108 675405 592109
rect 675339 592044 675340 592108
rect 675404 592044 675405 592108
rect 675339 592043 675405 592044
rect 676078 591701 676138 631347
rect 676814 619173 676874 694043
rect 676995 644332 677061 644333
rect 676995 644268 676996 644332
rect 677060 644268 677061 644332
rect 676995 644267 677061 644268
rect 676811 619172 676877 619173
rect 676811 619108 676812 619172
rect 676876 619108 676877 619172
rect 676811 619107 676877 619108
rect 676075 591700 676141 591701
rect 676075 591636 676076 591700
rect 676140 591636 676141 591700
rect 676075 591635 676141 591636
rect 676075 586260 676141 586261
rect 676075 586196 676076 586260
rect 676140 586196 676141 586260
rect 676075 586195 676141 586196
rect 675523 562732 675589 562733
rect 675523 562730 675524 562732
rect 675342 562670 675524 562730
rect 675155 550220 675221 550221
rect 675155 550156 675156 550220
rect 675220 550156 675221 550220
rect 675155 550155 675221 550156
rect 675158 547637 675218 550155
rect 675155 547636 675221 547637
rect 675155 547572 675156 547636
rect 675220 547572 675221 547636
rect 675155 547571 675221 547572
rect 675342 545597 675402 562670
rect 675523 562668 675524 562670
rect 675588 562668 675589 562732
rect 675523 562667 675589 562668
rect 675523 561236 675589 561237
rect 675523 561172 675524 561236
rect 675588 561172 675589 561236
rect 675523 561171 675589 561172
rect 675526 546141 675586 561171
rect 676078 547637 676138 586195
rect 676998 572797 677058 644267
rect 676995 572796 677061 572797
rect 676995 572732 676996 572796
rect 677060 572732 677061 572796
rect 676995 572731 677061 572732
rect 676811 557564 676877 557565
rect 676811 557500 676812 557564
rect 676876 557500 676877 557564
rect 676811 557499 676877 557500
rect 676075 547636 676141 547637
rect 676075 547572 676076 547636
rect 676140 547572 676141 547636
rect 676075 547571 676141 547572
rect 675523 546140 675589 546141
rect 675523 546076 675524 546140
rect 675588 546076 675589 546140
rect 675523 546075 675589 546076
rect 675339 545596 675405 545597
rect 675339 545532 675340 545596
rect 675404 545532 675405 545596
rect 675339 545531 675405 545532
rect 676814 492829 676874 557499
rect 676995 550356 677061 550357
rect 676995 550292 676996 550356
rect 677060 550292 677061 550356
rect 676995 550291 677061 550292
rect 676998 503709 677058 550291
rect 676995 503708 677061 503709
rect 676995 503644 676996 503708
rect 677060 503644 677061 503708
rect 676995 503643 677061 503644
rect 676811 492828 676877 492829
rect 676811 492764 676812 492828
rect 676876 492764 676877 492828
rect 676811 492763 676877 492764
rect 675891 488884 675957 488885
rect 675891 488820 675892 488884
rect 675956 488820 675957 488884
rect 675891 488819 675957 488820
rect 675894 488610 675954 488819
rect 675894 488550 676874 488610
rect 674603 475420 674669 475421
rect 674603 475356 674604 475420
rect 674668 475356 674669 475420
rect 674603 475355 674669 475356
rect 673867 455292 673933 455293
rect 673867 455228 673868 455292
rect 673932 455228 673933 455292
rect 673867 455227 673933 455228
rect 675339 453796 675405 453797
rect 675339 453732 675340 453796
rect 675404 453732 675405 453796
rect 675339 453731 675405 453732
rect 41827 425236 41893 425237
rect 41827 425172 41828 425236
rect 41892 425172 41893 425236
rect 41827 425171 41893 425172
rect 41830 424690 41890 425171
rect 42011 424828 42077 424829
rect 42011 424764 42012 424828
rect 42076 424764 42077 424828
rect 42011 424763 42077 424764
rect 41646 424630 41890 424690
rect 41459 418844 41525 418845
rect 41459 418780 41460 418844
rect 41524 418780 41525 418844
rect 41459 418779 41525 418780
rect 40723 418572 40789 418573
rect 40723 418508 40724 418572
rect 40788 418508 40789 418572
rect 40723 418507 40789 418508
rect 40539 418300 40605 418301
rect 40539 418236 40540 418300
rect 40604 418236 40605 418300
rect 40539 418235 40605 418236
rect 40542 403885 40602 418235
rect 40726 409461 40786 418507
rect 40723 409460 40789 409461
rect 40723 409396 40724 409460
rect 40788 409396 40789 409460
rect 40723 409395 40789 409396
rect 40539 403884 40605 403885
rect 40539 403820 40540 403884
rect 40604 403820 40605 403884
rect 40539 403819 40605 403820
rect 41462 398853 41522 418779
rect 41646 402990 41706 424630
rect 42014 424010 42074 424763
rect 41830 423950 42074 424010
rect 41830 406333 41890 423950
rect 42011 421972 42077 421973
rect 42011 421908 42012 421972
rect 42076 421908 42077 421972
rect 42011 421907 42077 421908
rect 42014 418301 42074 421907
rect 42011 418300 42077 418301
rect 42011 418236 42012 418300
rect 42076 418236 42077 418300
rect 42011 418235 42077 418236
rect 675342 410549 675402 453731
rect 675339 410548 675405 410549
rect 675339 410484 675340 410548
rect 675404 410484 675405 410548
rect 675339 410483 675405 410484
rect 41827 406332 41893 406333
rect 41827 406268 41828 406332
rect 41892 406268 41893 406332
rect 41827 406267 41893 406268
rect 41646 402930 41890 402990
rect 41830 401981 41890 402930
rect 41827 401980 41893 401981
rect 41827 401916 41828 401980
rect 41892 401916 41893 401980
rect 41827 401915 41893 401916
rect 676814 401301 676874 488550
rect 676811 401300 676877 401301
rect 676811 401236 676812 401300
rect 676876 401236 676877 401300
rect 676811 401235 676877 401236
rect 41459 398852 41525 398853
rect 41459 398788 41460 398852
rect 41524 398788 41525 398852
rect 41459 398787 41525 398788
rect 676075 398852 676141 398853
rect 676075 398788 676076 398852
rect 676140 398788 676141 398852
rect 676075 398787 676141 398788
rect 675891 389060 675957 389061
rect 675891 388996 675892 389060
rect 675956 388996 675957 389060
rect 675891 388995 675957 388996
rect 675707 387700 675773 387701
rect 675707 387636 675708 387700
rect 675772 387636 675773 387700
rect 675707 387635 675773 387636
rect 41459 381852 41525 381853
rect 41459 381788 41460 381852
rect 41524 381788 41525 381852
rect 41459 381787 41525 381788
rect 40539 378588 40605 378589
rect 40539 378524 40540 378588
rect 40604 378524 40605 378588
rect 40539 378523 40605 378524
rect 40355 375732 40421 375733
rect 40355 375668 40356 375732
rect 40420 375668 40421 375732
rect 40355 375667 40421 375668
rect 40358 368661 40418 375667
rect 40355 368660 40421 368661
rect 40355 368596 40356 368660
rect 40420 368596 40421 368660
rect 40355 368595 40421 368596
rect 40542 360093 40602 378523
rect 40723 378180 40789 378181
rect 40723 378116 40724 378180
rect 40788 378116 40789 378180
rect 40723 378115 40789 378116
rect 40726 363765 40786 378115
rect 40907 377772 40973 377773
rect 40907 377708 40908 377772
rect 40972 377708 40973 377772
rect 40907 377707 40973 377708
rect 40910 364309 40970 377707
rect 40907 364308 40973 364309
rect 40907 364244 40908 364308
rect 40972 364244 40973 364308
rect 40907 364243 40973 364244
rect 40723 363764 40789 363765
rect 40723 363700 40724 363764
rect 40788 363700 40789 363764
rect 40723 363699 40789 363700
rect 40539 360092 40605 360093
rect 40539 360028 40540 360092
rect 40604 360028 40605 360092
rect 40539 360027 40605 360028
rect 41462 358733 41522 381787
rect 675710 378725 675770 387635
rect 675707 378724 675773 378725
rect 675707 378660 675708 378724
rect 675772 378660 675773 378724
rect 675707 378659 675773 378660
rect 674787 378044 674853 378045
rect 674787 377980 674788 378044
rect 674852 377980 674853 378044
rect 674787 377979 674853 377980
rect 41643 376956 41709 376957
rect 41643 376892 41644 376956
rect 41708 376892 41709 376956
rect 41643 376891 41709 376892
rect 41646 360210 41706 376891
rect 674790 372605 674850 377979
rect 675894 373013 675954 388995
rect 676078 376957 676138 398787
rect 676627 396812 676693 396813
rect 676627 396748 676628 396812
rect 676692 396748 676693 396812
rect 676627 396747 676693 396748
rect 676259 395180 676325 395181
rect 676259 395116 676260 395180
rect 676324 395116 676325 395180
rect 676259 395115 676325 395116
rect 676262 377365 676322 395115
rect 676443 394772 676509 394773
rect 676443 394708 676444 394772
rect 676508 394708 676509 394772
rect 676443 394707 676509 394708
rect 676446 380629 676506 394707
rect 676630 384981 676690 396747
rect 676627 384980 676693 384981
rect 676627 384916 676628 384980
rect 676692 384916 676693 384980
rect 676627 384915 676693 384916
rect 676443 380628 676509 380629
rect 676443 380564 676444 380628
rect 676508 380564 676509 380628
rect 676443 380563 676509 380564
rect 676259 377364 676325 377365
rect 676259 377300 676260 377364
rect 676324 377300 676325 377364
rect 676259 377299 676325 377300
rect 676075 376956 676141 376957
rect 676075 376892 676076 376956
rect 676140 376892 676141 376956
rect 676075 376891 676141 376892
rect 675891 373012 675957 373013
rect 675891 372948 675892 373012
rect 675956 372948 675957 373012
rect 675891 372947 675957 372948
rect 674787 372604 674853 372605
rect 674787 372540 674788 372604
rect 674852 372540 674853 372604
rect 674787 372539 674853 372540
rect 41827 371380 41893 371381
rect 41827 371316 41828 371380
rect 41892 371316 41893 371380
rect 41827 371315 41893 371316
rect 41830 362949 41890 371315
rect 41827 362948 41893 362949
rect 41827 362884 41828 362948
rect 41892 362884 41893 362948
rect 41827 362883 41893 362884
rect 41646 360150 41890 360210
rect 41459 358732 41525 358733
rect 41459 358668 41460 358732
rect 41524 358668 41525 358732
rect 41459 358667 41525 358668
rect 41830 355741 41890 360150
rect 41827 355740 41893 355741
rect 41827 355676 41828 355740
rect 41892 355676 41893 355740
rect 41827 355675 41893 355676
rect 675339 354244 675405 354245
rect 675339 354180 675340 354244
rect 675404 354180 675405 354244
rect 675339 354179 675405 354180
rect 675155 349212 675221 349213
rect 675155 349148 675156 349212
rect 675220 349148 675221 349212
rect 675155 349147 675221 349148
rect 44219 342956 44285 342957
rect 44219 342892 44220 342956
rect 44284 342892 44285 342956
rect 44219 342891 44285 342892
rect 43667 340508 43733 340509
rect 43667 340444 43668 340508
rect 43732 340444 43733 340508
rect 43667 340443 43733 340444
rect 40723 338604 40789 338605
rect 40723 338540 40724 338604
rect 40788 338540 40789 338604
rect 40723 338539 40789 338540
rect 40539 336972 40605 336973
rect 40539 336908 40540 336972
rect 40604 336908 40605 336972
rect 40539 336907 40605 336908
rect 40542 316845 40602 336907
rect 40726 324730 40786 338539
rect 42931 337652 42997 337653
rect 42931 337588 42932 337652
rect 42996 337588 42997 337652
rect 42931 337587 42997 337588
rect 41827 336564 41893 336565
rect 41827 336500 41828 336564
rect 41892 336500 41893 336564
rect 41827 336499 41893 336500
rect 40907 333708 40973 333709
rect 40907 333644 40908 333708
rect 40972 333644 40973 333708
rect 40907 333643 40973 333644
rect 40910 325413 40970 333643
rect 41643 327724 41709 327725
rect 41643 327660 41644 327724
rect 41708 327660 41709 327724
rect 41643 327659 41709 327660
rect 40907 325412 40973 325413
rect 40907 325348 40908 325412
rect 40972 325348 40973 325412
rect 40907 325347 40973 325348
rect 40726 324670 41522 324730
rect 40539 316844 40605 316845
rect 40539 316780 40540 316844
rect 40604 316780 40605 316844
rect 40539 316779 40605 316780
rect 41462 315621 41522 324670
rect 41646 319970 41706 327659
rect 41830 324733 41890 336499
rect 42747 335476 42813 335477
rect 42747 335412 42748 335476
rect 42812 335412 42813 335476
rect 42747 335411 42813 335412
rect 42750 334661 42810 335411
rect 42747 334660 42813 334661
rect 42747 334596 42748 334660
rect 42812 334596 42813 334660
rect 42747 334595 42813 334596
rect 42011 329084 42077 329085
rect 42011 329020 42012 329084
rect 42076 329020 42077 329084
rect 42011 329019 42077 329020
rect 41827 324732 41893 324733
rect 41827 324668 41828 324732
rect 41892 324668 41893 324732
rect 41827 324667 41893 324668
rect 41827 319972 41893 319973
rect 41827 319970 41828 319972
rect 41646 319910 41828 319970
rect 41827 319908 41828 319910
rect 41892 319908 41893 319972
rect 41827 319907 41893 319908
rect 41459 315620 41525 315621
rect 41459 315556 41460 315620
rect 41524 315556 41525 315620
rect 41459 315555 41525 315556
rect 42014 312629 42074 329019
rect 42934 312765 42994 337587
rect 43299 337244 43365 337245
rect 43299 337180 43300 337244
rect 43364 337180 43365 337244
rect 43299 337179 43365 337180
rect 43115 336156 43181 336157
rect 43115 336092 43116 336156
rect 43180 336092 43181 336156
rect 43115 336091 43181 336092
rect 43118 334661 43178 336091
rect 43115 334660 43181 334661
rect 43115 334596 43116 334660
rect 43180 334596 43181 334660
rect 43115 334595 43181 334596
rect 43302 316050 43362 337179
rect 43118 316029 43362 316050
rect 43115 316028 43362 316029
rect 43115 315964 43116 316028
rect 43180 315990 43362 316028
rect 43180 315964 43181 315990
rect 43115 315963 43181 315964
rect 42931 312764 42997 312765
rect 42931 312700 42932 312764
rect 42996 312700 42997 312764
rect 42931 312699 42997 312700
rect 42011 312628 42077 312629
rect 42011 312564 42012 312628
rect 42076 312564 42077 312628
rect 42011 312563 42077 312564
rect 43670 297669 43730 340443
rect 43851 335748 43917 335749
rect 43851 335684 43852 335748
rect 43916 335684 43917 335748
rect 43851 335683 43917 335684
rect 43854 334661 43914 335683
rect 43851 334660 43917 334661
rect 43851 334596 43852 334660
rect 43916 334596 43917 334660
rect 43851 334595 43917 334596
rect 44222 311130 44282 342891
rect 44403 342140 44469 342141
rect 44403 342076 44404 342140
rect 44468 342076 44469 342140
rect 44403 342075 44469 342076
rect 44406 331230 44466 342075
rect 675158 340890 675218 349147
rect 675342 345130 675402 354179
rect 675707 353836 675773 353837
rect 675707 353772 675708 353836
rect 675772 353772 675773 353836
rect 675707 353771 675773 353772
rect 675710 345810 675770 353771
rect 675891 351932 675957 351933
rect 675891 351868 675892 351932
rect 675956 351930 675957 351932
rect 675956 351870 676322 351930
rect 675956 351868 675957 351870
rect 675891 351867 675957 351868
rect 676262 351250 676322 351870
rect 676262 351190 676690 351250
rect 675891 350980 675957 350981
rect 675891 350916 675892 350980
rect 675956 350916 675957 350980
rect 675891 350915 675957 350916
rect 675894 350570 675954 350915
rect 675894 350510 676506 350570
rect 675891 350164 675957 350165
rect 675891 350100 675892 350164
rect 675956 350100 675957 350164
rect 675891 350099 675957 350100
rect 675894 349890 675954 350099
rect 675894 349830 676322 349890
rect 675710 345750 676138 345810
rect 675342 345070 675770 345130
rect 675710 340890 675770 345070
rect 675158 340830 675586 340890
rect 675710 340830 675954 340890
rect 675526 337789 675586 340830
rect 675894 339421 675954 340830
rect 675891 339420 675957 339421
rect 675891 339356 675892 339420
rect 675956 339356 675957 339420
rect 675891 339355 675957 339356
rect 675523 337788 675589 337789
rect 675523 337724 675524 337788
rect 675588 337724 675589 337788
rect 675523 337723 675589 337724
rect 674787 336700 674853 336701
rect 674787 336636 674788 336700
rect 674852 336636 674853 336700
rect 674787 336635 674853 336636
rect 44406 331170 44650 331230
rect 44590 311405 44650 331170
rect 674790 326909 674850 336635
rect 676078 328405 676138 345750
rect 676262 332349 676322 349830
rect 676446 335341 676506 350510
rect 676630 340237 676690 351190
rect 676627 340236 676693 340237
rect 676627 340172 676628 340236
rect 676692 340172 676693 340236
rect 676627 340171 676693 340172
rect 676443 335340 676509 335341
rect 676443 335276 676444 335340
rect 676508 335276 676509 335340
rect 676443 335275 676509 335276
rect 676259 332348 676325 332349
rect 676259 332284 676260 332348
rect 676324 332284 676325 332348
rect 676259 332283 676325 332284
rect 676075 328404 676141 328405
rect 676075 328340 676076 328404
rect 676140 328340 676141 328404
rect 676075 328339 676141 328340
rect 674787 326908 674853 326909
rect 674787 326844 674788 326908
rect 674852 326844 674853 326908
rect 674787 326843 674853 326844
rect 44587 311404 44653 311405
rect 44587 311340 44588 311404
rect 44652 311340 44653 311404
rect 44587 311339 44653 311340
rect 44403 311132 44469 311133
rect 44403 311130 44404 311132
rect 44222 311070 44404 311130
rect 44403 311068 44404 311070
rect 44468 311068 44469 311132
rect 44403 311067 44469 311068
rect 675707 308820 675773 308821
rect 675707 308756 675708 308820
rect 675772 308756 675773 308820
rect 675707 308755 675773 308756
rect 675710 302250 675770 308755
rect 675891 306780 675957 306781
rect 675891 306716 675892 306780
rect 675956 306716 675957 306780
rect 675891 306715 675957 306716
rect 675894 306370 675954 306715
rect 675894 306310 676874 306370
rect 675891 305964 675957 305965
rect 675891 305900 675892 305964
rect 675956 305900 675957 305964
rect 675891 305899 675957 305900
rect 675894 305690 675954 305899
rect 675894 305630 676506 305690
rect 676029 305148 676095 305149
rect 676029 305084 676030 305148
rect 676094 305146 676095 305148
rect 676094 305084 676138 305146
rect 676029 305083 676138 305084
rect 676078 305010 676138 305083
rect 676078 304950 676322 305010
rect 675710 302190 676138 302250
rect 675707 299436 675773 299437
rect 675707 299372 675708 299436
rect 675772 299372 675773 299436
rect 675707 299371 675773 299372
rect 43667 297668 43733 297669
rect 43667 297604 43668 297668
rect 43732 297604 43733 297668
rect 43667 297603 43733 297604
rect 675523 297668 675589 297669
rect 675523 297604 675524 297668
rect 675588 297604 675589 297668
rect 675523 297603 675589 297604
rect 675339 296716 675405 296717
rect 675339 296652 675340 296716
rect 675404 296652 675405 296716
rect 675339 296651 675405 296652
rect 42011 296444 42077 296445
rect 42011 296380 42012 296444
rect 42076 296380 42077 296444
rect 42011 296379 42077 296380
rect 41827 295628 41893 295629
rect 41827 295564 41828 295628
rect 41892 295564 41893 295628
rect 41827 295563 41893 295564
rect 41830 294130 41890 295563
rect 40726 294070 41890 294130
rect 40539 292592 40605 292593
rect 40539 292528 40540 292592
rect 40604 292528 40605 292592
rect 40539 292527 40605 292528
rect 40542 274277 40602 292527
rect 40726 277677 40786 294070
rect 41827 292908 41893 292909
rect 41827 292844 41828 292908
rect 41892 292844 41893 292908
rect 41827 292843 41893 292844
rect 40907 292592 40973 292593
rect 40907 292528 40908 292592
rect 40972 292528 40973 292592
rect 41830 292590 41890 292843
rect 40907 292527 40973 292528
rect 41646 292530 41890 292590
rect 40910 277949 40970 292527
rect 41646 289830 41706 292530
rect 41827 292228 41893 292229
rect 41827 292164 41828 292228
rect 41892 292164 41893 292228
rect 41827 292163 41893 292164
rect 41462 289770 41706 289830
rect 40907 277948 40973 277949
rect 40907 277884 40908 277948
rect 40972 277884 40973 277948
rect 40907 277883 40973 277884
rect 40723 277676 40789 277677
rect 40723 277612 40724 277676
rect 40788 277612 40789 277676
rect 40723 277611 40789 277612
rect 40539 274276 40605 274277
rect 40539 274212 40540 274276
rect 40604 274212 40605 274276
rect 40539 274211 40605 274212
rect 41462 270469 41522 289770
rect 41459 270468 41525 270469
rect 41459 270404 41460 270468
rect 41524 270404 41525 270468
rect 41459 270403 41525 270404
rect 41830 269109 41890 292163
rect 42014 281485 42074 296379
rect 675342 292909 675402 296651
rect 675339 292908 675405 292909
rect 675339 292844 675340 292908
rect 675404 292844 675405 292908
rect 675339 292843 675405 292844
rect 675526 292093 675586 297603
rect 675523 292092 675589 292093
rect 675523 292028 675524 292092
rect 675588 292028 675589 292092
rect 675523 292027 675589 292028
rect 675710 282845 675770 299371
rect 675891 297396 675957 297397
rect 675891 297332 675892 297396
rect 675956 297332 675957 297396
rect 675891 297331 675957 297332
rect 675707 282844 675773 282845
rect 675707 282780 675708 282844
rect 675772 282780 675773 282844
rect 675707 282779 675773 282780
rect 42011 281484 42077 281485
rect 42011 281420 42012 281484
rect 42076 281420 42077 281484
rect 42011 281419 42077 281420
rect 675894 281213 675954 297331
rect 676078 283661 676138 302190
rect 676262 287061 676322 304950
rect 676446 291549 676506 305630
rect 676814 295221 676874 306310
rect 676811 295220 676877 295221
rect 676811 295156 676812 295220
rect 676876 295156 676877 295220
rect 676811 295155 676877 295156
rect 676443 291548 676509 291549
rect 676443 291484 676444 291548
rect 676508 291484 676509 291548
rect 676443 291483 676509 291484
rect 676259 287060 676325 287061
rect 676259 286996 676260 287060
rect 676324 286996 676325 287060
rect 676259 286995 676325 286996
rect 676075 283660 676141 283661
rect 676075 283596 676076 283660
rect 676140 283596 676141 283660
rect 676075 283595 676141 283596
rect 675891 281212 675957 281213
rect 675891 281148 675892 281212
rect 675956 281148 675957 281212
rect 675891 281147 675957 281148
rect 41827 269108 41893 269109
rect 41827 269044 41828 269108
rect 41892 269044 41893 269108
rect 41827 269043 41893 269044
rect 676075 263668 676141 263669
rect 676075 263604 676076 263668
rect 676140 263604 676141 263668
rect 676075 263603 676141 263604
rect 675891 261220 675957 261221
rect 675891 261156 675892 261220
rect 675956 261156 675957 261220
rect 675891 261155 675957 261156
rect 40539 251428 40605 251429
rect 40539 251364 40540 251428
rect 40604 251364 40605 251428
rect 40539 251363 40605 251364
rect 40542 240141 40602 251363
rect 40723 249796 40789 249797
rect 40723 249732 40724 249796
rect 40788 249732 40789 249796
rect 40723 249731 40789 249732
rect 40539 240140 40605 240141
rect 40539 240076 40540 240140
rect 40604 240076 40605 240140
rect 40539 240075 40605 240076
rect 40726 235925 40786 249731
rect 675894 249661 675954 261155
rect 676078 249661 676138 263603
rect 676995 261628 677061 261629
rect 676995 261564 676996 261628
rect 677060 261564 677061 261628
rect 676995 261563 677061 261564
rect 676811 259996 676877 259997
rect 676811 259932 676812 259996
rect 676876 259932 676877 259996
rect 676811 259931 676877 259932
rect 675891 249660 675957 249661
rect 675891 249596 675892 249660
rect 675956 249596 675957 249660
rect 675891 249595 675957 249596
rect 676075 249660 676141 249661
rect 676075 249596 676076 249660
rect 676140 249596 676141 249660
rect 676075 249595 676141 249596
rect 675339 245580 675405 245581
rect 675339 245516 675340 245580
rect 675404 245516 675405 245580
rect 675339 245515 675405 245516
rect 675342 238645 675402 245515
rect 676814 245309 676874 259931
rect 676998 250341 677058 261563
rect 676995 250340 677061 250341
rect 676995 250276 676996 250340
rect 677060 250276 677061 250340
rect 676995 250275 677061 250276
rect 676811 245308 676877 245309
rect 676811 245244 676812 245308
rect 676876 245244 676877 245308
rect 676811 245243 676877 245244
rect 675339 238644 675405 238645
rect 675339 238580 675340 238644
rect 675404 238580 675405 238644
rect 675339 238579 675405 238580
rect 42011 238100 42077 238101
rect 42011 238036 42012 238100
rect 42076 238036 42077 238100
rect 42011 238035 42077 238036
rect 40723 235924 40789 235925
rect 40723 235860 40724 235924
rect 40788 235860 40789 235924
rect 40723 235859 40789 235860
rect 42014 228989 42074 238035
rect 676811 236332 676877 236333
rect 676811 236268 676812 236332
rect 676876 236268 676877 236332
rect 676811 236267 676877 236268
rect 673499 236060 673565 236061
rect 673499 235996 673500 236060
rect 673564 235996 673565 236060
rect 673499 235995 673565 235996
rect 671291 234564 671357 234565
rect 671291 234500 671292 234564
rect 671356 234500 671357 234564
rect 671291 234499 671357 234500
rect 42011 228988 42077 228989
rect 42011 228924 42012 228988
rect 42076 228924 42077 228988
rect 42011 228923 42077 228924
rect 669819 220964 669885 220965
rect 669819 220900 669820 220964
rect 669884 220900 669885 220964
rect 669819 220899 669885 220900
rect 505050 218502 505054 218650
rect 553531 218652 553597 218653
rect 553531 218588 553532 218652
rect 553596 218650 553597 218652
rect 563102 218650 563162 219182
rect 553596 218590 553778 218650
rect 553596 218588 553597 218590
rect 553531 218587 553597 218588
rect 505050 218381 505110 218502
rect 493915 218380 493981 218381
rect 493915 218316 493916 218380
rect 493980 218316 493981 218380
rect 493915 218315 493981 218316
rect 505047 218380 505113 218381
rect 505047 218316 505048 218380
rect 505112 218316 505113 218380
rect 505047 218315 505113 218316
rect 493918 218058 493978 218315
rect 553718 217837 553778 218590
rect 562550 218590 563162 218650
rect 572486 218650 572546 219182
rect 572486 218590 572730 218650
rect 562550 217837 562610 218590
rect 572670 218381 572730 218590
rect 572667 218380 572733 218381
rect 572667 218316 572668 218380
rect 572732 218316 572733 218380
rect 572667 218315 572733 218316
rect 553715 217836 553781 217837
rect 493918 217701 493978 217822
rect 553715 217772 553716 217836
rect 553780 217772 553781 217836
rect 553715 217771 553781 217772
rect 562547 217836 562613 217837
rect 562547 217772 562548 217836
rect 562612 217772 562613 217836
rect 562547 217771 562613 217772
rect 493915 217700 493981 217701
rect 493915 217636 493916 217700
rect 493980 217636 493981 217700
rect 493915 217635 493981 217636
rect 576534 217290 576594 218502
rect 576807 217292 576873 217293
rect 576807 217290 576808 217292
rect 576534 217230 576808 217290
rect 576807 217228 576808 217230
rect 576872 217228 576873 217292
rect 576807 217227 576873 217228
rect 578190 213213 578250 217822
rect 666323 217292 666389 217293
rect 666323 217228 666324 217292
rect 666388 217228 666389 217292
rect 666323 217227 666389 217228
rect 578187 213212 578253 213213
rect 578187 213148 578188 213212
rect 578252 213148 578253 213212
rect 578187 213147 578253 213148
rect 666326 209790 666386 217227
rect 669822 215310 669882 220899
rect 670371 220692 670437 220693
rect 670371 220628 670372 220692
rect 670436 220690 670437 220692
rect 671107 220692 671173 220693
rect 671107 220690 671108 220692
rect 670436 220630 671108 220690
rect 670436 220628 670437 220630
rect 670371 220627 670437 220628
rect 671107 220628 671108 220630
rect 671172 220628 671173 220692
rect 671107 220627 671173 220628
rect 669454 215250 669882 215310
rect 666326 209730 666570 209790
rect 41643 209404 41709 209405
rect 41643 209340 41644 209404
rect 41708 209340 41709 209404
rect 41643 209339 41709 209340
rect 40539 208180 40605 208181
rect 40539 208116 40540 208180
rect 40604 208116 40605 208180
rect 40539 208115 40605 208116
rect 40542 197165 40602 208115
rect 41646 205650 41706 209339
rect 41827 207364 41893 207365
rect 41827 207300 41828 207364
rect 41892 207300 41893 207364
rect 41827 207299 41893 207300
rect 41462 205590 41706 205650
rect 40539 197164 40605 197165
rect 40539 197100 40540 197164
rect 40604 197100 40605 197164
rect 40539 197099 40605 197100
rect 41462 184109 41522 205590
rect 41643 204508 41709 204509
rect 41643 204444 41644 204508
rect 41708 204444 41709 204508
rect 41643 204443 41709 204444
rect 41646 190470 41706 204443
rect 41830 195261 41890 207299
rect 666510 202890 666570 209730
rect 667979 206548 668045 206549
rect 667979 206484 667980 206548
rect 668044 206484 668045 206548
rect 667979 206483 668045 206484
rect 666510 202830 666754 202890
rect 666694 198389 666754 202830
rect 666691 198388 666757 198389
rect 666691 198324 666692 198388
rect 666756 198324 666757 198388
rect 666691 198323 666757 198324
rect 41827 195260 41893 195261
rect 41827 195196 41828 195260
rect 41892 195196 41893 195260
rect 41827 195195 41893 195196
rect 41646 190410 41890 190470
rect 41830 185877 41890 190410
rect 41827 185876 41893 185877
rect 41827 185812 41828 185876
rect 41892 185812 41893 185876
rect 41827 185811 41893 185812
rect 41459 184108 41525 184109
rect 41459 184044 41460 184108
rect 41524 184044 41525 184108
rect 41459 184043 41525 184044
rect 667982 130661 668042 206483
rect 669083 206276 669149 206277
rect 669083 206212 669084 206276
rect 669148 206212 669149 206276
rect 669083 206211 669149 206212
rect 669086 202469 669146 206211
rect 669083 202468 669149 202469
rect 669083 202404 669084 202468
rect 669148 202404 669149 202468
rect 669083 202403 669149 202404
rect 669454 157350 669514 215250
rect 670739 211172 670805 211173
rect 670739 211108 670740 211172
rect 670804 211108 670805 211172
rect 670739 211107 670805 211108
rect 670742 164253 670802 211107
rect 670739 164252 670805 164253
rect 670739 164188 670740 164252
rect 670804 164188 670805 164252
rect 670739 164187 670805 164188
rect 669270 157290 669514 157350
rect 669270 137869 669330 157290
rect 671294 145349 671354 234499
rect 673502 232797 673562 235995
rect 673499 232796 673565 232797
rect 673499 232732 673500 232796
rect 673564 232732 673565 232796
rect 673499 232731 673565 232732
rect 673131 231844 673197 231845
rect 673131 231780 673132 231844
rect 673196 231780 673197 231844
rect 673131 231779 673197 231780
rect 673315 231844 673381 231845
rect 673315 231780 673316 231844
rect 673380 231780 673381 231844
rect 673315 231779 673381 231780
rect 674235 231844 674301 231845
rect 674235 231780 674236 231844
rect 674300 231780 674301 231844
rect 674235 231779 674301 231780
rect 671475 229396 671541 229397
rect 671475 229332 671476 229396
rect 671540 229332 671541 229396
rect 671475 229331 671541 229332
rect 671478 224909 671538 229331
rect 672947 228580 673013 228581
rect 672947 228516 672948 228580
rect 673012 228516 673013 228580
rect 672947 228515 673013 228516
rect 671843 227084 671909 227085
rect 671843 227020 671844 227084
rect 671908 227020 671909 227084
rect 671843 227019 671909 227020
rect 671659 226948 671725 226949
rect 671659 226884 671660 226948
rect 671724 226884 671725 226948
rect 671659 226883 671725 226884
rect 671475 224908 671541 224909
rect 671475 224844 671476 224908
rect 671540 224844 671541 224908
rect 671475 224843 671541 224844
rect 671662 224365 671722 226883
rect 671659 224364 671725 224365
rect 671659 224300 671660 224364
rect 671724 224300 671725 224364
rect 671659 224299 671725 224300
rect 671846 220421 671906 227019
rect 672763 225724 672829 225725
rect 672763 225660 672764 225724
rect 672828 225660 672829 225724
rect 672763 225659 672829 225660
rect 672766 223957 672826 225659
rect 672763 223956 672829 223957
rect 672763 223892 672764 223956
rect 672828 223892 672829 223956
rect 672763 223891 672829 223892
rect 671843 220420 671909 220421
rect 671843 220356 671844 220420
rect 671908 220356 671909 220420
rect 671843 220355 671909 220356
rect 672950 183565 673010 228515
rect 673134 222325 673194 231779
rect 673131 222324 673197 222325
rect 673131 222260 673132 222324
rect 673196 222260 673197 222324
rect 673131 222259 673197 222260
rect 673318 222210 673378 231779
rect 673318 222150 673562 222210
rect 673131 209676 673197 209677
rect 673131 209612 673132 209676
rect 673196 209612 673197 209676
rect 673131 209611 673197 209612
rect 672947 183564 673013 183565
rect 672947 183500 672948 183564
rect 673012 183500 673013 183564
rect 672947 183499 673013 183500
rect 671291 145348 671357 145349
rect 671291 145284 671292 145348
rect 671356 145284 671357 145348
rect 671291 145283 671357 145284
rect 669267 137868 669333 137869
rect 669267 137804 669268 137868
rect 669332 137804 669333 137868
rect 669267 137803 669333 137804
rect 673134 133925 673194 209611
rect 673131 133924 673197 133925
rect 673131 133860 673132 133924
rect 673196 133860 673197 133924
rect 673131 133859 673197 133860
rect 667979 130660 668045 130661
rect 667979 130596 667980 130660
rect 668044 130596 668045 130660
rect 667979 130595 668045 130596
rect 673502 128893 673562 222150
rect 674238 215310 674298 231779
rect 674971 228580 675037 228581
rect 674971 228516 674972 228580
rect 675036 228516 675037 228580
rect 674971 228515 675037 228516
rect 674974 217837 675034 228515
rect 675523 218652 675589 218653
rect 675523 218588 675524 218652
rect 675588 218588 675589 218652
rect 675523 218587 675589 218588
rect 674971 217836 675037 217837
rect 674971 217772 674972 217836
rect 675036 217772 675037 217836
rect 674971 217771 675037 217772
rect 673686 215250 674298 215310
rect 673686 141133 673746 215250
rect 674051 212124 674117 212125
rect 674051 212060 674052 212124
rect 674116 212060 674117 212124
rect 674051 212059 674117 212060
rect 673683 141132 673749 141133
rect 673683 141068 673684 141132
rect 673748 141068 673749 141132
rect 673683 141067 673749 141068
rect 673499 128892 673565 128893
rect 673499 128828 673500 128892
rect 673564 128828 673565 128892
rect 673499 128827 673565 128828
rect 674054 128349 674114 212059
rect 675526 210490 675586 218587
rect 675707 218108 675773 218109
rect 675707 218044 675708 218108
rect 675772 218044 675773 218108
rect 675707 218043 675773 218044
rect 675710 217834 675770 218043
rect 676078 217910 676506 217970
rect 676078 217834 676138 217910
rect 675710 217774 676138 217834
rect 675707 217020 675773 217021
rect 675707 216956 675708 217020
rect 675772 216956 675773 217020
rect 675707 216955 675773 216956
rect 675710 211170 675770 216955
rect 676259 215150 676325 215151
rect 676259 215086 676260 215150
rect 676324 215086 676325 215150
rect 676259 215085 676325 215086
rect 675710 211110 676138 211170
rect 675526 210430 675954 210490
rect 675707 207092 675773 207093
rect 675707 207028 675708 207092
rect 675772 207028 675773 207092
rect 675707 207027 675773 207028
rect 675710 204237 675770 207027
rect 675707 204236 675773 204237
rect 675707 204172 675708 204236
rect 675772 204172 675773 204236
rect 675707 204171 675773 204172
rect 675894 193221 675954 210430
rect 675891 193220 675957 193221
rect 675891 193156 675892 193220
rect 675956 193156 675957 193220
rect 675891 193155 675957 193156
rect 676078 191589 676138 211110
rect 676262 197165 676322 215085
rect 676446 205597 676506 217910
rect 676814 211445 676874 236267
rect 676811 211444 676877 211445
rect 676811 211380 676812 211444
rect 676876 211380 676877 211444
rect 676811 211379 676877 211380
rect 676995 211444 677061 211445
rect 676995 211380 676996 211444
rect 677060 211380 677061 211444
rect 676995 211379 677061 211380
rect 676443 205596 676509 205597
rect 676443 205532 676444 205596
rect 676508 205532 676509 205596
rect 676443 205531 676509 205532
rect 676998 200837 677058 211379
rect 676995 200836 677061 200837
rect 676995 200772 676996 200836
rect 677060 200772 677061 200836
rect 676995 200771 677061 200772
rect 676259 197164 676325 197165
rect 676259 197100 676260 197164
rect 676324 197100 676325 197164
rect 676259 197099 676325 197100
rect 676075 191588 676141 191589
rect 676075 191524 676076 191588
rect 676140 191524 676141 191588
rect 676075 191523 676141 191524
rect 675891 174044 675957 174045
rect 675891 173980 675892 174044
rect 675956 173980 675957 174044
rect 675891 173979 675957 173980
rect 675894 173770 675954 173979
rect 675894 173710 676506 173770
rect 675707 173636 675773 173637
rect 675707 173572 675708 173636
rect 675772 173572 675773 173636
rect 675707 173571 675773 173572
rect 675710 171050 675770 173571
rect 675891 172412 675957 172413
rect 675891 172348 675892 172412
rect 675956 172410 675957 172412
rect 675956 172350 676322 172410
rect 675956 172348 675957 172350
rect 675891 172347 675957 172348
rect 675710 170990 676138 171050
rect 675707 170372 675773 170373
rect 675707 170308 675708 170372
rect 675772 170308 675773 170372
rect 675707 170307 675773 170308
rect 675710 150381 675770 170307
rect 675891 167516 675957 167517
rect 675891 167452 675892 167516
rect 675956 167452 675957 167516
rect 675891 167451 675957 167452
rect 675707 150380 675773 150381
rect 675707 150316 675708 150380
rect 675772 150316 675773 150380
rect 675707 150315 675773 150316
rect 675894 147661 675954 167451
rect 676078 148477 676138 170990
rect 676262 151605 676322 172350
rect 676446 159357 676506 173710
rect 676627 166428 676693 166429
rect 676627 166364 676628 166428
rect 676692 166364 676693 166428
rect 676627 166363 676693 166364
rect 676443 159356 676509 159357
rect 676443 159292 676444 159356
rect 676508 159292 676509 159356
rect 676443 159291 676509 159292
rect 676630 156365 676690 166363
rect 676627 156364 676693 156365
rect 676627 156300 676628 156364
rect 676692 156300 676693 156364
rect 676627 156299 676693 156300
rect 676259 151604 676325 151605
rect 676259 151540 676260 151604
rect 676324 151540 676325 151604
rect 676259 151539 676325 151540
rect 676075 148476 676141 148477
rect 676075 148412 676076 148476
rect 676140 148412 676141 148476
rect 676075 148411 676141 148412
rect 675891 147660 675957 147661
rect 675891 147596 675892 147660
rect 675956 147596 675957 147660
rect 675891 147595 675957 147596
rect 676259 128620 676325 128621
rect 676259 128556 676260 128620
rect 676324 128556 676325 128620
rect 676259 128555 676325 128556
rect 674051 128348 674117 128349
rect 674051 128284 674052 128348
rect 674116 128284 674117 128348
rect 674051 128283 674117 128284
rect 676075 126988 676141 126989
rect 676075 126924 676076 126988
rect 676140 126924 676141 126988
rect 676075 126923 676141 126924
rect 675891 122364 675957 122365
rect 675891 122300 675892 122364
rect 675956 122300 675957 122364
rect 675891 122299 675957 122300
rect 675707 117332 675773 117333
rect 675707 117268 675708 117332
rect 675772 117268 675773 117332
rect 675707 117267 675773 117268
rect 675710 103189 675770 117267
rect 675707 103188 675773 103189
rect 675707 103124 675708 103188
rect 675772 103124 675773 103188
rect 675707 103123 675773 103124
rect 675894 102509 675954 122299
rect 676078 108221 676138 126923
rect 676262 113117 676322 128555
rect 676627 126580 676693 126581
rect 676627 126516 676628 126580
rect 676692 126516 676693 126580
rect 676627 126515 676693 126516
rect 676443 124540 676509 124541
rect 676443 124476 676444 124540
rect 676508 124476 676509 124540
rect 676443 124475 676509 124476
rect 676259 113116 676325 113117
rect 676259 113052 676260 113116
rect 676324 113052 676325 113116
rect 676259 113051 676325 113052
rect 676075 108220 676141 108221
rect 676075 108156 676076 108220
rect 676140 108156 676141 108220
rect 676075 108155 676141 108156
rect 676446 106181 676506 124475
rect 676443 106180 676509 106181
rect 676443 106116 676444 106180
rect 676508 106116 676509 106180
rect 676443 106115 676509 106116
rect 675891 102508 675957 102509
rect 675891 102444 675892 102508
rect 675956 102444 675957 102508
rect 675891 102443 675957 102444
rect 676630 101421 676690 126515
rect 676627 101420 676693 101421
rect 676627 101356 676628 101420
rect 676692 101356 676693 101420
rect 676627 101355 676693 101356
rect 637251 96932 637317 96933
rect 637251 96868 637252 96932
rect 637316 96868 637317 96932
rect 637251 96867 637317 96868
rect 633939 96116 634005 96117
rect 633939 96052 633940 96116
rect 634004 96052 634005 96116
rect 633939 96051 634005 96052
rect 633942 78573 634002 96051
rect 637254 84210 637314 96867
rect 647187 96116 647253 96117
rect 647187 96052 647188 96116
rect 647252 96052 647253 96116
rect 647187 96051 647253 96052
rect 647190 94298 647250 96051
rect 650318 93125 650378 93382
rect 650315 93124 650381 93125
rect 650315 93060 650316 93124
rect 650380 93060 650381 93124
rect 650315 93059 650381 93060
rect 637070 84150 637314 84210
rect 633939 78572 634005 78573
rect 633939 78508 633940 78572
rect 634004 78508 634005 78572
rect 633939 78507 634005 78508
rect 637070 77757 637130 84150
rect 637067 77756 637133 77757
rect 637067 77692 637068 77756
rect 637132 77692 637133 77756
rect 637067 77691 637133 77692
rect 194363 50284 194429 50285
rect 194363 50220 194364 50284
rect 194428 50220 194429 50284
rect 194363 50219 194429 50220
rect 141739 44028 141805 44029
rect 141739 43964 141740 44028
rect 141804 43964 141805 44028
rect 141739 43963 141805 43964
rect 141742 40493 141802 43963
rect 194366 42125 194426 50219
rect 522803 49468 522869 49469
rect 522803 49404 522804 49468
rect 522868 49404 522869 49468
rect 522803 49403 522869 49404
rect 518755 48924 518821 48925
rect 518755 48860 518756 48924
rect 518820 48860 518821 48924
rect 518755 48859 518821 48860
rect 515443 47020 515509 47021
rect 515443 46956 515444 47020
rect 515508 46956 515509 47020
rect 515443 46955 515509 46956
rect 463739 44436 463805 44437
rect 463739 44372 463740 44436
rect 463804 44372 463805 44436
rect 463739 44371 463805 44372
rect 440187 43892 440253 43893
rect 440187 43828 440188 43892
rect 440252 43890 440253 43892
rect 440923 43892 440989 43893
rect 440923 43890 440924 43892
rect 440252 43830 440924 43890
rect 440252 43828 440253 43830
rect 440187 43827 440253 43828
rect 440923 43828 440924 43830
rect 440988 43828 440989 43892
rect 440923 43827 440989 43828
rect 194363 42124 194429 42125
rect 194363 42060 194364 42124
rect 194428 42060 194429 42124
rect 194363 42059 194429 42060
rect 463742 41938 463802 44371
rect 464107 44300 464173 44301
rect 464107 44236 464108 44300
rect 464172 44236 464173 44300
rect 464107 44235 464173 44236
rect 365483 41852 365549 41853
rect 365483 41788 365484 41852
rect 365548 41788 365549 41852
rect 365483 41787 365549 41788
rect 365486 41258 365546 41787
rect 403019 41852 403085 41853
rect 403019 41850 403020 41852
rect 402802 41790 403020 41850
rect 403019 41788 403020 41790
rect 403084 41788 403085 41852
rect 403019 41787 403085 41788
rect 421971 41852 422037 41853
rect 421971 41788 421972 41852
rect 422036 41850 422037 41852
rect 422036 41790 422162 41850
rect 422036 41788 422037 41790
rect 421971 41787 422037 41788
rect 441843 41852 441909 41853
rect 441843 41850 441844 41852
rect 441626 41790 441844 41850
rect 441843 41788 441844 41790
rect 441908 41788 441909 41852
rect 441843 41787 441909 41788
rect 460795 41852 460861 41853
rect 460795 41788 460796 41852
rect 460860 41850 460861 41852
rect 460979 41852 461045 41853
rect 460979 41850 460980 41852
rect 460860 41790 460980 41850
rect 460860 41788 460861 41790
rect 460795 41787 460861 41788
rect 460979 41788 460980 41790
rect 461044 41788 461045 41852
rect 460979 41787 461045 41788
rect 464110 41853 464170 44235
rect 515446 42125 515506 46955
rect 518758 42805 518818 48859
rect 520963 47564 521029 47565
rect 520963 47500 520964 47564
rect 521028 47500 521029 47564
rect 520963 47499 521029 47500
rect 518755 42804 518821 42805
rect 518755 42740 518756 42804
rect 518820 42740 518821 42804
rect 518755 42739 518821 42740
rect 520966 42125 521026 47499
rect 522806 42125 522866 49403
rect 529795 49196 529861 49197
rect 529795 49132 529796 49196
rect 529860 49132 529861 49196
rect 529795 49131 529861 49132
rect 526483 47836 526549 47837
rect 526483 47772 526484 47836
rect 526548 47772 526549 47836
rect 526483 47771 526549 47772
rect 526486 42125 526546 47771
rect 529798 42125 529858 49131
rect 515443 42124 515509 42125
rect 515443 42060 515444 42124
rect 515508 42060 515509 42124
rect 515443 42059 515509 42060
rect 520963 42124 521029 42125
rect 520963 42060 520964 42124
rect 521028 42060 521029 42124
rect 520963 42059 521029 42060
rect 522803 42124 522869 42125
rect 522803 42060 522804 42124
rect 522868 42060 522869 42124
rect 522803 42059 522869 42060
rect 526483 42124 526549 42125
rect 526483 42060 526484 42124
rect 526548 42060 526549 42124
rect 526483 42059 526549 42060
rect 529795 42124 529861 42125
rect 529795 42060 529796 42124
rect 529860 42060 529861 42124
rect 529795 42059 529861 42060
rect 464107 41852 464173 41853
rect 464107 41788 464108 41852
rect 464172 41788 464173 41852
rect 464107 41787 464173 41788
rect 141739 40492 141805 40493
rect 141739 40428 141740 40492
rect 141804 40428 141805 40492
rect 141739 40427 141805 40428
<< via4 >>
rect 172382 997102 172618 997338
rect 245614 997252 245850 997338
rect 245614 997188 245700 997252
rect 245700 997188 245764 997252
rect 245764 997188 245850 997252
rect 245614 997102 245850 997188
rect 536702 993022 536938 993258
rect 572582 993022 572818 993258
rect 563014 219182 563250 219418
rect 572398 219182 572634 219418
rect 505054 218502 505290 218738
rect 493830 217822 494066 218058
rect 576446 218502 576682 218738
rect 578102 217822 578338 218058
rect 647102 94062 647338 94298
rect 650230 93382 650466 93618
rect 361902 41852 362138 41938
rect 361902 41788 361988 41852
rect 361988 41788 362052 41852
rect 362052 41788 362138 41852
rect 361902 41702 362138 41788
rect 402566 41702 402802 41938
rect 422162 41702 422398 41938
rect 441390 41702 441626 41938
rect 463654 41702 463890 41938
rect 365398 41022 365634 41258
<< metal5 >>
rect 78440 1018512 90960 1031002
rect 129840 1018512 142360 1031002
rect 181240 1018512 193760 1031002
rect 232640 1018512 245160 1031002
rect 284240 1018512 296760 1031002
rect 334810 1018624 346978 1030789
rect 386040 1018512 398560 1031002
rect 475040 1018512 487560 1031002
rect 526440 1018512 538960 1031002
rect 577010 1018624 589178 1030789
rect 628240 1018512 640760 1031002
rect 172340 997338 245892 997380
rect 172340 997102 172382 997338
rect 172618 997102 245614 997338
rect 245850 997102 245892 997338
rect 172340 997060 245892 997102
rect 536660 993258 572860 993300
rect 536660 993022 536702 993258
rect 536938 993022 572582 993258
rect 572818 993022 572860 993258
rect 536660 992980 572860 993022
rect 6598 956440 19088 968960
rect 698512 952840 711002 965360
rect 6167 914054 19620 924934
rect 697980 909666 711433 920546
rect 6811 871210 18976 883378
rect 698512 863640 711002 876160
rect 6811 829010 18976 841178
rect 698624 819822 710789 831990
rect 6598 786640 19088 799160
rect 698512 774440 711002 786960
rect 6598 743440 19088 755960
rect 698512 729440 711002 741960
rect 6598 700240 19088 712760
rect 698512 684440 711002 696960
rect 6598 657040 19088 669560
rect 698512 639240 711002 651760
rect 6598 613840 19088 626360
rect 698512 594240 711002 606760
rect 6598 570640 19088 583160
rect 698512 549040 711002 561560
rect 6598 527440 19088 539960
rect 698624 505222 710789 517390
rect 6811 484410 18976 496578
rect 697980 461866 711433 472746
rect 6167 442854 19620 453734
rect 698624 417022 710789 429190
rect 6598 399840 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 698512 326640 711002 339160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 6598 227040 19088 239560
rect 698512 236640 711002 249160
rect 562972 219418 572676 219460
rect 562972 219182 563014 219418
rect 563250 219182 572398 219418
rect 572634 219182 572676 219418
rect 562972 219140 572676 219182
rect 505012 218738 576724 218780
rect 505012 218502 505054 218738
rect 505290 218502 576446 218738
rect 576682 218502 576724 218738
rect 505012 218460 576724 218502
rect 493788 218058 578380 218100
rect 493788 217822 493830 218058
rect 494066 217822 578102 218058
rect 578338 217822 578380 218058
rect 493788 217780 578380 217822
rect 6598 183840 19088 196360
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 6811 111610 18976 123778
rect 698512 101240 711002 113760
rect 647060 94298 647748 94340
rect 647060 94062 647102 94298
rect 647338 94062 647748 94298
rect 647060 94020 647748 94062
rect 647428 93660 647748 94020
rect 647428 93618 650508 93660
rect 647428 93382 650230 93618
rect 650466 93382 650508 93618
rect 647428 93340 650508 93382
rect 6167 70054 19620 80934
rect 361860 41938 402844 41980
rect 361860 41702 361902 41938
rect 362138 41702 402566 41938
rect 402802 41702 402844 41938
rect 361860 41660 402844 41702
rect 403444 41660 412044 41980
rect 403444 41300 403764 41660
rect 365356 41258 403764 41300
rect 365356 41022 365398 41258
rect 365634 41022 403764 41258
rect 365356 40980 403764 41022
rect 411724 41300 412044 41660
rect 412460 41660 421796 41980
rect 422120 41938 441668 41980
rect 422120 41702 422162 41938
rect 422398 41702 441390 41938
rect 441626 41702 441668 41938
rect 422120 41660 441668 41702
rect 442084 41660 450684 41980
rect 412460 41300 412780 41660
rect 411724 40980 412780 41300
rect 421476 41300 421796 41660
rect 442084 41300 442404 41660
rect 421476 40980 442404 41300
rect 450364 41300 450684 41660
rect 451100 41660 461080 41980
rect 451100 41300 451420 41660
rect 450364 40980 451420 41300
rect 460760 41300 461080 41660
rect 461404 41938 463932 41980
rect 461404 41702 463654 41938
rect 463890 41702 463932 41938
rect 461404 41660 463932 41702
rect 461404 41300 461724 41660
rect 460760 40980 461724 41300
rect 80222 6811 92390 18976
rect 136713 7143 144150 18309
rect 187640 6598 200160 19088
rect 243266 6167 254146 19620
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 570422 6811 582590 18976
rect 624222 6811 636390 18976
use caravel_logo  caravel_logo
timestamp 0
transform 1 0 269370 0 1 5100
box 0 0 1 1
use caravel_motto  caravel_motto
timestamp 0
transform 1 0 -54372 0 1 -4446
box 0 0 1 1
use copyright_block  copyright_block
timestamp 0
transform 1 0 149582 0 1 16298
box 0 0 1 1
use open_source  open_source
timestamp 0
transform 1 0 206098 0 1 2054
box 0 0 1 1
use xres_buf  rstb_level
timestamp 1668092855
transform -1 0 145710 0 -1 50488
box 414 -400 3522 3800
use user_id_textblock  user_id_textblock
timestamp 0
transform 1 0 96272 0 1 6890
box 0 0 1 1
use caravel_clocking  clock_ctrl
timestamp 1668092855
transform 1 0 626764 0 1 55284
box 136 496 20000 20000
use buff_flash_clkrst  flash_clkrst_buffers
timestamp 1668092855
transform 1 0 458400 0 1 47600
box 330 0 7699 5000
use gpio_control_block  gpio_control_bidir_1\[0\]
timestamp 1668092855
transform -1 0 710203 0 1 121000
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_0
timestamp 1668092855
transform -1 0 709467 0 1 134000
box -38 0 6018 2224
use housekeeping  housekeeping
timestamp 1668092855
transform 1 0 592434 0 1 100002
box 0 0 74046 110190
use digital_pll  pll
timestamp 1668092855
transform 1 0 628146 0 1 80944
box 0 0 20000 15000
use simple_por  por
timestamp 1668092855
transform 1 0 650146 0 -1 55282
box -14 11 11344 8684
use user_id_programming  user_id_value
timestamp 1668092855
transform 1 0 656624 0 1 88126
box 0 0 7109 7077
use mgmt_core_wrapper  soc
timestamp 1668092855
transform 1 0 52034 0 1 53002
box -156 0 524096 164000
use gpio_control_block  gpio_control_bidir_1\[1\]
timestamp 1668092855
transform -1 0 710203 0 1 166200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_1
timestamp 1668092855
transform -1 0 709467 0 1 179200
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_2\[2\]
timestamp 1668092855
transform 1 0 7631 0 1 202600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[0\]
timestamp 1668092855
transform -1 0 710203 0 1 211200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_2
timestamp 1668092855
transform -1 0 709467 0 1 224200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_37
timestamp 1668092855
transform 1 0 8367 0 1 215600
box -38 0 6018 2224
use spare_logic_block  spare_logic\[2\]
timestamp 1668092855
transform 1 0 640874 0 1 220592
box 0 0 9000 9000
use gpio_control_block  gpio_control_bidir_2\[1\]
timestamp 1668092855
transform 1 0 7631 0 1 245800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[1\]
timestamp 1668092855
transform -1 0 710203 0 1 256400
box 872 416 34000 13000
use mgmt_protect  mgmt_buffers
timestamp 1668092855
transform 1 0 128180 0 1 232036
box 1066 -400 424400 32400
use spare_logic_block  spare_logic\[0\]
timestamp 1668092855
transform 1 0 88632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[1\]
timestamp 1668092855
transform 1 0 108632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[3\]
timestamp 1668092855
transform 1 0 578632 0 1 232528
box 0 0 9000 9000
use gpio_control_block  gpio_control_bidir_2\[0\]
timestamp 1668092855
transform 1 0 7631 0 1 289000
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_3
timestamp 1668092855
transform -1 0 709467 0 1 269400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_36
timestamp 1668092855
transform 1 0 8367 0 1 258800
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[2\]
timestamp 1668092855
transform -1 0 710203 0 1 301400
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_35
timestamp 1668092855
transform 1 0 8367 0 1 302000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_4
timestamp 1668092855
transform -1 0 709467 0 1 314400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[13\]
timestamp 1668092855
transform 1 0 7631 0 1 418600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[14\]
timestamp 1668092855
transform 1 0 7631 0 1 375400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[15\]
timestamp 1668092855
transform 1 0 7631 0 1 332200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_32
timestamp 1668092855
transform 1 0 8367 0 1 431600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_33
timestamp 1668092855
transform 1 0 8367 0 1 388400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_34
timestamp 1668092855
transform 1 0 8367 0 1 345200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[3\]
timestamp 1668092855
transform -1 0 710203 0 1 346400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[4\]
timestamp 1668092855
transform -1 0 710203 0 1 391600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[5\]
timestamp 1668092855
transform -1 0 710203 0 1 479800
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_5
timestamp 1668092855
transform -1 0 709467 0 1 359400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_6
timestamp 1668092855
transform -1 0 709467 0 1 404600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_7
timestamp 1668092855
transform -1 0 709467 0 1 492800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_31
timestamp 1668092855
transform 1 0 8367 0 1 559200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_30
timestamp 1668092855
transform 1 0 8367 0 1 602400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[12\]
timestamp 1668092855
transform 1 0 7631 0 1 546200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[11\]
timestamp 1668092855
transform 1 0 7631 0 1 589400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[1\]
timestamp 1668092855
transform -1 0 710203 0 1 568800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[0\]
timestamp 1668092855
transform -1 0 710203 0 1 523800
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_9
timestamp 1668092855
transform -1 0 709467 0 1 581800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_8
timestamp 1668092855
transform -1 0 709467 0 1 536800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_29
timestamp 1668092855
transform 1 0 8367 0 1 645600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_28
timestamp 1668092855
transform 1 0 8367 0 1 688800
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[9\]
timestamp 1668092855
transform 1 0 7631 0 1 675800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[10\]
timestamp 1668092855
transform 1 0 7631 0 1 632600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[3\]
timestamp 1668092855
transform -1 0 710203 0 1 659000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[2\]
timestamp 1668092855
transform -1 0 710203 0 1 614000
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_11
timestamp 1668092855
transform -1 0 709467 0 1 672000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_10
timestamp 1668092855
transform -1 0 709467 0 1 627000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_27
timestamp 1668092855
transform 1 0 8367 0 1 732000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_26
timestamp 1668092855
transform 1 0 8367 0 1 775200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[8\]
timestamp 1668092855
transform 1 0 7631 0 1 719000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[7\]
timestamp 1668092855
transform 1 0 7631 0 1 762200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[5\]
timestamp 1668092855
transform -1 0 710203 0 1 749200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[4\]
timestamp 1668092855
transform -1 0 710203 0 1 704200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_13
timestamp 1668092855
transform -1 0 709467 0 1 762200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_12
timestamp 1668092855
transform -1 0 709467 0 1 717200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_25
timestamp 1668092855
transform 1 0 8367 0 1 818400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[6\]
timestamp 1668092855
transform 1 0 7631 0 1 805400
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_24
timestamp 1668092855
transform 1 0 8367 0 1 944200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[5\]
timestamp 1668092855
transform 1 0 7631 0 1 931200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[6\]
timestamp 1668092855
transform -1 0 710203 0 1 927600
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_14
timestamp 1668092855
transform -1 0 709467 0 1 940600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_23
timestamp 1668092855
transform 0 1 110194 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[4\]
timestamp 1668092855
transform 0 1 97200 -1 0 1030077
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_22
timestamp 1668092855
transform 0 1 161594 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_21
timestamp 1668092855
transform 0 1 212994 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[3\]
timestamp 1668092855
transform 0 1 148600 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[2\]
timestamp 1668092855
transform 0 1 200000 -1 0 1030077
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_20
timestamp 1668092855
transform 0 1 264394 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[1\]
timestamp 1668092855
transform 0 1 251400 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[0\]
timestamp 1668092855
transform 0 1 303000 -1 0 1030077
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_19
timestamp 1668092855
transform 0 1 315994 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_18
timestamp 1668092855
transform 0 1 366394 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[10\]
timestamp 1668092855
transform 0 1 353400 -1 0 1030077
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_17
timestamp 1668092855
transform 0 1 433794 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[9\]
timestamp 1668092855
transform 0 1 420800 -1 0 1030077
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_16
timestamp 1668092855
transform 0 1 510794 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_15
timestamp 1668092855
transform 0 1 562194 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[8\]
timestamp 1668092855
transform 0 1 497800 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[7\]
timestamp 1668092855
transform 0 1 549200 -1 0 1030077
box 872 416 34000 13000
use caravel_power_routing  caravel_power_routing
timestamp 1668092855
transform 1 0 0 0 1 0
box 6022 30806 711814 1031696
use user_project_wrapper  mprj
timestamp 1668092855
transform 1 0 65308 0 1 278718
box -8726 -7654 592650 711590
use chip_io  padframe
timestamp 1668092855
transform 1 0 0 0 1 0
box 0 0 717600 1037600
use gpio_signal_buffering  sigbuf
timestamp 1668092855
transform 1 0 0 0 1 0
box 39992 41960 677583 997915
<< labels >>
rlabel metal5 s 187640 6598 200160 19088 6 clock
port 0 nsew signal input
rlabel metal5 s 351040 6598 363560 19088 6 flash_clk
port 1 nsew signal tristate
rlabel metal5 s 296240 6598 308760 19088 6 flash_csb
port 2 nsew signal tristate
rlabel metal5 s 405840 6598 418360 19088 6 flash_io0
port 3 nsew signal tristate
rlabel metal5 s 460640 6598 473160 19088 6 flash_io1
port 4 nsew signal tristate
rlabel metal5 s 515440 6598 527960 19088 6 gpio
port 5 nsew signal bidirectional
rlabel metal5 s 698512 101240 711002 113760 6 mprj_io[0]
port 6 nsew signal bidirectional
rlabel metal5 s 698512 684440 711002 696960 6 mprj_io[10]
port 7 nsew signal bidirectional
rlabel metal5 s 698512 729440 711002 741960 6 mprj_io[11]
port 8 nsew signal bidirectional
rlabel metal5 s 698512 774440 711002 786960 6 mprj_io[12]
port 9 nsew signal bidirectional
rlabel metal5 s 698512 863640 711002 876160 6 mprj_io[13]
port 10 nsew signal bidirectional
rlabel metal5 s 698512 952840 711002 965360 6 mprj_io[14]
port 11 nsew signal bidirectional
rlabel metal5 s 628240 1018512 640760 1031002 6 mprj_io[15]
port 12 nsew signal bidirectional
rlabel metal5 s 526440 1018512 538960 1031002 6 mprj_io[16]
port 13 nsew signal bidirectional
rlabel metal5 s 475040 1018512 487560 1031002 6 mprj_io[17]
port 14 nsew signal bidirectional
rlabel metal5 s 386040 1018512 398560 1031002 6 mprj_io[18]
port 15 nsew signal bidirectional
rlabel metal5 s 284240 1018512 296760 1031002 6 mprj_io[19]
port 16 nsew signal bidirectional
rlabel metal5 s 698512 146440 711002 158960 6 mprj_io[1]
port 17 nsew signal bidirectional
rlabel metal5 s 232640 1018512 245160 1031002 6 mprj_io[20]
port 18 nsew signal bidirectional
rlabel metal5 s 181240 1018512 193760 1031002 6 mprj_io[21]
port 19 nsew signal bidirectional
rlabel metal5 s 129840 1018512 142360 1031002 6 mprj_io[22]
port 20 nsew signal bidirectional
rlabel metal5 s 78440 1018512 90960 1031002 6 mprj_io[23]
port 21 nsew signal bidirectional
rlabel metal5 s 6598 956440 19088 968960 6 mprj_io[24]
port 22 nsew signal bidirectional
rlabel metal5 s 6598 786640 19088 799160 6 mprj_io[25]
port 23 nsew signal bidirectional
rlabel metal5 s 6598 743440 19088 755960 6 mprj_io[26]
port 24 nsew signal bidirectional
rlabel metal5 s 6598 700240 19088 712760 6 mprj_io[27]
port 25 nsew signal bidirectional
rlabel metal5 s 6598 657040 19088 669560 6 mprj_io[28]
port 26 nsew signal bidirectional
rlabel metal5 s 6598 613840 19088 626360 6 mprj_io[29]
port 27 nsew signal bidirectional
rlabel metal5 s 698512 191440 711002 203960 6 mprj_io[2]
port 28 nsew signal bidirectional
rlabel metal5 s 6598 570640 19088 583160 6 mprj_io[30]
port 29 nsew signal bidirectional
rlabel metal5 s 6598 527440 19088 539960 6 mprj_io[31]
port 30 nsew signal bidirectional
rlabel metal5 s 6598 399840 19088 412360 6 mprj_io[32]
port 31 nsew signal bidirectional
rlabel metal5 s 6598 356640 19088 369160 6 mprj_io[33]
port 32 nsew signal bidirectional
rlabel metal5 s 6598 313440 19088 325960 6 mprj_io[34]
port 33 nsew signal bidirectional
rlabel metal5 s 6598 270240 19088 282760 6 mprj_io[35]
port 34 nsew signal bidirectional
rlabel metal5 s 6598 227040 19088 239560 6 mprj_io[36]
port 35 nsew signal bidirectional
rlabel metal5 s 6598 183840 19088 196360 6 mprj_io[37]
port 36 nsew signal bidirectional
rlabel metal5 s 698512 236640 711002 249160 6 mprj_io[3]
port 37 nsew signal bidirectional
rlabel metal5 s 698512 281640 711002 294160 6 mprj_io[4]
port 38 nsew signal bidirectional
rlabel metal5 s 698512 326640 711002 339160 6 mprj_io[5]
port 39 nsew signal bidirectional
rlabel metal5 s 698512 371840 711002 384360 6 mprj_io[6]
port 40 nsew signal bidirectional
rlabel metal5 s 698512 549040 711002 561560 6 mprj_io[7]
port 41 nsew signal bidirectional
rlabel metal5 s 698512 594240 711002 606760 6 mprj_io[8]
port 42 nsew signal bidirectional
rlabel metal5 s 698512 639240 711002 651760 6 mprj_io[9]
port 43 nsew signal bidirectional
rlabel metal5 s 136713 7143 144150 18309 6 resetb
port 44 nsew signal input
rlabel metal5 s 6167 70054 19620 80934 6 vccd
port 45 nsew signal bidirectional
rlabel metal5 s 697980 909666 711433 920546 6 vccd1
port 46 nsew signal bidirectional
rlabel metal5 s 6167 914054 19620 924934 6 vccd2
port 47 nsew signal bidirectional
rlabel metal5 s 624222 6811 636390 18976 6 vdda
port 48 nsew signal bidirectional
rlabel metal5 s 698624 819822 710789 831990 6 vdda1
port 49 nsew signal bidirectional
rlabel metal5 s 698624 505222 710789 517390 6 vdda1_2
port 50 nsew signal bidirectional
rlabel metal5 s 6811 484410 18976 496578 6 vdda2
port 51 nsew signal bidirectional
rlabel metal5 s 6811 111610 18976 123778 6 vddio
port 52 nsew signal bidirectional
rlabel metal5 s 6811 871210 18976 883378 6 vddio_2
port 53 nsew signal bidirectional
rlabel metal5 s 80222 6811 92390 18976 6 vssa
port 54 nsew signal bidirectional
rlabel metal5 s 577010 1018624 589178 1030789 6 vssa1
port 55 nsew signal bidirectional
rlabel metal5 s 698624 417022 710789 429190 6 vssa1_2
port 56 nsew signal bidirectional
rlabel metal5 s 6811 829010 18976 841178 6 vssa2
port 57 nsew signal bidirectional
rlabel metal5 s 243266 6167 254146 19620 6 vssd
port 58 nsew signal bidirectional
rlabel metal5 s 697980 461866 711433 472746 6 vssd1
port 59 nsew signal bidirectional
rlabel metal5 s 6167 442854 19620 453734 6 vssd2
port 60 nsew signal bidirectional
rlabel metal5 s 570422 6811 582590 18976 6 vssio
port 61 nsew signal bidirectional
rlabel metal5 s 334810 1018624 346978 1030789 6 vssio_2
port 62 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
