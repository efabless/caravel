* NGSPICE file created from gpio_logic_high.ext - technology: sky130A

.subckt sky130_fd_sc_hd__decap_6 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.97e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.97e+06u
.ends

.subckt sky130_fd_sc_hd__decap_8 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=2.89e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=2.89e+06u
.ends

.subckt sky130_fd_sc_hd__decap_3 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=590000u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=590000u
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=870000u l=1.05e+06u
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=550000u l=1.05e+06u
.ends

.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
R0 HI VPWR sky130_fd_pr__res_generic_po w=480000u l=45000u
R1 VGND LO sky130_fd_pr__res_generic_po w=480000u l=45000u
.ends

.subckt gpio_logic_high gpio_logic1 vccd1 vssd1
XFILLER_3_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_0 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_7 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_8 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_9 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
Xgpio_logic_high vssd1 vssd1 vccd1 vccd1 gpio_logic1 gpio_logic_high/LO sky130_fd_sc_hd__conb_1
XFILLER_4_9 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_9 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9 vssd1 vccd1 vssd1 vccd1 sky130_fd_sc_hd__decap_3
.ends

