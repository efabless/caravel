* NGSPICE file created from housekeeping.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtn_1 abstract view
.subckt sky130_fd_sc_hd__dfrtn_1 CLK_N D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_1 abstract view
.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_1 abstract view
.subckt sky130_fd_sc_hd__o32ai_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

.subckt housekeeping VGND VPWR debug_in debug_mode debug_oeb debug_out irq[0] irq[1]
+ irq[2] mask_rev_in[0] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13]
+ mask_rev_in[14] mask_rev_in[15] mask_rev_in[16] mask_rev_in[17] mask_rev_in[18]
+ mask_rev_in[19] mask_rev_in[1] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23]
+ mask_rev_in[24] mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28]
+ mask_rev_in[29] mask_rev_in[2] mask_rev_in[30] mask_rev_in[31] mask_rev_in[3] mask_rev_in[4]
+ mask_rev_in[5] mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9] mgmt_gpio_in[0]
+ mgmt_gpio_in[10] mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14]
+ mgmt_gpio_in[15] mgmt_gpio_in[16] mgmt_gpio_in[17] mgmt_gpio_in[18] mgmt_gpio_in[19]
+ mgmt_gpio_in[1] mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23]
+ mgmt_gpio_in[24] mgmt_gpio_in[25] mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28]
+ mgmt_gpio_in[29] mgmt_gpio_in[2] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32]
+ mgmt_gpio_in[33] mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37]
+ mgmt_gpio_in[3] mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7]
+ mgmt_gpio_in[8] mgmt_gpio_in[9] mgmt_gpio_oeb[0] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11]
+ mgmt_gpio_oeb[12] mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16]
+ mgmt_gpio_oeb[17] mgmt_gpio_oeb[18] mgmt_gpio_oeb[19] mgmt_gpio_oeb[1] mgmt_gpio_oeb[20]
+ mgmt_gpio_oeb[21] mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25]
+ mgmt_gpio_oeb[26] mgmt_gpio_oeb[27] mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[2]
+ mgmt_gpio_oeb[30] mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34]
+ mgmt_gpio_oeb[35] mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_oeb[3] mgmt_gpio_oeb[4]
+ mgmt_gpio_oeb[5] mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9]
+ mgmt_gpio_out[0] mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13]
+ mgmt_gpio_out[14] mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18]
+ mgmt_gpio_out[19] mgmt_gpio_out[1] mgmt_gpio_out[20] mgmt_gpio_out[21] mgmt_gpio_out[22]
+ mgmt_gpio_out[23] mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27]
+ mgmt_gpio_out[28] mgmt_gpio_out[29] mgmt_gpio_out[2] mgmt_gpio_out[30] mgmt_gpio_out[31]
+ mgmt_gpio_out[32] mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36]
+ mgmt_gpio_out[37] mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5] mgmt_gpio_out[6]
+ mgmt_gpio_out[7] mgmt_gpio_out[8] mgmt_gpio_out[9] pad_flash_clk pad_flash_clk_oeb
+ pad_flash_csb pad_flash_csb_oeb pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ieb
+ pad_flash_io0_oeb pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ieb pad_flash_io1_oeb
+ pll90_sel[0] pll90_sel[1] pll90_sel[2] pll_bypass pll_dco_ena pll_div[0] pll_div[1]
+ pll_div[2] pll_div[3] pll_div[4] pll_ena pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0]
+ pll_trim[10] pll_trim[11] pll_trim[12] pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16]
+ pll_trim[17] pll_trim[18] pll_trim[19] pll_trim[1] pll_trim[20] pll_trim[21] pll_trim[22]
+ pll_trim[23] pll_trim[24] pll_trim[25] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5]
+ pll_trim[6] pll_trim[7] pll_trim[8] pll_trim[9] porb pwr_ctrl_out[0] pwr_ctrl_out[1]
+ pwr_ctrl_out[2] pwr_ctrl_out[3] qspi_enabled reset ser_rx ser_tx serial_clock serial_data_1
+ serial_data_2 serial_load serial_resetn spi_csb spi_enabled spi_sck spi_sdi spi_sdo
+ spi_sdoenb spimemio_flash_clk spimemio_flash_csb spimemio_flash_io0_di spimemio_flash_io0_do
+ spimemio_flash_io0_oeb spimemio_flash_io1_di spimemio_flash_io1_do spimemio_flash_io1_oeb
+ spimemio_flash_io2_di spimemio_flash_io2_do spimemio_flash_io2_oeb spimemio_flash_io3_di
+ spimemio_flash_io3_do spimemio_flash_io3_oeb trap uart_enabled user_clock usr1_vcc_pwrgood
+ usr1_vdd_pwrgood usr2_vcc_pwrgood usr2_vdd_pwrgood wb_ack_o wb_adr_i[0] wb_adr_i[10]
+ wb_adr_i[11] wb_adr_i[12] wb_adr_i[13] wb_adr_i[14] wb_adr_i[15] wb_adr_i[16] wb_adr_i[17]
+ wb_adr_i[18] wb_adr_i[19] wb_adr_i[1] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22] wb_adr_i[23]
+ wb_adr_i[24] wb_adr_i[25] wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[2]
+ wb_adr_i[30] wb_adr_i[31] wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6] wb_adr_i[7]
+ wb_adr_i[8] wb_adr_i[9] wb_clk_i wb_cyc_i wb_dat_i[0] wb_dat_i[10] wb_dat_i[11]
+ wb_dat_i[12] wb_dat_i[13] wb_dat_i[14] wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18]
+ wb_dat_i[19] wb_dat_i[1] wb_dat_i[20] wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24]
+ wb_dat_i[25] wb_dat_i[26] wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[2] wb_dat_i[30]
+ wb_dat_i[31] wb_dat_i[3] wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7] wb_dat_i[8]
+ wb_dat_i[9] wb_dat_o[0] wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14]
+ wb_dat_o[15] wb_dat_o[16] wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[1] wb_dat_o[20]
+ wb_dat_o[21] wb_dat_o[22] wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27]
+ wb_dat_o[28] wb_dat_o[29] wb_dat_o[2] wb_dat_o[30] wb_dat_o[31] wb_dat_o[3] wb_dat_o[4]
+ wb_dat_o[5] wb_dat_o[6] wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_rstn_i wb_sel_i[0]
+ wb_sel_i[1] wb_sel_i[2] wb_sel_i[3] wb_stb_i wb_we_i
XFILLER_39_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6914_ clknet_leaf_15_csclk net1790 net513 VGND VGND VPWR VPWR gpio_configure\[9\]\[0\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6845_ clknet_leaf_65_csclk net739 net505 VGND VGND VPWR VPWR gpio_configure\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6776_ clknet_3_7_0_wb_clk_i _0379_ net528 VGND VGND VPWR VPWR wbbd_addr\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_168_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3988_ net1019 net443 _1470_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__mux2_1
XFILLER_148_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5727_ gpio_configure\[22\]\[1\] _2498_ _2513_ gpio_configure\[28\]\[1\] _2560_ VGND
+ VGND VPWR VPWR _2561_ sky130_fd_sc_hd__a221o_1
XFILLER_109_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5658_ pad_count_1\[3\] pad_count_1\[2\] VGND VGND VPWR VPWR _2493_ sky130_fd_sc_hd__and2_2
X_4609_ _1750_ _1769_ _1772_ VGND VGND VPWR VPWR _1821_ sky130_fd_sc_hd__nor3_2
XFILLER_190_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5589_ xfer_state\[0\] _0823_ serial_busy VGND VGND VPWR VPWR _2442_ sky130_fd_sc_hd__a21o_1
XFILLER_151_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold340 _0510_ VGND VGND VPWR VPWR net873 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold351 gpio_configure\[5\]\[1\] VGND VGND VPWR VPWR net884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 _0251_ VGND VGND VPWR VPWR net895 sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 gpio_configure\[34\]\[1\] VGND VGND VPWR VPWR net906 sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 _0312_ VGND VGND VPWR VPWR net917 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold395 gpio_configure\[28\]\[7\] VGND VGND VPWR VPWR net928 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1040 _0172_ VGND VGND VPWR VPWR net1573 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1051 gpio_configure\[7\]\[0\] VGND VGND VPWR VPWR net1584 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1062 _0329_ VGND VGND VPWR VPWR net1595 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1073 gpio_configure\[11\]\[0\] VGND VGND VPWR VPWR net1606 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1084 _0461_ VGND VGND VPWR VPWR net1617 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_202 _2497_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1095 _0738_ VGND VGND VPWR VPWR net1628 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_213 serial_data_staging_1\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_224 net373 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_235 net463 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_246 _2512_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_257 net471 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4960_ _2156_ _2164_ _2169_ VGND VGND VPWR VPWR _2170_ sky130_fd_sc_hd__or3b_1
XFILLER_17_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3911_ _0818_ net431 _0820_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__o21ai_1
X_4891_ _1652_ _2082_ _2091_ _2101_ VGND VGND VPWR VPWR _2102_ sky130_fd_sc_hd__a211o_1
XFILLER_149_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6630_ clknet_3_4_0_wb_clk_i _0243_ VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__dfxtp_1
X_3842_ hkspi.readmode _1378_ hkspi.rdstb VGND VGND VPWR VPWR _1412_ sky130_fd_sc_hd__a21oi_1
XFILLER_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6561_ clknet_leaf_57_csclk net1507 net504 VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__dfrtp_4
X_3773_ gpio_configure\[28\]\[0\] _0888_ _1086_ gpio_configure\[29\]\[8\] VGND VGND
+ VPWR VPWR _1359_ sky130_fd_sc_hd__a22o_1
XFILLER_192_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5512_ net469 net1598 _2433_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__mux2_1
X_6492_ clknet_leaf_73_csclk net1990 net488 VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__dfstp_1
XFILLER_172_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5443_ net452 net962 _2425_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__mux2_1
XFILLER_105_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5374_ net439 net852 _2417_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__mux2_1
X_7113_ clknet_leaf_26_csclk net1733 net519 VGND VGND VPWR VPWR gpio_configure\[34\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_4325_ net1816 net467 _1546_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__mux2_1
XFILLER_114_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7044_ clknet_leaf_64_csclk net843 net501 VGND VGND VPWR VPWR gpio_configure\[25\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_4256_ net916 net450 _1534_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__mux2_1
XFILLER_113_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3207_ gpio_configure\[27\]\[3\] VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__inv_2
XFILLER_74_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4187_ net2013 _1004_ _1519_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__mux2_1
XFILLER_27_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6828_ clknet_leaf_29_csclk net1615 net520 VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__dfrtp_1
XFILLER_50_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6759_ clknet_leaf_73_csclk net1036 net489 VGND VGND VPWR VPWR gpio_configure\[33\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_109_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold170 _0232_ VGND VGND VPWR VPWR net703 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold181 gpio_configure\[5\]\[11\] VGND VGND VPWR VPWR net714 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 _0416_ VGND VGND VPWR VPWR net725 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_120_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4110_ net660 net706 _1508_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__mux2_1
X_5090_ _2011_ _2194_ _2298_ VGND VGND VPWR VPWR _2299_ sky130_fd_sc_hd__or3b_1
X_4041_ net468 net1785 _1478_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__mux2_1
XFILLER_56_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5992_ _2469_ _2796_ _2809_ VGND VGND VPWR VPWR _2814_ sky130_fd_sc_hd__and3_4
XFILLER_24_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4943_ _1607_ _2152_ _2044_ VGND VGND VPWR VPWR _2153_ sky130_fd_sc_hd__a21o_1
XFILLER_17_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4874_ _1622_ _1642_ _1937_ VGND VGND VPWR VPWR _2085_ sky130_fd_sc_hd__and3_1
XFILLER_177_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6613_ clknet_leaf_3_csclk net1341 net493 VGND VGND VPWR VPWR gpio_configure\[3\]\[10\]
+ sky130_fd_sc_hd__dfrtp_4
X_3825_ _1402_ net2085 _1388_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__mux2_1
XFILLER_193_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6544_ clknet_2_1__leaf_mgmt_gpio_in[4] _0007_ _0055_ VGND VGND VPWR VPWR hkspi.state\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_158_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3756_ gpio_configure\[33\]\[0\] _0938_ _1007_ net61 _1325_ VGND VGND VPWR VPWR _1342_
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_5_0_csclk clknet_2_2_0_csclk VGND VGND VPWR VPWR clknet_3_5_0_csclk sky130_fd_sc_hd__clkbuf_8
XFILLER_145_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6475_ clknet_leaf_72_csclk net1719 net490 VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__dfstp_1
XFILLER_145_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3687_ gpio_configure\[19\]\[1\] _0896_ _1073_ gpio_configure\[24\]\[9\] _1274_ VGND
+ VGND VPWR VPWR _1275_ sky130_fd_sc_hd__a221o_1
XFILLER_106_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5426_ net445 net720 _2423_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__mux2_1
XFILLER_118_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput220 net220 VGND VGND VPWR VPWR mgmt_gpio_out[16] sky130_fd_sc_hd__buf_12
Xoutput231 net231 VGND VGND VPWR VPWR mgmt_gpio_out[26] sky130_fd_sc_hd__buf_12
Xoutput242 net242 VGND VGND VPWR VPWR mgmt_gpio_out[36] sky130_fd_sc_hd__buf_12
Xoutput253 net253 VGND VGND VPWR VPWR pad_flash_csb sky130_fd_sc_hd__buf_12
XFILLER_133_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput264 net264 VGND VGND VPWR VPWR pll_bypass sky130_fd_sc_hd__buf_12
X_5357_ net434 net1037 _2415_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__mux2_1
XFILLER_99_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput275 net275 VGND VGND VPWR VPWR pll_trim[0] sky130_fd_sc_hd__buf_12
XFILLER_87_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput286 net286 VGND VGND VPWR VPWR pll_trim[1] sky130_fd_sc_hd__buf_12
Xoutput297 net297 VGND VGND VPWR VPWR pll_trim[6] sky130_fd_sc_hd__buf_12
X_4308_ net462 net1481 _1543_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__mux2_1
XFILLER_99_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5288_ net542 net1922 net565 VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__mux2_1
XFILLER_59_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7027_ clknet_leaf_22_csclk net875 net515 VGND VGND VPWR VPWR gpio_configure\[23\]\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_4239_ net446 net910 net592 VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__mux2_1
XFILLER_28_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_199 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout491 net527 VGND VGND VPWR VPWR net491 sky130_fd_sc_hd__buf_6
XFILLER_171_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3610_ gpio_configure\[4\]\[10\] _1093_ _1110_ gpio_configure\[2\]\[10\] VGND VGND
+ VPWR VPWR _1199_ sky130_fd_sc_hd__a22o_1
XFILLER_159_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4590_ net424 _1801_ VGND VGND VPWR VPWR _1802_ sky130_fd_sc_hd__nor2_1
X_3541_ _1120_ _1124_ _1128_ _1131_ VGND VGND VPWR VPWR _1132_ sky130_fd_sc_hd__or4_1
XFILLER_190_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold906 net2136 VGND VGND VPWR VPWR net1439 sky130_fd_sc_hd__dlygate4sd3_1
Xhold917 _0102_ VGND VGND VPWR VPWR net1450 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold928 gpio_configure\[1\]\[1\] VGND VGND VPWR VPWR net1461 sky130_fd_sc_hd__dlygate4sd3_1
Xhold939 _0611_ VGND VGND VPWR VPWR net1472 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6260_ gpio_configure\[9\]\[9\] net412 _2838_ gpio_configure\[12\]\[9\] VGND VGND
+ VPWR VPWR _3073_ sky130_fd_sc_hd__a22o_1
X_3472_ net389 _0973_ VGND VGND VPWR VPWR _1063_ sky130_fd_sc_hd__nor2_1
X_5211_ net466 net1767 _2395_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__mux2_1
X_6191_ gpio_configure\[29\]\[6\] _2816_ _2852_ gpio_configure\[19\]\[6\] _3006_ VGND
+ VGND VPWR VPWR _3007_ sky130_fd_sc_hd__a221o_1
XFILLER_170_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5142_ _2175_ _2307_ _2348_ VGND VGND VPWR VPWR _2349_ sky130_fd_sc_hd__or3b_1
XFILLER_111_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1606 wbbd_state\[0\] VGND VGND VPWR VPWR net2139 sky130_fd_sc_hd__dlygate4sd3_1
X_5073_ _1821_ _2230_ _2281_ VGND VGND VPWR VPWR _2282_ sky130_fd_sc_hd__or3b_1
X_4024_ net1674 net461 _1475_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__mux2_1
XFILLER_65_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5975_ pad_count_2\[4\] pad_count_2\[5\] VGND VGND VPWR VPWR _2797_ sky130_fd_sc_hd__or2_4
X_4926_ _1704_ _1933_ VGND VGND VPWR VPWR _2137_ sky130_fd_sc_hd__nand2_1
XFILLER_21_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4857_ _2046_ _2065_ _2066_ _2067_ VGND VGND VPWR VPWR _2068_ sky130_fd_sc_hd__and4_1
XFILLER_165_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3808_ hkspi.addr\[3\] _1389_ VGND VGND VPWR VPWR _1390_ sky130_fd_sc_hd__and2_1
XFILLER_165_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4788_ _1655_ _1745_ net424 _1836_ VGND VGND VPWR VPWR _1999_ sky130_fd_sc_hd__o22ai_1
X_6527_ clknet_leaf_76_csclk net1655 net484 VGND VGND VPWR VPWR gpio_configure\[25\]\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_118_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3739_ gpio_configure\[6\]\[0\] net357 net352 gpio_configure\[36\]\[0\] VGND VGND
+ VPWR VPWR _1325_ sky130_fd_sc_hd__a22o_1
X_6458_ clknet_2_1__leaf_mgmt_gpio_in[4] _0080_ _0036_ VGND VGND VPWR VPWR hkspi.rdstb
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_134_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5409_ net440 net1554 _2421_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__mux2_1
XFILLER_134_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6389_ wbbd_state\[8\] net166 _3179_ VGND VGND VPWR VPWR _3180_ sky130_fd_sc_hd__a21o_1
XFILLER_87_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5760_ gpio_configure\[28\]\[3\] _2513_ _2517_ gpio_configure\[30\]\[3\] _2591_ VGND
+ VGND VPWR VPWR _2592_ sky130_fd_sc_hd__a221o_1
XFILLER_15_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4711_ net477 _1684_ _1685_ _1901_ _1922_ VGND VGND VPWR VPWR _1923_ sky130_fd_sc_hd__o311a_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5691_ _0831_ net419 VGND VGND VPWR VPWR _2526_ sky130_fd_sc_hd__nand2_8
XFILLER_147_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4642_ _1830_ _1846_ _1849_ _1853_ VGND VGND VPWR VPWR _1854_ sky130_fd_sc_hd__and4_1
XFILLER_163_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4573_ _1679_ _1758_ VGND VGND VPWR VPWR _1785_ sky130_fd_sc_hd__nand2b_2
Xmax_cap400 _2806_ VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__buf_8
XFILLER_162_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap411 _2836_ VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__buf_12
Xhold703 gpio_configure\[13\]\[11\] VGND VGND VPWR VPWR net1236 sky130_fd_sc_hd__dlygate4sd3_1
Xhold714 _0368_ VGND VGND VPWR VPWR net1247 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap422 _2496_ VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__buf_8
X_6312_ gpio_configure\[13\]\[11\] net417 _2862_ gpio_configure\[25\]\[11\] VGND VGND
+ VPWR VPWR _3123_ sky130_fd_sc_hd__a22o_1
Xmax_cap433 _1526_ VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__clkbuf_2
X_3524_ _1108_ _1111_ _1112_ _1114_ VGND VGND VPWR VPWR _1115_ sky130_fd_sc_hd__or4_2
Xhold725 net290 VGND VGND VPWR VPWR net1258 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold736 _0593_ VGND VGND VPWR VPWR net1269 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold747 gpio_configure\[28\]\[11\] VGND VGND VPWR VPWR net1280 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold758 _0684_ VGND VGND VPWR VPWR net1291 sky130_fd_sc_hd__dlygate4sd3_1
X_6243_ gpio_configure\[0\]\[8\] _2851_ _3046_ _3056_ net473 VGND VGND VPWR VPWR _3057_
+ sky130_fd_sc_hd__o221a_1
Xhold769 gpio_configure\[7\]\[4\] VGND VGND VPWR VPWR net1302 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3455_ net590 net388 VGND VGND VPWR VPWR _1046_ sky130_fd_sc_hd__nor2_4
XFILLER_115_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6174_ gpio_configure\[7\]\[6\] _2811_ net413 gpio_configure\[3\]\[6\] VGND VGND
+ VPWR VPWR _2990_ sky130_fd_sc_hd__a22o_1
XFILLER_130_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3386_ gpio_configure\[13\]\[6\] _0906_ _0932_ gpio_configure\[35\]\[6\] _0975_ VGND
+ VGND VPWR VPWR _0980_ sky130_fd_sc_hd__a221o_1
XFILLER_57_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5125_ _2273_ _2332_ VGND VGND VPWR VPWR _2333_ sky130_fd_sc_hd__nor2_1
Xhold1403 gpio_configure\[12\]\[10\] VGND VGND VPWR VPWR net1936 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1414 net337 VGND VGND VPWR VPWR net1947 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1425 net320 VGND VGND VPWR VPWR net1958 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1436 net334 VGND VGND VPWR VPWR net1969 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1447 _0541_ VGND VGND VPWR VPWR net1980 sky130_fd_sc_hd__dlygate4sd3_1
X_5056_ _1588_ _1801_ _2158_ _1697_ VGND VGND VPWR VPWR _2265_ sky130_fd_sc_hd__o211a_1
Xhold1458 wbbd_addr\[2\] VGND VGND VPWR VPWR net1991 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1469 _0391_ VGND VGND VPWR VPWR net2002 sky130_fd_sc_hd__dlygate4sd3_1
X_4007_ net440 net1558 _1472_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__mux2_1
XTAP_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_1_0_1_wb_clk_i clknet_1_0_0_wb_clk_i VGND VGND VPWR VPWR clknet_1_0_1_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_80_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5958_ gpio_configure\[17\]\[12\] _2537_ _2541_ gpio_configure\[31\]\[12\] VGND VGND
+ VPWR VPWR _2781_ sky130_fd_sc_hd__a22o_1
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4909_ _2119_ VGND VGND VPWR VPWR _2120_ sky130_fd_sc_hd__inv_2
X_5889_ gpio_configure\[17\]\[9\] _2537_ _2541_ gpio_configure\[31\]\[9\] VGND VGND
+ VPWR VPWR _2715_ sky130_fd_sc_hd__a22o_1
XFILLER_187_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_2_2_0_csclk clknet_1_1_1_csclk VGND VGND VPWR VPWR clknet_2_2_0_csclk sky130_fd_sc_hd__clkbuf_8
XFILLER_181_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold30 _0935_ VGND VGND VPWR VPWR net563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 _0200_ VGND VGND VPWR VPWR net574 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold52 _0290_ VGND VGND VPWR VPWR net585 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold63 _0296_ VGND VGND VPWR VPWR net596 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 _0854_ VGND VGND VPWR VPWR net607 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 net448 VGND VGND VPWR VPWR net618 sky130_fd_sc_hd__buf_6
Xhold96 net379 VGND VGND VPWR VPWR net629 sky130_fd_sc_hd__buf_6
XFILLER_29_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_5 _0908_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3240_ net125 VGND VGND VPWR VPWR _0836_ sky130_fd_sc_hd__clkinv_2
XFILLER_100_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6930_ clknet_leaf_27_csclk net1607 net519 VGND VGND VPWR VPWR gpio_configure\[11\]\[0\]
+ sky130_fd_sc_hd__dfstp_4
XFILLER_35_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6861_ clknet_leaf_50_csclk net695 net507 VGND VGND VPWR VPWR gpio_configure\[2\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_6_csclk clknet_3_1_0_csclk VGND VGND VPWR VPWR clknet_leaf_6_csclk sky130_fd_sc_hd__clkbuf_16
XFILLER_34_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5812_ gpio_configure\[6\]\[5\] _2490_ _2523_ gpio_configure\[2\]\[5\] _2641_ VGND
+ VGND VPWR VPWR _2642_ sky130_fd_sc_hd__a221o_1
X_6792_ clknet_leaf_77_csclk net1593 net484 VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__dfstp_1
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5743_ gpio_configure\[16\]\[2\] _0831_ VGND VGND VPWR VPWR _2576_ sky130_fd_sc_hd__or2_1
XFILLER_148_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5674_ gpio_configure\[11\]\[0\] _2505_ _2508_ VGND VGND VPWR VPWR _2509_ sky130_fd_sc_hd__a21o_1
X_4625_ net432 _1836_ VGND VGND VPWR VPWR _1837_ sky130_fd_sc_hd__nor2_1
XFILLER_148_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold500 gpio_configure\[33\]\[7\] VGND VGND VPWR VPWR net1033 sky130_fd_sc_hd__dlygate4sd3_1
Xhold511 _0460_ VGND VGND VPWR VPWR net1044 sky130_fd_sc_hd__dlygate4sd3_1
X_4556_ _1767_ VGND VGND VPWR VPWR _1768_ sky130_fd_sc_hd__inv_2
Xhold522 gpio_configure\[27\]\[11\] VGND VGND VPWR VPWR net1055 sky130_fd_sc_hd__dlygate4sd3_1
Xhold533 _0490_ VGND VGND VPWR VPWR net1066 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3507_ _0885_ net384 VGND VGND VPWR VPWR _1098_ sky130_fd_sc_hd__nor2_4
Xhold544 gpio_configure\[1\]\[3\] VGND VGND VPWR VPWR net1077 sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 _0500_ VGND VGND VPWR VPWR net1088 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold566 _0409_ VGND VGND VPWR VPWR net1099 sky130_fd_sc_hd__dlygate4sd3_1
X_4487_ _1598_ _1675_ VGND VGND VPWR VPWR _1699_ sky130_fd_sc_hd__nand2_2
Xhold577 gpio_configure\[37\]\[11\] VGND VGND VPWR VPWR net1110 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold588 _0530_ VGND VGND VPWR VPWR net1121 sky130_fd_sc_hd__dlygate4sd3_1
X_6226_ gpio_configure\[29\]\[8\] _2816_ _2820_ gpio_configure\[21\]\[8\] _3037_ VGND
+ VGND VPWR VPWR _3040_ sky130_fd_sc_hd__a221o_1
XFILLER_103_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3438_ gpio_configure\[6\]\[5\] net357 _0888_ gpio_configure\[28\]\[5\] _1017_ VGND
+ VGND VPWR VPWR _1030_ sky130_fd_sc_hd__a221o_1
Xhold599 gpio_configure\[29\]\[5\] VGND VGND VPWR VPWR net1132 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6157_ gpio_configure\[37\]\[5\] net400 net416 gpio_configure\[32\]\[5\] _2964_ VGND
+ VGND VPWR VPWR _2974_ sky130_fd_sc_hd__a221o_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3369_ gpio_configure\[5\]\[7\] _0914_ _0921_ gpio_configure\[12\]\[7\] VGND VGND
+ VPWR VPWR _0965_ sky130_fd_sc_hd__a22o_1
Xhold1200 _0716_ VGND VGND VPWR VPWR net1733 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1211 net266 VGND VGND VPWR VPWR net1744 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5108_ _1805_ _2285_ VGND VGND VPWR VPWR _2316_ sky130_fd_sc_hd__nor2_1
Xhold1222 gpio_configure\[4\]\[8\] VGND VGND VPWR VPWR net1755 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1233 _0557_ VGND VGND VPWR VPWR net1766 sky130_fd_sc_hd__dlygate4sd3_1
X_6088_ gpio_configure\[27\]\[2\] net406 net391 gpio_configure\[17\]\[2\] VGND VGND
+ VPWR VPWR _2908_ sky130_fd_sc_hd__a22o_1
Xhold1244 gpio_configure\[16\]\[0\] VGND VGND VPWR VPWR net1777 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1255 _0234_ VGND VGND VPWR VPWR net1788 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1266 _0685_ VGND VGND VPWR VPWR net1799 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1277 gpio_configure\[30\]\[8\] VGND VGND VPWR VPWR net1810 sky130_fd_sc_hd__dlygate4sd3_1
X_5039_ _1944_ _2210_ _2247_ VGND VGND VPWR VPWR _2248_ sky130_fd_sc_hd__or3b_1
XTAP_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1288 _0096_ VGND VGND VPWR VPWR net1821 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1299 net299 VGND VGND VPWR VPWR net1832 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_578 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput120 wb_adr_i[29] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_1
Xinput131 wb_cyc_i VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_1
XFILLER_163_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput142 wb_dat_i[19] VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_1
Xinput153 wb_dat_i[29] VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_1
Xinput164 wb_rstn_i VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_4
XFILLER_48_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4410_ _1621_ _1619_ VGND VGND VPWR VPWR _1622_ sky130_fd_sc_hd__and2b_1
XFILLER_184_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5390_ net447 net1298 _2419_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__mux2_1
X_4341_ net126 net125 VGND VGND VPWR VPWR _1553_ sky130_fd_sc_hd__and2_2
XFILLER_113_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7060_ clknet_leaf_23_csclk net1351 net515 VGND VGND VPWR VPWR gpio_configure\[27\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_4272_ net830 net465 _1537_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__mux2_1
XFILLER_140_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6011_ gpio_configure\[20\]\[0\] _2828_ _2829_ gpio_configure\[33\]\[0\] _2832_ VGND
+ VGND VPWR VPWR _2833_ sky130_fd_sc_hd__a221o_1
XFILLER_140_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3223_ gpio_configure\[11\]\[3\] VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__inv_2
XFILLER_79_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6913_ clknet_leaf_29_csclk net909 net524 VGND VGND VPWR VPWR gpio_configure\[8\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_35_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6844_ clknet_leaf_50_csclk net751 net505 VGND VGND VPWR VPWR gpio_configure\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6775_ clknet_leaf_70_csclk net1064 net491 VGND VGND VPWR VPWR gpio_configure\[22\]\[12\]
+ sky130_fd_sc_hd__dfrtp_4
X_3987_ net1124 net449 _1470_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__mux2_1
X_5726_ gpio_configure\[13\]\[1\] _2501_ _2523_ gpio_configure\[2\]\[1\] VGND VGND
+ VPWR VPWR _2560_ sky130_fd_sc_hd__a22o_1
XFILLER_109_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5657_ gpio_configure\[6\]\[0\] _2490_ _2491_ gpio_configure\[19\]\[0\] VGND VGND
+ VPWR VPWR _2492_ sky130_fd_sc_hd__a22o_1
XFILLER_136_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4608_ _1752_ _1771_ _1819_ VGND VGND VPWR VPWR _1820_ sky130_fd_sc_hd__a21o_1
XFILLER_184_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5588_ net573 net1908 net603 VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__mux2_1
Xhold330 _0203_ VGND VGND VPWR VPWR net863 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_163_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold341 gpio_configure\[23\]\[1\] VGND VGND VPWR VPWR net874 sky130_fd_sc_hd__dlygate4sd3_1
X_4539_ _1554_ _1749_ VGND VGND VPWR VPWR _1751_ sky130_fd_sc_hd__and2_1
Xhold352 _0486_ VGND VGND VPWR VPWR net885 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold363 gpio_configure\[9\]\[12\] VGND VGND VPWR VPWR net896 sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 _0715_ VGND VGND VPWR VPWR net907 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold385 gpio_configure\[7\]\[11\] VGND VGND VPWR VPWR net918 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold396 _0676_ VGND VGND VPWR VPWR net929 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6209_ gpio_configure\[34\]\[7\] net393 _2852_ gpio_configure\[19\]\[7\] _3023_ VGND
+ VGND VPWR VPWR _3024_ sky130_fd_sc_hd__a221o_1
X_7189_ clknet_3_4_0_wb_clk_i _0791_ VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__dfxtp_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1030 _0714_ VGND VGND VPWR VPWR net1563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1041 gpio_configure\[31\]\[0\] VGND VGND VPWR VPWR net1574 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1052 _0501_ VGND VGND VPWR VPWR net1585 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1063 gpio_configure\[23\]\[0\] VGND VGND VPWR VPWR net1596 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1074 _0533_ VGND VGND VPWR VPWR net1607 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1085 net1986 VGND VGND VPWR VPWR net1618 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_203 _2534_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1096 gpio_configure\[26\]\[10\] VGND VGND VPWR VPWR net1629 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_214 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_225 net392 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_236 net471 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_247 _2520_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_258 clknet_3_6_0_wb_clk_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_71_csclk clknet_3_0_0_csclk VGND VGND VPWR VPWR clknet_leaf_71_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_64_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3910_ _1451_ _1453_ xfer_state\[3\] _1442_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_32_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4890_ _2090_ _2098_ _2099_ _2100_ VGND VGND VPWR VPWR _2101_ sky130_fd_sc_hd__or4_1
X_3841_ net2097 _1380_ hkspi.pass_thru_mgmt VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__a21o_1
XFILLER_60_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3772_ net266 _1117_ _1353_ _1355_ _1357_ VGND VGND VPWR VPWR _1358_ sky130_fd_sc_hd__a2111o_1
X_6560_ clknet_leaf_78_csclk net943 net486 VGND VGND VPWR VPWR mgmt_gpio_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_9_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5511_ _0917_ net427 VGND VGND VPWR VPWR _2433_ sky130_fd_sc_hd__nand2_8
X_6491_ clknet_leaf_73_csclk net1950 net488 VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__dfstp_2
XFILLER_118_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5442_ net457 net778 _2425_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__mux2_1
XFILLER_145_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5373_ net441 net1102 _2417_ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__mux2_1
XFILLER_114_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_24_csclk clknet_3_7_0_csclk VGND VGND VPWR VPWR clknet_leaf_24_csclk
+ sky130_fd_sc_hd__clkbuf_16
X_7112_ clknet_leaf_64_csclk net907 net501 VGND VGND VPWR VPWR gpio_configure\[34\]\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_4324_ _1101_ net427 VGND VGND VPWR VPWR _1546_ sky130_fd_sc_hd__and2_2
XFILLER_160_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7043_ clknet_leaf_21_csclk net1378 net514 VGND VGND VPWR VPWR gpio_configure\[25\]\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_4255_ net1362 net456 _1534_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__mux2_1
X_3206_ gpio_configure\[28\]\[3\] VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__inv_2
X_4186_ net2024 _1039_ _1519_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_39_csclk clknet_3_6_0_csclk VGND VGND VPWR VPWR clknet_leaf_39_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_95_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_1_0_csclk clknet_2_0_0_csclk VGND VGND VPWR VPWR clknet_3_1_0_csclk sky130_fd_sc_hd__clkbuf_8
XFILLER_82_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6827_ clknet_leaf_28_csclk net737 net520 VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__dfrtp_1
XFILLER_50_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6758_ clknet_leaf_72_csclk net1283 net490 VGND VGND VPWR VPWR gpio_configure\[33\]\[10\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_149_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5709_ gpio_configure\[0\]\[0\] _2526_ _2543_ _2516_ _2485_ VGND VGND VPWR VPWR _2544_
+ sky130_fd_sc_hd__o221a_1
XFILLER_148_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6689_ clknet_leaf_5_csclk net1237 net494 VGND VGND VPWR VPWR gpio_configure\[13\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_109_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold160 _0680_ VGND VGND VPWR VPWR net693 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold171 gpio_configure\[36\]\[4\] VGND VGND VPWR VPWR net704 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold182 _0237_ VGND VGND VPWR VPWR net715 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold193 net2128 VGND VGND VPWR VPWR net726 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_120_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4040_ _1046_ net426 VGND VGND VPWR VPWR _1478_ sky130_fd_sc_hd__nand2_2
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5991_ _1447_ _2793_ _2800_ VGND VGND VPWR VPWR _2813_ sky130_fd_sc_hd__and3b_2
XFILLER_91_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4942_ _1663_ _1684_ VGND VGND VPWR VPWR _2152_ sky130_fd_sc_hd__nand2_1
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_735 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4873_ _1708_ _1929_ VGND VGND VPWR VPWR _2084_ sky130_fd_sc_hd__nand2_1
XFILLER_178_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6612_ clknet_leaf_78_csclk net1673 net486 VGND VGND VPWR VPWR gpio_configure\[3\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_3824_ hkspi.addr\[2\] hkspi.state\[3\] _1396_ _1401_ VGND VGND VPWR VPWR _1402_
+ sky130_fd_sc_hd__a22o_1
XFILLER_177_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6543_ clknet_2_1__leaf_mgmt_gpio_in[4] _0006_ _0054_ VGND VGND VPWR VPWR hkspi.state\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_3755_ _1337_ _1338_ _1339_ _1340_ VGND VGND VPWR VPWR _1341_ sky130_fd_sc_hd__or4_1
XFILLER_192_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3686_ gpio_configure\[20\]\[1\] _0928_ _1098_ gpio_configure\[25\]\[9\] VGND VGND
+ VPWR VPWR _1274_ sky130_fd_sc_hd__a22o_1
X_6474_ clknet_leaf_71_csclk net1821 net490 VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__dfstp_1
XFILLER_145_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5425_ net451 net812 _2423_ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__mux2_1
Xoutput210 net210 VGND VGND VPWR VPWR mgmt_gpio_oeb[7] sky130_fd_sc_hd__buf_12
Xoutput221 net221 VGND VGND VPWR VPWR mgmt_gpio_out[17] sky130_fd_sc_hd__buf_12
XFILLER_133_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput232 net232 VGND VGND VPWR VPWR mgmt_gpio_out[27] sky130_fd_sc_hd__buf_12
Xoutput243 net243 VGND VGND VPWR VPWR mgmt_gpio_out[37] sky130_fd_sc_hd__buf_12
Xoutput254 net254 VGND VGND VPWR VPWR pad_flash_csb_oeb sky130_fd_sc_hd__buf_12
X_5356_ net438 net1365 _2415_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__mux2_1
Xoutput265 net265 VGND VGND VPWR VPWR pll_dco_ena sky130_fd_sc_hd__buf_12
Xoutput276 net276 VGND VGND VPWR VPWR pll_trim[10] sky130_fd_sc_hd__buf_12
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput287 net287 VGND VGND VPWR VPWR pll_trim[20] sky130_fd_sc_hd__buf_12
X_4307_ net467 net1493 _1543_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__mux2_1
Xoutput298 net298 VGND VGND VPWR VPWR pll_trim[7] sky130_fd_sc_hd__buf_12
X_5287_ net1098 net1308 net565 VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__mux2_1
XFILLER_102_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7026_ clknet_leaf_63_csclk net1597 net501 VGND VGND VPWR VPWR gpio_configure\[23\]\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_87_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4238_ net569 net1915 net592 VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__mux2_1
XFILLER_28_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4169_ net2014 _1191_ _1517_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__mux2_1
XFILLER_83_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire359 net365 VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__clkbuf_2
XFILLER_136_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout470 net471 VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__buf_6
XFILLER_59_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout481 net482 VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__buf_4
XFILLER_120_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout492 net493 VGND VGND VPWR VPWR net492 sky130_fd_sc_hd__buf_4
XFILLER_65_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3540_ net30 _0900_ net353 net39 _1130_ VGND VGND VPWR VPWR _1131_ sky130_fd_sc_hd__a221o_2
Xhold907 _0744_ VGND VGND VPWR VPWR net1440 sky130_fd_sc_hd__dlygate4sd3_1
Xhold918 mgmt_gpio_data_buf\[8\] VGND VGND VPWR VPWR net1451 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3471_ net385 net1972 VGND VGND VPWR VPWR _1062_ sky130_fd_sc_hd__nor2_4
Xhold929 _0454_ VGND VGND VPWR VPWR net1462 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5210_ _1317_ net425 VGND VGND VPWR VPWR _2395_ sky130_fd_sc_hd__nand2_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6190_ gpio_configure\[13\]\[6\] net417 _2831_ gpio_configure\[16\]\[6\] VGND VGND
+ VPWR VPWR _3006_ sky130_fd_sc_hd__a22o_1
XFILLER_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5141_ _1657_ _1940_ _1826_ _1824_ VGND VGND VPWR VPWR _2348_ sky130_fd_sc_hd__o211a_1
XFILLER_69_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5072_ _1857_ _1876_ _1880_ _1602_ VGND VGND VPWR VPWR _2281_ sky130_fd_sc_hd__a31o_1
Xhold1607 mgmt_gpio_data_buf\[13\] VGND VGND VPWR VPWR net2140 sky130_fd_sc_hd__dlygate4sd3_1
X_4023_ net1828 net466 _1475_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__mux2_1
XFILLER_65_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5974_ pad_count_2\[4\] pad_count_2\[5\] VGND VGND VPWR VPWR _2796_ sky130_fd_sc_hd__nor2_4
XFILLER_80_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4925_ _1821_ _2116_ _2135_ VGND VGND VPWR VPWR _2136_ sky130_fd_sc_hd__or3b_1
XFILLER_100_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4856_ _1598_ _1607_ _1661_ _2044_ VGND VGND VPWR VPWR _2067_ sky130_fd_sc_hd__a211oi_1
XFILLER_178_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3807_ hkspi.addr\[2\] hkspi.addr\[1\] hkspi.addr\[0\] VGND VGND VPWR VPWR _1389_
+ sky130_fd_sc_hd__and3_1
XFILLER_119_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4787_ net424 _1850_ _1946_ VGND VGND VPWR VPWR _1998_ sky130_fd_sc_hd__o21bai_2
XFILLER_119_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6526_ clknet_leaf_76_csclk net1837 net484 VGND VGND VPWR VPWR gpio_configure\[25\]\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_3738_ gpio_configure\[2\]\[0\] _0908_ _0920_ gpio_configure\[10\]\[0\] VGND VGND
+ VPWR VPWR _1324_ sky130_fd_sc_hd__a22o_1
XFILLER_109_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6457_ clknet_2_0__leaf_mgmt_gpio_in[4] _0079_ _0035_ VGND VGND VPWR VPWR hkspi.writemode
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_161_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3669_ _1251_ _1252_ _1254_ _1256_ VGND VGND VPWR VPWR _1257_ sky130_fd_sc_hd__or4_1
XFILLER_118_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5408_ net446 net1170 _2421_ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__mux2_1
XFILLER_192_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6388_ wbbd_state\[9\] net168 net167 wbbd_state\[7\] VGND VGND VPWR VPWR _3179_ sky130_fd_sc_hd__a22o_1
X_5339_ net435 net1039 _2413_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__mux2_1
XFILLER_102_554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7009_ clknet_leaf_59_csclk net1313 net502 VGND VGND VPWR VPWR gpio_configure\[20\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_75_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_719 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4710_ _1678_ _1798_ _1850_ _1581_ _1921_ VGND VGND VPWR VPWR _1922_ sky130_fd_sc_hd__o221a_1
XFILLER_30_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5690_ net472 _2459_ _2466_ VGND VGND VPWR VPWR _2525_ sky130_fd_sc_hd__and3_4
XFILLER_147_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4641_ _1791_ _1833_ _1850_ net424 _1852_ VGND VGND VPWR VPWR _1853_ sky130_fd_sc_hd__o221a_1
X_4572_ _1592_ _1599_ _1783_ VGND VGND VPWR VPWR _1784_ sky130_fd_sc_hd__o21ai_1
Xmax_cap401 _2802_ VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__buf_12
XFILLER_116_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold704 _0302_ VGND VGND VPWR VPWR net1237 sky130_fd_sc_hd__dlygate4sd3_1
X_6311_ gpio_configure\[10\]\[11\] net414 net394 gpio_configure\[6\]\[11\] _3121_
+ VGND VGND VPWR VPWR _3122_ sky130_fd_sc_hd__a221o_1
Xmax_cap423 _2480_ VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__buf_12
Xhold715 gpio_configure\[24\]\[12\] VGND VGND VPWR VPWR net1248 sky130_fd_sc_hd__dlygate4sd3_1
X_3523_ gpio_configure\[31\]\[4\] net375 net355 gpio_configure\[5\]\[4\] _1113_ VGND
+ VGND VPWR VPWR _1114_ sky130_fd_sc_hd__a221o_1
Xhold726 _0103_ VGND VGND VPWR VPWR net1259 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold737 gpio_configure\[31\]\[7\] VGND VGND VPWR VPWR net1270 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold748 _0156_ VGND VGND VPWR VPWR net1281 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6242_ net359 _3048_ _3050_ _3055_ VGND VGND VPWR VPWR _3056_ sky130_fd_sc_hd__or4_1
Xhold759 gpio_configure\[3\]\[11\] VGND VGND VPWR VPWR net1292 sky130_fd_sc_hd__dlygate4sd3_1
X_3454_ _0899_ net582 VGND VGND VPWR VPWR _1045_ sky130_fd_sc_hd__nor2_4
Xmax_cap478 _1591_ VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__clkbuf_2
XFILLER_130_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3385_ gpio_configure\[29\]\[6\] _0917_ _0928_ gpio_configure\[20\]\[6\] VGND VGND
+ VPWR VPWR _0979_ sky130_fd_sc_hd__a22o_1
X_6173_ gpio_configure\[15\]\[6\] net407 net404 gpio_configure\[25\]\[6\] _2988_ VGND
+ VGND VPWR VPWR _2989_ sky130_fd_sc_hd__a221o_1
XFILLER_97_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5124_ _1729_ _2061_ _2147_ _1903_ VGND VGND VPWR VPWR _2332_ sky130_fd_sc_hd__or4b_1
Xhold1404 net341 VGND VGND VPWR VPWR net1937 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1415 net342 VGND VGND VPWR VPWR net1948 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1426 net330 VGND VGND VPWR VPWR net1959 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1437 wbbd_addr\[3\] VGND VGND VPWR VPWR net1970 sky130_fd_sc_hd__dlygate4sd3_1
X_5055_ _2041_ _2052_ _2151_ _2263_ VGND VGND VPWR VPWR _2264_ sky130_fd_sc_hd__or4_1
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1448 gpio_configure\[15\]\[10\] VGND VGND VPWR VPWR net1981 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1459 _0422_ VGND VGND VPWR VPWR net1992 sky130_fd_sc_hd__dlygate4sd3_1
X_4006_ net618 net700 _1472_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__mux2_1
XFILLER_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5957_ _2773_ _2775_ _2777_ _2779_ VGND VGND VPWR VPWR _2780_ sky130_fd_sc_hd__or4_1
X_4908_ _1678_ _1805_ net432 _1798_ VGND VGND VPWR VPWR _2119_ sky130_fd_sc_hd__o22ai_1
XFILLER_21_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5888_ gpio_configure\[24\]\[9\] net418 _2713_ VGND VGND VPWR VPWR _2714_ sky130_fd_sc_hd__a21o_1
XFILLER_178_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4839_ _1681_ _1685_ VGND VGND VPWR VPWR _2050_ sky130_fd_sc_hd__nor2_1
XFILLER_138_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6509_ clknet_leaf_3_csclk net1275 net493 VGND VGND VPWR VPWR gpio_configure\[23\]\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_134_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold20 _0875_ VGND VGND VPWR VPWR net553 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold31 net350 VGND VGND VPWR VPWR net564 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold42 hkspi.odata\[2\] VGND VGND VPWR VPWR net575 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 hkspi.addr\[1\] VGND VGND VPWR VPWR net586 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold64 hkspi.addr\[2\] VGND VGND VPWR VPWR net597 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 _0872_ VGND VGND VPWR VPWR net608 sky130_fd_sc_hd__buf_6
Xhold86 net1910 VGND VGND VPWR VPWR net619 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 _1509_ VGND VGND VPWR VPWR net630 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_6 _0909_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6860_ clknet_leaf_28_csclk net1571 net520 VGND VGND VPWR VPWR gpio_configure\[2\]\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_35_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5811_ gpio_configure\[9\]\[5\] _2512_ _2529_ gpio_configure\[29\]\[5\] VGND VGND
+ VPWR VPWR _2641_ sky130_fd_sc_hd__a22o_1
XFILLER_62_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6791_ clknet_leaf_77_csclk net1601 net484 VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__dfrtp_2
XFILLER_50_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5742_ gpio_configure\[21\]\[2\] _2521_ net418 gpio_configure\[24\]\[2\] _2574_ VGND
+ VGND VPWR VPWR _2575_ sky130_fd_sc_hd__a221o_1
XFILLER_50_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5673_ gpio_configure\[27\]\[0\] _2506_ net421 gpio_configure\[10\]\[0\] VGND VGND
+ VPWR VPWR _2508_ sky130_fd_sc_hd__a22o_1
XFILLER_148_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4624_ net477 _1833_ VGND VGND VPWR VPWR _1836_ sky130_fd_sc_hd__or2_4
XFILLER_163_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold501 _0713_ VGND VGND VPWR VPWR net1034 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4555_ _1759_ _1766_ VGND VGND VPWR VPWR _1767_ sky130_fd_sc_hd__nor2_1
Xhold512 gpio_configure\[17\]\[7\] VGND VGND VPWR VPWR net1045 sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 _0812_ VGND VGND VPWR VPWR net1056 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold534 net269 VGND VGND VPWR VPWR net1067 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3506_ gpio_configure\[2\]\[4\] _0908_ _1093_ gpio_configure\[4\]\[12\] _1096_ VGND
+ VGND VPWR VPWR _1097_ sky130_fd_sc_hd__a221o_1
Xhold545 _0456_ VGND VGND VPWR VPWR net1078 sky130_fd_sc_hd__dlygate4sd3_1
Xhold556 gpio_configure\[20\]\[3\] VGND VGND VPWR VPWR net1089 sky130_fd_sc_hd__dlygate4sd3_1
X_4486_ _1651_ _1663_ VGND VGND VPWR VPWR _1698_ sky130_fd_sc_hd__nor2_1
Xhold567 gpio_configure\[2\]\[7\] VGND VGND VPWR VPWR net1100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 _0322_ VGND VGND VPWR VPWR net1111 sky130_fd_sc_hd__dlygate4sd3_1
X_6225_ gpio_configure\[3\]\[8\] _2830_ _2842_ gpio_configure\[15\]\[8\] VGND VGND
+ VPWR VPWR _3039_ sky130_fd_sc_hd__a22o_1
Xhold589 gpio_configure\[2\]\[5\] VGND VGND VPWR VPWR net1122 sky130_fd_sc_hd__dlygate4sd3_1
X_3437_ gpio_configure\[14\]\[5\] _0916_ _0933_ net68 _1028_ VGND VGND VPWR VPWR _1029_
+ sky130_fd_sc_hd__a221o_1
XFILLER_106_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3368_ gpio_configure\[27\]\[7\] net370 _0934_ gpio_configure\[1\]\[7\] _0942_ VGND
+ VGND VPWR VPWR _0964_ sky130_fd_sc_hd__a221o_1
X_6156_ _2967_ _2968_ _2970_ _2972_ VGND VGND VPWR VPWR _2973_ sky130_fd_sc_hd__or4_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1201 gpio_configure\[21\]\[9\] VGND VGND VPWR VPWR net1734 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1212 _0396_ VGND VGND VPWR VPWR net1745 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5107_ _1829_ _2292_ _1885_ _1888_ VGND VGND VPWR VPWR _2315_ sky130_fd_sc_hd__or4b_1
Xhold1223 _0229_ VGND VGND VPWR VPWR net1756 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1234 reset_reg VGND VGND VPWR VPWR net1767 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6087_ gpio_configure\[18\]\[2\] net399 net411 gpio_configure\[14\]\[2\] _2906_ VGND
+ VGND VPWR VPWR _2907_ sky130_fd_sc_hd__a221o_1
X_3299_ _0857_ net2006 VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__nand2_8
Xhold1245 _0573_ VGND VGND VPWR VPWR net1778 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1256 gpio_configure\[9\]\[0\] VGND VGND VPWR VPWR net1789 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1267 gpio_configure\[1\]\[8\] VGND VGND VPWR VPWR net1800 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1278 _0133_ VGND VGND VPWR VPWR net1811 sky130_fd_sc_hd__dlygate4sd3_1
X_5038_ _1608_ _1880_ _2047_ _1618_ VGND VGND VPWR VPWR _2247_ sky130_fd_sc_hd__a31o_1
Xhold1289 gpio_configure\[31\]\[8\] VGND VGND VPWR VPWR net1822 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6989_ clknet_leaf_36_csclk net1153 net523 VGND VGND VPWR VPWR gpio_configure\[18\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_41_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput110 wb_adr_i[1] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__buf_6
Xinput121 wb_adr_i[2] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_2
Xinput132 wb_dat_i[0] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput143 wb_dat_i[1] VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_1
XFILLER_49_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput154 wb_dat_i[2] VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_1
Xinput165 wb_sel_i[0] VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4340_ _1549_ _1550_ _1551_ VGND VGND VPWR VPWR _1552_ sky130_fd_sc_hd__and3_1
XFILLER_125_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4271_ net1779 net470 _1537_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__mux2_1
XFILLER_141_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6010_ gpio_configure\[3\]\[0\] _2830_ _2831_ gpio_configure\[16\]\[0\] VGND VGND
+ VPWR VPWR _2832_ sky130_fd_sc_hd__a22o_1
X_3222_ gpio_configure\[12\]\[3\] VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__inv_2
XFILLER_140_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6912_ clknet_leaf_33_csclk net536 net524 VGND VGND VPWR VPWR gpio_configure\[8\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_35_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6843_ clknet_leaf_67_csclk net881 net505 VGND VGND VPWR VPWR gpio_configure\[0\]\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_62_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6774_ clknet_leaf_71_csclk net993 net498 VGND VGND VPWR VPWR gpio_configure\[22\]\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_3986_ net1692 net455 _1470_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__mux2_1
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5725_ gpio_configure\[19\]\[1\] _2491_ _2496_ gpio_configure\[5\]\[1\] _2558_ VGND
+ VGND VPWR VPWR _2559_ sky130_fd_sc_hd__a221o_1
XFILLER_148_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5656_ pad_count_1\[4\] _2461_ _2466_ VGND VGND VPWR VPWR _2491_ sky130_fd_sc_hd__and3_4
XFILLER_191_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4607_ _1785_ _0834_ _1584_ _1818_ VGND VGND VPWR VPWR _1819_ sky130_fd_sc_hd__and4b_1
X_5587_ net437 net1439 net603 VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__mux2_1
Xhold320 _0555_ VGND VGND VPWR VPWR net853 sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 net303 VGND VGND VPWR VPWR net864 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4538_ net99 _1610_ VGND VGND VPWR VPWR _1750_ sky130_fd_sc_hd__nand2_8
XFILLER_190_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold342 _0630_ VGND VGND VPWR VPWR net875 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold353 gpio_configure\[2\]\[1\] VGND VGND VPWR VPWR net886 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold364 _0282_ VGND VGND VPWR VPWR net897 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold375 gpio_configure\[8\]\[7\] VGND VGND VPWR VPWR net908 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold386 _0271_ VGND VGND VPWR VPWR net919 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4469_ _1564_ _1678_ VGND VGND VPWR VPWR _1681_ sky130_fd_sc_hd__or2_1
Xhold397 gpio_configure\[4\]\[7\] VGND VGND VPWR VPWR net930 sky130_fd_sc_hd__dlygate4sd3_1
X_6208_ gpio_configure\[37\]\[7\] net400 net416 gpio_configure\[32\]\[7\] _3012_ VGND
+ VGND VPWR VPWR _3023_ sky130_fd_sc_hd__a221o_1
X_7188_ clknet_3_7_0_wb_clk_i _0790_ net528 VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__dfrtp_4
XFILLER_58_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6139_ gpio_configure\[2\]\[4\] _2823_ net392 gpio_configure\[5\]\[4\] _2956_ VGND
+ VGND VPWR VPWR _2957_ sky130_fd_sc_hd__a221o_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1020 _0506_ VGND VGND VPWR VPWR net1553 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1031 gpio_configure\[6\]\[0\] VGND VGND VPWR VPWR net1564 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1042 _0120_ VGND VGND VPWR VPWR net1575 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_133_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1053 gpio_configure\[10\]\[2\] VGND VGND VPWR VPWR net1586 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1064 _0629_ VGND VGND VPWR VPWR net1597 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1075 gpio_configure\[17\]\[0\] VGND VGND VPWR VPWR net1608 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1086 gpio_configure\[26\]\[9\] VGND VGND VPWR VPWR net1619 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1097 _0160_ VGND VGND VPWR VPWR net1630 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_204 _2804_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_215 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_226 net394 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_237 net471 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_248 _2528_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_259 net569 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_5_csclk clknet_3_1_0_csclk VGND VGND VPWR VPWR clknet_leaf_5_csclk sky130_fd_sc_hd__clkbuf_16
XFILLER_150_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3840_ hkspi.pass_thru_mgmt_delay hkspi.pre_pass_thru_mgmt _1411_ VGND VGND VPWR
+ VPWR _0082_ sky130_fd_sc_hd__mux2_1
XFILLER_32_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3771_ gpio_configure\[27\]\[0\] _0925_ _1046_ gpio_configure\[28\]\[8\] _1356_ VGND
+ VGND VPWR VPWR _1357_ sky130_fd_sc_hd__a221o_1
XFILLER_158_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5510_ net435 net928 _2432_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__mux2_1
XFILLER_157_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6490_ clknet_leaf_73_csclk net1827 net488 VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__dfstp_2
XFILLER_9_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5441_ net464 net1330 _2425_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__mux2_1
XFILLER_172_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5372_ net446 net1190 _2417_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__mux2_1
X_7111_ clknet_leaf_15_csclk net1563 net527 VGND VGND VPWR VPWR gpio_configure\[34\]\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_4323_ net1246 net443 _1545_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__mux2_1
XFILLER_153_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7042_ clknet_leaf_69_csclk net1815 net497 VGND VGND VPWR VPWR gpio_configure\[25\]\[0\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_101_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4254_ net1475 net462 _1534_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__mux2_1
XFILLER_141_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3205_ gpio_configure\[29\]\[3\] VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__inv_2
XFILLER_101_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4185_ net321 clknet_1_1__leaf__1134_ _1519_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__mux2_1
XFILLER_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6826_ clknet_leaf_28_csclk net1505 net520 VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__dfrtp_1
XFILLER_51_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6757_ clknet_leaf_73_csclk net1339 net488 VGND VGND VPWR VPWR gpio_configure\[33\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_149_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3969_ net537 net540 net474 VGND VGND VPWR VPWR _1463_ sky130_fd_sc_hd__mux2_8
XFILLER_50_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5708_ _2522_ _2530_ _2536_ _2542_ VGND VGND VPWR VPWR _2543_ sky130_fd_sc_hd__or4_1
XFILLER_109_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6688_ clknet_leaf_5_csclk net1323 net496 VGND VGND VPWR VPWR gpio_configure\[13\]\[10\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_148_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5639_ _2474_ _2477_ _2476_ VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__a21oi_1
XFILLER_164_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold150 gpio_configure\[35\]\[11\] VGND VGND VPWR VPWR net683 sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 gpio_configure\[2\]\[3\] VGND VGND VPWR VPWR net694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 _0734_ VGND VGND VPWR VPWR net705 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold183 gpio_configure\[14\]\[7\] VGND VGND VPWR VPWR net716 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 _0206_ VGND VGND VPWR VPWR net727 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5990_ gpio_configure\[26\]\[0\] _2810_ _2811_ gpio_configure\[7\]\[0\] VGND VGND
+ VPWR VPWR _2812_ sky130_fd_sc_hd__a22o_1
XFILLER_64_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4941_ _1631_ _1658_ _2043_ _2150_ VGND VGND VPWR VPWR _2151_ sky130_fd_sc_hd__a211o_1
X_4872_ _1657_ _2081_ VGND VGND VPWR VPWR _2083_ sky130_fd_sc_hd__nor2_1
XFILLER_178_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6611_ clknet_leaf_78_csclk net1679 net486 VGND VGND VPWR VPWR gpio_configure\[3\]\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_3823_ hkspi.addr\[3\] _1389_ VGND VGND VPWR VPWR _1401_ sky130_fd_sc_hd__or2_1
X_6542_ clknet_2_1__leaf_mgmt_gpio_in[4] _0005_ _0053_ VGND VGND VPWR VPWR hkspi.state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3754_ gpio_configure\[13\]\[0\] _0906_ _1102_ gpio_configure\[15\]\[8\] _1324_ VGND
+ VGND VPWR VPWR _1340_ sky130_fd_sc_hd__a221o_1
XFILLER_158_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6473_ clknet_2_1__leaf_mgmt_gpio_in[4] _0095_ _0051_ VGND VGND VPWR VPWR hkspi.count\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_3685_ gpio_configure\[23\]\[1\] _0922_ _1093_ gpio_configure\[4\]\[9\] _1272_ VGND
+ VGND VPWR VPWR _1273_ sky130_fd_sc_hd__a221o_2
X_5424_ net457 net772 _2423_ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__mux2_1
XFILLER_161_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput200 net200 VGND VGND VPWR VPWR mgmt_gpio_oeb[32] sky130_fd_sc_hd__buf_12
Xoutput211 net211 VGND VGND VPWR VPWR mgmt_gpio_oeb[8] sky130_fd_sc_hd__buf_12
Xoutput222 net222 VGND VGND VPWR VPWR mgmt_gpio_out[18] sky130_fd_sc_hd__buf_12
Xoutput233 net233 VGND VGND VPWR VPWR mgmt_gpio_out[28] sky130_fd_sc_hd__buf_12
Xoutput244 net244 VGND VGND VPWR VPWR mgmt_gpio_out[3] sky130_fd_sc_hd__buf_12
XFILLER_160_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5355_ net440 net1522 _2415_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__mux2_1
Xoutput255 net255 VGND VGND VPWR VPWR pad_flash_io0_do sky130_fd_sc_hd__buf_12
Xoutput266 net266 VGND VGND VPWR VPWR pll_div[0] sky130_fd_sc_hd__buf_12
Xoutput277 net277 VGND VGND VPWR VPWR pll_trim[11] sky130_fd_sc_hd__buf_12
X_4306_ _1053_ net425 VGND VGND VPWR VPWR _1543_ sky130_fd_sc_hd__nand2_4
Xoutput288 net288 VGND VGND VPWR VPWR pll_trim[21] sky130_fd_sc_hd__buf_12
XFILLER_160_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput299 net299 VGND VGND VPWR VPWR pll_trim[8] sky130_fd_sc_hd__buf_12
XFILLER_99_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5286_ net564 net428 VGND VGND VPWR VPWR _2408_ sky130_fd_sc_hd__nand2_4
XFILLER_141_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7025_ clknet_leaf_50_csclk net653 net507 VGND VGND VPWR VPWR gpio_configure\[22\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_4237_ net577 net1936 net592 VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__mux2_1
XFILLER_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4168_ net1960 _1249_ _1517_ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__mux2_1
XFILLER_95_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4099_ net1373 _1505_ _1499_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__mux2_1
XFILLER_43_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6809_ clknet_leaf_57_csclk net865 net503 VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__dfrtp_4
XFILLER_11_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_70_csclk clknet_3_0_0_csclk VGND VGND VPWR VPWR clknet_leaf_70_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_124_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout460 net576 VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__buf_4
XFILLER_93_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout471 net1098 VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__buf_8
Xfanout482 net483 VGND VGND VPWR VPWR net482 sky130_fd_sc_hd__buf_4
XFILLER_46_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout493 net496 VGND VGND VPWR VPWR net493 sky130_fd_sc_hd__buf_6
XFILLER_58_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_23_csclk clknet_3_4_0_csclk VGND VGND VPWR VPWR clknet_leaf_23_csclk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_38_csclk clknet_3_7_0_csclk VGND VGND VPWR VPWR clknet_leaf_38_csclk
+ sky130_fd_sc_hd__clkbuf_16
Xhold908 gpio_configure\[13\]\[9\] VGND VGND VPWR VPWR net1441 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold919 _0437_ VGND VGND VPWR VPWR net1452 sky130_fd_sc_hd__dlygate4sd3_1
X_3470_ gpio_configure\[10\]\[4\] _0920_ _0939_ gpio_configure\[8\]\[4\] _1060_ VGND
+ VGND VPWR VPWR _1061_ sky130_fd_sc_hd__a221o_1
XFILLER_127_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5140_ _2180_ _2320_ _2327_ VGND VGND VPWR VPWR _2347_ sky130_fd_sc_hd__or3b_1
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1608 pad_count_2\[3\] VGND VGND VPWR VPWR net2141 sky130_fd_sc_hd__dlygate4sd3_1
X_5071_ _1529_ _2222_ _2241_ VGND VGND VPWR VPWR _2280_ sky130_fd_sc_hd__or3_1
XFILLER_96_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4022_ _1073_ net426 VGND VGND VPWR VPWR _1475_ sky130_fd_sc_hd__and2_2
XFILLER_84_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5973_ _1447_ _2794_ VGND VGND VPWR VPWR _2795_ sky130_fd_sc_hd__nor2_2
XFILLER_64_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4924_ _2126_ _2134_ VGND VGND VPWR VPWR _2135_ sky130_fd_sc_hd__nor2_1
XFILLER_178_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4855_ _1606_ net432 _1863_ _1777_ _2048_ VGND VGND VPWR VPWR _2066_ sky130_fd_sc_hd__o221a_1
X_3806_ hkspi.state\[0\] _1387_ VGND VGND VPWR VPWR _1388_ sky130_fd_sc_hd__nand2b_4
XFILLER_166_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4786_ _1635_ _1744_ _1802_ VGND VGND VPWR VPWR _1997_ sky130_fd_sc_hd__a21oi_1
XFILLER_165_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6525_ clknet_leaf_3_csclk net1255 net495 VGND VGND VPWR VPWR gpio_configure\[29\]\[12\]
+ sky130_fd_sc_hd__dfrtp_4
X_3737_ gpio_configure\[9\]\[8\] _1057_ _1119_ gpio_configure\[5\]\[8\] VGND VGND
+ VPWR VPWR _1323_ sky130_fd_sc_hd__a22o_2
XFILLER_118_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6456_ clknet_2_0__leaf_mgmt_gpio_in[4] _0078_ _0034_ VGND VGND VPWR VPWR hkspi.readmode
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_146_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3668_ gpio_configure\[37\]\[1\] _0902_ _0927_ gpio_configure\[25\]\[1\] _1255_ VGND
+ VGND VPWR VPWR _1256_ sky130_fd_sc_hd__a221o_1
XFILLER_133_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5407_ net453 net1136 _2421_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__mux2_1
X_6387_ clknet_1_0__leaf_wbbd_sck _1528_ _1529_ _0820_ VGND VGND VPWR VPWR _0807_
+ sky130_fd_sc_hd__o211a_2
X_3599_ gpio_configure\[30\]\[3\] _0892_ _1125_ gpio_configure\[22\]\[11\] _1188_
+ VGND VGND VPWR VPWR _1189_ sky130_fd_sc_hd__a221o_1
XFILLER_88_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5338_ net438 net1342 _2413_ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__mux2_1
XFILLER_102_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5269_ net469 net1616 _2406_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__mux2_1
X_7008_ clknet_leaf_59_csclk net1472 net502 VGND VGND VPWR VPWR gpio_configure\[20\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4640_ _1798_ _1805_ net424 VGND VGND VPWR VPWR _1852_ sky130_fd_sc_hd__a21o_1
XFILLER_30_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4571_ _1774_ _1777_ _1780_ _1609_ VGND VGND VPWR VPWR _1783_ sky130_fd_sc_hd__o211a_1
XFILLER_190_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap402 _2798_ VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__buf_8
X_6310_ gpio_configure\[9\]\[11\] net412 _2838_ gpio_configure\[12\]\[11\] VGND VGND
+ VPWR VPWR _3121_ sky130_fd_sc_hd__a22o_1
Xmax_cap413 _2830_ VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__buf_8
X_3522_ gpio_configure\[30\]\[4\] _0892_ _0925_ gpio_configure\[27\]\[4\] VGND VGND
+ VPWR VPWR _1113_ sky130_fd_sc_hd__a22o_1
Xhold705 gpio_configure\[16\]\[4\] VGND VGND VPWR VPWR net1238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold716 _0142_ VGND VGND VPWR VPWR net1249 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold727 gpio_configure\[14\]\[11\] VGND VGND VPWR VPWR net1260 sky130_fd_sc_hd__dlygate4sd3_1
Xhold738 _0127_ VGND VGND VPWR VPWR net1271 sky130_fd_sc_hd__dlygate4sd3_1
X_6241_ _3038_ _3039_ _3052_ _3054_ VGND VGND VPWR VPWR _3055_ sky130_fd_sc_hd__or4_1
Xhold749 gpio_configure\[33\]\[10\] VGND VGND VPWR VPWR net1282 sky130_fd_sc_hd__dlygate4sd3_1
X_3453_ gpio_configure\[7\]\[4\] _0913_ _1041_ gpio_configure\[31\]\[12\] _1043_ VGND
+ VGND VPWR VPWR _1044_ sky130_fd_sc_hd__a221o_1
XFILLER_170_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap479 net480 VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__clkbuf_2
X_6172_ gpio_configure\[26\]\[6\] _2810_ net409 gpio_configure\[12\]\[6\] VGND VGND
+ VPWR VPWR _2988_ sky130_fd_sc_hd__a22o_1
X_3384_ gpio_configure\[17\]\[6\] _0937_ _0940_ net280 VGND VGND VPWR VPWR _0978_
+ sky130_fd_sc_hd__a22o_1
XFILLER_97_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5123_ _2165_ _2266_ _2330_ VGND VGND VPWR VPWR _2331_ sky130_fd_sc_hd__and3_1
Xhold1405 net333 VGND VGND VPWR VPWR net1938 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1416 net286 VGND VGND VPWR VPWR net1949 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1427 net327 VGND VGND VPWR VPWR net1960 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1438 _0857_ VGND VGND VPWR VPWR net1971 sky130_fd_sc_hd__dlygate4sd3_1
X_5054_ _1733_ _1889_ VGND VGND VPWR VPWR _2263_ sky130_fd_sc_hd__nand2_1
Xhold1449 _0311_ VGND VGND VPWR VPWR net1982 sky130_fd_sc_hd__dlygate4sd3_1
X_4005_ net452 net1023 _1472_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__mux2_1
XFILLER_65_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5956_ gpio_configure\[20\]\[12\] _2499_ _2505_ gpio_configure\[11\]\[12\] _2778_
+ VGND VGND VPWR VPWR _2779_ sky130_fd_sc_hd__a221o_1
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4907_ _1794_ _1806_ _1831_ _2117_ VGND VGND VPWR VPWR _2118_ sky130_fd_sc_hd__or4_1
XFILLER_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5887_ gpio_configure\[22\]\[9\] _2498_ _2502_ gpio_configure\[4\]\[9\] VGND VGND
+ VPWR VPWR _2713_ sky130_fd_sc_hd__a22o_1
XFILLER_138_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4838_ _1587_ net380 VGND VGND VPWR VPWR _2049_ sky130_fd_sc_hd__and2_1
XFILLER_138_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4769_ _1658_ _1706_ _1953_ _1954_ _1980_ VGND VGND VPWR VPWR _1981_ sky130_fd_sc_hd__a2111o_1
XFILLER_107_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6508_ clknet_leaf_78_csclk net1647 net486 VGND VGND VPWR VPWR gpio_configure\[23\]\[10\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_193_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6439_ net495 net482 VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__and2_1
XFILLER_162_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold10 _0425_ VGND VGND VPWR VPWR net543 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 net377 VGND VGND VPWR VPWR net554 sky130_fd_sc_hd__buf_8
XFILLER_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold32 _2408_ VGND VGND VPWR VPWR net565 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 net595 VGND VGND VPWR VPWR net576 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold54 _0858_ VGND VGND VPWR VPWR net587 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 _0855_ VGND VGND VPWR VPWR net598 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 _0926_ VGND VGND VPWR VPWR net609 sky130_fd_sc_hd__buf_8
XFILLER_188_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold87 gpio_configure\[11\]\[9\] VGND VGND VPWR VPWR net620 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold98 _0199_ VGND VGND VPWR VPWR net631 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_7 _0913_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5810_ gpio_configure\[7\]\[5\] _2528_ _2538_ gpio_configure\[1\]\[5\] _2639_ VGND
+ VGND VPWR VPWR _2640_ sky130_fd_sc_hd__a221o_1
X_6790_ clknet_2_1__leaf_mgmt_gpio_in[4] _0393_ _0064_ VGND VGND VPWR VPWR hkspi.SDO
+ sky130_fd_sc_hd__dfrtn_1
X_5741_ gpio_configure\[15\]\[2\] _2510_ _2537_ gpio_configure\[17\]\[2\] VGND VGND
+ VPWR VPWR _2574_ sky130_fd_sc_hd__a22o_1
XFILLER_148_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5672_ net472 _2489_ _2504_ VGND VGND VPWR VPWR _2507_ sky130_fd_sc_hd__and3_4
XFILLER_187_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4623_ _1795_ _1833_ VGND VGND VPWR VPWR _1835_ sky130_fd_sc_hd__nor2_1
XFILLER_148_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4554_ _1752_ _1765_ _1764_ VGND VGND VPWR VPWR _1766_ sky130_fd_sc_hd__o21bai_1
Xhold502 gpio_configure\[33\]\[11\] VGND VGND VPWR VPWR net1035 sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 _0588_ VGND VGND VPWR VPWR net1046 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold524 gpio_configure\[5\]\[7\] VGND VGND VPWR VPWR net1057 sky130_fd_sc_hd__dlygate4sd3_1
X_3505_ gpio_configure\[7\]\[12\] _1094_ _1095_ gpio_configure\[3\]\[12\] VGND VGND
+ VPWR VPWR _1096_ sky130_fd_sc_hd__a22o_1
Xhold535 _0399_ VGND VGND VPWR VPWR net1068 sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 gpio_configure\[1\]\[11\] VGND VGND VPWR VPWR net1079 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4485_ _1635_ _1662_ VGND VGND VPWR VPWR _1697_ sky130_fd_sc_hd__nand2_1
XFILLER_116_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold557 _0608_ VGND VGND VPWR VPWR net1090 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold568 _0468_ VGND VGND VPWR VPWR net1101 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6224_ gpio_configure\[26\]\[8\] _2810_ _2811_ gpio_configure\[7\]\[8\] VGND VGND
+ VPWR VPWR _3038_ sky130_fd_sc_hd__a22o_1
Xhold579 gpio_configure\[34\]\[12\] VGND VGND VPWR VPWR net1112 sky130_fd_sc_hd__dlygate4sd3_1
X_3436_ gpio_configure\[12\]\[5\] _0921_ net352 gpio_configure\[36\]\[5\] VGND VGND
+ VPWR VPWR _1028_ sky130_fd_sc_hd__a22o_1
XFILLER_131_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6155_ gpio_configure\[16\]\[5\] _2831_ net391 gpio_configure\[17\]\[5\] _2971_ VGND
+ VGND VPWR VPWR _2972_ sky130_fd_sc_hd__a221o_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3367_ gpio_configure\[19\]\[7\] _0896_ _0919_ gpio_configure\[24\]\[7\] _0941_ VGND
+ VGND VPWR VPWR _0963_ sky130_fd_sc_hd__a221o_2
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1202 _0365_ VGND VGND VPWR VPWR net1735 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5106_ _1695_ _2228_ _2288_ _2313_ VGND VGND VPWR VPWR _2314_ sky130_fd_sc_hd__or4b_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1213 gpio_configure\[28\]\[10\] VGND VGND VPWR VPWR net1746 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6086_ gpio_configure\[16\]\[2\] _2831_ _2852_ gpio_configure\[19\]\[2\] VGND VGND
+ VPWR VPWR _2906_ sky130_fd_sc_hd__a22o_1
Xhold1224 gpio_configure\[3\]\[0\] VGND VGND VPWR VPWR net1757 sky130_fd_sc_hd__dlygate4sd3_1
X_3298_ _0873_ net385 VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__nor2_8
Xhold1235 _0414_ VGND VGND VPWR VPWR net1768 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1246 gpio_configure\[17\]\[8\] VGND VGND VPWR VPWR net1779 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1257 _0517_ VGND VGND VPWR VPWR net1790 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5037_ _1635_ _2244_ _2245_ _1629_ VGND VGND VPWR VPWR _2246_ sky130_fd_sc_hd__a22o_1
Xhold1268 _0214_ VGND VGND VPWR VPWR net1801 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1279 gpio_configure\[9\]\[8\] VGND VGND VPWR VPWR net1812 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6988_ clknet_leaf_64_csclk net851 net501 VGND VGND VPWR VPWR gpio_configure\[18\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_15_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5939_ gpio_configure\[9\]\[11\] _2512_ _2524_ _2762_ VGND VGND VPWR VPWR _2763_
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput100 wb_adr_i[10] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput111 wb_adr_i[20] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_4
XFILLER_49_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput122 wb_adr_i[30] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput133 wb_dat_i[10] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_1
Xinput144 wb_dat_i[20] VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__clkbuf_1
Xinput155 wb_dat_i[30] VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput166 wb_sel_i[1] VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4270_ _1121_ net429 VGND VGND VPWR VPWR _1537_ sky130_fd_sc_hd__and2_2
XFILLER_113_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3221_ gpio_configure\[13\]\[3\] VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__inv_2
XFILLER_79_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6911_ clknet_leaf_32_csclk net1529 net524 VGND VGND VPWR VPWR gpio_configure\[8\]\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_63_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6842_ clknet_leaf_65_csclk net1643 net501 VGND VGND VPWR VPWR gpio_configure\[0\]\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_62_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6773_ clknet_leaf_70_csclk net1703 net491 VGND VGND VPWR VPWR gpio_configure\[22\]\[10\]
+ sky130_fd_sc_hd__dfstp_1
X_3985_ net1715 net461 _1470_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__mux2_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5724_ gpio_configure\[6\]\[1\] _2490_ _2502_ gpio_configure\[4\]\[1\] VGND VGND
+ VPWR VPWR _2558_ sky130_fd_sc_hd__a22o_1
X_5655_ net472 _2488_ _2489_ VGND VGND VPWR VPWR _2490_ sky130_fd_sc_hd__and3_4
XFILLER_148_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4606_ _1766_ _1816_ _1817_ _1762_ VGND VGND VPWR VPWR _1818_ sky130_fd_sc_hd__and4b_1
X_5586_ net440 net1532 net603 VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__mux2_1
XFILLER_190_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold310 _0647_ VGND VGND VPWR VPWR net843 sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 net292 VGND VGND VPWR VPWR net854 sky130_fd_sc_hd__dlygate4sd3_1
X_4537_ net110 net99 net124 net530 VGND VGND VPWR VPWR _1749_ sky130_fd_sc_hd__and4_4
Xhold332 _0412_ VGND VGND VPWR VPWR net865 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold343 gpio_configure\[36\]\[9\] VGND VGND VPWR VPWR net876 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold354 _0462_ VGND VGND VPWR VPWR net887 sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 gpio_configure\[7\]\[12\] VGND VGND VPWR VPWR net898 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold376 _0516_ VGND VGND VPWR VPWR net909 sky130_fd_sc_hd__dlygate4sd3_1
X_4468_ _1575_ _1679_ _1563_ VGND VGND VPWR VPWR _1680_ sky130_fd_sc_hd__or3b_2
Xhold387 gpio_configure\[9\]\[11\] VGND VGND VPWR VPWR net920 sky130_fd_sc_hd__dlygate4sd3_1
Xhold398 _0484_ VGND VGND VPWR VPWR net931 sky130_fd_sc_hd__dlygate4sd3_1
X_6207_ gpio_configure\[28\]\[7\] _2861_ _3017_ _3019_ _3021_ VGND VGND VPWR VPWR
+ _3022_ sky130_fd_sc_hd__a2111o_1
XFILLER_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3419_ gpio_configure\[2\]\[5\] _0908_ _0920_ gpio_configure\[10\]\[5\] VGND VGND
+ VPWR VPWR _1011_ sky130_fd_sc_hd__a22o_1
X_7187_ clknet_3_1_0_wb_clk_i _0789_ net490 VGND VGND VPWR VPWR serial_data_staging_2\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_4399_ _0832_ _1555_ VGND VGND VPWR VPWR _1611_ sky130_fd_sc_hd__or2_2
XFILLER_98_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6138_ gpio_configure\[13\]\[4\] net417 net404 gpio_configure\[25\]\[4\] VGND VGND
+ VPWR VPWR _2956_ sky130_fd_sc_hd__a22o_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1010 _0522_ VGND VGND VPWR VPWR net1543 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1021 gpio_configure\[17\]\[5\] VGND VGND VPWR VPWR net1554 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1032 _0493_ VGND VGND VPWR VPWR net1565 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1043 net291 VGND VGND VPWR VPWR net1576 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6069_ net363 _2879_ _2881_ _2889_ VGND VGND VPWR VPWR _2890_ sky130_fd_sc_hd__or4_1
XFILLER_100_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1054 _0527_ VGND VGND VPWR VPWR net1587 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1065 gpio_configure\[29\]\[0\] VGND VGND VPWR VPWR net1598 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_133_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1076 _0581_ VGND VGND VPWR VPWR net1609 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1087 _0159_ VGND VGND VPWR VPWR net1620 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1098 net1984 VGND VGND VPWR VPWR net1631 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_205 _2810_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_216 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_227 net405 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_238 net542 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_249 _2540_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3770_ gpio_configure\[1\]\[8\] _1103_ _1137_ net98 VGND VGND VPWR VPWR _1356_ sky130_fd_sc_hd__a22o_1
XFILLER_118_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5440_ net1098 net1214 _2425_ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__mux2_1
XFILLER_173_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5371_ net453 net1130 _2417_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__mux2_1
X_7110_ clknet_leaf_50_csclk net1034 net507 VGND VGND VPWR VPWR gpio_configure\[33\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_4322_ net1244 net449 _1545_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__mux2_1
XFILLER_113_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7041_ clknet_leaf_58_csclk net1267 net503 VGND VGND VPWR VPWR gpio_configure\[24\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_113_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4253_ net1802 net468 _1534_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__mux2_1
XFILLER_87_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3204_ gpio_configure\[30\]\[3\] VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__inv_2
X_4184_ net1958 _1191_ _1519_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__mux2_1
XFILLER_95_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_7_0_wb_clk_i clknet_2_3_0_wb_clk_i VGND VGND VPWR VPWR clknet_3_7_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_6825_ clknet_leaf_71_csclk net1613 net491 VGND VGND VPWR VPWR irq_2_inputsrc sky130_fd_sc_hd__dfrtp_1
XFILLER_50_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3968_ net1820 net467 _1461_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__mux2_1
X_6756_ clknet_leaf_73_csclk net1825 net488 VGND VGND VPWR VPWR gpio_configure\[33\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_149_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5707_ gpio_configure\[12\]\[0\] _2540_ _2541_ gpio_configure\[31\]\[0\] _2539_ VGND
+ VGND VPWR VPWR _2542_ sky130_fd_sc_hd__a221o_1
XFILLER_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6687_ clknet_leaf_5_csclk net1442 net494 VGND VGND VPWR VPWR gpio_configure\[13\]\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_109_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3899_ net307 _1444_ xfer_count\[2\] xfer_count\[3\] VGND VGND VPWR VPWR _1445_ sky130_fd_sc_hd__and4b_1
XFILLER_149_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5638_ pad_count_2\[4\] _2462_ VGND VGND VPWR VPWR _2477_ sky130_fd_sc_hd__nor2_1
XFILLER_164_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5569_ net439 net1916 net648 VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__mux2_1
XFILLER_2_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold140 net279 VGND VGND VPWR VPWR net673 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 _0342_ VGND VGND VPWR VPWR net684 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold162 _0464_ VGND VGND VPWR VPWR net695 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold173 net2106 VGND VGND VPWR VPWR net706 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 _0564_ VGND VGND VPWR VPWR net717 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 gpio_configure\[10\]\[3\] VGND VGND VPWR VPWR net728 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4940_ _1680_ _1684_ VGND VGND VPWR VPWR _2150_ sky130_fd_sc_hd__nor2_1
XFILLER_64_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4871_ _1643_ _1707_ VGND VGND VPWR VPWR _2082_ sky130_fd_sc_hd__nand2_1
XFILLER_33_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3822_ _1400_ hkspi.addr\[4\] _1388_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__mux2_1
X_6610_ clknet_leaf_8_csclk net1119 net509 VGND VGND VPWR VPWR gpio_configure\[2\]\[12\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_177_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6541_ clknet_2_0__leaf_mgmt_gpio_in[4] _0004_ _0052_ VGND VGND VPWR VPWR hkspi.state\[0\]
+ sky130_fd_sc_hd__dfstp_4
XFILLER_193_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3753_ gpio_configure\[35\]\[8\] _1051_ _1313_ hkspi_disable _1318_ VGND VGND VPWR
+ VPWR _1339_ sky130_fd_sc_hd__a221o_1
XFILLER_146_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6472_ clknet_2_0__leaf_mgmt_gpio_in[4] _0094_ _0050_ VGND VGND VPWR VPWR hkspi.count\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_146_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3684_ gpio_configure\[29\]\[1\] _0917_ net371 gpio_configure\[26\]\[1\] VGND VGND
+ VPWR VPWR _1272_ sky130_fd_sc_hd__a22o_1
X_5423_ net463 net940 _2423_ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__mux2_1
XFILLER_146_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput201 net201 VGND VGND VPWR VPWR mgmt_gpio_oeb[33] sky130_fd_sc_hd__buf_12
Xoutput212 net212 VGND VGND VPWR VPWR mgmt_gpio_oeb[9] sky130_fd_sc_hd__buf_12
Xoutput223 net223 VGND VGND VPWR VPWR mgmt_gpio_out[19] sky130_fd_sc_hd__buf_12
X_5354_ net618 net710 _2415_ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__mux2_1
Xoutput234 net234 VGND VGND VPWR VPWR mgmt_gpio_out[29] sky130_fd_sc_hd__buf_12
Xoutput245 net245 VGND VGND VPWR VPWR mgmt_gpio_out[4] sky130_fd_sc_hd__buf_12
XFILLER_114_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput256 net256 VGND VGND VPWR VPWR pad_flash_io0_ieb sky130_fd_sc_hd__buf_12
Xoutput267 net267 VGND VGND VPWR VPWR pll_div[1] sky130_fd_sc_hd__buf_12
X_4305_ net446 net1112 _1542_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__mux2_1
Xoutput278 net278 VGND VGND VPWR VPWR pll_trim[12] sky130_fd_sc_hd__buf_12
Xoutput289 net289 VGND VGND VPWR VPWR pll_trim[22] sky130_fd_sc_hd__buf_12
X_5285_ net435 net1051 _2407_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__mux2_1
XFILLER_59_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7024_ clknet_leaf_59_csclk net1470 net502 VGND VGND VPWR VPWR gpio_configure\[22\]\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4236_ net465 net622 net592 VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__mux2_1
X_4167_ net2007 _1311_ _1517_ VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__mux2_1
X_4098_ net974 net441 net354 VGND VGND VPWR VPWR _1505_ sky130_fd_sc_hd__mux2_1
XFILLER_43_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_4_csclk clknet_opt_1_0_csclk VGND VGND VPWR VPWR clknet_leaf_4_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6808_ clknet_leaf_57_csclk net925 net503 VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__dfrtp_4
XFILLER_168_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6739_ clknet_leaf_8_csclk net684 net510 VGND VGND VPWR VPWR gpio_configure\[35\]\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_99_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout450 net451 VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__clkbuf_4
Xfanout461 net462 VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__buf_6
XFILLER_171_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout472 _0831_ VGND VGND VPWR VPWR net472 sky130_fd_sc_hd__buf_6
XFILLER_59_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout483 _1427_ VGND VGND VPWR VPWR net483 sky130_fd_sc_hd__clkbuf_16
XFILLER_120_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout494 net496 VGND VGND VPWR VPWR net494 sky130_fd_sc_hd__buf_8
XFILLER_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold909 _0300_ VGND VGND VPWR VPWR net1442 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5070_ _1529_ _2222_ _2241_ VGND VGND VPWR VPWR _2279_ sky130_fd_sc_hd__nor3_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1609 pad_count_1\[2\] VGND VGND VPWR VPWR net2142 sky130_fd_sc_hd__dlygate4sd3_1
X_4021_ net443 net1093 _1474_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__mux2_1
XFILLER_84_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5972_ _1449_ _2793_ VGND VGND VPWR VPWR _2794_ sky130_fd_sc_hd__nand2_2
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4923_ _2127_ _2128_ _2129_ _2133_ VGND VGND VPWR VPWR _2134_ sky130_fd_sc_hd__or4_1
XFILLER_178_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4854_ _1605_ _1684_ _1800_ _1630_ VGND VGND VPWR VPWR _2065_ sky130_fd_sc_hd__o31a_1
X_3805_ hkspi.state\[2\] _1384_ _1386_ hkspi.state\[3\] VGND VGND VPWR VPWR _1387_
+ sky130_fd_sc_hd__a31o_1
XFILLER_178_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4785_ _1598_ _1635_ _1995_ VGND VGND VPWR VPWR _1996_ sky130_fd_sc_hd__a21o_1
X_3736_ gpio_configure\[29\]\[0\] _0917_ _0923_ gpio_configure\[22\]\[0\] VGND VGND
+ VPWR VPWR _1322_ sky130_fd_sc_hd__a22o_1
X_6524_ clknet_leaf_3_csclk net1277 net493 VGND VGND VPWR VPWR gpio_configure\[29\]\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_174_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6455_ clknet_2_0__leaf_mgmt_gpio_in[4] net2093 _0033_ VGND VGND VPWR VPWR hkspi.fixed\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3667_ gpio_configure\[10\]\[1\] _0920_ _1067_ gpio_configure\[23\]\[9\] VGND VGND
+ VPWR VPWR _1255_ sky130_fd_sc_hd__a22o_1
XFILLER_109_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5406_ net457 net780 _2421_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__mux2_1
XFILLER_133_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6386_ _3178_ net2036 _3162_ VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__mux2_1
X_3598_ net67 net351 _1065_ gpio_configure\[37\]\[11\] _1187_ VGND VGND VPWR VPWR
+ _1188_ sky130_fd_sc_hd__a221o_1
XFILLER_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5337_ net440 net1542 _2413_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__mux2_1
XFILLER_142_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5268_ _0908_ net646 VGND VGND VPWR VPWR _2406_ sky130_fd_sc_hd__nand2_8
X_4219_ net577 net1926 _1524_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__mux2_1
XFILLER_102_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7007_ clknet_leaf_45_csclk net1211 net526 VGND VGND VPWR VPWR gpio_configure\[20\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_28_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5199_ net660 net708 _2391_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__mux2_1
XFILLER_141_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4570_ net110 net99 net124 net530 VGND VGND VPWR VPWR _1782_ sky130_fd_sc_hd__or4_4
X_3521_ gpio_configure\[9\]\[4\] net368 _0932_ gpio_configure\[35\]\[4\] VGND VGND
+ VPWR VPWR _1112_ sky130_fd_sc_hd__a22o_1
XFILLER_156_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap403 _2795_ VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__buf_8
Xmax_cap414 _2825_ VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__buf_12
Xhold706 _0577_ VGND VGND VPWR VPWR net1239 sky130_fd_sc_hd__dlygate4sd3_1
Xhold717 gpio_configure\[3\]\[12\] VGND VGND VPWR VPWR net1250 sky130_fd_sc_hd__dlygate4sd3_1
Xhold728 _0307_ VGND VGND VPWR VPWR net1261 sky130_fd_sc_hd__dlygate4sd3_1
X_6240_ gpio_configure\[1\]\[8\] _2802_ _2858_ gpio_configure\[24\]\[8\] _3053_ VGND
+ VGND VPWR VPWR _3054_ sky130_fd_sc_hd__a221o_1
Xhold739 gpio_configure\[26\]\[7\] VGND VGND VPWR VPWR net1272 sky130_fd_sc_hd__dlygate4sd3_1
X_3452_ gpio_configure\[23\]\[4\] _0922_ _1042_ gpio_configure\[6\]\[12\] VGND VGND
+ VPWR VPWR _1043_ sky130_fd_sc_hd__a22o_1
XFILLER_170_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6171_ net2042 _2987_ _2486_ VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__mux2_1
XFILLER_131_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3383_ gpio_configure\[31\]\[6\] _0883_ _0911_ gpio_configure\[21\]\[6\] VGND VGND
+ VPWR VPWR _0977_ sky130_fd_sc_hd__a22o_1
X_5122_ _1793_ _1872_ _1637_ _1669_ VGND VGND VPWR VPWR _2330_ sky130_fd_sc_hd__o211a_1
Xhold1406 net319 VGND VGND VPWR VPWR net1939 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1417 _0113_ VGND VGND VPWR VPWR net1950 sky130_fd_sc_hd__dlygate4sd3_1
X_5053_ _1713_ _2153_ _2261_ VGND VGND VPWR VPWR _2262_ sky130_fd_sc_hd__or3b_1
Xhold1428 net340 VGND VGND VPWR VPWR net1961 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1439 _0899_ VGND VGND VPWR VPWR net1972 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4004_ net458 net1726 _1472_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__mux2_1
XFILLER_38_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_665 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5955_ gpio_configure\[10\]\[12\] net421 _2540_ gpio_configure\[12\]\[12\] VGND VGND
+ VPWR VPWR _2778_ sky130_fd_sc_hd__a22o_1
XFILLER_40_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4906_ _1592_ _1778_ _1866_ VGND VGND VPWR VPWR _2117_ sky130_fd_sc_hd__nor3_1
X_5886_ gpio_configure\[5\]\[9\] _2496_ _2532_ gpio_configure\[18\]\[9\] _2711_ VGND
+ VGND VPWR VPWR _2712_ sky130_fd_sc_hd__a221o_1
XFILLER_139_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4837_ _1864_ _2047_ _1605_ VGND VGND VPWR VPWR _2048_ sky130_fd_sc_hd__a21o_1
XFILLER_178_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4768_ _1584_ _1667_ _1960_ _1961_ _1979_ VGND VGND VPWR VPWR _1980_ sky130_fd_sc_hd__a2111o_1
XFILLER_107_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6507_ clknet_leaf_2_csclk net1468 net492 VGND VGND VPWR VPWR gpio_configure\[23\]\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_134_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3719_ gpio_configure\[21\]\[1\] _0911_ _1062_ gpio_configure\[21\]\[9\] VGND VGND
+ VPWR VPWR _1307_ sky130_fd_sc_hd__a22o_1
XFILLER_106_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4699_ _1894_ _1895_ _1896_ _1910_ VGND VGND VPWR VPWR _1911_ sky130_fd_sc_hd__and4_1
XFILLER_134_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6438_ net495 net482 VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__and2_1
XFILLER_106_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6369_ wbbd_state\[7\] net141 net133 wbbd_state\[8\] VGND VGND VPWR VPWR _3167_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_22_csclk clknet_3_4_0_csclk VGND VGND VPWR VPWR clknet_leaf_22_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold11 hkspi.wrstb VGND VGND VPWR VPWR net544 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold22 _0913_ VGND VGND VPWR VPWR net555 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold33 _0478_ VGND VGND VPWR VPWR net566 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold44 net460 VGND VGND VPWR VPWR net577 sky130_fd_sc_hd__buf_4
Xhold55 _0859_ VGND VGND VPWR VPWR net588 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 _0856_ VGND VGND VPWR VPWR net599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 _0927_ VGND VGND VPWR VPWR net610 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 _0289_ VGND VGND VPWR VPWR net621 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 wbbd_data\[6\] VGND VGND VPWR VPWR net632 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_37_csclk clknet_3_7_0_csclk VGND VGND VPWR VPWR clknet_leaf_37_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_16_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_mgmt_gpio_in[4] mgmt_gpio_in[4] VGND VGND VPWR VPWR clknet_0_mgmt_gpio_in[4]
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_8 _0915_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_719 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_270 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5740_ _2566_ _2568_ _2570_ _2572_ VGND VGND VPWR VPWR _2573_ sky130_fd_sc_hd__or4_1
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5671_ pad_count_1\[4\] _2461_ _2504_ VGND VGND VPWR VPWR _2506_ sky130_fd_sc_hd__and3_4
XFILLER_188_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4622_ _1833_ VGND VGND VPWR VPWR _1834_ sky130_fd_sc_hd__inv_2
XFILLER_128_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4553_ net128 _1751_ VGND VGND VPWR VPWR _1765_ sky130_fd_sc_hd__nor2_1
XFILLER_190_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold503 _0362_ VGND VGND VPWR VPWR net1036 sky130_fd_sc_hd__dlygate4sd3_1
Xhold514 gpio_configure\[13\]\[7\] VGND VGND VPWR VPWR net1047 sky130_fd_sc_hd__dlygate4sd3_1
X_3504_ net554 _0973_ VGND VGND VPWR VPWR _1095_ sky130_fd_sc_hd__nor2_8
Xhold525 _0492_ VGND VGND VPWR VPWR net1058 sky130_fd_sc_hd__dlygate4sd3_1
Xhold536 gpio_configure\[7\]\[7\] VGND VGND VPWR VPWR net1069 sky130_fd_sc_hd__dlygate4sd3_1
X_4484_ _1609_ _1679_ _1563_ VGND VGND VPWR VPWR _1696_ sky130_fd_sc_hd__or3b_1
Xhold547 _0217_ VGND VGND VPWR VPWR net1080 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold558 gpio_configure\[4\]\[12\] VGND VGND VPWR VPWR net1091 sky130_fd_sc_hd__dlygate4sd3_1
X_6223_ gpio_configure\[30\]\[8\] _2799_ net408 gpio_configure\[35\]\[8\] VGND VGND
+ VPWR VPWR _3037_ sky130_fd_sc_hd__a22o_1
XFILLER_116_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold569 gpio_configure\[13\]\[5\] VGND VGND VPWR VPWR net1102 sky130_fd_sc_hd__dlygate4sd3_1
X_3435_ gpio_configure\[16\]\[5\] _0912_ _0915_ gpio_configure\[3\]\[5\] _1026_ VGND
+ VGND VPWR VPWR _1027_ sky130_fd_sc_hd__a221o_1
XFILLER_171_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6154_ gpio_configure\[14\]\[5\] net411 net406 gpio_configure\[27\]\[5\] VGND VGND
+ VPWR VPWR _2971_ sky130_fd_sc_hd__a22o_1
X_3366_ gpio_configure\[2\]\[7\] _0908_ _0940_ net281 _0961_ VGND VGND VPWR VPWR _0962_
+ sky130_fd_sc_hd__a221o_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1203 gpio_configure\[9\]\[9\] VGND VGND VPWR VPWR net1736 sky130_fd_sc_hd__dlygate4sd3_1
X_5105_ _1689_ _1750_ _1778_ _1693_ _1870_ VGND VGND VPWR VPWR _2313_ sky130_fd_sc_hd__o221a_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1214 _0155_ VGND VGND VPWR VPWR net1747 sky130_fd_sc_hd__dlygate4sd3_1
X_6085_ _2895_ _2904_ VGND VGND VPWR VPWR _2905_ sky130_fd_sc_hd__or2_2
XFILLER_58_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3297_ net627 net638 net551 VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__or3b_4
Xhold1225 _0469_ VGND VGND VPWR VPWR net1758 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1236 gpio_configure\[22\]\[8\] VGND VGND VPWR VPWR net1769 sky130_fd_sc_hd__dlygate4sd3_1
X_5036_ _1750_ _2203_ VGND VGND VPWR VPWR _2245_ sky130_fd_sc_hd__nand2_1
Xhold1247 _0324_ VGND VGND VPWR VPWR net1780 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1258 net1976 VGND VGND VPWR VPWR net1791 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1269 gpio_configure\[15\]\[8\] VGND VGND VPWR VPWR net1802 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6987_ clknet_leaf_25_csclk net1398 net518 VGND VGND VPWR VPWR gpio_configure\[18\]\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_179_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5938_ gpio_configure\[16\]\[11\] net472 VGND VGND VPWR VPWR _2762_ sky130_fd_sc_hd__or2_1
XFILLER_179_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5869_ _2689_ _2691_ _2693_ _2695_ VGND VGND VPWR VPWR _2696_ sky130_fd_sc_hd__or4_1
XFILLER_139_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput101 wb_adr_i[11] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_1
XFILLER_103_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput112 wb_adr_i[21] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_1
XFILLER_163_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput123 wb_adr_i[31] VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_1
Xinput134 wb_dat_i[11] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_1
Xinput145 wb_dat_i[21] VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput156 wb_dat_i[31] VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_1
Xinput167 wb_sel_i[2] VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3220_ gpio_configure\[14\]\[3\] VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__inv_2
XFILLER_97_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6910_ clknet_leaf_15_csclk net1167 net513 VGND VGND VPWR VPWR gpio_configure\[8\]\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6841_ clknet_leaf_36_csclk net615 net522 VGND VGND VPWR VPWR mgmt_gpio_data_buf\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_62_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6772_ clknet_leaf_70_csclk net1406 net501 VGND VGND VPWR VPWR gpio_configure\[22\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_3984_ net1832 net467 _1470_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__mux2_1
XFILLER_50_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5723_ gpio_configure\[21\]\[1\] _2521_ _2538_ gpio_configure\[1\]\[1\] _2556_ VGND
+ VGND VPWR VPWR _2557_ sky130_fd_sc_hd__a221o_1
XFILLER_188_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5654_ pad_count_1\[0\] pad_count_1\[1\] VGND VGND VPWR VPWR _2489_ sky130_fd_sc_hd__and2b_2
X_4605_ net126 _0836_ _1750_ VGND VGND VPWR VPWR _1817_ sky130_fd_sc_hd__or3_1
XFILLER_117_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5585_ net618 net698 net603 VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__mux2_1
XFILLER_163_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold300 _0350_ VGND VGND VPWR VPWR net833 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold311 gpio_configure\[16\]\[6\] VGND VGND VPWR VPWR net844 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_191_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4536_ _1704_ _1705_ _1743_ _1747_ _1582_ VGND VGND VPWR VPWR _1748_ sky130_fd_sc_hd__a41oi_1
Xhold322 _0408_ VGND VGND VPWR VPWR net855 sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 gpio_configure\[5\]\[9\] VGND VGND VPWR VPWR net866 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold344 _0330_ VGND VGND VPWR VPWR net877 sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 serial_bb_enable VGND VGND VPWR VPWR net888 sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 _0272_ VGND VGND VPWR VPWR net899 sky130_fd_sc_hd__dlygate4sd3_1
X_4467_ _1434_ _1435_ _1600_ VGND VGND VPWR VPWR _1679_ sky130_fd_sc_hd__or3_2
Xhold377 gpio_configure\[12\]\[12\] VGND VGND VPWR VPWR net910 sky130_fd_sc_hd__dlygate4sd3_1
Xhold388 _0281_ VGND VGND VPWR VPWR net921 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6206_ gpio_configure\[16\]\[7\] _2831_ net391 gpio_configure\[17\]\[7\] _3020_ VGND
+ VGND VPWR VPWR _3021_ sky130_fd_sc_hd__a221o_1
Xhold399 net237 VGND VGND VPWR VPWR net932 sky130_fd_sc_hd__dlygate4sd3_1
X_3418_ gpio_configure\[13\]\[5\] _0906_ net355 gpio_configure\[5\]\[5\] VGND VGND
+ VPWR VPWR _1010_ sky130_fd_sc_hd__a22o_1
X_7186_ clknet_3_1_0_wb_clk_i _0788_ net490 VGND VGND VPWR VPWR serial_data_staging_2\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_4398_ net110 net124 net530 VGND VGND VPWR VPWR _1610_ sky130_fd_sc_hd__and3_4
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3349_ gpio_configure\[31\]\[7\] net375 _0900_ net33 VGND VGND VPWR VPWR _0945_ sky130_fd_sc_hd__a22o_1
XFILLER_98_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6137_ gpio_configure\[10\]\[4\] _2825_ net394 gpio_configure\[6\]\[4\] _2954_ VGND
+ VGND VPWR VPWR _2955_ sky130_fd_sc_hd__a221o_1
Xhold1000 _0743_ VGND VGND VPWR VPWR net1533 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1011 gpio_configure\[16\]\[5\] VGND VGND VPWR VPWR net1544 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1022 _0586_ VGND VGND VPWR VPWR net1555 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1033 gpio_configure\[35\]\[0\] VGND VGND VPWR VPWR net1566 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1044 _0407_ VGND VGND VPWR VPWR net1577 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6068_ _2883_ _2885_ _2886_ _2888_ VGND VGND VPWR VPWR _2889_ sky130_fd_sc_hd__or4_1
Xhold1055 gpio_configure\[5\]\[2\] VGND VGND VPWR VPWR net1588 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1066 _0677_ VGND VGND VPWR VPWR net1599 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1077 net2048 VGND VGND VPWR VPWR net1610 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1088 gpio_configure\[26\]\[8\] VGND VGND VPWR VPWR net1621 sky130_fd_sc_hd__dlygate4sd3_1
X_5019_ _1828_ _2225_ _2227_ _2228_ VGND VGND VPWR VPWR _2229_ sky130_fd_sc_hd__or4_1
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1099 gpio_configure\[19\]\[10\] VGND VGND VPWR VPWR net1632 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_206 _2816_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_217 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_228 net412 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_239 net569 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5370_ net458 net1740 _2417_ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__mux2_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4321_ net1729 net455 _1545_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__mux2_1
XFILLER_113_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7040_ clknet_leaf_58_csclk net1444 net503 VGND VGND VPWR VPWR gpio_configure\[24\]\[6\]
+ sky130_fd_sc_hd__dfrtp_2
X_4252_ _1102_ net426 VGND VGND VPWR VPWR _1534_ sky130_fd_sc_hd__and2_2
XFILLER_113_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3203_ gpio_configure\[31\]\[3\] VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__inv_2
X_4183_ net2080 _1249_ _1519_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__mux2_1
XFILLER_55_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6824_ clknet_leaf_71_csclk net1611 net491 VGND VGND VPWR VPWR irq_1_inputsrc sky130_fd_sc_hd__dfrtp_1
X_6755_ clknet_leaf_6_csclk net1301 net497 VGND VGND VPWR VPWR gpio_configure\[20\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_3967_ net58 net1097 net669 VGND VGND VPWR VPWR _1462_ sky130_fd_sc_hd__mux2_8
X_5706_ pad_count_1\[4\] _2461_ _2493_ VGND VGND VPWR VPWR _2541_ sky130_fd_sc_hd__and3_4
XFILLER_148_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6686_ clknet_leaf_5_csclk net1774 net494 VGND VGND VPWR VPWR gpio_configure\[13\]\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_3898_ xfer_count\[0\] xfer_count\[1\] VGND VGND VPWR VPWR _1444_ sky130_fd_sc_hd__nor2_1
XFILLER_109_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5637_ pad_count_2\[4\] _2470_ _2473_ VGND VGND VPWR VPWR _2476_ sky130_fd_sc_hd__and3_1
XFILLER_148_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5568_ net440 net1520 net648 VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__mux2_1
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold130 _0180_ VGND VGND VPWR VPWR net663 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_191_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold141 _0109_ VGND VGND VPWR VPWR net674 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_163_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4519_ _1643_ _1653_ _1727_ _1728_ _1730_ VGND VGND VPWR VPWR _1731_ sky130_fd_sc_hd__o2111a_1
Xhold152 mgmt_gpio_data_buf\[12\] VGND VGND VPWR VPWR net685 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold163 gpio_configure\[34\]\[11\] VGND VGND VPWR VPWR net696 sky130_fd_sc_hd__dlygate4sd3_1
X_5499_ net440 net1536 net641 VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__mux2_1
Xhold174 _0192_ VGND VGND VPWR VPWR net707 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold185 gpio_configure\[36\]\[11\] VGND VGND VPWR VPWR net718 sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 _0528_ VGND VGND VPWR VPWR net729 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7169_ clknet_3_2_0_wb_clk_i _0771_ net498 VGND VGND VPWR VPWR serial_data_staging_1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4870_ _1642_ _1706_ VGND VGND VPWR VPWR _2081_ sky130_fd_sc_hd__nor2_1
XTAP_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3821_ _0845_ _0844_ _1390_ VGND VGND VPWR VPWR _1400_ sky130_fd_sc_hd__mux2_1
XFILLER_32_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6540_ clknet_leaf_1_csclk net1199 net493 VGND VGND VPWR VPWR gpio_configure\[26\]\[12\]
+ sky130_fd_sc_hd__dfrtp_2
X_3752_ gpio_configure\[7\]\[8\] _1094_ _1319_ VGND VGND VPWR VPWR _1338_ sky130_fd_sc_hd__a21o_1
XFILLER_146_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6471_ clknet_2_1__leaf_mgmt_gpio_in[4] _0093_ _0049_ VGND VGND VPWR VPWR hkspi.count\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_185_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3683_ gpio_configure\[6\]\[9\] _1042_ _1117_ net267 _1270_ VGND VGND VPWR VPWR _1271_
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5422_ net469 net1724 _2423_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__mux2_1
Xoutput202 net202 VGND VGND VPWR VPWR mgmt_gpio_oeb[34] sky130_fd_sc_hd__buf_12
Xoutput213 net213 VGND VGND VPWR VPWR mgmt_gpio_out[0] sky130_fd_sc_hd__buf_12
Xoutput224 net224 VGND VGND VPWR VPWR mgmt_gpio_out[1] sky130_fd_sc_hd__buf_12
Xoutput235 net235 VGND VGND VPWR VPWR mgmt_gpio_out[2] sky130_fd_sc_hd__buf_12
X_5353_ net453 net1242 _2415_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__mux2_1
Xoutput246 net246 VGND VGND VPWR VPWR mgmt_gpio_out[5] sky130_fd_sc_hd__buf_12
Xoutput257 net257 VGND VGND VPWR VPWR pad_flash_io0_oeb sky130_fd_sc_hd__buf_12
XFILLER_160_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput268 net268 VGND VGND VPWR VPWR pll_div[2] sky130_fd_sc_hd__buf_12
X_4304_ net569 net696 _1542_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__mux2_1
Xoutput279 net279 VGND VGND VPWR VPWR pll_trim[13] sky130_fd_sc_hd__buf_12
X_5284_ net439 net756 _2407_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__mux2_1
XFILLER_99_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7023_ clknet_leaf_59_csclk net825 net502 VGND VGND VPWR VPWR gpio_configure\[22\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_99_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4235_ net470 net1497 net592 VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__mux2_1
XFILLER_102_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4166_ net1953 _1376_ _1517_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__mux2_1
XFILLER_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4097_ net912 _1504_ _1499_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__mux2_1
XFILLER_36_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6807_ clknet_leaf_58_csclk net1705 net503 VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__dfrtp_4
XFILLER_168_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4999_ net478 _1596_ VGND VGND VPWR VPWR _2209_ sky130_fd_sc_hd__nand2_1
XFILLER_139_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6738_ clknet_leaf_18_csclk net787 net510 VGND VGND VPWR VPWR gpio_configure\[35\]\[10\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_23_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6669_ clknet_leaf_4_csclk net897 net494 VGND VGND VPWR VPWR gpio_configure\[9\]\[12\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_109_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout440 net441 VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__buf_4
XFILLER_48_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout451 net568 VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__buf_8
XFILLER_120_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout462 net463 VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__buf_6
XFILLER_171_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout473 _0824_ VGND VGND VPWR VPWR net473 sky130_fd_sc_hd__buf_12
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout484 net487 VGND VGND VPWR VPWR net484 sky130_fd_sc_hd__buf_6
XFILLER_59_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout495 net496 VGND VGND VPWR VPWR net495 sky130_fd_sc_hd__buf_4
XFILLER_58_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4020_ net449 net1150 _1474_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__mux2_1
XFILLER_96_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5971_ pad_count_2\[1\] pad_count_2\[0\] VGND VGND VPWR VPWR _2793_ sky130_fd_sc_hd__nor2_2
XFILLER_64_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4922_ _1837_ _2132_ _1867_ _2131_ VGND VGND VPWR VPWR _2133_ sky130_fd_sc_hd__or4b_1
XFILLER_45_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4853_ _1757_ _1863_ _1659_ VGND VGND VPWR VPWR _2064_ sky130_fd_sc_hd__o21a_1
XFILLER_193_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3804_ hkspi.fixed\[2\] hkspi.fixed\[1\] hkspi.fixed\[0\] VGND VGND VPWR VPWR _1386_
+ sky130_fd_sc_hd__or3b_1
X_4784_ _1777_ _1795_ VGND VGND VPWR VPWR _1995_ sky130_fd_sc_hd__nor2_1
XFILLER_119_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_opt_2_0_csclk clknet_3_4_0_csclk VGND VGND VPWR VPWR clknet_opt_2_0_csclk
+ sky130_fd_sc_hd__clkbuf_16
X_6523_ clknet_leaf_2_csclk net1364 net492 VGND VGND VPWR VPWR gpio_configure\[29\]\[10\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_20_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3735_ net299 _0940_ net305 _1317_ VGND VGND VPWR VPWR _1321_ sky130_fd_sc_hd__a22o_1
XFILLER_146_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6454_ clknet_2_1__leaf_mgmt_gpio_in[4] _0076_ _0032_ VGND VGND VPWR VPWR hkspi.fixed\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_118_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3666_ gpio_configure\[13\]\[1\] _0906_ _0921_ gpio_configure\[12\]\[1\] _1253_ VGND
+ VGND VPWR VPWR _1254_ sky130_fd_sc_hd__a221o_1
XFILLER_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5405_ net465 net868 _2421_ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__mux2_1
XFILLER_134_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6385_ wbbd_state\[7\] net147 net161 net433 _3177_ VGND VGND VPWR VPWR _3178_ sky130_fd_sc_hd__a221o_1
X_3597_ gpio_configure\[36\]\[3\] net352 _1122_ gpio_configure\[8\]\[11\] VGND VGND
+ VPWR VPWR _1187_ sky130_fd_sc_hd__a22o_1
XFILLER_133_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5336_ net447 net1174 _2413_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__mux2_1
XFILLER_0_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5267_ net435 net1043 _2405_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__mux2_1
X_7006_ clknet_leaf_20_csclk net1183 net514 VGND VGND VPWR VPWR gpio_configure\[20\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_4218_ net462 net1427 _1524_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__mux2_1
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5198_ net443 net1085 _2391_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__mux2_1
X_4149_ net461 net1672 _1514_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__mux2_1
XFILLER_16_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3520_ gpio_configure\[36\]\[12\] _1109_ _1110_ gpio_configure\[2\]\[12\] VGND VGND
+ VPWR VPWR _1111_ sky130_fd_sc_hd__a22o_1
Xmax_cap404 _2862_ VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__buf_8
XFILLER_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap415 _2814_ VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__buf_12
Xhold707 gpio_configure\[21\]\[4\] VGND VGND VPWR VPWR net1240 sky130_fd_sc_hd__dlygate4sd3_1
Xhold718 _0228_ VGND VGND VPWR VPWR net1251 sky130_fd_sc_hd__dlygate4sd3_1
Xhold729 gpio_configure\[32\]\[7\] VGND VGND VPWR VPWR net1262 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3451_ net554 _1006_ VGND VGND VPWR VPWR _1042_ sky130_fd_sc_hd__nor2_8
XFILLER_143_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3382_ net289 _0886_ _0924_ gpio_configure\[26\]\[6\] VGND VGND VPWR VPWR _0976_
+ sky130_fd_sc_hd__a22o_1
X_6170_ xfer_state\[1\] serial_data_staging_2\[4\] _2986_ VGND VGND VPWR VPWR _2987_
+ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_3_csclk clknet_3_1_0_csclk VGND VGND VPWR VPWR clknet_leaf_3_csclk sky130_fd_sc_hd__clkbuf_16
X_5121_ _2320_ _2328_ VGND VGND VPWR VPWR _2329_ sky130_fd_sc_hd__and2b_1
XFILLER_69_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1407 net345 VGND VGND VPWR VPWR net1940 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1418 net344 VGND VGND VPWR VPWR net1951 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5052_ _1606_ net432 _1822_ _1873_ VGND VGND VPWR VPWR _2261_ sky130_fd_sc_hd__o22a_1
Xhold1429 net335 VGND VGND VPWR VPWR net1962 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4003_ net464 net1431 _1472_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__mux2_1
XFILLER_65_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5954_ gpio_configure\[18\]\[12\] _2532_ _2776_ VGND VGND VPWR VPWR _2777_ sky130_fd_sc_hd__a21o_1
XFILLER_80_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4905_ _2112_ _2115_ VGND VGND VPWR VPWR _2116_ sky130_fd_sc_hd__nand2_1
XFILLER_21_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5885_ gpio_configure\[28\]\[9\] _2513_ _2517_ gpio_configure\[30\]\[9\] VGND VGND
+ VPWR VPWR _2711_ sky130_fd_sc_hd__a22o_1
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4836_ _1641_ _1670_ VGND VGND VPWR VPWR _2047_ sky130_fd_sc_hd__nand2_1
XFILLER_178_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4767_ _1584_ _1666_ _1948_ _1962_ _1978_ VGND VGND VPWR VPWR _1979_ sky130_fd_sc_hd__a2111o_1
X_6506_ clknet_leaf_78_csclk net1831 net486 VGND VGND VPWR VPWR gpio_configure\[23\]\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_3718_ gpio_configure\[35\]\[1\] _0932_ _1007_ net62 _1305_ VGND VGND VPWR VPWR _1306_
+ sky130_fd_sc_hd__a221o_1
XFILLER_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4698_ _1881_ _1905_ _1907_ _1909_ VGND VGND VPWR VPWR _1910_ sky130_fd_sc_hd__and4b_1
XFILLER_106_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6437_ net495 net482 VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__and2_1
X_3649_ gpio_configure\[31\]\[2\] net375 _1137_ net97 VGND VGND VPWR VPWR _1238_ sky130_fd_sc_hd__a22o_1
XFILLER_136_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6368_ _3166_ net2059 _3162_ VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__mux2_1
XFILLER_0_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5319_ net440 net1552 net556 VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__mux2_1
XFILLER_130_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6299_ gpio_configure\[30\]\[11\] _2799_ net408 gpio_configure\[35\]\[11\] VGND VGND
+ VPWR VPWR _3110_ sky130_fd_sc_hd__a22o_1
Xhold12 net476 VGND VGND VPWR VPWR net545 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold23 _2411_ VGND VGND VPWR VPWR net556 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold34 hkspi.odata\[3\] VGND VGND VPWR VPWR net567 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 _0285_ VGND VGND VPWR VPWR net578 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 _0862_ VGND VGND VPWR VPWR net589 sky130_fd_sc_hd__buf_6
Xhold67 _0869_ VGND VGND VPWR VPWR net600 sky130_fd_sc_hd__buf_6
Xhold78 net369 VGND VGND VPWR VPWR net611 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold89 gpio_configure\[12\]\[9\] VGND VGND VPWR VPWR net622 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_9 _0919_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5670_ net472 _2461_ _2504_ VGND VGND VPWR VPWR _2505_ sky130_fd_sc_hd__and3_4
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4621_ _0835_ net125 _1755_ VGND VGND VPWR VPWR _1833_ sky130_fd_sc_hd__or3_4
XFILLER_175_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4552_ _1751_ _1763_ VGND VGND VPWR VPWR _1764_ sky130_fd_sc_hd__nor2_1
XFILLER_116_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold504 gpio_configure\[11\]\[7\] VGND VGND VPWR VPWR net1037 sky130_fd_sc_hd__dlygate4sd3_1
X_3503_ net376 _0903_ VGND VGND VPWR VPWR _1094_ sky130_fd_sc_hd__nor2_4
Xhold515 _0556_ VGND VGND VPWR VPWR net1048 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold526 net294 VGND VGND VPWR VPWR net1059 sky130_fd_sc_hd__dlygate4sd3_1
X_4483_ _1694_ VGND VGND VPWR VPWR _1695_ sky130_fd_sc_hd__inv_2
Xhold537 _0508_ VGND VGND VPWR VPWR net1070 sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 gpio_configure\[19\]\[11\] VGND VGND VPWR VPWR net1081 sky130_fd_sc_hd__dlygate4sd3_1
X_6222_ gpio_configure\[28\]\[8\] _2861_ VGND VGND VPWR VPWR _3036_ sky130_fd_sc_hd__and2_1
XFILLER_131_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold559 _0233_ VGND VGND VPWR VPWR net1092 sky130_fd_sc_hd__dlygate4sd3_1
X_3434_ gpio_configure\[30\]\[5\] _0892_ _0907_ gpio_configure\[11\]\[5\] VGND VGND
+ VPWR VPWR _1026_ sky130_fd_sc_hd__a22o_1
XFILLER_171_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6153_ gpio_configure\[18\]\[5\] net399 net410 gpio_configure\[8\]\[5\] _2969_ VGND
+ VGND VPWR VPWR _2970_ sky130_fd_sc_hd__a221o_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3365_ gpio_configure\[13\]\[7\] _0906_ _0920_ gpio_configure\[10\]\[7\] VGND VGND
+ VPWR VPWR _0961_ sky130_fd_sc_hd__a22o_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5104_ _2260_ _2278_ _2297_ _2312_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__or4_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1204 _0279_ VGND VGND VPWR VPWR net1737 sky130_fd_sc_hd__dlygate4sd3_1
X_6084_ _2897_ _2899_ _2901_ _2903_ VGND VGND VPWR VPWR _2904_ sky130_fd_sc_hd__or4_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3296_ _0870_ net388 VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__nor2_8
Xhold1215 net1979 VGND VGND VPWR VPWR net1748 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1226 mgmt_gpio_data\[8\] VGND VGND VPWR VPWR net1759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1237 _0374_ VGND VGND VPWR VPWR net1770 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1248 gpio_configure\[18\]\[0\] VGND VGND VPWR VPWR net1781 sky130_fd_sc_hd__dlygate4sd3_1
X_5035_ _1597_ _1671_ VGND VGND VPWR VPWR _2244_ sky130_fd_sc_hd__nand2_1
Xhold1259 gpio_configure\[22\]\[0\] VGND VGND VPWR VPWR net1792 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6986_ clknet_leaf_70_csclk net1782 net491 VGND VGND VPWR VPWR gpio_configure\[18\]\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_25_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5937_ gpio_configure\[6\]\[11\] _2490_ _2528_ gpio_configure\[7\]\[11\] _2760_ VGND
+ VGND VPWR VPWR _2761_ sky130_fd_sc_hd__a221o_1
XFILLER_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5868_ gpio_configure\[11\]\[8\] _2505_ _2511_ gpio_configure\[25\]\[8\] _2694_ VGND
+ VGND VPWR VPWR _2695_ sky130_fd_sc_hd__a221o_1
XFILLER_179_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4819_ _1756_ _1785_ _1554_ _1749_ VGND VGND VPWR VPWR _2030_ sky130_fd_sc_hd__and4bb_1
XFILLER_166_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5799_ gpio_configure\[20\]\[5\] _2499_ _2517_ gpio_configure\[30\]\[5\] _2628_ VGND
+ VGND VPWR VPWR _2629_ sky130_fd_sc_hd__a221o_1
XFILLER_119_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput102 wb_adr_i[12] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_1
Xinput113 wb_adr_i[22] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_130_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput124 wb_adr_i[3] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_16
Xinput135 wb_dat_i[12] VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_1
XFILLER_193_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput146 wb_dat_i[22] VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput157 wb_dat_i[3] VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_1
Xinput168 wb_sel_i[3] VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6840_ clknet_leaf_32_csclk net657 net524 VGND VGND VPWR VPWR mgmt_gpio_data_buf\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_63_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6771_ clknet_leaf_71_csclk net1770 net491 VGND VGND VPWR VPWR gpio_configure\[22\]\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_3983_ _0940_ net425 VGND VGND VPWR VPWR _1470_ sky130_fd_sc_hd__and2_2
XFILLER_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5722_ gpio_configure\[25\]\[1\] net420 net419 gpio_configure\[16\]\[1\] _2525_ VGND
+ VGND VPWR VPWR _2556_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_21_csclk clknet_3_4_0_csclk VGND VGND VPWR VPWR clknet_leaf_21_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_31_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5653_ pad_count_1\[3\] pad_count_1\[2\] VGND VGND VPWR VPWR _2488_ sky130_fd_sc_hd__and2b_2
XFILLER_176_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4604_ net125 _1749_ _0835_ VGND VGND VPWR VPWR _1816_ sky130_fd_sc_hd__a21o_1
X_5584_ net452 net980 net603 VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__mux2_1
XFILLER_175_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_36_csclk clknet_3_7_0_csclk VGND VGND VPWR VPWR clknet_leaf_36_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_163_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold301 net2145 VGND VGND VPWR VPWR net834 sky130_fd_sc_hd__dlygate4sd3_1
X_4535_ _1576_ _1745_ VGND VGND VPWR VPWR _1747_ sky130_fd_sc_hd__or2_1
Xhold312 _0579_ VGND VGND VPWR VPWR net845 sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 gpio_configure\[37\]\[2\] VGND VGND VPWR VPWR net856 sky130_fd_sc_hd__dlygate4sd3_1
Xhold334 _0235_ VGND VGND VPWR VPWR net867 sky130_fd_sc_hd__dlygate4sd3_1
Xhold345 gpio_configure\[6\]\[1\] VGND VGND VPWR VPWR net878 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold356 _0421_ VGND VGND VPWR VPWR net889 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4466_ _0834_ net479 VGND VGND VPWR VPWR _1678_ sky130_fd_sc_hd__nand2_8
Xhold367 gpio_configure\[4\]\[9\] VGND VGND VPWR VPWR net900 sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 _0298_ VGND VGND VPWR VPWR net911 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6205_ gpio_configure\[14\]\[7\] net411 net406 gpio_configure\[27\]\[7\] VGND VGND
+ VPWR VPWR _3020_ sky130_fd_sc_hd__a22o_1
XFILLER_171_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold389 gpio_configure\[21\]\[7\] VGND VGND VPWR VPWR net922 sky130_fd_sc_hd__dlygate4sd3_1
X_3417_ net383 _1008_ VGND VGND VPWR VPWR _1009_ sky130_fd_sc_hd__nor2_8
X_7185_ clknet_3_1_0_wb_clk_i _0787_ net490 VGND VGND VPWR VPWR serial_data_staging_2\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_4397_ _1580_ _1591_ VGND VGND VPWR VPWR _1609_ sky130_fd_sc_hd__nand2_1
XFILLER_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6136_ gpio_configure\[9\]\[4\] net412 net409 gpio_configure\[12\]\[4\] VGND VGND
+ VPWR VPWR _2954_ sky130_fd_sc_hd__a22o_1
X_3348_ gpio_configure\[18\]\[7\] net374 _0924_ gpio_configure\[26\]\[7\] _0943_ VGND
+ VGND VPWR VPWR _0944_ sky130_fd_sc_hd__a221o_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1001 gpio_configure\[15\]\[5\] VGND VGND VPWR VPWR net1534 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_133_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1012 _0578_ VGND VGND VPWR VPWR net1545 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1023 gpio_configure\[26\]\[5\] VGND VGND VPWR VPWR net1556 sky130_fd_sc_hd__dlygate4sd3_1
X_6067_ gpio_configure\[3\]\[1\] net413 net407 gpio_configure\[15\]\[1\] _2887_ VGND
+ VGND VPWR VPWR _2888_ sky130_fd_sc_hd__a221o_1
Xhold1034 _0722_ VGND VGND VPWR VPWR net1567 sky130_fd_sc_hd__dlygate4sd3_1
X_3279_ net581 net552 VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__or2_2
Xhold1045 gpio_configure\[12\]\[2\] VGND VGND VPWR VPWR net1578 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1056 _0487_ VGND VGND VPWR VPWR net1589 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1067 net271 VGND VGND VPWR VPWR net1600 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5018_ _1590_ _1778_ _1797_ VGND VGND VPWR VPWR _2228_ sky130_fd_sc_hd__nor3_1
Xhold1078 _0427_ VGND VGND VPWR VPWR net1611 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1089 _0158_ VGND VGND VPWR VPWR net1622 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_207 _2825_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_218 net263 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_229 net439 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6969_ clknet_leaf_54_csclk net1135 net506 VGND VGND VPWR VPWR gpio_configure\[15\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_186_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold890 gpio_configure\[26\]\[6\] VGND VGND VPWR VPWR net1423 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_95_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1590 serial_data_staging_1\[7\] VGND VGND VPWR VPWR net2123 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4320_ net1734 net461 _1545_ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__mux2_1
XFILLER_160_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4251_ net444 net1310 _1533_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__mux2_1
X_3202_ gpio_configure\[32\]\[3\] VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__inv_2
XFILLER_113_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4182_ net2046 _1311_ _1519_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__mux2_1
XFILLER_79_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6823_ clknet_leaf_29_csclk net1513 net520 VGND VGND VPWR VPWR trap_output_dest sky130_fd_sc_hd__dfrtp_4
XFILLER_168_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6754_ clknet_leaf_6_csclk net1253 net497 VGND VGND VPWR VPWR gpio_configure\[20\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_3966_ _0886_ net427 VGND VGND VPWR VPWR _1461_ sky130_fd_sc_hd__and2_2
X_5705_ net472 _2459_ _2493_ VGND VGND VPWR VPWR _2540_ sky130_fd_sc_hd__and3_4
X_6685_ clknet_leaf_4_csclk net911 net511 VGND VGND VPWR VPWR gpio_configure\[12\]\[12\]
+ sky130_fd_sc_hd__dfrtp_2
X_3897_ _0822_ serial_xfer _1443_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__o21ai_1
XFILLER_176_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5636_ net2141 _2463_ _2474_ _2475_ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__a31o_1
XFILLER_164_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5567_ net447 net1188 net648 VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__mux2_1
Xhold120 _0628_ VGND VGND VPWR VPWR net653 sky130_fd_sc_hd__dlygate4sd3_1
X_4518_ _1729_ VGND VGND VPWR VPWR _1730_ sky130_fd_sc_hd__inv_2
Xhold131 wbbd_data\[5\] VGND VGND VPWR VPWR net664 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold142 gpio_configure\[29\]\[4\] VGND VGND VPWR VPWR net675 sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 _0441_ VGND VGND VPWR VPWR net686 sky130_fd_sc_hd__dlygate4sd3_1
X_5498_ net618 net654 net641 VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__mux2_1
XFILLER_132_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold164 _0352_ VGND VGND VPWR VPWR net697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 net263 VGND VGND VPWR VPWR net708 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold186 _0332_ VGND VGND VPWR VPWR net719 sky130_fd_sc_hd__dlygate4sd3_1
X_4449_ _1605_ _1612_ _1641_ VGND VGND VPWR VPWR _1661_ sky130_fd_sc_hd__and3b_1
XFILLER_104_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold197 mgmt_gpio_data_buf\[11\] VGND VGND VPWR VPWR net730 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7168_ clknet_3_2_0_wb_clk_i net2018 net502 VGND VGND VPWR VPWR serial_data_staging_1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6119_ net362 _2931_ _2933_ _2937_ VGND VGND VPWR VPWR _2938_ sky130_fd_sc_hd__or4_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7099_ clknet_leaf_62_csclk net793 net501 VGND VGND VPWR VPWR gpio_configure\[32\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3820_ hkspi.state\[3\] _1389_ VGND VGND VPWR VPWR _1399_ sky130_fd_sc_hd__nor2_1
XFILLER_177_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3751_ net71 net353 net351 net36 _1336_ VGND VGND VPWR VPWR _1337_ sky130_fd_sc_hd__a221o_1
XFILLER_32_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6470_ clknet_2_1__leaf_mgmt_gpio_in[4] _0092_ _0048_ VGND VGND VPWR VPWR hkspi.addr\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_146_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3682_ net12 _0864_ _0936_ net21 VGND VGND VPWR VPWR _1270_ sky130_fd_sc_hd__a22o_2
XFILLER_145_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5421_ net1967 net427 VGND VGND VPWR VPWR _2423_ sky130_fd_sc_hd__nand2_8
XFILLER_173_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput203 net203 VGND VGND VPWR VPWR mgmt_gpio_oeb[35] sky130_fd_sc_hd__buf_12
XFILLER_126_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput214 net214 VGND VGND VPWR VPWR mgmt_gpio_out[10] sky130_fd_sc_hd__buf_12
X_5352_ net458 net1550 _2415_ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__mux2_1
Xoutput225 net225 VGND VGND VPWR VPWR mgmt_gpio_out[20] sky130_fd_sc_hd__buf_12
Xoutput236 net236 VGND VGND VPWR VPWR mgmt_gpio_out[30] sky130_fd_sc_hd__buf_12
Xoutput247 net247 VGND VGND VPWR VPWR mgmt_gpio_out[6] sky130_fd_sc_hd__buf_12
XFILLER_114_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput258 net258 VGND VGND VPWR VPWR pad_flash_io1_do sky130_fd_sc_hd__buf_12
X_4303_ net577 net758 _1542_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__mux2_1
Xoutput269 net269 VGND VGND VPWR VPWR pll_div[3] sky130_fd_sc_hd__buf_12
X_5283_ net440 net1548 _2407_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__mux2_1
X_7022_ clknet_leaf_16_csclk net1305 net518 VGND VGND VPWR VPWR gpio_configure\[22\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_4234_ net591 net429 VGND VGND VPWR VPWR _1531_ sky130_fd_sc_hd__nand2_2
XFILLER_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4165_ wbbd_state\[4\] net528 VGND VGND VPWR VPWR _1517_ sky130_fd_sc_hd__and2_4
XFILLER_114_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4096_ net685 net618 net354 VGND VGND VPWR VPWR _1504_ sky130_fd_sc_hd__mux2_1
XFILLER_82_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6806_ clknet_leaf_63_csclk net1099 net501 VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__dfstp_2
XFILLER_168_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4998_ net478 _1662_ _1943_ _1946_ _2083_ VGND VGND VPWR VPWR _2208_ sky130_fd_sc_hd__a311o_1
XFILLER_11_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3949_ hkspi.pass_thru_mgmt net88 VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__or2_1
X_6737_ clknet_leaf_18_csclk net861 net510 VGND VGND VPWR VPWR gpio_configure\[35\]\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_23_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6668_ clknet_leaf_4_csclk net921 net494 VGND VGND VPWR VPWR gpio_configure\[9\]\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_139_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5619_ _2464_ VGND VGND VPWR VPWR _2465_ sky130_fd_sc_hd__inv_2
X_6599_ clknet_leaf_73_csclk net1032 net489 VGND VGND VPWR VPWR gpio_configure\[0\]\[11\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_192_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout441 net660 VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__buf_6
Xfanout452 net569 VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__buf_6
XFILLER_59_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout463 net542 VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__buf_6
XFILLER_120_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout474 net668 VGND VGND VPWR VPWR net474 sky130_fd_sc_hd__buf_12
XFILLER_171_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout485 net487 VGND VGND VPWR VPWR net485 sky130_fd_sc_hd__buf_4
Xfanout496 net497 VGND VGND VPWR VPWR net496 sky130_fd_sc_hd__buf_6
XFILLER_59_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5970_ net2070 _2792_ _2486_ VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__mux2_1
XFILLER_18_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4921_ _1601_ _1677_ _1834_ _1847_ VGND VGND VPWR VPWR _2132_ sky130_fd_sc_hd__a31o_1
XFILLER_52_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4852_ _1601_ _1677_ _1756_ _1718_ VGND VGND VPWR VPWR _2063_ sky130_fd_sc_hd__a31o_1
XFILLER_178_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3803_ hkspi.count\[0\] _1382_ VGND VGND VPWR VPWR _1385_ sky130_fd_sc_hd__nand2_1
XFILLER_21_748 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4783_ _1768_ _1993_ VGND VGND VPWR VPWR _1994_ sky130_fd_sc_hd__nor2_1
X_6522_ clknet_leaf_2_csclk net1474 net492 VGND VGND VPWR VPWR gpio_configure\[29\]\[9\]
+ sky130_fd_sc_hd__dfrtp_2
X_3734_ gpio_configure\[23\]\[0\] net372 _1316_ net264 VGND VGND VPWR VPWR _1320_
+ sky130_fd_sc_hd__a22o_1
XFILLER_186_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6453_ clknet_2_1__leaf_mgmt_gpio_in[4] _0075_ _0031_ VGND VGND VPWR VPWR hkspi.fixed\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3665_ gpio_configure\[32\]\[9\] _1101_ _1125_ gpio_configure\[22\]\[9\] VGND VGND
+ VPWR VPWR _1253_ sky130_fd_sc_hd__a22o_2
XFILLER_174_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5404_ net471 net1608 _2421_ VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__mux2_1
X_6384_ wbbd_state\[9\] net156 net138 wbbd_state\[8\] VGND VGND VPWR VPWR _3177_ sky130_fd_sc_hd__a22o_1
X_3596_ gpio_configure\[21\]\[3\] _0911_ _1067_ gpio_configure\[23\]\[11\] _1147_
+ VGND VGND VPWR VPWR _1186_ sky130_fd_sc_hd__a221o_1
X_5335_ net453 net1138 _2413_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__mux2_1
XFILLER_87_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5266_ net438 net1356 _2405_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__mux2_1
XFILLER_125_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7005_ clknet_leaf_23_csclk net1090 net526 VGND VGND VPWR VPWR gpio_configure\[20\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_4217_ net470 net1487 _1524_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__mux2_1
XFILLER_75_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5197_ net449 net1126 _2391_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__mux2_1
XFILLER_56_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4148_ net467 net1678 _1514_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__mux2_1
XFILLER_110_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4079_ net742 net445 net351 VGND VGND VPWR VPWR _1495_ sky130_fd_sc_hd__mux2_1
XFILLER_71_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_723 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap405 _2858_ VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__buf_12
XFILLER_128_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap416 _2813_ VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__buf_8
XFILLER_116_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold708 _0617_ VGND VGND VPWR VPWR net1241 sky130_fd_sc_hd__dlygate4sd3_1
Xhold719 gpio_configure\[20\]\[11\] VGND VGND VPWR VPWR net1252 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3450_ net388 _0903_ VGND VGND VPWR VPWR _1041_ sky130_fd_sc_hd__nor2_4
XFILLER_170_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3381_ gpio_configure\[16\]\[6\] _0912_ net350 gpio_configure\[4\]\[6\] VGND VGND
+ VPWR VPWR _0975_ sky130_fd_sc_hd__a22o_1
XFILLER_97_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5120_ _2322_ _2324_ _2327_ VGND VGND VPWR VPWR _2328_ sky130_fd_sc_hd__or3b_1
XFILLER_124_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5051_ _2253_ _2257_ _2259_ VGND VGND VPWR VPWR _2260_ sky130_fd_sc_hd__o21a_1
Xhold1408 net346 VGND VGND VPWR VPWR net1941 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1419 net329 VGND VGND VPWR VPWR net1952 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4002_ net469 net1574 _1472_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__mux2_1
XFILLER_38_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5953_ gpio_configure\[6\]\[12\] _2490_ _2494_ gpio_configure\[14\]\[12\] VGND VGND
+ VPWR VPWR _2776_ sky130_fd_sc_hd__a22o_1
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4904_ _1791_ _1800_ _2113_ _1602_ _2114_ VGND VGND VPWR VPWR _2115_ sky130_fd_sc_hd__o221a_1
X_5884_ gpio_configure\[15\]\[9\] _2510_ _2518_ gpio_configure\[3\]\[9\] _2709_ VGND
+ VGND VPWR VPWR _2710_ sky130_fd_sc_hd__a221o_1
XFILLER_33_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4835_ _1605_ _2045_ VGND VGND VPWR VPWR _2046_ sky130_fd_sc_hd__or2_1
XFILLER_178_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4766_ _1584_ _1652_ _1942_ _1963_ _1977_ VGND VGND VPWR VPWR _1978_ sky130_fd_sc_hd__a2111o_1
X_6505_ clknet_leaf_58_csclk net1271 net502 VGND VGND VPWR VPWR gpio_configure\[31\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_3717_ net283 _0886_ _0940_ net300 VGND VGND VPWR VPWR _1305_ sky130_fd_sc_hd__a22o_4
XFILLER_162_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4697_ _1777_ _1874_ _1908_ _1865_ VGND VGND VPWR VPWR _1909_ sky130_fd_sc_hd__o211a_1
XFILLER_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3648_ gpio_configure\[31\]\[10\] _1041_ _1087_ gpio_configure\[0\]\[10\] _1236_
+ VGND VGND VPWR VPWR _1237_ sky130_fd_sc_hd__a221o_1
X_6436_ net495 net482 VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__and2_1
XFILLER_161_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6367_ wbbd_state\[7\] net140 net143 net433 _3165_ VGND VGND VPWR VPWR _3166_ sky130_fd_sc_hd__a221o_1
XFILLER_88_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3579_ net55 _0871_ _1080_ gpio_configure\[16\]\[11\] _1168_ VGND VGND VPWR VPWR
+ _1169_ sky130_fd_sc_hd__a221o_1
XFILLER_161_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5318_ net447 net1302 net556 VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__mux2_1
X_6298_ gpio_configure\[31\]\[11\] _2480_ _2814_ gpio_configure\[11\]\[11\] VGND VGND
+ VPWR VPWR _3109_ sky130_fd_sc_hd__a22o_1
XFILLER_0_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_718 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold13 _1460_ VGND VGND VPWR VPWR net546 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 _0502_ VGND VGND VPWR VPWR net557 sky130_fd_sc_hd__dlygate4sd3_1
X_5249_ net573 net614 net547 VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__mux2_1
XFILLER_29_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold35 net692 VGND VGND VPWR VPWR net568 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 hkspi.addr\[6\] VGND VGND VPWR VPWR net579 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold57 _0863_ VGND VGND VPWR VPWR net590 sky130_fd_sc_hd__clkbuf_8
XFILLER_75_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold68 _0901_ VGND VGND VPWR VPWR net601 sky130_fd_sc_hd__clkbuf_16
XFILLER_29_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold79 _2429_ VGND VGND VPWR VPWR net612 sky130_fd_sc_hd__clkbuf_16
XFILLER_90_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4620_ _1805_ net432 VGND VGND VPWR VPWR _1832_ sky130_fd_sc_hd__nor2_1
XFILLER_175_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4551_ _1553_ _1749_ net127 VGND VGND VPWR VPWR _1763_ sky130_fd_sc_hd__a21oi_1
XFILLER_144_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3502_ net590 net554 VGND VGND VPWR VPWR _1093_ sky130_fd_sc_hd__nor2_2
XFILLER_156_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold505 _0540_ VGND VGND VPWR VPWR net1038 sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 net295 VGND VGND VPWR VPWR net1049 sky130_fd_sc_hd__dlygate4sd3_1
X_4482_ _1555_ _1693_ VGND VGND VPWR VPWR _1694_ sky130_fd_sc_hd__or2_2
Xhold527 _0115_ VGND VGND VPWR VPWR net1060 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold538 gpio_configure\[16\]\[7\] VGND VGND VPWR VPWR net1071 sky130_fd_sc_hd__dlygate4sd3_1
X_6221_ gpio_configure\[36\]\[8\] net403 net402 gpio_configure\[4\]\[8\] VGND VGND
+ VPWR VPWR _3035_ sky130_fd_sc_hd__a22o_2
XFILLER_171_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold549 _0347_ VGND VGND VPWR VPWR net1082 sky130_fd_sc_hd__dlygate4sd3_1
X_3433_ gpio_configure\[31\]\[5\] net375 net367 gpio_configure\[17\]\[5\] _1024_ VGND
+ VGND VPWR VPWR _1025_ sky130_fd_sc_hd__a221o_1
XFILLER_131_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6152_ gpio_configure\[22\]\[5\] net397 net395 gpio_configure\[33\]\[5\] VGND VGND
+ VPWR VPWR _2969_ sky130_fd_sc_hd__a22o_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ gpio_configure\[22\]\[7\] _0923_ _0938_ gpio_configure\[33\]\[7\] _0959_ VGND
+ VGND VPWR VPWR _0960_ sky130_fd_sc_hd__a221o_1
XFILLER_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ _2174_ _2311_ VGND VGND VPWR VPWR _2312_ sky130_fd_sc_hd__nor2_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6083_ gpio_configure\[13\]\[2\] net417 net393 gpio_configure\[34\]\[2\] _2902_ VGND
+ VGND VPWR VPWR _2903_ sky130_fd_sc_hd__a221o_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3295_ net390 _0887_ VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__nor2_8
XFILLER_57_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1205 gpio_configure\[15\]\[0\] VGND VGND VPWR VPWR net1738 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1216 net272 VGND VGND VPWR VPWR net1749 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_112_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _2172_ _2201_ _2243_ _1530_ net1991 VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__o32a_1
Xhold1227 _0179_ VGND VGND VPWR VPWR net1760 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1238 hkspi_disable VGND VGND VPWR VPWR net1771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1249 _0589_ VGND VGND VPWR VPWR net1782 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_65_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6985_ clknet_leaf_41_csclk net1046 net517 VGND VGND VPWR VPWR gpio_configure\[17\]\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5936_ gpio_configure\[5\]\[11\] _2496_ _2511_ gpio_configure\[25\]\[11\] VGND VGND
+ VPWR VPWR _2760_ sky130_fd_sc_hd__a22o_1
XFILLER_34_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5867_ gpio_configure\[15\]\[8\] _2510_ _2532_ gpio_configure\[18\]\[8\] VGND VGND
+ VPWR VPWR _2694_ sky130_fd_sc_hd__a22o_1
XFILLER_139_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4818_ _2028_ _1960_ _1824_ VGND VGND VPWR VPWR _2029_ sky130_fd_sc_hd__or3b_1
X_5798_ gpio_configure\[28\]\[5\] _2513_ _2521_ gpio_configure\[21\]\[5\] _2627_ VGND
+ VGND VPWR VPWR _2628_ sky130_fd_sc_hd__a221o_1
XFILLER_135_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4749_ _1692_ _1749_ _1771_ VGND VGND VPWR VPWR _1961_ sky130_fd_sc_hd__and3b_2
XFILLER_147_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6419_ net495 net482 VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__and2_1
XFILLER_162_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput103 wb_adr_i[13] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput114 wb_adr_i[23] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput125 wb_adr_i[4] VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__buf_6
XFILLER_130_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput136 wb_dat_i[13] VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_1
XFILLER_103_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput147 wb_dat_i[23] VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput158 wb_dat_i[4] VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_1
Xinput169 wb_stb_i VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_4
XFILLER_186_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_2_csclk clknet_3_1_0_csclk VGND VGND VPWR VPWR clknet_leaf_2_csclk sky130_fd_sc_hd__clkbuf_16
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6770_ clknet_leaf_71_csclk net987 net490 VGND VGND VPWR VPWR gpio_configure\[32\]\[12\]
+ sky130_fd_sc_hd__dfrtp_2
X_3982_ net1258 net434 _1461_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__mux2_1
XFILLER_16_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5721_ gpio_configure\[8\]\[1\] _2520_ net418 gpio_configure\[24\]\[1\] _2554_ VGND
+ VGND VPWR VPWR _2555_ sky130_fd_sc_hd__a221o_1
XFILLER_175_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5652_ net366 VGND VGND VPWR VPWR _2487_ sky130_fd_sc_hd__inv_2
XFILLER_176_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4603_ _1576_ _1684_ VGND VGND VPWR VPWR _1815_ sky130_fd_sc_hd__nor2_2
X_5583_ net457 net856 net603 VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__mux2_1
XFILLER_129_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4534_ _1576_ _1745_ VGND VGND VPWR VPWR _1746_ sky130_fd_sc_hd__nor2_1
Xhold302 _0370_ VGND VGND VPWR VPWR net835 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold313 gpio_configure\[24\]\[2\] VGND VGND VPWR VPWR net846 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold324 _0740_ VGND VGND VPWR VPWR net857 sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 gpio_configure\[17\]\[1\] VGND VGND VPWR VPWR net868 sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 _0494_ VGND VGND VPWR VPWR net879 sky130_fd_sc_hd__dlygate4sd3_1
X_4465_ _0834_ net479 VGND VGND VPWR VPWR _1677_ sky130_fd_sc_hd__and2_4
Xhold357 gpio_configure\[20\]\[1\] VGND VGND VPWR VPWR net890 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold368 _0230_ VGND VGND VPWR VPWR net901 sky130_fd_sc_hd__dlygate4sd3_1
X_6204_ gpio_configure\[22\]\[7\] net397 net395 gpio_configure\[33\]\[7\] _3018_ VGND
+ VGND VPWR VPWR _3019_ sky130_fd_sc_hd__a221o_1
X_3416_ net589 net608 VGND VGND VPWR VPWR _1008_ sky130_fd_sc_hd__nand2_8
XFILLER_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold379 net216 VGND VGND VPWR VPWR net912 sky130_fd_sc_hd__dlygate4sd3_1
X_7184_ clknet_3_1_0_wb_clk_i _0786_ net490 VGND VGND VPWR VPWR serial_data_staging_2\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_4396_ net110 _1555_ _1592_ VGND VGND VPWR VPWR _1608_ sky130_fd_sc_hd__or3_2
X_6135_ gpio_configure\[34\]\[4\] _2841_ _2852_ gpio_configure\[19\]\[4\] _2952_ VGND
+ VGND VPWR VPWR _2953_ sky130_fd_sc_hd__a221o_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3347_ net19 _0864_ _0898_ gpio_configure\[0\]\[7\] VGND VGND VPWR VPWR _0943_ sky130_fd_sc_hd__a22o_1
XFILLER_100_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1002 _0570_ VGND VGND VPWR VPWR net1535 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1013 gpio_configure\[12\]\[5\] VGND VGND VPWR VPWR net1546 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6066_ gpio_configure\[26\]\[1\] _2810_ _2811_ gpio_configure\[7\]\[1\] VGND VGND
+ VPWR VPWR _2887_ sky130_fd_sc_hd__a22o_1
Xhold1024 _0658_ VGND VGND VPWR VPWR net1557 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1035 gpio_configure\[20\]\[0\] VGND VGND VPWR VPWR net1568 sky130_fd_sc_hd__dlygate4sd3_1
X_3278_ net378 _0873_ VGND VGND VPWR VPWR _0874_ sky130_fd_sc_hd__nor2_8
Xhold1046 _0543_ VGND VGND VPWR VPWR net1579 sky130_fd_sc_hd__dlygate4sd3_1
X_5017_ _1841_ _2226_ VGND VGND VPWR VPWR _2227_ sky130_fd_sc_hd__nor2_1
Xhold1057 clk1_output_dest VGND VGND VPWR VPWR net1590 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1068 _0394_ VGND VGND VPWR VPWR net1601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1079 net2077 VGND VGND VPWR VPWR net1612 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_208 _2843_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_219 net280 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6968_ clknet_leaf_54_csclk net1370 net506 VGND VGND VPWR VPWR gpio_configure\[15\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_13_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5919_ gpio_configure\[20\]\[10\] _2499_ _2505_ gpio_configure\[11\]\[10\] VGND VGND
+ VPWR VPWR _2744_ sky130_fd_sc_hd__a22o_1
XFILLER_22_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6899_ clknet_leaf_25_csclk net557 net518 VGND VGND VPWR VPWR gpio_configure\[7\]\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_179_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold880 gpio_configure\[33\]\[1\] VGND VGND VPWR VPWR net1413 sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 _0659_ VGND VGND VPWR VPWR net1424 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_67_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1580 xfer_state\[0\] VGND VGND VPWR VPWR net2113 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1591 mgmt_gpio_data\[35\] VGND VGND VPWR VPWR net2124 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_724 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4250_ net450 net1260 _1533_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__mux2_1
XFILLER_113_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3201_ gpio_configure\[33\]\[3\] VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__inv_2
X_4181_ net2079 _1376_ _1519_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__mux2_1
XFILLER_121_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6822_ clknet_leaf_29_csclk net543 net520 VGND VGND VPWR VPWR clk2_output_dest sky130_fd_sc_hd__dfrtp_4
X_6753_ clknet_3_0_0_csclk net1762 net491 VGND VGND VPWR VPWR gpio_configure\[20\]\[10\]
+ sky130_fd_sc_hd__dfstp_1
X_3965_ net545 net474 net644 VGND VGND VPWR VPWR _1460_ sky130_fd_sc_hd__o21ai_4
X_5704_ gpio_configure\[17\]\[0\] _2537_ _2538_ gpio_configure\[1\]\[0\] VGND VGND
+ VPWR VPWR _2539_ sky130_fd_sc_hd__a22o_2
X_3896_ _0823_ _1442_ VGND VGND VPWR VPWR _1443_ sky130_fd_sc_hd__or2_1
X_6684_ clknet_leaf_4_csclk net593 net495 VGND VGND VPWR VPWR gpio_configure\[12\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_148_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5635_ xfer_state\[2\] _1449_ _2469_ VGND VGND VPWR VPWR _2475_ sky130_fd_sc_hd__and3_1
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5566_ net452 net976 net648 VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__mux2_1
Xhold110 wbbd_write VGND VGND VPWR VPWR net643 sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 gpio_configure\[27\]\[4\] VGND VGND VPWR VPWR net654 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_163_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4517_ _1663_ _1665_ VGND VGND VPWR VPWR _1729_ sky130_fd_sc_hd__nor2_2
Xhold132 _1467_ VGND VGND VPWR VPWR net665 sky130_fd_sc_hd__dlygate4sd3_1
X_5497_ net452 net968 net641 VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__mux2_1
XFILLER_117_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold143 _0681_ VGND VGND VPWR VPWR net676 sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 gpio_configure\[19\]\[5\] VGND VGND VPWR VPWR net687 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 gpio_configure\[37\]\[4\] VGND VGND VPWR VPWR net698 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 _0406_ VGND VGND VPWR VPWR net709 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4448_ _1612_ _1650_ VGND VGND VPWR VPWR _1660_ sky130_fd_sc_hd__nand2_1
XFILLER_171_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold187 gpio_configure\[19\]\[4\] VGND VGND VPWR VPWR net720 sky130_fd_sc_hd__dlygate4sd3_1
Xhold198 _0440_ VGND VGND VPWR VPWR net731 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7167_ clknet_3_3_0_wb_clk_i net2050 net502 VGND VGND VPWR VPWR serial_data_staging_1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_113_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4379_ net127 net128 net126 net125 VGND VGND VPWR VPWR _1591_ sky130_fd_sc_hd__nor4_4
XFILLER_86_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6118_ gpio_configure\[15\]\[3\] net407 _2934_ _2936_ VGND VGND VPWR VPWR _2937_
+ sky130_fd_sc_hd__a211o_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7098_ clknet_leaf_51_csclk net741 net506 VGND VGND VPWR VPWR gpio_configure\[32\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6049_ gpio_configure\[23\]\[1\] _2822_ VGND VGND VPWR VPWR _2870_ sky130_fd_sc_hd__and2_1
XFILLER_37_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_20_csclk clknet_3_4_0_csclk VGND VGND VPWR VPWR clknet_leaf_20_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_64_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_35_csclk clknet_3_7_0_csclk VGND VGND VPWR VPWR clknet_leaf_35_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_91_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3750_ gpio_configure\[37\]\[8\] _1065_ _1122_ gpio_configure\[8\]\[8\] VGND VGND
+ VPWR VPWR _1336_ sky130_fd_sc_hd__a22o_1
XFILLER_118_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3681_ gpio_configure\[30\]\[1\] _0892_ _1086_ gpio_configure\[29\]\[9\] _1268_ VGND
+ VGND VPWR VPWR _1269_ sky130_fd_sc_hd__a221o_1
XFILLER_158_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5420_ net434 net1314 _2422_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__mux2_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5351_ net464 net1668 _2415_ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__mux2_1
Xoutput204 net204 VGND VGND VPWR VPWR mgmt_gpio_oeb[36] sky130_fd_sc_hd__buf_12
Xoutput215 net215 VGND VGND VPWR VPWR mgmt_gpio_out[11] sky130_fd_sc_hd__buf_12
XFILLER_160_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput226 net226 VGND VGND VPWR VPWR mgmt_gpio_out[21] sky130_fd_sc_hd__buf_12
XFILLER_99_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput237 net237 VGND VGND VPWR VPWR mgmt_gpio_out[31] sky130_fd_sc_hd__buf_12
Xoutput248 net248 VGND VGND VPWR VPWR mgmt_gpio_out[7] sky130_fd_sc_hd__buf_12
X_4302_ net465 net832 _1542_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__mux2_1
Xoutput259 net259 VGND VGND VPWR VPWR pad_flash_io1_ieb sky130_fd_sc_hd__buf_12
XFILLER_114_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5282_ net447 net1306 _2407_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__mux2_1
XFILLER_153_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4233_ _0818_ net474 net2103 _1528_ _1530_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__a2111o_1
X_7021_ clknet_leaf_28_csclk net961 net521 VGND VGND VPWR VPWR gpio_configure\[22\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_114_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4164_ net1202 net446 _1516_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__mux2_1
XFILLER_114_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4095_ net946 _1503_ _1499_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__mux2_1
XFILLER_55_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6805_ clknet_leaf_61_csclk net855 net498 VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__dfstp_2
XFILLER_169_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4997_ _1668_ _2203_ VGND VGND VPWR VPWR _2207_ sky130_fd_sc_hd__nor2_1
XFILLER_23_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6736_ clknet_leaf_19_csclk net1691 net510 VGND VGND VPWR VPWR gpio_configure\[35\]\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_3948_ net256 VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__inv_2
XFILLER_176_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6667_ clknet_leaf_1_csclk net1390 net493 VGND VGND VPWR VPWR gpio_configure\[9\]\[10\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_109_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3879_ net130 net129 _1430_ VGND VGND VPWR VPWR _1431_ sky130_fd_sc_hd__or3_1
XFILLER_192_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5618_ pad_count_1\[2\] _2460_ VGND VGND VPWR VPWR _2464_ sky130_fd_sc_hd__or2_1
XFILLER_137_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6598_ clknet_leaf_73_csclk net1635 net489 VGND VGND VPWR VPWR gpio_configure\[0\]\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_124_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5549_ net446 net1186 _2437_ VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__mux2_1
XFILLER_145_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout442 net666 VGND VGND VPWR VPWR net442 sky130_fd_sc_hd__clkbuf_16
Xfanout453 net569 VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__clkbuf_4
Xfanout464 net465 VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__buf_6
Xfanout475 xfer_state\[1\] VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__buf_8
XFILLER_59_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout486 net487 VGND VGND VPWR VPWR net486 sky130_fd_sc_hd__buf_6
XFILLER_19_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout497 net527 VGND VGND VPWR VPWR net497 sky130_fd_sc_hd__buf_4
XFILLER_58_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_554 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_6_0_wb_clk_i clknet_2_3_0_wb_clk_i VGND VGND VPWR VPWR clknet_3_6_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_97_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4920_ _1807_ net432 _1886_ _1790_ _2130_ VGND VGND VPWR VPWR _2131_ sky130_fd_sc_hd__o221a_1
XFILLER_45_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4851_ _1833_ _1886_ _1721_ VGND VGND VPWR VPWR _2062_ sky130_fd_sc_hd__o21ai_1
XTAP_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3802_ hkspi.count\[2\] hkspi.count\[1\] hkspi.count\[0\] VGND VGND VPWR VPWR _1384_
+ sky130_fd_sc_hd__and3_2
X_4782_ _1816_ _1817_ _1762_ VGND VGND VPWR VPWR _1993_ sky130_fd_sc_hd__a21bo_1
X_6521_ clknet_leaf_2_csclk net1809 net492 VGND VGND VPWR VPWR gpio_configure\[29\]\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_3733_ gpio_configure\[16\]\[0\] _0912_ _0930_ gpio_configure\[9\]\[0\] VGND VGND
+ VPWR VPWR _1319_ sky130_fd_sc_hd__a22o_1
XFILLER_146_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6452_ clknet_2_3__leaf_mgmt_gpio_in[4] net2022 _0030_ VGND VGND VPWR VPWR hkspi.odata\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_3664_ gpio_configure\[6\]\[1\] _0876_ _1054_ gpio_configure\[19\]\[9\] VGND VGND
+ VPWR VPWR _1252_ sky130_fd_sc_hd__a22o_1
XFILLER_106_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5403_ net367 net647 VGND VGND VPWR VPWR _2421_ sky130_fd_sc_hd__nand2_8
X_3595_ net14 _0864_ _0896_ gpio_configure\[19\]\[3\] _1146_ VGND VGND VPWR VPWR _1185_
+ sky130_fd_sc_hd__a221o_2
X_6383_ _3176_ net2062 _3162_ VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__mux2_1
X_5334_ net459 net1447 _2413_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__mux2_1
XFILLER_114_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5265_ net440 net1530 _2405_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__mux2_1
X_7004_ clknet_leaf_24_csclk net1665 net526 VGND VGND VPWR VPWR gpio_configure\[20\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_4216_ _1068_ net429 VGND VGND VPWR VPWR _1524_ sky130_fd_sc_hd__nand2_2
X_5196_ net455 net1696 _2391_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__mux2_1
XFILLER_68_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4147_ _1095_ net425 VGND VGND VPWR VPWR _1514_ sky130_fd_sc_hd__nand2_4
XFILLER_95_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4078_ net964 _1494_ _1490_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__mux2_1
XFILLER_36_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6719_ clknet_leaf_63_csclk net1111 net501 VGND VGND VPWR VPWR gpio_configure\[37\]\[11\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_177_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap406 _2855_ VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__buf_12
XFILLER_7_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap417 _2804_ VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__buf_12
XFILLER_115_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold709 gpio_configure\[11\]\[3\] VGND VGND VPWR VPWR net1242 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3380_ serial_data_staging_2\[12\] serial_bb_data_2 serial_bb_enable VGND VGND VPWR
+ VPWR net309 sky130_fd_sc_hd__mux2_4
XFILLER_156_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5050_ _1708_ _1929_ _2202_ VGND VGND VPWR VPWR _2259_ sky130_fd_sc_hd__and3_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1409 net322 VGND VGND VPWR VPWR net1942 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4001_ _0883_ net427 VGND VGND VPWR VPWR _1472_ sky130_fd_sc_hd__nand2_8
XFILLER_77_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5952_ gpio_configure\[25\]\[12\] _2511_ _2538_ gpio_configure\[1\]\[12\] _2774_
+ VGND VGND VPWR VPWR _2775_ sky130_fd_sc_hd__a221o_1
XFILLER_18_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4903_ _1693_ _1779_ _1992_ _1689_ VGND VGND VPWR VPWR _2114_ sky130_fd_sc_hd__o22a_1
X_5883_ gpio_configure\[27\]\[9\] _2506_ _2511_ gpio_configure\[25\]\[9\] VGND VGND
+ VPWR VPWR _2709_ sky130_fd_sc_hd__a22o_1
XFILLER_61_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4834_ _1638_ _1639_ _1671_ _1678_ _1777_ VGND VGND VPWR VPWR _2045_ sky130_fd_sc_hd__o32a_1
XFILLER_60_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4765_ _1584_ _1654_ _1958_ _1959_ _1976_ VGND VGND VPWR VPWR _1977_ sky130_fd_sc_hd__a2111o_1
XFILLER_193_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6504_ clknet_leaf_57_csclk net1454 net502 VGND VGND VPWR VPWR gpio_configure\[31\]\[6\]
+ sky130_fd_sc_hd__dfrtp_2
X_3716_ gpio_configure\[27\]\[1\] _0925_ _0934_ gpio_configure\[1\]\[1\] _1303_ VGND
+ VGND VPWR VPWR _1304_ sky130_fd_sc_hd__a221o_1
XFILLER_147_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4696_ _1581_ _1801_ _1863_ _1776_ VGND VGND VPWR VPWR _1908_ sky130_fd_sc_hd__o22a_1
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6435_ net495 net481 VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__and2_1
X_3647_ net13 _0864_ _1196_ clk1_output_dest VGND VGND VPWR VPWR _1236_ sky130_fd_sc_hd__a22o_1
XFILLER_146_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6366_ wbbd_state\[9\] net149 net163 wbbd_state\[8\] VGND VGND VPWR VPWR _3165_ sky130_fd_sc_hd__a22o_1
X_3578_ gpio_configure\[34\]\[3\] net358 _1109_ gpio_configure\[36\]\[11\] VGND VGND
+ VPWR VPWR _1168_ sky130_fd_sc_hd__a22o_1
XFILLER_161_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5317_ net453 net1178 net556 VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__mux2_1
XFILLER_130_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6297_ gpio_configure\[3\]\[11\] _2830_ _2842_ gpio_configure\[15\]\[11\] VGND VGND
+ VPWR VPWR _3108_ sky130_fd_sc_hd__a22o_1
XFILLER_142_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold14 _2403_ VGND VGND VPWR VPWR net547 sky130_fd_sc_hd__dlygate4sd3_1
X_5248_ net439 net656 net547 VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__mux2_1
Xhold25 hkspi.addr\[0\] VGND VGND VPWR VPWR net558 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold36 net454 VGND VGND VPWR VPWR net569 sky130_fd_sc_hd__buf_8
XFILLER_29_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold47 _0842_ VGND VGND VPWR VPWR net580 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 _1056_ VGND VGND VPWR VPWR net591 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold69 _0902_ VGND VGND VPWR VPWR net602 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5179_ _1588_ _1836_ _1891_ _1660_ _1682_ VGND VGND VPWR VPWR _2385_ sky130_fd_sc_hd__o2111a_1
XFILLER_29_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4550_ net125 _1749_ VGND VGND VPWR VPWR _1762_ sky130_fd_sc_hd__xnor2_1
XFILLER_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3501_ gpio_configure\[34\]\[4\] _0874_ _0974_ serial_bb_clock _1091_ VGND VGND VPWR
+ VPWR _1092_ sky130_fd_sc_hd__a221o_2
XFILLER_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold506 gpio_configure\[9\]\[7\] VGND VGND VPWR VPWR net1039 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4481_ _1590_ _1692_ VGND VGND VPWR VPWR _1693_ sky130_fd_sc_hd__or2_4
XFILLER_156_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold517 _0116_ VGND VGND VPWR VPWR net1050 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold528 net285 VGND VGND VPWR VPWR net1061 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6220_ net2068 _3034_ net366 VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__mux2_1
Xhold539 _0580_ VGND VGND VPWR VPWR net1072 sky130_fd_sc_hd__dlygate4sd3_1
X_3432_ gpio_configure\[27\]\[5\] net370 _0974_ net308 VGND VGND VPWR VPWR _1024_
+ sky130_fd_sc_hd__a22o_1
XFILLER_103_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3363_ gpio_configure\[30\]\[7\] _0892_ _0913_ gpio_configure\[7\]\[7\] _0958_ VGND
+ VGND VPWR VPWR _0959_ sky130_fd_sc_hd__a221o_1
X_6151_ gpio_configure\[23\]\[5\] _2822_ net396 gpio_configure\[20\]\[5\] _2965_ VGND
+ VGND VPWR VPWR _2968_ sky130_fd_sc_hd__a221o_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _2301_ _2310_ VGND VGND VPWR VPWR _2311_ sky130_fd_sc_hd__nor2_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3294_ net387 _0889_ VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__nor2_8
XFILLER_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6082_ gpio_configure\[12\]\[2\] net409 net392 gpio_configure\[5\]\[2\] VGND VGND
+ VPWR VPWR _2902_ sky130_fd_sc_hd__a22o_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1206 _0565_ VGND VGND VPWR VPWR net1739 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1217 _0401_ VGND VGND VPWR VPWR net1750 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1228 gpio_configure\[20\]\[10\] VGND VGND VPWR VPWR net1761 sky130_fd_sc_hd__dlygate4sd3_1
X_5033_ _1529_ _2221_ _2242_ VGND VGND VPWR VPWR _2243_ sky130_fd_sc_hd__or3_1
Xhold1239 _0423_ VGND VGND VPWR VPWR net1772 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6984_ clknet_leaf_56_csclk net1434 net504 VGND VGND VPWR VPWR gpio_configure\[17\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_53_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5935_ _2752_ _2754_ _2756_ _2758_ VGND VGND VPWR VPWR _2759_ sky130_fd_sc_hd__or4_1
XFILLER_80_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5866_ gpio_configure\[8\]\[8\] _2520_ _2692_ VGND VGND VPWR VPWR _2693_ sky130_fd_sc_hd__a21o_1
XFILLER_33_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4817_ _2000_ _2014_ _2026_ _2027_ VGND VGND VPWR VPWR _2028_ sky130_fd_sc_hd__or4b_1
X_5797_ gpio_configure\[11\]\[5\] _2505_ _2506_ gpio_configure\[27\]\[5\] VGND VGND
+ VPWR VPWR _2627_ sky130_fd_sc_hd__a22o_1
XFILLER_178_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4748_ _1599_ _1657_ VGND VGND VPWR VPWR _1960_ sky130_fd_sc_hd__nor2_1
XFILLER_135_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4679_ _1684_ _1836_ VGND VGND VPWR VPWR _1891_ sky130_fd_sc_hd__or2_1
X_6418_ net495 net482 VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__and2_1
XFILLER_162_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6349_ net1969 _1376_ _3156_ VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__mux2_1
XFILLER_88_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_759 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput104 wb_adr_i[14] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput115 wb_adr_i[24] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput126 wb_adr_i[5] VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__buf_6
Xinput137 wb_dat_i[14] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_1
Xinput148 wb_dat_i[24] VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_1
Xinput159 wb_dat_i[5] VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_1
XFILLER_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3981_ net571 net1002 net668 VGND VGND VPWR VPWR _1469_ sky130_fd_sc_hd__mux2_1
XFILLER_16_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5720_ gpio_configure\[10\]\[1\] net421 _2528_ gpio_configure\[7\]\[1\] VGND VGND
+ VPWR VPWR _2554_ sky130_fd_sc_hd__a22o_1
XFILLER_43_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5651_ _1452_ _2443_ VGND VGND VPWR VPWR _2486_ sky130_fd_sc_hd__nor2_4
XFILLER_30_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4602_ net110 net99 net530 _1770_ _1813_ VGND VGND VPWR VPWR _1814_ sky130_fd_sc_hd__a41o_1
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5582_ net542 gpio_configure\[37\]\[1\] net603 VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__mux2_1
XFILLER_175_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4533_ _0834_ _1584_ VGND VGND VPWR VPWR _1745_ sky130_fd_sc_hd__nand2_8
XFILLER_116_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold303 gpio_configure\[36\]\[10\] VGND VGND VPWR VPWR net836 sky130_fd_sc_hd__dlygate4sd3_1
Xhold314 _0639_ VGND VGND VPWR VPWR net847 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold325 gpio_configure\[3\]\[1\] VGND VGND VPWR VPWR net858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold336 _0582_ VGND VGND VPWR VPWR net869 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4464_ net380 VGND VGND VPWR VPWR _1676_ sky130_fd_sc_hd__inv_2
Xhold347 gpio_configure\[0\]\[1\] VGND VGND VPWR VPWR net880 sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 _0606_ VGND VGND VPWR VPWR net891 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6203_ gpio_configure\[18\]\[7\] net399 net410 gpio_configure\[8\]\[7\] VGND VGND
+ VPWR VPWR _3018_ sky130_fd_sc_hd__a22o_1
Xhold369 gpio_configure\[23\]\[12\] VGND VGND VPWR VPWR net902 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3415_ net628 _1006_ VGND VGND VPWR VPWR _1007_ sky130_fd_sc_hd__nor2_8
X_7183_ clknet_3_0_0_wb_clk_i _0785_ net490 VGND VGND VPWR VPWR serial_data_staging_2\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_98_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4395_ _1606_ VGND VGND VPWR VPWR _1607_ sky130_fd_sc_hd__inv_2
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6134_ gpio_configure\[37\]\[4\] net400 net416 gpio_configure\[32\]\[4\] _2941_ VGND
+ VGND VPWR VPWR _2952_ sky130_fd_sc_hd__a221o_4
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3346_ gpio_configure\[11\]\[7\] _0907_ net368 gpio_configure\[9\]\[7\] VGND VGND
+ VPWR VPWR _0942_ sky130_fd_sc_hd__a22o_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1003 gpio_configure\[27\]\[5\] VGND VGND VPWR VPWR net1536 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6065_ gpio_configure\[1\]\[1\] net401 net405 gpio_configure\[24\]\[1\] _2869_ VGND
+ VGND VPWR VPWR _2886_ sky130_fd_sc_hd__a221o_1
Xhold1014 _0546_ VGND VGND VPWR VPWR net1547 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3277_ net561 net608 VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__nand2_8
Xhold1025 gpio_configure\[31\]\[5\] VGND VGND VPWR VPWR net1558 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1036 _0605_ VGND VGND VPWR VPWR net1569 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1047 gpio_configure\[35\]\[2\] VGND VGND VPWR VPWR net1580 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5016_ _1779_ _1872_ VGND VGND VPWR VPWR _2226_ sky130_fd_sc_hd__and2_1
Xhold1058 _0424_ VGND VGND VPWR VPWR net1591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1069 gpio_configure\[33\]\[0\] VGND VGND VPWR VPWR net1602 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_209 _2852_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6967_ clknet_leaf_31_csclk net1535 net523 VGND VGND VPWR VPWR gpio_configure\[15\]\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_5918_ gpio_configure\[15\]\[10\] _2510_ _2535_ gpio_configure\[23\]\[10\] _2742_
+ VGND VGND VPWR VPWR _2743_ sky130_fd_sc_hd__a221o_1
X_6898_ clknet_leaf_25_csclk net1585 net518 VGND VGND VPWR VPWR gpio_configure\[7\]\[0\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_179_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5849_ gpio_configure\[15\]\[7\] _2510_ _2535_ gpio_configure\[23\]\[7\] _2676_ VGND
+ VGND VPWR VPWR _2677_ sky130_fd_sc_hd__a221o_1
XFILLER_166_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold870 gpio_configure\[30\]\[10\] VGND VGND VPWR VPWR net1403 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold881 _0707_ VGND VGND VPWR VPWR net1414 sky130_fd_sc_hd__dlygate4sd3_1
Xhold892 gpio_configure\[19\]\[6\] VGND VGND VPWR VPWR net1425 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1570 wbbd_state\[6\] VGND VGND VPWR VPWR net2103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1581 serial_bb_data_2 VGND VGND VPWR VPWR net2114 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_83_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1592 gpio_configure\[32\]\[6\] VGND VGND VPWR VPWR net2125 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3200_ gpio_configure\[34\]\[3\] VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__inv_2
X_4180_ wbbd_state\[2\] net528 VGND VGND VPWR VPWR _1519_ sky130_fd_sc_hd__and2_4
XFILLER_79_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6821_ clknet_leaf_28_csclk net1591 net520 VGND VGND VPWR VPWR clk1_output_dest sky130_fd_sc_hd__dfrtp_4
XFILLER_35_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6752_ clknet_leaf_6_csclk net1482 net497 VGND VGND VPWR VPWR gpio_configure\[20\]\[9\]
+ sky130_fd_sc_hd__dfrtp_2
X_3964_ net545 net669 net644 VGND VGND VPWR VPWR _1459_ sky130_fd_sc_hd__o21a_4
X_5703_ net472 _2466_ _2495_ VGND VGND VPWR VPWR _2538_ sky130_fd_sc_hd__and3_4
XFILLER_176_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6683_ clknet_leaf_11_csclk net596 net511 VGND VGND VPWR VPWR gpio_configure\[12\]\[10\]
+ sky130_fd_sc_hd__dfstp_1
X_3895_ xfer_count\[0\] xfer_count\[2\] xfer_count\[3\] xfer_count\[1\] VGND VGND
+ VPWR VPWR _1442_ sky130_fd_sc_hd__or4b_1
X_5634_ _2470_ _2473_ VGND VGND VPWR VPWR _2474_ sky130_fd_sc_hd__nand2_1
XFILLER_136_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5565_ net458 net1580 net648 VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__mux2_1
XFILLER_191_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold100 net1994 VGND VGND VPWR VPWR net633 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold111 _1458_ VGND VGND VPWR VPWR net644 sky130_fd_sc_hd__dlygate4sd3_1
X_4516_ _1612_ _1652_ VGND VGND VPWR VPWR _1728_ sky130_fd_sc_hd__nand2_1
Xhold122 _0665_ VGND VGND VPWR VPWR net655 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5496_ net459 net1350 net641 VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__mux2_1
Xhold133 net659 VGND VGND VPWR VPWR net666 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 net288 VGND VGND VPWR VPWR net677 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold155 _0602_ VGND VGND VPWR VPWR net688 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 _0742_ VGND VGND VPWR VPWR net699 sky130_fd_sc_hd__dlygate4sd3_1
X_4447_ _1612_ _1645_ VGND VGND VPWR VPWR _1659_ sky130_fd_sc_hd__nand2_1
Xhold177 gpio_configure\[11\]\[4\] VGND VGND VPWR VPWR net710 sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 _0601_ VGND VGND VPWR VPWR net721 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold199 gpio_configure\[6\]\[3\] VGND VGND VPWR VPWR net732 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7166_ clknet_3_2_0_wb_clk_i _0768_ net500 VGND VGND VPWR VPWR serial_data_staging_1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_98_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4378_ _0817_ _1548_ VGND VGND VPWR VPWR _1590_ sky130_fd_sc_hd__or2_4
XFILLER_86_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_1_csclk clknet_3_1_0_csclk VGND VGND VPWR VPWR clknet_leaf_1_csclk sky130_fd_sc_hd__clkbuf_16
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6117_ gpio_configure\[37\]\[3\] net400 net416 gpio_configure\[32\]\[3\] _2935_ VGND
+ VGND VPWR VPWR _2936_ sky130_fd_sc_hd__a221o_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3329_ net388 _0895_ VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__nor2_4
XFILLER_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7097_ clknet_leaf_51_csclk net799 net505 VGND VGND VPWR VPWR gpio_configure\[32\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_85_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6048_ gpio_configure\[31\]\[1\] net423 net415 gpio_configure\[11\]\[1\] VGND VGND
+ VPWR VPWR _2869_ sky130_fd_sc_hd__a22o_1
XTAP_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3680_ gpio_configure\[15\]\[9\] _1102_ _1122_ gpio_configure\[8\]\[9\] VGND VGND
+ VPWR VPWR _1268_ sky130_fd_sc_hd__a22o_1
XFILLER_158_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5350_ net471 net1606 _2415_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__mux2_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput205 net205 VGND VGND VPWR VPWR mgmt_gpio_oeb[37] sky130_fd_sc_hd__buf_12
Xoutput216 net216 VGND VGND VPWR VPWR mgmt_gpio_out[12] sky130_fd_sc_hd__buf_12
XFILLER_160_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput227 net227 VGND VGND VPWR VPWR mgmt_gpio_out[22] sky130_fd_sc_hd__buf_12
Xoutput238 net238 VGND VGND VPWR VPWR mgmt_gpio_out[32] sky130_fd_sc_hd__buf_12
X_4301_ net470 net1648 _1542_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__mux2_1
XFILLER_141_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput249 net249 VGND VGND VPWR VPWR mgmt_gpio_out[8] sky130_fd_sc_hd__buf_12
X_5281_ net453 net1200 _2407_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__mux2_1
XFILLER_153_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7020_ clknet_leaf_60_csclk net821 net499 VGND VGND VPWR VPWR gpio_configure\[22\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_114_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4232_ wbbd_state\[5\] _1527_ VGND VGND VPWR VPWR _1530_ sky130_fd_sc_hd__or2_2
XFILLER_141_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4163_ net714 net569 _1516_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__mux2_1
XFILLER_110_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4094_ net730 net569 net354 VGND VGND VPWR VPWR _1503_ sky130_fd_sc_hd__mux2_1
XFILLER_55_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6804_ clknet_leaf_61_csclk net1577 net498 VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__dfstp_1
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4996_ _1651_ _2203_ VGND VGND VPWR VPWR _2206_ sky130_fd_sc_hd__nor2_1
X_6735_ clknet_leaf_73_csclk net989 net489 VGND VGND VPWR VPWR gpio_configure\[18\]\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_23_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3947_ hkspi.pass_thru_mgmt_delay net86 VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__nand2b_1
XFILLER_149_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6666_ clknet_leaf_0_csclk net1737 net487 VGND VGND VPWR VPWR gpio_configure\[9\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_3878_ net101 net100 net103 net102 VGND VGND VPWR VPWR _1430_ sky130_fd_sc_hd__or4_1
XFILLER_109_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5617_ _0825_ _2459_ _2461_ net2135 _2458_ VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__o32a_1
XFILLER_164_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6597_ clknet_leaf_75_csclk net1699 net489 VGND VGND VPWR VPWR gpio_configure\[0\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_136_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5548_ net452 net970 _2437_ VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__mux2_1
XFILLER_191_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5479_ net452 net1025 net612 VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__mux2_1
XFILLER_78_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout432 _1808_ VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__buf_8
Xfanout443 net445 VGND VGND VPWR VPWR net443 sky130_fd_sc_hd__buf_8
X_7149_ clknet_3_0_0_wb_clk_i _0752_ net499 VGND VGND VPWR VPWR pad_count_1\[1\] sky130_fd_sc_hd__dfstp_1
Xfanout454 net568 VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__buf_8
XFILLER_101_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout465 net542 VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__buf_8
Xfanout487 net527 VGND VGND VPWR VPWR net487 sky130_fd_sc_hd__buf_6
Xfanout498 net500 VGND VGND VPWR VPWR net498 sky130_fd_sc_hd__buf_8
XFILLER_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4850_ _1728_ _1919_ VGND VGND VPWR VPWR _2061_ sky130_fd_sc_hd__nand2_1
XTAP_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3801_ net2127 _1379_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__xor2_1
XFILLER_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4781_ _1557_ _1583_ VGND VGND VPWR VPWR _1992_ sky130_fd_sc_hd__nand2_2
X_6520_ clknet_leaf_3_csclk net1249 net494 VGND VGND VPWR VPWR gpio_configure\[24\]\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_119_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3732_ net52 _0871_ _0902_ gpio_configure\[37\]\[0\] VGND VGND VPWR VPWR _1318_ sky130_fd_sc_hd__a22o_2
XFILLER_9_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6451_ clknet_2_3__leaf_mgmt_gpio_in[4] net2055 _0029_ VGND VGND VPWR VPWR hkspi.odata\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_3663_ gpio_configure\[18\]\[1\] _0894_ _0912_ gpio_configure\[16\]\[1\] VGND VGND
+ VPWR VPWR _1251_ sky130_fd_sc_hd__a22o_1
X_5402_ net1071 net434 _2420_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__mux2_1
X_6382_ wbbd_state\[7\] net146 net160 net433 _3175_ VGND VGND VPWR VPWR _3176_ sky130_fd_sc_hd__a221o_1
X_3594_ gpio_configure\[27\]\[3\] _0925_ _1041_ gpio_configure\[31\]\[11\] _1145_
+ VGND VGND VPWR VPWR _1184_ sky130_fd_sc_hd__a221o_1
XFILLER_127_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5333_ net464 net1421 _2413_ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__mux2_1
XFILLER_114_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5264_ net447 net1264 _2405_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__mux2_1
X_7003_ clknet_leaf_60_csclk net891 net499 VGND VGND VPWR VPWR gpio_configure\[20\]\[1\]
+ sky130_fd_sc_hd__dfstp_4
X_4215_ net896 net444 _1523_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__mux2_1
X_5195_ net461 net1720 _2391_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__mux2_1
XFILLER_68_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4146_ net446 net1118 net671 VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__mux2_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4077_ net828 net451 net351 VGND VGND VPWR VPWR _1494_ sky130_fd_sc_hd__mux2_1
XFILLER_56_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4979_ _2175_ _2179_ _2183_ _2188_ VGND VGND VPWR VPWR _2189_ sky130_fd_sc_hd__or4_1
X_6718_ clknet_leaf_63_csclk net745 net501 VGND VGND VPWR VPWR gpio_configure\[37\]\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_50_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6649_ clknet_3_1_0_wb_clk_i _0262_ VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__dfxtp_1
XFILLER_109_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_34_csclk clknet_3_7_0_csclk VGND VGND VPWR VPWR clknet_leaf_34_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_117_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_49_csclk clknet_3_3_0_csclk VGND VGND VPWR VPWR clknet_leaf_49_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_87_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap407 _2842_ VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__buf_12
Xmax_cap418 _2531_ VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__buf_12
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4000_ net1116 net434 _1471_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__mux2_1
XFILLER_111_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5951_ gpio_configure\[22\]\[12\] _2498_ _2506_ gpio_configure\[27\]\[12\] VGND VGND
+ VPWR VPWR _2774_ sky130_fd_sc_hd__a22o_1
XFILLER_52_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4902_ _1684_ _1800_ _2111_ _1776_ _1880_ VGND VGND VPWR VPWR _2113_ sky130_fd_sc_hd__o221a_1
X_5882_ net2063 _2708_ net366 VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__mux2_1
XFILLER_178_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4833_ _1606_ _1678_ _1696_ VGND VGND VPWR VPWR _2044_ sky130_fd_sc_hd__o21ai_1
XFILLER_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4764_ _1955_ _1964_ _1975_ VGND VGND VPWR VPWR _1976_ sky130_fd_sc_hd__or3_1
XFILLER_193_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6503_ clknet_leaf_38_csclk net1559 net523 VGND VGND VPWR VPWR gpio_configure\[31\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_159_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3715_ gpio_configure\[18\]\[9\] _1047_ _1302_ irq_2_inputsrc VGND VGND VPWR VPWR
+ _1303_ sky130_fd_sc_hd__a22o_2
XFILLER_174_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4695_ _1581_ _1793_ _1801_ _1872_ _1906_ VGND VGND VPWR VPWR _1907_ sky130_fd_sc_hd__o221a_1
X_6434_ net495 net481 VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__and2_1
X_3646_ net284 _0886_ _0919_ gpio_configure\[24\]\[2\] _1234_ VGND VGND VPWR VPWR
+ _1235_ sky130_fd_sc_hd__a221o_1
XFILLER_162_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6365_ _3164_ net2052 _3162_ VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__mux2_1
XFILLER_115_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3577_ gpio_configure\[5\]\[3\] net355 _0939_ gpio_configure\[8\]\[3\] _1166_ VGND
+ VGND VPWR VPWR _1167_ sky130_fd_sc_hd__a221o_1
X_5316_ net458 net1676 net556 VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__mux2_1
XFILLER_115_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6296_ gpio_configure\[36\]\[11\] net403 net402 gpio_configure\[4\]\[11\] VGND VGND
+ VPWR VPWR _3107_ sky130_fd_sc_hd__a22o_2
XFILLER_130_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5247_ net441 net974 net547 VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__mux2_1
Xhold15 net1907 VGND VGND VPWR VPWR net548 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 _0860_ VGND VGND VPWR VPWR net559 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 _0291_ VGND VGND VPWR VPWR net570 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold48 _0843_ VGND VGND VPWR VPWR net581 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold59 _1531_ VGND VGND VPWR VPWR net592 sky130_fd_sc_hd__dlygate4sd3_1
X_5178_ _2287_ _2315_ _2362_ _2383_ VGND VGND VPWR VPWR _2384_ sky130_fd_sc_hd__or4_1
XFILLER_56_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4129_ _1087_ net425 VGND VGND VPWR VPWR _1511_ sky130_fd_sc_hd__and2_1
XFILLER_29_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3500_ net7 _0891_ _0896_ gpio_configure\[19\]\[4\] VGND VGND VPWR VPWR _1091_ sky130_fd_sc_hd__a22o_1
XFILLER_190_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4480_ net127 net128 _0835_ net125 VGND VGND VPWR VPWR _1692_ sky130_fd_sc_hd__or4_4
Xhold507 _0524_ VGND VGND VPWR VPWR net1040 sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 gpio_configure\[3\]\[7\] VGND VGND VPWR VPWR net1051 sky130_fd_sc_hd__dlygate4sd3_1
Xhold529 _0099_ VGND VGND VPWR VPWR net1062 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3431_ _1019_ _1020_ _1021_ _1022_ VGND VGND VPWR VPWR _1023_ sky130_fd_sc_hd__or4_1
X_6150_ gpio_configure\[29\]\[5\] _2816_ _2820_ gpio_configure\[21\]\[5\] _2966_ VGND
+ VGND VPWR VPWR _2967_ sky130_fd_sc_hd__a221o_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3362_ gpio_configure\[6\]\[7\] net357 _0939_ gpio_configure\[8\]\[7\] VGND VGND
+ VPWR VPWR _0958_ sky130_fd_sc_hd__a22o_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5101_ _2302_ _2304_ _2306_ _2309_ VGND VGND VPWR VPWR _2310_ sky130_fd_sc_hd__or4_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6081_ gpio_configure\[1\]\[2\] net401 net415 gpio_configure\[11\]\[2\] _2900_ VGND
+ VGND VPWR VPWR _2901_ sky130_fd_sc_hd__a221o_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ net561 _0879_ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__nand2_8
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1207 gpio_configure\[13\]\[2\] VGND VGND VPWR VPWR net1740 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _2222_ _2240_ _2241_ VGND VGND VPWR VPWR _2242_ sky130_fd_sc_hd__o21ba_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1218 gpio_configure\[6\]\[8\] VGND VGND VPWR VPWR net1751 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1229 _0356_ VGND VGND VPWR VPWR net1762 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6983_ clknet_leaf_38_csclk net1555 net523 VGND VGND VPWR VPWR gpio_configure\[17\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_80_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5934_ gpio_configure\[8\]\[11\] _2520_ net418 gpio_configure\[24\]\[11\] _2757_
+ VGND VGND VPWR VPWR _2758_ sky130_fd_sc_hd__a221o_1
X_5865_ gpio_configure\[9\]\[8\] _2512_ net418 gpio_configure\[24\]\[8\] VGND VGND
+ VPWR VPWR _2692_ sky130_fd_sc_hd__a22o_1
XFILLER_33_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4816_ _1668_ _1745_ net424 _1798_ VGND VGND VPWR VPWR _2027_ sky130_fd_sc_hd__o22a_1
X_5796_ gpio_configure\[16\]\[5\] _0831_ net419 VGND VGND VPWR VPWR _2626_ sky130_fd_sc_hd__o21a_1
XFILLER_193_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4747_ _1655_ _1750_ VGND VGND VPWR VPWR _1959_ sky130_fd_sc_hd__nor2_1
XFILLER_147_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4678_ _1797_ _1886_ VGND VGND VPWR VPWR _1890_ sky130_fd_sc_hd__or2_2
XFILLER_162_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6417_ net492 net481 VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__and2_1
XFILLER_107_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3629_ net37 net353 _1122_ gpio_configure\[8\]\[10\] _1195_ VGND VGND VPWR VPWR _1218_
+ sky130_fd_sc_hd__a221o_1
XFILLER_150_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6348_ wbbd_state\[1\] net528 VGND VGND VPWR VPWR _3156_ sky130_fd_sc_hd__and2_4
XFILLER_1_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6279_ gpio_configure\[16\]\[10\] _2831_ _2860_ gpio_configure\[17\]\[10\] _3085_
+ VGND VGND VPWR VPWR _3091_ sky130_fd_sc_hd__a221o_1
Xinput105 wb_adr_i[15] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_1
Xinput116 wb_adr_i[25] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput127 wb_adr_i[6] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__buf_4
XFILLER_48_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput138 wb_dat_i[15] VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_1
Xinput149 wb_dat_i[25] VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_1
XFILLER_57_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3980_ net1449 net437 _1461_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__mux2_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5650_ net475 _0825_ VGND VGND VPWR VPWR _2485_ sky130_fd_sc_hd__nor2_4
XFILLER_188_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4601_ _1771_ _1784_ _1812_ _1594_ _1586_ VGND VGND VPWR VPWR _1813_ sky130_fd_sc_hd__a2111o_1
X_5581_ net471 net1627 net603 VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__mux2_1
XFILLER_163_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4532_ net530 _1585_ VGND VGND VPWR VPWR _1744_ sky130_fd_sc_hd__nor2_2
XFILLER_191_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold304 _0331_ VGND VGND VPWR VPWR net837 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold315 gpio_configure\[15\]\[1\] VGND VGND VPWR VPWR net848 sky130_fd_sc_hd__dlygate4sd3_1
Xhold326 _0470_ VGND VGND VPWR VPWR net859 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4463_ _1564_ _1568_ _1674_ VGND VGND VPWR VPWR _1675_ sky130_fd_sc_hd__nor3b_4
Xhold337 gpio_configure\[14\]\[1\] VGND VGND VPWR VPWR net870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 _0446_ VGND VGND VPWR VPWR net881 sky130_fd_sc_hd__dlygate4sd3_1
X_6202_ gpio_configure\[23\]\[7\] _2822_ net396 gpio_configure\[20\]\[7\] VGND VGND
+ VPWR VPWR _3017_ sky130_fd_sc_hd__a22o_1
XFILLER_171_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold359 gpio_configure\[24\]\[1\] VGND VGND VPWR VPWR net892 sky130_fd_sc_hd__dlygate4sd3_1
X_3414_ net589 net600 VGND VGND VPWR VPWR _1006_ sky130_fd_sc_hd__nand2_8
X_7182_ clknet_3_2_0_wb_clk_i _0784_ net499 VGND VGND VPWR VPWR serial_data_staging_2\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_4394_ _1575_ _1605_ VGND VGND VPWR VPWR _1606_ sky130_fd_sc_hd__or2_2
XFILLER_98_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6133_ gpio_configure\[28\]\[4\] _2861_ _2946_ _2948_ _2950_ VGND VGND VPWR VPWR
+ _2951_ sky130_fd_sc_hd__a2111o_2
X_3345_ net298 _0910_ _0917_ gpio_configure\[29\]\[7\] VGND VGND VPWR VPWR _0941_
+ sky130_fd_sc_hd__a22o_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6064_ gpio_configure\[2\]\[1\] net398 _2843_ gpio_configure\[5\]\[1\] _2884_ VGND
+ VGND VPWR VPWR _2885_ sky130_fd_sc_hd__a221o_1
XFILLER_100_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1004 _0666_ VGND VGND VPWR VPWR net1537 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3276_ net607 net599 VGND VGND VPWR VPWR _0872_ sky130_fd_sc_hd__nor2_8
Xhold1015 gpio_configure\[3\]\[5\] VGND VGND VPWR VPWR net1548 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1026 _0125_ VGND VGND VPWR VPWR net1559 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _1885_ _1995_ _2224_ VGND VGND VPWR VPWR _2225_ sky130_fd_sc_hd__or3_1
Xhold1037 gpio_configure\[2\]\[2\] VGND VGND VPWR VPWR net1570 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1048 _0724_ VGND VGND VPWR VPWR net1581 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1059 net265 VGND VGND VPWR VPWR net1592 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6966_ clknet_leaf_16_csclk net1299 net512 VGND VGND VPWR VPWR gpio_configure\[15\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_41_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5917_ gpio_configure\[22\]\[10\] _2498_ _2524_ _2741_ VGND VGND VPWR VPWR _2742_
+ sky130_fd_sc_hd__a22o_1
X_6897_ clknet_leaf_43_csclk net1088 net517 VGND VGND VPWR VPWR gpio_configure\[6\]\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_167_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5848_ gpio_configure\[20\]\[7\] _2499_ net420 gpio_configure\[25\]\[7\] VGND VGND
+ VPWR VPWR _2676_ sky130_fd_sc_hd__a22o_1
X_5779_ gpio_configure\[13\]\[4\] _2501_ _2520_ gpio_configure\[8\]\[4\] VGND VGND
+ VPWR VPWR _2610_ sky130_fd_sc_hd__a22o_1
XFILLER_166_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold860 gpio_configure\[33\]\[6\] VGND VGND VPWR VPWR net1393 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_174_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold871 _0135_ VGND VGND VPWR VPWR net1404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 gpio_configure\[23\]\[6\] VGND VGND VPWR VPWR net1415 sky130_fd_sc_hd__dlygate4sd3_1
Xhold893 _0603_ VGND VGND VPWR VPWR net1426 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1560 _0077_ VGND VGND VPWR VPWR net2093 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1571 mgmt_gpio_data_buf\[18\] VGND VGND VPWR VPWR net2104 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1582 mgmt_gpio_data_buf\[6\] VGND VGND VPWR VPWR net2115 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1593 hkspi.addr\[6\] VGND VGND VPWR VPWR net2126 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6820_ clknet_3_4_0_csclk net1772 net511 VGND VGND VPWR VPWR hkspi_disable sky130_fd_sc_hd__dfrtp_1
XFILLER_51_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6751_ clknet_leaf_73_csclk net1494 net489 VGND VGND VPWR VPWR gpio_configure\[20\]\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_3963_ net643 net474 VGND VGND VPWR VPWR _1458_ sky130_fd_sc_hd__nand2b_1
X_5702_ pad_count_1\[4\] _2466_ _2495_ VGND VGND VPWR VPWR _2537_ sky130_fd_sc_hd__and3_4
Xclkbuf_1_1_0_wb_clk_i clknet_0_wb_clk_i VGND VGND VPWR VPWR clknet_1_1_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_6682_ clknet_leaf_11_csclk net623 net511 VGND VGND VPWR VPWR gpio_configure\[12\]\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_31_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3894_ wbbd_state\[9\] _1428_ net2025 VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__a21o_1
X_5633_ pad_count_2\[3\] pad_count_2\[2\] VGND VGND VPWR VPWR _2473_ sky130_fd_sc_hd__and2_2
XFILLER_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5564_ net464 net1411 net648 VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__mux2_1
XFILLER_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4515_ _1723_ _1724_ _1725_ _1726_ VGND VGND VPWR VPWR _1727_ sky130_fd_sc_hd__and4_1
Xhold101 net535 VGND VGND VPWR VPWR net634 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 net670 VGND VGND VPWR VPWR net645 sky130_fd_sc_hd__buf_6
X_5495_ net464 net1383 net641 VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__mux2_1
Xhold123 net2111 VGND VGND VPWR VPWR net656 sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 _0117_ VGND VGND VPWR VPWR net667 sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 _0101_ VGND VGND VPWR VPWR net678 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 gpio_configure\[0\]\[4\] VGND VGND VPWR VPWR net689 sky130_fd_sc_hd__dlygate4sd3_1
X_4446_ _1657_ VGND VGND VPWR VPWR _1658_ sky130_fd_sc_hd__inv_2
Xhold167 gpio_configure\[31\]\[4\] VGND VGND VPWR VPWR net700 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold178 _0537_ VGND VGND VPWR VPWR net711 sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 gpio_configure\[4\]\[4\] VGND VGND VPWR VPWR net722 sky130_fd_sc_hd__dlygate4sd3_1
X_7165_ clknet_3_0_0_wb_clk_i net2035 net500 VGND VGND VPWR VPWR serial_data_staging_1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_98_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4377_ _0817_ _1548_ VGND VGND VPWR VPWR _1589_ sky130_fd_sc_hd__nor2_2
XFILLER_98_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6116_ gpio_configure\[16\]\[3\] _2831_ _2852_ gpio_configure\[19\]\[3\] VGND VGND
+ VPWR VPWR _2935_ sky130_fd_sc_hd__a22o_1
X_3328_ _0873_ net387 VGND VGND VPWR VPWR _0924_ sky130_fd_sc_hd__nor2_4
X_7096_ clknet_leaf_64_csclk net905 net501 VGND VGND VPWR VPWR gpio_configure\[32\]\[1\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6047_ _2485_ _2867_ _2868_ _2487_ net2040 VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__a32o_1
X_3259_ net597 net586 net605 VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__mux2_1
XTAP_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6949_ clknet_leaf_36_csclk net1131 net522 VGND VGND VPWR VPWR gpio_configure\[13\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold690 _0286_ VGND VGND VPWR VPWR net1223 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1390 gpio_configure\[27\]\[6\] VGND VGND VPWR VPWR net1923 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_691 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput206 net206 VGND VGND VPWR VPWR mgmt_gpio_oeb[3] sky130_fd_sc_hd__buf_12
Xoutput217 net217 VGND VGND VPWR VPWR mgmt_gpio_out[13] sky130_fd_sc_hd__buf_12
X_4300_ _1081_ net429 VGND VGND VPWR VPWR _1542_ sky130_fd_sc_hd__nand2_2
Xoutput228 net228 VGND VGND VPWR VPWR mgmt_gpio_out[23] sky130_fd_sc_hd__buf_12
XFILLER_99_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5280_ net459 net1344 _2407_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__mux2_1
Xoutput239 net239 VGND VGND VPWR VPWR mgmt_gpio_out[33] sky130_fd_sc_hd__buf_12
XFILLER_141_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4231_ wbbd_state\[5\] _1527_ VGND VGND VPWR VPWR _1529_ sky130_fd_sc_hd__nor2_8
XFILLER_141_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4162_ net806 net577 _1516_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__mux2_1
XFILLER_68_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4093_ net1540 _1502_ _1499_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__mux2_1
XFILLER_82_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6803_ clknet_leaf_76_csclk net709 net488 VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__dfrtp_4
XFILLER_169_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4995_ _1646_ _2203_ VGND VGND VPWR VPWR _2205_ sky130_fd_sc_hd__nor2_1
X_6734_ clknet_leaf_75_csclk net1074 net489 VGND VGND VPWR VPWR gpio_configure\[18\]\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_149_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3946_ hkspi.pass_thru_mgmt net487 VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__nor2_1
XFILLER_51_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6665_ clknet_leaf_0_csclk net1813 net487 VGND VGND VPWR VPWR gpio_configure\[9\]\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_137_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3877_ hkspi.rdstb net476 net483 VGND VGND VPWR VPWR _1429_ sky130_fd_sc_hd__o21ai_1
XFILLER_192_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5616_ xfer_state\[0\] _0825_ VGND VGND VPWR VPWR _2463_ sky130_fd_sc_hd__nand2_1
XFILLER_176_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6596_ clknet_leaf_73_csclk net1797 net489 VGND VGND VPWR VPWR gpio_configure\[0\]\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_164_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5547_ net458 net1680 _2437_ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__mux2_1
XFILLER_105_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5478_ net457 net842 net612 VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__mux2_1
XFILLER_3_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4429_ _1639_ _1640_ VGND VGND VPWR VPWR _1641_ sky130_fd_sc_hd__nor2_1
XFILLER_48_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7148_ clknet_3_3_0_wb_clk_i _0751_ net499 VGND VGND VPWR VPWR pad_count_1\[0\] sky130_fd_sc_hd__dfrtp_2
Xfanout444 net445 VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__clkbuf_4
Xfanout455 net456 VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__buf_6
Xfanout466 net467 VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__buf_6
Xfanout477 _1602_ VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__buf_6
Xfanout488 net491 VGND VGND VPWR VPWR net488 sky130_fd_sc_hd__buf_6
X_7079_ clknet_leaf_39_csclk net1133 net517 VGND VGND VPWR VPWR gpio_configure\[29\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout499 net500 VGND VGND VPWR VPWR net499 sky130_fd_sc_hd__buf_8
XFILLER_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3800_ _1381_ _1383_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__nor2_1
XFILLER_178_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4780_ _1753_ _1785_ VGND VGND VPWR VPWR _1991_ sky130_fd_sc_hd__nor2_1
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3731_ net389 _0903_ VGND VGND VPWR VPWR _1317_ sky130_fd_sc_hd__nor2_1
XFILLER_159_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_0_csclk clknet_3_1_0_csclk VGND VGND VPWR VPWR clknet_leaf_0_csclk sky130_fd_sc_hd__clkbuf_16
XFILLER_158_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_119_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3662_ _1250_ net1997 _0970_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__mux2_1
XFILLER_158_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6450_ clknet_2_3__leaf_mgmt_gpio_in[4] _0072_ _0028_ VGND VGND VPWR VPWR hkspi.odata\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_5401_ net844 net439 _2420_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__mux2_1
X_6381_ wbbd_state\[9\] net155 net137 wbbd_state\[8\] VGND VGND VPWR VPWR _3175_ sky130_fd_sc_hd__a22o_1
X_3593_ _1179_ _1180_ _1181_ _1182_ VGND VGND VPWR VPWR _1183_ sky130_fd_sc_hd__or4_1
XFILLER_126_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5332_ net470 net1789 _2413_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__mux2_1
XFILLER_126_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5263_ net452 net1077 _2405_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__mux2_1
XFILLER_114_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7002_ clknet_leaf_61_csclk net1569 net500 VGND VGND VPWR VPWR gpio_configure\[20\]\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_4214_ net920 net450 _1523_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__mux2_1
X_5194_ net466 net1749 _2391_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__mux2_1
X_4145_ net569 net1918 net671 VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__mux2_1
XFILLER_95_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4076_ net1083 _1493_ _1490_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__mux2_1
XFILLER_55_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4978_ _1706_ _1994_ _2185_ _2187_ VGND VGND VPWR VPWR _2188_ sky130_fd_sc_hd__a211o_1
X_6717_ clknet_leaf_62_csclk net939 net501 VGND VGND VPWR VPWR gpio_configure\[37\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_3929_ mgmt_gpio_data\[6\] net77 net94 VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__mux2_4
XFILLER_20_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6648_ clknet_3_1_0_wb_clk_i _0261_ VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__dfxtp_1
XFILLER_166_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6579_ clknet_leaf_14_csclk net707 net513 VGND VGND VPWR VPWR mgmt_gpio_data\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_117_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap408 _2839_ VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__buf_12
XFILLER_171_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap419 _2524_ VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__buf_12
XFILLER_143_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_694 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5950_ gpio_configure\[9\]\[12\] _2512_ _2523_ gpio_configure\[2\]\[12\] _2772_ VGND
+ VGND VPWR VPWR _2773_ sky130_fd_sc_hd__a221o_1
XFILLER_46_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4901_ _1788_ _1798_ _1836_ _1850_ _2111_ VGND VGND VPWR VPWR _2112_ sky130_fd_sc_hd__a41o_1
X_5881_ xfer_state\[1\] serial_data_staging_1\[7\] _2707_ VGND VGND VPWR VPWR _2708_
+ sky130_fd_sc_hd__a21o_1
XFILLER_61_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4832_ _1605_ _1678_ _1685_ VGND VGND VPWR VPWR _2043_ sky130_fd_sc_hd__nor3_1
XANTENNA_190 _0904_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4763_ _1584_ _1650_ _1965_ _1974_ VGND VGND VPWR VPWR _1975_ sky130_fd_sc_hd__a211o_1
XFILLER_159_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6502_ clknet_leaf_25_csclk net701 net518 VGND VGND VPWR VPWR gpio_configure\[31\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_3714_ _0881_ net383 VGND VGND VPWR VPWR _1302_ sky130_fd_sc_hd__nor2_1
X_4694_ _1678_ _1801_ VGND VGND VPWR VPWR _1906_ sky130_fd_sc_hd__or2_1
X_6433_ net492 net481 VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__and2_1
X_3645_ gpio_configure\[23\]\[2\] _0922_ _1116_ gpio_configure\[26\]\[10\] VGND VGND
+ VPWR VPWR _1234_ sky130_fd_sc_hd__a22o_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3576_ gpio_configure\[6\]\[3\] net357 _1042_ gpio_configure\[6\]\[11\] VGND VGND
+ VPWR VPWR _1166_ sky130_fd_sc_hd__a22o_1
XFILLER_136_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6364_ wbbd_state\[9\] net148 net162 wbbd_state\[8\] _3163_ VGND VGND VPWR VPWR _3164_
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5315_ net542 net1921 net556 VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__mux2_1
X_6295_ net2094 net366 _3105_ _3106_ VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__o22a_1
XFILLER_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5246_ net618 net685 net547 VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__mux2_1
XFILLER_29_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold16 hkspi.addr\[3\] VGND VGND VPWR VPWR net549 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 _0861_ VGND VGND VPWR VPWR net560 sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 hkspi.odata\[7\] VGND VGND VPWR VPWR net571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 _0905_ VGND VGND VPWR VPWR net582 sky130_fd_sc_hd__dlygate4sd3_1
X_5177_ _1837_ _1867_ _2382_ VGND VGND VPWR VPWR _2383_ sky130_fd_sc_hd__or3b_1
XFILLER_68_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4128_ net434 net1288 _1510_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__mux2_1
XFILLER_84_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4059_ net1508 _1484_ _1481_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__mux2_1
XFILLER_37_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold508 gpio_configure\[12\]\[7\] VGND VGND VPWR VPWR net1041 sky130_fd_sc_hd__dlygate4sd3_1
Xhold519 _0476_ VGND VGND VPWR VPWR net1052 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3430_ net57 _0871_ _0902_ gpio_configure\[37\]\[5\] _1010_ VGND VGND VPWR VPWR _1022_
+ sky130_fd_sc_hd__a221o_1
XFILLER_143_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3361_ net290 _0886_ _0935_ gpio_configure\[4\]\[7\] _0956_ VGND VGND VPWR VPWR _0957_
+ sky130_fd_sc_hd__a221o_1
XFILLER_112_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5100_ _2178_ _2180_ _2307_ _2308_ VGND VGND VPWR VPWR _2309_ sky130_fd_sc_hd__or4_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6080_ gpio_configure\[31\]\[2\] net423 _2810_ gpio_configure\[26\]\[2\] VGND VGND
+ VPWR VPWR _2900_ sky130_fd_sc_hd__a22o_1
X_3292_ net388 net562 VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__nor2_8
XFILLER_112_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _1861_ _1928_ _2137_ VGND VGND VPWR VPWR _2241_ sky130_fd_sc_hd__or3_2
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1208 _0551_ VGND VGND VPWR VPWR net1741 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1219 _0247_ VGND VGND VPWR VPWR net1752 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6982_ clknet_leaf_19_csclk net1171 net510 VGND VGND VPWR VPWR gpio_configure\[17\]\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_5933_ gpio_configure\[14\]\[11\] _2494_ _2534_ gpio_configure\[26\]\[11\] VGND VGND
+ VPWR VPWR _2757_ sky130_fd_sc_hd__a22o_1
XFILLER_34_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_33_csclk clknet_3_7_0_csclk VGND VGND VPWR VPWR clknet_leaf_33_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_178_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5864_ gpio_configure\[17\]\[8\] _2537_ _2538_ gpio_configure\[1\]\[8\] _2690_ VGND
+ VGND VPWR VPWR _2691_ sky130_fd_sc_hd__a221o_1
X_4815_ _1942_ _2002_ _2024_ _2025_ VGND VGND VPWR VPWR _2026_ sky130_fd_sc_hd__or4b_1
XFILLER_166_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5795_ net2056 _2625_ net366 VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__mux2_1
XFILLER_119_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_48_csclk clknet_3_6_0_csclk VGND VGND VPWR VPWR clknet_leaf_48_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_119_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4746_ _1599_ _1653_ VGND VGND VPWR VPWR _1958_ sky130_fd_sc_hd__nor2_1
XFILLER_193_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4677_ _1588_ _1798_ VGND VGND VPWR VPWR _1889_ sky130_fd_sc_hd__or2_1
XFILLER_134_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6416_ net492 net481 VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__and2_1
X_3628_ gpio_configure\[10\]\[10\] _1068_ _1119_ gpio_configure\[5\]\[10\] _1198_
+ VGND VGND VPWR VPWR _1217_ sky130_fd_sc_hd__a221o_1
XFILLER_115_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6347_ net2081 _1440_ _3155_ _3154_ VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__a31o_1
XFILLER_0_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3559_ gpio_configure\[31\]\[3\] net375 _1101_ gpio_configure\[32\]\[11\] VGND VGND
+ VPWR VPWR _1149_ sky130_fd_sc_hd__a22o_1
XFILLER_88_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6278_ gpio_configure\[22\]\[10\] _2824_ _2829_ gpio_configure\[33\]\[10\] _3089_
+ VGND VGND VPWR VPWR _3090_ sky130_fd_sc_hd__a221o_1
XFILLER_103_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput106 wb_adr_i[16] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_1
Xinput117 wb_adr_i[26] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_1
Xinput128 wb_adr_i[7] VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__buf_6
X_5229_ _1302_ net425 VGND VGND VPWR VPWR _2401_ sky130_fd_sc_hd__nand2_1
XFILLER_76_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput139 wb_dat_i[16] VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_1
XFILLER_56_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_90 hkspi.pass_thru_user VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_3_0_wb_clk_i clknet_1_1_1_wb_clk_i VGND VGND VPWR VPWR clknet_2_3_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_121_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4600_ _1578_ _1695_ _1786_ _1811_ _1691_ VGND VGND VPWR VPWR _1812_ sky130_fd_sc_hd__a2111o_1
XFILLER_30_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5580_ net602 net429 VGND VGND VPWR VPWR _2441_ sky130_fd_sc_hd__nand2_8
XFILLER_30_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4531_ _0834_ _1577_ _1676_ _1708_ _1742_ VGND VGND VPWR VPWR _1743_ sky130_fd_sc_hd__o311a_1
XFILLER_129_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold305 gpio_configure\[23\]\[2\] VGND VGND VPWR VPWR net838 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold316 _0566_ VGND VGND VPWR VPWR net849 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4462_ net126 _1572_ VGND VGND VPWR VPWR _1674_ sky130_fd_sc_hd__nor2_1
Xhold327 gpio_configure\[35\]\[9\] VGND VGND VPWR VPWR net860 sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 _0558_ VGND VGND VPWR VPWR net871 sky130_fd_sc_hd__dlygate4sd3_1
X_6201_ gpio_configure\[29\]\[7\] _2816_ _2820_ gpio_configure\[21\]\[7\] _3013_ VGND
+ VGND VPWR VPWR _3016_ sky130_fd_sc_hd__a221o_1
Xhold349 net2133 VGND VGND VPWR VPWR net882 sky130_fd_sc_hd__dlygate4sd3_1
X_3413_ serial_data_staging_1\[12\] serial_bb_data_1 serial_bb_enable VGND VGND VPWR
+ VPWR net308 sky130_fd_sc_hd__mux2_8
XFILLER_144_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7181_ clknet_3_3_0_wb_clk_i _0783_ net505 VGND VGND VPWR VPWR serial_data_staging_2\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_171_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4393_ _1561_ _1562_ _1603_ VGND VGND VPWR VPWR _1605_ sky130_fd_sc_hd__a21o_4
XFILLER_98_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3344_ net389 _0889_ VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__nor2_8
X_6132_ gpio_configure\[16\]\[4\] _2831_ net391 gpio_configure\[17\]\[4\] _2949_ VGND
+ VGND VPWR VPWR _2950_ sky130_fd_sc_hd__a221o_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3275_ net378 _0870_ VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__nor2_8
X_6063_ gpio_configure\[13\]\[1\] net417 _2862_ gpio_configure\[25\]\[1\] VGND VGND
+ VPWR VPWR _2884_ sky130_fd_sc_hd__a22o_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1005 gpio_configure\[14\]\[5\] VGND VGND VPWR VPWR net1538 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1016 _0474_ VGND VGND VPWR VPWR net1549 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1027 gpio_configure\[36\]\[5\] VGND VGND VPWR VPWR net1560 sky130_fd_sc_hd__dlygate4sd3_1
X_5014_ _1611_ _1775_ _1693_ VGND VGND VPWR VPWR _2224_ sky130_fd_sc_hd__a21oi_1
Xhold1038 _0463_ VGND VGND VPWR VPWR net1571 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 gpio_configure\[13\]\[0\] VGND VGND VPWR VPWR net1582 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_521 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6965_ clknet_leaf_36_csclk net1141 net522 VGND VGND VPWR VPWR gpio_configure\[15\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_53_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5916_ gpio_configure\[16\]\[10\] net472 VGND VGND VPWR VPWR _2741_ sky130_fd_sc_hd__or2_1
XFILLER_81_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6896_ clknet_leaf_54_csclk net1380 net506 VGND VGND VPWR VPWR gpio_configure\[6\]\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_22_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5847_ _2668_ _2670_ _2672_ _2674_ VGND VGND VPWR VPWR _2675_ sky130_fd_sc_hd__or4_1
XFILLER_21_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5778_ gpio_configure\[10\]\[4\] net421 _2535_ gpio_configure\[23\]\[4\] _2608_ VGND
+ VGND VPWR VPWR _2609_ sky130_fd_sc_hd__a221o_1
XFILLER_154_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4729_ _1599_ _1707_ VGND VGND VPWR VPWR _1941_ sky130_fd_sc_hd__nand2_1
XFILLER_135_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold850 gpio_configure\[27\]\[1\] VGND VGND VPWR VPWR net1383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold861 _0712_ VGND VGND VPWR VPWR net1394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold872 gpio_configure\[22\]\[9\] VGND VGND VPWR VPWR net1405 sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 _0635_ VGND VGND VPWR VPWR net1416 sky130_fd_sc_hd__dlygate4sd3_1
Xhold894 gpio_configure\[10\]\[9\] VGND VGND VPWR VPWR net1427 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1550 hkspi.state\[1\] VGND VGND VPWR VPWR net2083 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1561 serial_data_staging_2\[10\] VGND VGND VPWR VPWR net2094 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1572 mgmt_gpio_data\[36\] VGND VGND VPWR VPWR net2105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1583 hkspi.addr\[2\] VGND VGND VPWR VPWR net2116 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1594 hkspi.count\[0\] VGND VGND VPWR VPWR net2127 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6750_ clknet_leaf_8_csclk net1113 net509 VGND VGND VPWR VPWR gpio_configure\[34\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_3962_ wbbd_state\[9\] _1429_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__and2_1
XFILLER_189_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5701_ gpio_configure\[26\]\[0\] _2534_ _2535_ gpio_configure\[23\]\[0\] _2533_ VGND
+ VGND VPWR VPWR _2536_ sky130_fd_sc_hd__a221o_1
XFILLER_188_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6681_ clknet_leaf_11_csclk net1498 net511 VGND VGND VPWR VPWR gpio_configure\[12\]\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_3893_ wbbd_state\[8\] _1428_ net2020 VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__a21o_1
XFILLER_31_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5632_ net2084 _2470_ _2472_ VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__a21oi_1
XFILLER_129_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5563_ net471 net1566 net648 VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__mux2_1
XFILLER_8_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4514_ _1652_ _1670_ VGND VGND VPWR VPWR _1726_ sky130_fd_sc_hd__nand2_1
Xhold102 _0435_ VGND VGND VPWR VPWR net635 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold113 net430 VGND VGND VPWR VPWR net646 sky130_fd_sc_hd__buf_8
X_5494_ net471 net1618 net641 VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__mux2_1
Xhold124 _0443_ VGND VGND VPWR VPWR net657 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 wbbd_busy VGND VGND VPWR VPWR net668 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold146 gpio_configure\[17\]\[11\] VGND VGND VPWR VPWR net679 sky130_fd_sc_hd__dlygate4sd3_1
X_4445_ _1623_ _1656_ VGND VGND VPWR VPWR _1657_ sky130_fd_sc_hd__or2_4
Xhold157 _0449_ VGND VGND VPWR VPWR net690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 _0124_ VGND VGND VPWR VPWR net701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold179 net2010 VGND VGND VPWR VPWR net712 sky130_fd_sc_hd__dlygate4sd3_1
X_7164_ clknet_3_0_0_wb_clk_i net2038 net500 VGND VGND VPWR VPWR serial_data_staging_1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_144_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4376_ net530 net480 VGND VGND VPWR VPWR _1588_ sky130_fd_sc_hd__nand2_8
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6115_ gpio_configure\[31\]\[3\] net423 net412 gpio_configure\[9\]\[3\] VGND VGND
+ VPWR VPWR _2934_ sky130_fd_sc_hd__a22o_1
X_3327_ _0870_ net386 VGND VGND VPWR VPWR _0923_ sky130_fd_sc_hd__nor2_8
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7095_ clknet_leaf_64_csclk net1714 net501 VGND VGND VPWR VPWR gpio_configure\[32\]\[0\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ gpio_configure\[0\]\[0\] _2851_ VGND VGND VPWR VPWR _2868_ sky130_fd_sc_hd__or2_1
X_3258_ net606 net1970 net474 VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__mux2_2
XFILLER_39_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3189_ gpio_configure\[3\]\[3\] VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__inv_2
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6948_ clknet_leaf_26_csclk net1741 net526 VGND VGND VPWR VPWR gpio_configure\[13\]\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_169_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6879_ clknet_leaf_32_csclk net1525 net523 VGND VGND VPWR VPWR gpio_configure\[4\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_139_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold680 _0674_ VGND VGND VPWR VPWR net1213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold691 gpio_configure\[36\]\[3\] VGND VGND VPWR VPWR net1224 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1380 _0739_ VGND VGND VPWR VPWR net1913 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1391 gpio_configure\[29\]\[3\] VGND VGND VPWR VPWR net1924 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput207 net207 VGND VGND VPWR VPWR mgmt_gpio_oeb[4] sky130_fd_sc_hd__buf_12
XFILLER_99_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput218 net218 VGND VGND VPWR VPWR mgmt_gpio_out[14] sky130_fd_sc_hd__clkbuf_1
XFILLER_153_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput229 net229 VGND VGND VPWR VPWR mgmt_gpio_out[24] sky130_fd_sc_hd__buf_12
XFILLER_99_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4230_ wbbd_state\[1\] wbbd_state\[2\] wbbd_state\[4\] wbbd_state\[3\] VGND VGND
+ VPWR VPWR _1528_ sky130_fd_sc_hd__or4_1
XFILLER_141_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4161_ net866 net465 _1516_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__mux2_1
XFILLER_122_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4092_ net1401 net459 net354 VGND VGND VPWR VPWR _1502_ sky130_fd_sc_hd__mux2_1
XFILLER_55_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6802_ clknet_leaf_76_csclk net1086 net488 VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__dfstp_1
XFILLER_51_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4994_ _1653_ _2203_ VGND VGND VPWR VPWR _2204_ sky130_fd_sc_hd__nor2_1
XFILLER_90_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6733_ clknet_leaf_75_csclk net1667 net489 VGND VGND VPWR VPWR gpio_configure\[18\]\[10\]
+ sky130_fd_sc_hd__dfstp_2
X_3945_ net83 clknet_2_1__leaf_mgmt_gpio_in[4] hkspi.pass_thru_mgmt VGND VGND VPWR
+ VPWR net251 sky130_fd_sc_hd__mux2_1
XFILLER_176_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6664_ clknet_leaf_78_csclk net995 net487 VGND VGND VPWR VPWR gpio_configure\[8\]\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_31_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3876_ hkspi.rdstb net476 net483 VGND VGND VPWR VPWR _1428_ sky130_fd_sc_hd__o21a_1
XFILLER_177_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5615_ _0822_ xfer_state\[2\] VGND VGND VPWR VPWR _2462_ sky130_fd_sc_hd__nor2_1
XFILLER_136_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6595_ clknet_leaf_57_csclk net1289 net504 VGND VGND VPWR VPWR mgmt_gpio_data_buf\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_192_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5546_ net464 net1413 _2437_ VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__mux2_1
XFILLER_145_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5477_ net464 net1377 net612 VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__mux2_1
XFILLER_155_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4428_ net126 _1571_ VGND VGND VPWR VPWR _1640_ sky130_fd_sc_hd__nand2_1
Xclkbuf_2_3__f_mgmt_gpio_in[4] clknet_0_mgmt_gpio_in[4] VGND VGND VPWR VPWR clknet_2_3__leaf_mgmt_gpio_in[4]
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_48_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7147_ clknet_3_3_0_wb_clk_i _0750_ net502 VGND VGND VPWR VPWR xfer_count\[3\] sky130_fd_sc_hd__dfrtp_1
Xfanout434 net573 VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__buf_8
Xfanout445 net617 VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__buf_6
XFILLER_101_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4359_ _0836_ _1557_ VGND VGND VPWR VPWR _1571_ sky130_fd_sc_hd__xnor2_2
XFILLER_86_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout456 net457 VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__buf_4
Xfanout467 net468 VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__clkbuf_8
Xfanout489 net491 VGND VGND VPWR VPWR net489 sky130_fd_sc_hd__buf_4
X_7078_ clknet_leaf_22_csclk net676 net515 VGND VGND VPWR VPWR gpio_configure\[29\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6029_ _2478_ _2813_ _2848_ _2849_ VGND VGND VPWR VPWR _2851_ sky130_fd_sc_hd__or4_4
XFILLER_100_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3730_ hkspi.pass_thru_mgmt_delay hkspi.pre_pass_thru_mgmt reset_reg VGND VGND VPWR
+ VPWR net305 sky130_fd_sc_hd__or3_4
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3661_ _1249_ hkspi.ldata\[1\] _0837_ VGND VGND VPWR VPWR _1250_ sky130_fd_sc_hd__mux2_1
XFILLER_118_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5400_ net1544 net440 _2420_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__mux2_1
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6380_ _3174_ net2061 _3162_ VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__mux2_1
X_3592_ net6 _0891_ _0900_ net29 _1144_ VGND VGND VPWR VPWR _1182_ sky130_fd_sc_hd__a221o_2
XFILLER_127_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5331_ net368 net647 VGND VGND VPWR VPWR _2413_ sky130_fd_sc_hd__nand2_8
XFILLER_161_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5262_ net458 net1660 _2405_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__mux2_1
X_7001_ clknet_leaf_58_csclk net1257 net503 VGND VGND VPWR VPWR gpio_configure\[19\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_4213_ net1389 net456 _1523_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__mux2_1
XFILLER_142_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5193_ _1009_ net425 VGND VGND VPWR VPWR _2391_ sky130_fd_sc_hd__nand2_2
XFILLER_68_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4144_ net577 net774 net671 VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__mux2_1
XFILLER_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4075_ net862 net457 net351 VGND VGND VPWR VPWR _1493_ sky130_fd_sc_hd__mux2_1
XFILLER_83_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_4_0_csclk clknet_2_2_0_csclk VGND VGND VPWR VPWR clknet_3_4_0_csclk sky130_fd_sc_hd__clkbuf_8
XFILLER_64_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4977_ _2005_ _2181_ _2186_ VGND VGND VPWR VPWR _2187_ sky130_fd_sc_hd__o21ai_1
X_6716_ clknet_leaf_63_csclk net1819 net501 VGND VGND VPWR VPWR gpio_configure\[37\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_3928_ mgmt_gpio_data\[8\] net67 hkspi.pass_thru_user_delay VGND VGND VPWR VPWR net249
+ sky130_fd_sc_hd__mux2_1
XFILLER_165_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6647_ clknet_3_1_0_wb_clk_i _0260_ VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__dfxtp_1
X_3859_ net58 _1416_ _1419_ net2096 _1423_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__a221o_1
XFILLER_165_746 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6578_ clknet_leaf_14_csclk net1333 net513 VGND VGND VPWR VPWR mgmt_gpio_data\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_124_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5529_ _1041_ net425 VGND VGND VPWR VPWR _2435_ sky130_fd_sc_hd__and2_2
XFILLER_3_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_693 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_74 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap409 _2838_ VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__buf_12
XFILLER_40_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4900_ _1684_ _1779_ VGND VGND VPWR VPWR _2111_ sky130_fd_sc_hd__and2_1
XFILLER_46_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5880_ gpio_configure\[0\]\[8\] _2526_ _2696_ _2706_ net473 VGND VGND VPWR VPWR _2707_
+ sky130_fd_sc_hd__o221a_1
XFILLER_73_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4831_ _1684_ _1850_ _1736_ VGND VGND VPWR VPWR _2042_ sky130_fd_sc_hd__o21ai_1
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_180 clknet_2_0__leaf_mgmt_gpio_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_191 _0933_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4762_ _1584_ _1645_ _1966_ _1973_ VGND VGND VPWR VPWR _1974_ sky130_fd_sc_hd__a211o_1
XFILLER_159_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6501_ clknet_leaf_31_csclk net1024 net523 VGND VGND VPWR VPWR gpio_configure\[31\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_3713_ gpio_configure\[2\]\[1\] _0908_ _0914_ gpio_configure\[5\]\[1\] _1300_ VGND
+ VGND VPWR VPWR _1301_ sky130_fd_sc_hd__a221o_1
XFILLER_146_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4693_ _1602_ _1678_ _1777_ VGND VGND VPWR VPWR _1905_ sky130_fd_sc_hd__or3_1
X_6432_ net493 net481 VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__and2_1
X_3644_ net274 _1009_ _1083_ gpio_configure\[30\]\[10\] _1232_ VGND VGND VPWR VPWR
+ _1233_ sky130_fd_sc_hd__a221o_1
XFILLER_134_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6363_ wbbd_state\[7\] net139 net132 net433 VGND VGND VPWR VPWR _3163_ sky130_fd_sc_hd__a22o_1
X_3575_ gpio_configure\[1\]\[3\] _0934_ _1110_ gpio_configure\[2\]\[11\] _1164_ VGND
+ VGND VPWR VPWR _1165_ sky130_fd_sc_hd__a221o_1
X_5314_ net471 net1584 net556 VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__mux2_1
XFILLER_115_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6294_ serial_data_staging_2\[9\] _2444_ _2485_ VGND VGND VPWR VPWR _3106_ sky130_fd_sc_hd__o21ba_1
XFILLER_114_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5245_ net569 net730 net547 VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__mux2_1
XFILLER_69_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold17 _0845_ VGND VGND VPWR VPWR net550 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold28 _0868_ VGND VGND VPWR VPWR net561 sky130_fd_sc_hd__buf_6
XFILLER_102_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5176_ _1807_ _2233_ _2285_ _1836_ VGND VGND VPWR VPWR _2382_ sky130_fd_sc_hd__o22a_1
XFILLER_152_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold39 net1003 VGND VGND VPWR VPWR net572 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4127_ net439 net760 _1510_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__mux2_1
XFILLER_28_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4058_ net1316 net459 net356 VGND VGND VPWR VPWR _1484_ sky130_fd_sc_hd__mux2_1
XFILLER_45_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_5_0_wb_clk_i clknet_2_2_0_wb_clk_i VGND VGND VPWR VPWR clknet_3_5_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_726 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold509 _0548_ VGND VGND VPWR VPWR net1042 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_440 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3360_ gpio_configure\[32\]\[7\] _0890_ _0953_ _0955_ VGND VGND VPWR VPWR _0956_
+ sky130_fd_sc_hd__a211o_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3291_ net1971 net561 VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__nand2_8
XFILLER_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5030_ _2229_ _2230_ _2232_ _2239_ VGND VGND VPWR VPWR _2240_ sky130_fd_sc_hd__or4b_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1209 net2143 VGND VGND VPWR VPWR net1742 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6981_ clknet_leaf_36_csclk net1137 net522 VGND VGND VPWR VPWR gpio_configure\[17\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_19_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5932_ gpio_configure\[18\]\[11\] _2532_ _2755_ VGND VGND VPWR VPWR _2756_ sky130_fd_sc_hd__a21o_1
XFILLER_80_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5863_ gpio_configure\[10\]\[8\] net421 _2523_ gpio_configure\[2\]\[8\] VGND VGND
+ VPWR VPWR _2690_ sky130_fd_sc_hd__a22o_1
XFILLER_178_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4814_ net477 _1782_ _1787_ VGND VGND VPWR VPWR _2025_ sky130_fd_sc_hd__or3_1
XFILLER_21_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5794_ net475 net2034 _2624_ VGND VGND VPWR VPWR _2625_ sky130_fd_sc_hd__a21o_1
XFILLER_119_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4745_ _1576_ _1643_ VGND VGND VPWR VPWR _1957_ sky130_fd_sc_hd__nor2_1
XFILLER_193_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4676_ _1790_ _1874_ _1886_ _1800_ VGND VGND VPWR VPWR _1888_ sky130_fd_sc_hd__o22a_1
XFILLER_107_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6415_ net486 net481 VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__and2_1
X_3627_ _1212_ _1213_ _1214_ _1215_ VGND VGND VPWR VPWR _1216_ sky130_fd_sc_hd__or4_1
XFILLER_134_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6346_ _0818_ wbbd_state\[6\] VGND VGND VPWR VPWR _3155_ sky130_fd_sc_hd__nand2_1
X_3558_ gpio_configure\[10\]\[3\] _0920_ _1102_ gpio_configure\[15\]\[11\] VGND VGND
+ VPWR VPWR _1148_ sky130_fd_sc_hd__a22o_1
XFILLER_1_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6277_ gpio_configure\[18\]\[10\] _2819_ _2837_ gpio_configure\[8\]\[10\] VGND VGND
+ VPWR VPWR _3089_ sky130_fd_sc_hd__a22o_1
XFILLER_130_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3489_ net382 _0909_ VGND VGND VPWR VPWR _1080_ sky130_fd_sc_hd__nor2_4
Xinput107 wb_adr_i[17] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput118 wb_adr_i[27] VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_1
X_5228_ net1512 net471 _2400_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__mux2_1
Xinput129 wb_adr_i[8] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_1
XFILLER_56_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5159_ _2268_ _2335_ _2365_ VGND VGND VPWR VPWR _2366_ sky130_fd_sc_hd__nand3_1
XFILLER_84_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_2_1_0_csclk clknet_1_0_1_csclk VGND VGND VPWR VPWR clknet_2_1_0_csclk sky130_fd_sc_hd__clkbuf_8
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_80 _2986_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_91 hkspi.pass_thru_user VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4530_ _1687_ _1699_ _1740_ _1741_ VGND VGND VPWR VPWR _1742_ sky130_fd_sc_hd__and4_1
XFILLER_7_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold306 _0631_ VGND VGND VPWR VPWR net839 sky130_fd_sc_hd__dlygate4sd3_1
X_4461_ _1581_ _1606_ VGND VGND VPWR VPWR _1673_ sky130_fd_sc_hd__nor2_1
Xhold317 gpio_configure\[18\]\[2\] VGND VGND VPWR VPWR net850 sky130_fd_sc_hd__dlygate4sd3_1
Xhold328 _0340_ VGND VGND VPWR VPWR net861 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6200_ gpio_configure\[7\]\[7\] _2811_ net407 gpio_configure\[15\]\[7\] VGND VGND
+ VPWR VPWR _3015_ sky130_fd_sc_hd__a22o_1
Xhold339 gpio_configure\[8\]\[1\] VGND VGND VPWR VPWR net872 sky130_fd_sc_hd__dlygate4sd3_1
X_3412_ _1005_ net2004 _0970_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__mux2_1
X_7180_ clknet_3_3_0_wb_clk_i net2043 net506 VGND VGND VPWR VPWR serial_data_staging_2\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_4392_ net114 net113 _1434_ _1601_ VGND VGND VPWR VPWR _1604_ sky130_fd_sc_hd__a31o_2
XFILLER_171_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6131_ gpio_configure\[14\]\[4\] net411 net406 gpio_configure\[27\]\[4\] VGND VGND
+ VPWR VPWR _2949_ sky130_fd_sc_hd__a22o_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ net376 _0889_ VGND VGND VPWR VPWR _0939_ sky130_fd_sc_hd__nor2_8
XFILLER_97_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6062_ gpio_configure\[10\]\[1\] net414 net394 gpio_configure\[6\]\[1\] _2882_ VGND
+ VGND VPWR VPWR _2883_ sky130_fd_sc_hd__a221o_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ net561 net600 VGND VGND VPWR VPWR _0870_ sky130_fd_sc_hd__nand2_8
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1006 _0562_ VGND VGND VPWR VPWR net1539 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1017 gpio_configure\[11\]\[2\] VGND VGND VPWR VPWR net1550 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _1693_ net424 VGND VGND VPWR VPWR _2223_ sky130_fd_sc_hd__or2_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1028 _0735_ VGND VGND VPWR VPWR net1561 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1039 net2095 VGND VGND VPWR VPWR net1572 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6964_ clknet_leaf_23_csclk net1349 net514 VGND VGND VPWR VPWR gpio_configure\[15\]\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_5915_ gpio_configure\[13\]\[10\] _2501_ _2532_ gpio_configure\[18\]\[10\] _2739_
+ VGND VGND VPWR VPWR _2740_ sky130_fd_sc_hd__a221o_1
X_6895_ clknet_leaf_39_csclk net1107 net516 VGND VGND VPWR VPWR gpio_configure\[6\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5846_ gpio_configure\[5\]\[7\] net422 _2501_ gpio_configure\[13\]\[7\] _2673_ VGND
+ VGND VPWR VPWR _2674_ sky130_fd_sc_hd__a221o_1
XFILLER_42_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5777_ gpio_configure\[24\]\[4\] _2531_ _2532_ gpio_configure\[18\]\[4\] VGND VGND
+ VPWR VPWR _2608_ sky130_fd_sc_hd__a22o_1
X_4728_ _1598_ _1706_ VGND VGND VPWR VPWR _1940_ sky130_fd_sc_hd__nor2_1
XFILLER_147_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4659_ _1588_ _1807_ VGND VGND VPWR VPWR _1871_ sky130_fd_sc_hd__nor2_1
XFILLER_162_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold840 mgmt_gpio_data\[13\] VGND VGND VPWR VPWR net1373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold851 _0662_ VGND VGND VPWR VPWR net1384 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_107_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold862 gpio_configure\[30\]\[1\] VGND VGND VPWR VPWR net1395 sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 _0375_ VGND VGND VPWR VPWR net1406 sky130_fd_sc_hd__dlygate4sd3_1
Xhold884 gpio_configure\[14\]\[6\] VGND VGND VPWR VPWR net1417 sky130_fd_sc_hd__dlygate4sd3_1
X_6329_ gpio_configure\[8\]\[12\] net410 net405 gpio_configure\[24\]\[12\] VGND VGND
+ VPWR VPWR _3139_ sky130_fd_sc_hd__a22o_1
XFILLER_115_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold895 _0284_ VGND VGND VPWR VPWR net1428 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_107_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1540 serial_data_staging_1\[10\] VGND VGND VPWR VPWR net2073 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1551 pad_count_2\[2\] VGND VGND VPWR VPWR net2084 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1562 mgmt_gpio_data\[1\] VGND VGND VPWR VPWR net2095 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1573 mgmt_gpio_data\[37\] VGND VGND VPWR VPWR net2106 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1584 serial_data_staging_2\[12\] VGND VGND VPWR VPWR net2117 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_177_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1595 mgmt_gpio_data_buf\[5\] VGND VGND VPWR VPWR net2128 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_32_csclk clknet_3_7_0_csclk VGND VGND VPWR VPWR clknet_leaf_32_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_79_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_47_csclk clknet_3_6_0_csclk VGND VGND VPWR VPWR clknet_leaf_47_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_36_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3961_ irq_2_inputsrc net39 VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__and2_2
XFILLER_189_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5700_ pad_count_1\[4\] _2461_ _2488_ VGND VGND VPWR VPWR _2535_ sky130_fd_sc_hd__and3_4
XFILLER_50_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6680_ clknet_3_7_0_wb_clk_i _0293_ net528 VGND VGND VPWR VPWR wbbd_busy sky130_fd_sc_hd__dfrtp_4
X_3892_ wbbd_state\[7\] _1428_ net2032 VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__a21o_1
XFILLER_176_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5631_ pad_count_2\[2\] _2463_ _2470_ VGND VGND VPWR VPWR _2472_ sky130_fd_sc_hd__a21oi_1
XFILLER_148_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5562_ _0932_ net647 VGND VGND VPWR VPWR _2439_ sky130_fd_sc_hd__nand2_4
XFILLER_129_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4513_ _1652_ _1662_ VGND VGND VPWR VPWR _1725_ sky130_fd_sc_hd__nand2_1
XFILLER_191_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold103 hkspi.addr\[4\] VGND VGND VPWR VPWR net636 sky130_fd_sc_hd__dlygate4sd3_1
X_5493_ net370 net647 VGND VGND VPWR VPWR _2431_ sky130_fd_sc_hd__nand2_8
Xhold114 net428 VGND VGND VPWR VPWR net647 sky130_fd_sc_hd__buf_12
Xhold125 hkspi.odata\[5\] VGND VGND VPWR VPWR net658 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4444_ _1625_ _1627_ VGND VGND VPWR VPWR _1656_ sky130_fd_sc_hd__nand2b_2
Xhold136 net474 VGND VGND VPWR VPWR net669 sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 _0327_ VGND VGND VPWR VPWR net680 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 wbbd_data\[3\] VGND VGND VPWR VPWR net691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold169 gpio_configure\[4\]\[11\] VGND VGND VPWR VPWR net702 sky130_fd_sc_hd__dlygate4sd3_1
X_7163_ clknet_3_0_0_wb_clk_i net2030 net508 VGND VGND VPWR VPWR serial_data_staging_1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_113_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4375_ net110 net124 net99 VGND VGND VPWR VPWR _1587_ sky130_fd_sc_hd__nor3b_2
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6114_ gpio_configure\[10\]\[3\] _2825_ net394 gpio_configure\[6\]\[3\] _2932_ VGND
+ VGND VPWR VPWR _2933_ sky130_fd_sc_hd__a221o_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3326_ _0881_ net386 VGND VGND VPWR VPWR _0922_ sky130_fd_sc_hd__nor2_8
XFILLER_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7094_ clknet_leaf_5_csclk net1229 net494 VGND VGND VPWR VPWR gpio_configure\[31\]\[12\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _2808_ _2834_ _2866_ VGND VGND VPWR VPWR _2867_ sky130_fd_sc_hd__or3_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3257_ net549 net597 net605 VGND VGND VPWR VPWR _0853_ sky130_fd_sc_hd__mux2_1
XTAP_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3188_ net2086 VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__inv_2
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6947_ clknet_leaf_21_csclk net1372 net514 VGND VGND VPWR VPWR gpio_configure\[13\]\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_41_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6878_ clknet_leaf_26_csclk net723 net519 VGND VGND VPWR VPWR gpio_configure\[4\]\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_5829_ gpio_configure\[9\]\[6\] _2512_ net419 _2657_ VGND VGND VPWR VPWR _2658_ sky130_fd_sc_hd__a22o_1
XFILLER_139_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold670 _0238_ VGND VGND VPWR VPWR net1203 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold681 gpio_configure\[21\]\[0\] VGND VGND VPWR VPWR net1214 sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 _0733_ VGND VGND VPWR VPWR net1225 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1370 mgmt_gpio_data_buf\[21\] VGND VGND VPWR VPWR net1903 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1381 clk2_output_dest VGND VGND VPWR VPWR net1914 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1392 wbbd_data\[4\] VGND VGND VPWR VPWR net1925 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput208 net208 VGND VGND VPWR VPWR mgmt_gpio_oeb[5] sky130_fd_sc_hd__buf_12
XFILLER_154_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput219 net219 VGND VGND VPWR VPWR mgmt_gpio_out[15] sky130_fd_sc_hd__clkbuf_1
XFILLER_5_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4160_ net1787 net470 _1516_ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__mux2_1
XFILLER_4_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4091_ net662 _1501_ _1499_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__mux2_1
XFILLER_83_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6801_ clknet_leaf_76_csclk net1127 net488 VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__dfrtp_4
XFILLER_90_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4993_ _1584_ _1703_ VGND VGND VPWR VPWR _2203_ sky130_fd_sc_hd__nor2_4
XFILLER_23_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6732_ clknet_leaf_75_csclk net1695 net489 VGND VGND VPWR VPWR gpio_configure\[18\]\[9\]
+ sky130_fd_sc_hd__dfrtp_2
X_3944_ hkspi.pass_thru_mgmt_delay net487 VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__nor2_1
X_6663_ clknet_leaf_78_csclk net1028 net485 VGND VGND VPWR VPWR gpio_configure\[8\]\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_3875_ serial_clock_pre serial_bb_clock serial_bb_enable VGND VGND VPWR VPWR net307
+ sky130_fd_sc_hd__mux2_4
XFILLER_139_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5614_ pad_count_1\[1\] pad_count_1\[0\] VGND VGND VPWR VPWR _2461_ sky130_fd_sc_hd__and2_2
X_6594_ clknet_leaf_78_csclk net761 net486 VGND VGND VPWR VPWR mgmt_gpio_data_buf\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_164_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5545_ net471 net1602 _2437_ VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__mux2_1
XFILLER_145_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_0_0_csclk clknet_2_0_0_csclk VGND VGND VPWR VPWR clknet_3_0_0_csclk sky130_fd_sc_hd__clkbuf_8
X_5476_ net468 net1814 net612 VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__mux2_1
XFILLER_144_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7215_ net66 VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__buf_2
X_4427_ _1558_ _1565_ _1567_ _1559_ VGND VGND VPWR VPWR _1639_ sky130_fd_sc_hd__a211o_2
XFILLER_160_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7146_ clknet_3_3_0_wb_clk_i _0749_ net502 VGND VGND VPWR VPWR xfer_count\[2\] sky130_fd_sc_hd__dfrtp_1
Xfanout424 _1775_ VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__buf_6
X_4358_ net125 _1557_ VGND VGND VPWR VPWR _1570_ sky130_fd_sc_hd__and2_1
Xfanout435 net573 VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__buf_6
Xfanout446 net618 VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__buf_6
XFILLER_58_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout457 net576 VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__buf_8
X_3309_ net581 net551 net638 VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__or3b_4
Xfanout468 net469 VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__clkbuf_4
XFILLER_100_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7077_ clknet_leaf_50_csclk net693 net506 VGND VGND VPWR VPWR gpio_configure\[29\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_4289_ net470 net1690 _1540_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__mux2_1
XFILLER_86_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6028_ _2478_ _2813_ _2848_ _2849_ VGND VGND VPWR VPWR _2850_ sky130_fd_sc_hd__nor4_1
XFILLER_39_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3660_ _1222_ _1231_ _1248_ VGND VGND VPWR VPWR _1249_ sky130_fd_sc_hd__or3_4
X_3591_ net285 _0886_ _0910_ net294 _1150_ VGND VGND VPWR VPWR _1181_ sky130_fd_sc_hd__a221o_1
XFILLER_127_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5330_ net908 net435 _2412_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__mux2_1
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5261_ net464 net1461 _2405_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__mux2_1
XFILLER_88_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7000_ clknet_leaf_58_csclk net1426 net503 VGND VGND VPWR VPWR gpio_configure\[19\]\[6\]
+ sky130_fd_sc_hd__dfrtp_2
X_4212_ net1736 net461 _1523_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__mux2_1
X_5192_ net443 net1011 _2390_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__mux2_1
XFILLER_68_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4143_ net465 net822 net671 VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__mux2_1
XFILLER_68_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4074_ net1572 _1492_ _1490_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__mux2_1
XFILLER_71_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4976_ net424 _1779_ _1823_ VGND VGND VPWR VPWR _2186_ sky130_fd_sc_hd__a21o_1
X_6715_ clknet_leaf_8_csclk net1149 net509 VGND VGND VPWR VPWR gpio_configure\[16\]\[12\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_189_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3927_ mgmt_gpio_data\[9\] clknet_2_0__leaf_mgmt_gpio_in[4] hkspi.pass_thru_user
+ VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__mux2_1
XFILLER_20_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3858_ hkspi.state\[0\] _1420_ VGND VGND VPWR VPWR _1423_ sky130_fd_sc_hd__and2b_1
X_6646_ clknet_3_5_0_wb_clk_i _0259_ VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__dfxtp_1
XFILLER_149_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3789_ _1352_ _1358_ _1367_ _1374_ VGND VGND VPWR VPWR _1375_ sky130_fd_sc_hd__or4_1
X_6577_ clknet_leaf_0_csclk net1233 net486 VGND VGND VPWR VPWR mgmt_gpio_data\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_164_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5528_ net435 net948 _2434_ VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__mux2_1
X_5459_ net465 net874 _2427_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__mux2_1
XFILLER_59_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7129_ clknet_leaf_24_csclk net1653 net518 VGND VGND VPWR VPWR gpio_configure\[36\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_47_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_170 net458 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4830_ _1581_ _1678_ _1680_ VGND VGND VPWR VPWR _2041_ sky130_fd_sc_hd__a21oi_1
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_181 clknet_2_0__leaf_mgmt_gpio_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_192 _0972_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4761_ _1945_ _1968_ _1969_ _1972_ VGND VGND VPWR VPWR _1973_ sky130_fd_sc_hd__or4b_1
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3712_ net96 _1137_ _1299_ net292 VGND VGND VPWR VPWR _1300_ sky130_fd_sc_hd__a22o_1
X_6500_ clknet_leaf_25_csclk net1727 net518 VGND VGND VPWR VPWR gpio_configure\[31\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_119_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4692_ _1787_ _1886_ VGND VGND VPWR VPWR _1904_ sky130_fd_sc_hd__or2_1
XFILLER_174_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3643_ gpio_configure\[27\]\[10\] _1076_ _1117_ net268 VGND VGND VPWR VPWR _1232_
+ sky130_fd_sc_hd__a22o_1
X_6431_ net493 net481 VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__and2_1
XFILLER_147_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6362_ _1529_ _3161_ _3159_ _3160_ VGND VGND VPWR VPWR _3162_ sky130_fd_sc_hd__or4b_4
X_3574_ gpio_configure\[12\]\[11\] _1056_ _1069_ gpio_configure\[14\]\[11\] VGND VGND
+ VPWR VPWR _1164_ sky130_fd_sc_hd__a22o_1
X_5313_ net555 net428 VGND VGND VPWR VPWR _2411_ sky130_fd_sc_hd__nand2_4
XFILLER_114_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6293_ gpio_configure\[0\]\[10\] _2851_ _3092_ _3104_ net473 VGND VGND VPWR VPWR
+ _3105_ sky130_fd_sc_hd__o221a_1
XFILLER_115_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5244_ net459 net1401 net547 VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__mux2_1
XFILLER_102_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold18 _0847_ VGND VGND VPWR VPWR net551 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 _0887_ VGND VGND VPWR VPWR net562 sky130_fd_sc_hd__buf_6
XFILLER_130_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5175_ _2344_ _2380_ _2355_ VGND VGND VPWR VPWR _2381_ sky130_fd_sc_hd__o21a_1
XFILLER_69_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4126_ net660 net726 _1510_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__mux2_1
XFILLER_84_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4057_ net958 _1483_ _1481_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__mux2_1
XFILLER_83_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4959_ _2165_ _2166_ _2168_ VGND VGND VPWR VPWR _2169_ sky130_fd_sc_hd__and3_1
XFILLER_177_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6629_ clknet_3_5_0_wb_clk_i _0242_ VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__dfxtp_1
XFILLER_192_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3290_ net389 _0885_ VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__nor2_8
XFILLER_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_704 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6980_ clknet_leaf_67_csclk net781 net505 VGND VGND VPWR VPWR gpio_configure\[17\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_80_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5931_ gpio_configure\[3\]\[11\] _2518_ _2535_ gpio_configure\[23\]\[11\] VGND VGND
+ VPWR VPWR _2755_ sky130_fd_sc_hd__a22o_1
XFILLER_179_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5862_ gpio_configure\[27\]\[8\] _2506_ _2517_ gpio_configure\[30\]\[8\] _2688_ VGND
+ VGND VPWR VPWR _2689_ sky130_fd_sc_hd__a221o_1
XFILLER_61_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4813_ _1999_ _2012_ _2015_ _2023_ VGND VGND VPWR VPWR _2024_ sky130_fd_sc_hd__or4_1
X_5793_ gpio_configure\[0\]\[4\] _2526_ _2616_ _2623_ _0824_ VGND VGND VPWR VPWR _2624_
+ sky130_fd_sc_hd__o221a_4
XFILLER_21_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4744_ _1617_ _1628_ _1648_ VGND VGND VPWR VPWR _1956_ sky130_fd_sc_hd__and3_1
XFILLER_159_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4675_ _1800_ _1886_ VGND VGND VPWR VPWR _1887_ sky130_fd_sc_hd__nor2_1
XFILLER_147_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6414_ net486 net481 VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__and2_1
X_3626_ net54 _0871_ _1081_ gpio_configure\[34\]\[10\] _1203_ VGND VGND VPWR VPWR
+ _1215_ sky130_fd_sc_hd__a221o_1
XFILLER_147_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3557_ gpio_configure\[23\]\[3\] _0922_ net367 gpio_configure\[17\]\[3\] VGND VGND
+ VPWR VPWR _1147_ sky130_fd_sc_hd__a22o_1
X_6345_ _0818_ net431 wbbd_state\[1\] VGND VGND VPWR VPWR _3154_ sky130_fd_sc_hd__o21a_1
X_6276_ gpio_configure\[23\]\[10\] _2822_ _2828_ gpio_configure\[20\]\[10\] _3084_
+ VGND VGND VPWR VPWR _3088_ sky130_fd_sc_hd__a221o_1
XFILLER_115_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3488_ gpio_configure\[4\]\[4\] net350 _1007_ net65 VGND VGND VPWR VPWR _1079_ sky130_fd_sc_hd__a22o_1
XFILLER_130_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5227_ net1914 net542 _2400_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__mux2_1
Xinput108 wb_adr_i[18] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_1
Xinput119 wb_adr_i[28] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_1
XFILLER_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5158_ _1883_ _1988_ _2163_ VGND VGND VPWR VPWR _2365_ sky130_fd_sc_hd__nor3_1
XFILLER_84_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4109_ net447 net1332 _1508_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__mux2_1
X_5089_ _1651_ _1707_ _1807_ net432 VGND VGND VPWR VPWR _2298_ sky130_fd_sc_hd__o22a_1
XFILLER_71_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_70 _2537_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_81 _3107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_92 mask_rev_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4460_ _1645_ _1670_ VGND VGND VPWR VPWR _1672_ sky130_fd_sc_hd__nand2_1
Xhold307 gpio_configure\[29\]\[2\] VGND VGND VPWR VPWR net840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold318 _0591_ VGND VGND VPWR VPWR net851 sky130_fd_sc_hd__dlygate4sd3_1
Xhold329 mgmt_gpio_data_buf\[2\] VGND VGND VPWR VPWR net862 sky130_fd_sc_hd__dlygate4sd3_1
X_3411_ _1004_ net2001 _0837_ VGND VGND VPWR VPWR _1005_ sky130_fd_sc_hd__mux2_1
XFILLER_144_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4391_ net114 net113 _1434_ _1601_ VGND VGND VPWR VPWR _1603_ sky130_fd_sc_hd__a31oi_2
XFILLER_98_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6130_ gpio_configure\[22\]\[4\] net397 _2829_ gpio_configure\[33\]\[4\] _2947_ VGND
+ VGND VPWR VPWR _2948_ sky130_fd_sc_hd__a221o_1
X_3342_ net378 net609 VGND VGND VPWR VPWR _0938_ sky130_fd_sc_hd__nor2_8
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ gpio_configure\[9\]\[1\] net412 net409 gpio_configure\[12\]\[1\] VGND VGND
+ VPWR VPWR _2882_ sky130_fd_sc_hd__a22o_1
X_3273_ net599 net607 VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__and2b_4
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1007 net2131 VGND VGND VPWR VPWR net1540 sky130_fd_sc_hd__dlygate4sd3_1
X_5012_ _1589_ net478 _1596_ _2110_ VGND VGND VPWR VPWR _2222_ sky130_fd_sc_hd__a31o_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1018 _0535_ VGND VGND VPWR VPWR net1551 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 gpio_configure\[34\]\[0\] VGND VGND VPWR VPWR net1562 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6963_ clknet_leaf_8_csclk net849 net509 VGND VGND VPWR VPWR gpio_configure\[15\]\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_5914_ gpio_configure\[27\]\[10\] _2506_ _2541_ gpio_configure\[31\]\[10\] VGND VGND
+ VPWR VPWR _2739_ sky130_fd_sc_hd__a22o_1
XFILLER_62_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6894_ clknet_leaf_15_csclk net1197 net513 VGND VGND VPWR VPWR gpio_configure\[6\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_5845_ gpio_configure\[3\]\[7\] _2518_ _2538_ gpio_configure\[1\]\[7\] VGND VGND
+ VPWR VPWR _2673_ sky130_fd_sc_hd__a22o_1
XFILLER_22_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5776_ gpio_configure\[9\]\[4\] _2512_ _2529_ gpio_configure\[29\]\[4\] VGND VGND
+ VPWR VPWR _2607_ sky130_fd_sc_hd__a22o_1
XFILLER_158_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4727_ _1613_ _1644_ _1938_ wbbd_state\[7\] VGND VGND VPWR VPWR _1939_ sky130_fd_sc_hd__o31a_1
XFILLER_175_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4658_ _1592_ _1795_ VGND VGND VPWR VPWR _1870_ sky130_fd_sc_hd__or2_1
XFILLER_135_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput90 spimemio_flash_io2_oeb VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_2
Xhold830 gpio_configure\[29\]\[10\] VGND VGND VPWR VPWR net1363 sky130_fd_sc_hd__dlygate4sd3_1
X_3609_ gpio_configure\[9\]\[2\] _0930_ _1129_ gpio_configure\[11\]\[10\] VGND VGND
+ VPWR VPWR _1198_ sky130_fd_sc_hd__a22o_1
Xhold841 _0184_ VGND VGND VPWR VPWR net1374 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold852 gpio_configure\[30\]\[6\] VGND VGND VPWR VPWR net1385 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4589_ net477 _1800_ VGND VGND VPWR VPWR _1801_ sky130_fd_sc_hd__or2_4
XFILLER_150_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold863 _0686_ VGND VGND VPWR VPWR net1396 sky130_fd_sc_hd__dlygate4sd3_1
Xhold874 gpio_configure\[14\]\[10\] VGND VGND VPWR VPWR net1407 sky130_fd_sc_hd__dlygate4sd3_1
X_6328_ gpio_configure\[1\]\[12\] _2802_ _2860_ gpio_configure\[17\]\[12\] _3137_
+ VGND VGND VPWR VPWR _3138_ sky130_fd_sc_hd__a221o_1
Xhold885 _0563_ VGND VGND VPWR VPWR net1418 sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 gpio_configure\[36\]\[1\] VGND VGND VPWR VPWR net1429 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6259_ gpio_configure\[34\]\[9\] net393 _2852_ gpio_configure\[19\]\[9\] _3071_ VGND
+ VGND VPWR VPWR _3072_ sky130_fd_sc_hd__a221o_1
XFILLER_29_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1530 serial_data_staging_1\[8\] VGND VGND VPWR VPWR net2063 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1541 serial_load_pre VGND VGND VPWR VPWR net2074 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1552 hkspi.addr\[3\] VGND VGND VPWR VPWR net2085 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_91_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1563 hkspi.fixed\[0\] VGND VGND VPWR VPWR net2096 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1574 pad_count_2\[1\] VGND VGND VPWR VPWR net2107 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1585 gpio_configure\[32\]\[2\] VGND VGND VPWR VPWR net2118 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1596 gpio_configure\[34\]\[6\] VGND VGND VPWR VPWR net2129 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3960_ irq_1_inputsrc net70 VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__and2_2
XFILLER_51_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3891_ hkspi.state\[0\] _1385_ _1441_ hkspi.state\[2\] VGND VGND VPWR VPWR _0004_
+ sky130_fd_sc_hd__a22o_1
XFILLER_189_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5630_ _0825_ _1448_ _2471_ _2458_ net2107 VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__o32a_1
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5561_ net435 net966 _2438_ VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__mux2_1
XFILLER_117_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4512_ _1612_ _1654_ VGND VGND VPWR VPWR _1724_ sky130_fd_sc_hd__nand2_1
X_5492_ net434 net1272 _2430_ VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__mux2_1
XFILLER_184_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold104 _0849_ VGND VGND VPWR VPWR net637 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_156_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold115 _2439_ VGND VGND VPWR VPWR net648 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_105_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold126 net665 VGND VGND VPWR VPWR net659 sky130_fd_sc_hd__dlygate4sd3_1
X_4443_ _1623_ _1647_ VGND VGND VPWR VPWR _1655_ sky130_fd_sc_hd__or2_4
XFILLER_171_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold137 _1459_ VGND VGND VPWR VPWR net670 sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 gpio_configure\[16\]\[11\] VGND VGND VPWR VPWR net681 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold159 _1465_ VGND VGND VPWR VPWR net692 sky130_fd_sc_hd__dlygate4sd3_1
X_7162_ clknet_3_0_0_wb_clk_i _0764_ net508 VGND VGND VPWR VPWR serial_data_staging_1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_4374_ _1576_ _1585_ VGND VGND VPWR VPWR _1586_ sky130_fd_sc_hd__nor2_1
XFILLER_171_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3325_ net562 net381 VGND VGND VPWR VPWR _0921_ sky130_fd_sc_hd__nor2_8
X_6113_ gpio_configure\[12\]\[3\] net409 net405 gpio_configure\[24\]\[3\] VGND VGND
+ VPWR VPWR _2932_ sky130_fd_sc_hd__a22o_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7093_ clknet_leaf_1_csclk net1325 net496 VGND VGND VPWR VPWR gpio_configure\[31\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3256_ net389 VGND VGND VPWR VPWR _0852_ sky130_fd_sc_hd__inv_2
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6044_ net360 _2854_ _2857_ _2865_ VGND VGND VPWR VPWR _2866_ sky130_fd_sc_hd__or4_4
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3187_ net111 VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__clkinv_2
XFILLER_94_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6946_ clknet_leaf_25_csclk net1583 net518 VGND VGND VPWR VPWR gpio_configure\[13\]\[0\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_41_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6877_ clknet_leaf_29_csclk net991 net520 VGND VGND VPWR VPWR gpio_configure\[4\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_22_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5828_ gpio_configure\[16\]\[6\] _0831_ VGND VGND VPWR VPWR _2657_ sky130_fd_sc_hd__or2_1
XFILLER_167_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5759_ gpio_configure\[20\]\[3\] _2499_ _2523_ gpio_configure\[2\]\[3\] VGND VGND
+ VPWR VPWR _2591_ sky130_fd_sc_hd__a22o_1
XFILLER_135_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold660 _0576_ VGND VGND VPWR VPWR net1193 sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 gpio_configure\[28\]\[12\] VGND VGND VPWR VPWR net1204 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold682 _0613_ VGND VGND VPWR VPWR net1215 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold693 gpio_configure\[6\]\[11\] VGND VGND VPWR VPWR net1226 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_618 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1360 net1893 VGND VGND VPWR VPWR wb_dat_o[20] sky130_fd_sc_hd__buf_12
XFILLER_45_523 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1371 mgmt_gpio_data_buf\[23\] VGND VGND VPWR VPWR net1904 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1382 gpio_configure\[12\]\[11\] VGND VGND VPWR VPWR net1915 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1393 gpio_configure\[10\]\[10\] VGND VGND VPWR VPWR net1926 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput209 net209 VGND VGND VPWR VPWR mgmt_gpio_oeb[6] sky130_fd_sc_hd__buf_12
XFILLER_5_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4090_ net1906 net542 net354 VGND VGND VPWR VPWR _1501_ sky130_fd_sc_hd__mux2_1
XFILLER_95_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6800_ clknet_leaf_76_csclk net1697 net484 VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__dfrtp_2
XFILLER_91_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4992_ _2086_ _1933_ _1939_ VGND VGND VPWR VPWR _2202_ sky130_fd_sc_hd__and3b_1
X_6731_ clknet_leaf_75_csclk net1712 net489 VGND VGND VPWR VPWR gpio_configure\[18\]\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_3943_ net84 net67 hkspi.pass_thru_mgmt_delay VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__mux2_2
XFILLER_16_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6662_ clknet_leaf_78_csclk net1985 net487 VGND VGND VPWR VPWR gpio_configure\[8\]\[10\]
+ sky130_fd_sc_hd__dfstp_4
XFILLER_31_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3874_ hkspi.writemode net2015 hkspi.state\[2\] _1384_ VGND VGND VPWR VPWR _0065_
+ sky130_fd_sc_hd__o211a_1
XFILLER_149_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5613_ xfer_state\[2\] _2459_ VGND VGND VPWR VPWR _2460_ sky130_fd_sc_hd__nand2_1
X_6593_ clknet_leaf_54_csclk net727 net506 VGND VGND VPWR VPWR mgmt_gpio_data_buf\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_191_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5544_ _0938_ net647 VGND VGND VPWR VPWR _2437_ sky130_fd_sc_hd__nand2_8
XFILLER_145_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5475_ net611 net647 VGND VGND VPWR VPWR _2429_ sky130_fd_sc_hd__nand2_8
XFILLER_117_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7214_ net65 VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__clkbuf_1
XFILLER_160_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4426_ _1572_ _1573_ VGND VGND VPWR VPWR _1638_ sky130_fd_sc_hd__nand2_1
X_7145_ clknet_3_2_0_wb_clk_i _0748_ net502 VGND VGND VPWR VPWR xfer_count\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_99_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout425 net426 VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__buf_12
XFILLER_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4357_ net125 _1557_ VGND VGND VPWR VPWR _1569_ sky130_fd_sc_hd__nor2_1
Xfanout436 net572 VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__buf_6
XFILLER_86_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout447 net618 VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__buf_4
X_3308_ net629 _0903_ VGND VGND VPWR VPWR _0904_ sky130_fd_sc_hd__nor2_8
Xfanout458 net459 VGND VGND VPWR VPWR net458 sky130_fd_sc_hd__clkbuf_8
X_7076_ clknet_leaf_64_csclk net841 net501 VGND VGND VPWR VPWR gpio_configure\[29\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout469 net1098 VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__buf_8
XFILLER_86_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4288_ _1051_ net429 VGND VGND VPWR VPWR _1540_ sky130_fd_sc_hd__nand2_2
XFILLER_100_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6027_ net401 _2825_ _2835_ net392 VGND VGND VPWR VPWR _2849_ sky130_fd_sc_hd__or4_1
X_3239_ net126 VGND VGND VPWR VPWR _0835_ sky130_fd_sc_hd__inv_2
XFILLER_86_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6929_ clknet_leaf_41_csclk net1054 net517 VGND VGND VPWR VPWR gpio_configure\[10\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_31_csclk clknet_3_7_0_csclk VGND VGND VPWR VPWR clknet_leaf_31_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_168_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_46_csclk clknet_3_6_0_csclk VGND VGND VPWR VPWR clknet_leaf_46_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold490 gpio_configure\[31\]\[3\] VGND VGND VPWR VPWR net1023 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_1_0_0_wb_clk_i clknet_0_wb_clk_i VGND VGND VPWR VPWR clknet_1_0_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_150_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1190 _0163_ VGND VGND VPWR VPWR net1723 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3590_ gpio_configure\[29\]\[3\] _0917_ _1087_ gpio_configure\[0\]\[11\] _1151_ VGND
+ VGND VPWR VPWR _1180_ sky130_fd_sc_hd__a221o_1
XFILLER_139_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5260_ net470 net1763 _2405_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__mux2_1
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4211_ net1812 net466 _1523_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__mux2_1
X_5191_ net449 net1067 _2390_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__mux2_1
XFILLER_142_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4142_ net470 net1700 net671 VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__mux2_1
XFILLER_96_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4073_ net1455 net462 _0933_ VGND VGND VPWR VPWR _1492_ sky130_fd_sc_hd__mux2_1
XFILLER_49_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4975_ _1744_ _1771_ _1818_ _2184_ _1786_ VGND VGND VPWR VPWR _2185_ sky130_fd_sc_hd__a311o_1
X_6714_ clknet_leaf_9_csclk net682 net509 VGND VGND VPWR VPWR gpio_configure\[16\]\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_51_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3926_ mgmt_gpio_data\[10\] net58 hkspi.pass_thru_user_delay VGND VGND VPWR VPWR
+ net214 sky130_fd_sc_hd__mux2_1
XFILLER_20_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6645_ clknet_3_5_0_wb_clk_i _0258_ VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__dfxtp_1
X_3857_ _1420_ _1422_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__xnor2_1
XFILLER_165_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6576_ clknet_leaf_27_csclk net815 net519 VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__dfrtp_2
X_3788_ _1368_ _1370_ _1372_ _1373_ VGND VGND VPWR VPWR _1374_ sky130_fd_sc_hd__or4_1
XFILLER_152_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5527_ net438 net1385 _2434_ VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__mux2_1
XFILLER_192_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_634 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5458_ net469 net1596 _2427_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__mux2_1
XFILLER_172_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4409_ _1553_ _1610_ _1620_ VGND VGND VPWR VPWR _1621_ sky130_fd_sc_hd__a21o_1
X_5389_ net453 net1140 _2419_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__mux2_1
X_7128_ clknet_leaf_47_csclk net1430 net514 VGND VGND VPWR VPWR gpio_configure\[36\]\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_101_531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7059_ clknet_leaf_22_csclk net1384 net515 VGND VGND VPWR VPWR gpio_configure\[27\]\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_131_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_160 net391 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_171 net462 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_182 clknet_2_0__leaf_mgmt_gpio_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_193 _1073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4760_ _1599_ _1646_ _1745_ _1636_ _1970_ VGND VGND VPWR VPWR _1972_ sky130_fd_sc_hd__o221a_1
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_193_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3711_ net383 net609 VGND VGND VPWR VPWR _1299_ sky130_fd_sc_hd__nor2_2
XFILLER_147_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4691_ _1803_ _1873_ VGND VGND VPWR VPWR _1903_ sky130_fd_sc_hd__or2_1
XFILLER_119_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6430_ net492 net481 VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__and2_1
XFILLER_146_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3642_ _1224_ _1226_ _1228_ _1230_ VGND VGND VPWR VPWR _1231_ sky130_fd_sc_hd__or4_1
XFILLER_174_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6361_ net170 net166 wbbd_state\[8\] VGND VGND VPWR VPWR _3161_ sky130_fd_sc_hd__a21boi_1
X_3573_ _1156_ _1158_ _1160_ _1162_ VGND VGND VPWR VPWR _1163_ sky130_fd_sc_hd__or4_1
XFILLER_161_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5312_ net435 net1087 _2410_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__mux2_1
XFILLER_161_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6292_ net359 _3094_ _3103_ VGND VGND VPWR VPWR _3104_ sky130_fd_sc_hd__or3_1
XFILLER_114_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5243_ net542 net1906 net547 VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__mux2_1
Xhold19 _0866_ VGND VGND VPWR VPWR net552 sky130_fd_sc_hd__dlygate4sd3_1
X_5174_ _2090_ _2252_ _2357_ _2379_ VGND VGND VPWR VPWR _2380_ sky130_fd_sc_hd__or4b_1
XFILLER_68_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4125_ net445 net742 _1510_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__mux2_1
XFILLER_84_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4056_ net770 net465 net356 VGND VGND VPWR VPWR _1483_ sky130_fd_sc_hd__mux2_1
XFILLER_83_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_418 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4958_ _1665_ _1671_ _1678_ _1805_ _2167_ VGND VGND VPWR VPWR _2168_ sky130_fd_sc_hd__o221a_1
XFILLER_184_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3909_ net475 _1445_ _1451_ serial_xfer xfer_state\[0\] VGND VGND VPWR VPWR _0016_
+ sky130_fd_sc_hd__a32o_1
XFILLER_177_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4889_ _1651_ _1655_ _2081_ VGND VGND VPWR VPWR _2100_ sky130_fd_sc_hd__a21oi_1
XFILLER_137_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6628_ clknet_3_4_0_wb_clk_i _0241_ VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__dfxtp_1
XFILLER_165_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6559_ clknet_leaf_54_csclk net937 net506 VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__dfrtp_1
XFILLER_118_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire431 _1439_ VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__clkbuf_2
XFILLER_156_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5930_ gpio_configure\[20\]\[11\] _2499_ _2537_ gpio_configure\[17\]\[11\] _2753_
+ VGND VGND VPWR VPWR _2754_ sky130_fd_sc_hd__a221o_1
XFILLER_80_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5861_ gpio_configure\[14\]\[8\] _2494_ _2528_ gpio_configure\[7\]\[8\] VGND VGND
+ VPWR VPWR _2688_ sky130_fd_sc_hd__a22o_1
XFILLER_179_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4812_ _2009_ _2011_ _2016_ _2022_ VGND VGND VPWR VPWR _2023_ sky130_fd_sc_hd__or4bb_1
XFILLER_61_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5792_ _2618_ _2620_ _2622_ VGND VGND VPWR VPWR _2623_ sky130_fd_sc_hd__or3_1
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4743_ _1599_ _1655_ VGND VGND VPWR VPWR _1955_ sky130_fd_sc_hd__nor2_1
XFILLER_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4674_ _1601_ _1677_ VGND VGND VPWR VPWR _1886_ sky130_fd_sc_hd__nand2_8
X_6413_ net492 net482 VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__and2_1
X_3625_ gpio_configure\[16\]\[2\] _0912_ _1102_ gpio_configure\[15\]\[10\] _1202_
+ VGND VGND VPWR VPWR _1214_ sky130_fd_sc_hd__a221o_1
XFILLER_135_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6344_ net2117 net366 _3152_ _3153_ VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__o22a_1
X_3556_ gpio_configure\[1\]\[11\] _1103_ _1127_ gpio_configure\[33\]\[11\] VGND VGND
+ VPWR VPWR _1146_ sky130_fd_sc_hd__a22o_1
XFILLER_103_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6275_ gpio_configure\[29\]\[10\] _2816_ _2820_ gpio_configure\[21\]\[10\] _3086_
+ VGND VGND VPWR VPWR _3087_ sky130_fd_sc_hd__a221o_1
XFILLER_163_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3487_ gpio_configure\[26\]\[4\] net371 _0933_ clknet_2_2__leaf_mgmt_gpio_in[4] _1077_
+ VGND VGND VPWR VPWR _1078_ sky130_fd_sc_hd__a221o_2
XFILLER_115_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5226_ net1590 net458 _2400_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__mux2_1
Xinput109 wb_adr_i[19] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_1
XFILLER_130_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5157_ _2317_ _2360_ _2362_ _2363_ VGND VGND VPWR VPWR _2364_ sky130_fd_sc_hd__o31a_1
XFILLER_56_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4108_ net449 net1232 _1508_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__mux2_1
XFILLER_84_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5088_ wbbd_addr\[3\] _1529_ _2279_ _2296_ VGND VGND VPWR VPWR _2297_ sky130_fd_sc_hd__a22o_1
X_4039_ net1000 net443 _1477_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__mux2_1
XFILLER_71_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_60 _2498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_71 _2538_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_82 _3130_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_93 mask_rev_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold308 _0679_ VGND VGND VPWR VPWR net841 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold319 gpio_configure\[13\]\[6\] VGND VGND VPWR VPWR net852 sky130_fd_sc_hd__dlygate4sd3_1
X_3410_ _0986_ _1003_ VGND VGND VPWR VPWR _1004_ sky130_fd_sc_hd__or2_4
XFILLER_109_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4390_ net112 net111 net114 net113 VGND VGND VPWR VPWR _1602_ sky130_fd_sc_hd__or4_4
XFILLER_98_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3341_ net386 net609 VGND VGND VPWR VPWR _0937_ sky130_fd_sc_hd__nor2_2
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ gpio_configure\[34\]\[1\] net393 _2852_ gpio_configure\[19\]\[1\] _2880_ VGND
+ VGND VPWR VPWR _2881_ sky130_fd_sc_hd__a221o_1
XFILLER_140_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ net560 net588 VGND VGND VPWR VPWR _0868_ sky130_fd_sc_hd__and2b_4
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1008 _0181_ VGND VGND VPWR VPWR net1541 sky130_fd_sc_hd__dlygate4sd3_1
X_5011_ _2084_ _2110_ _2220_ _2202_ VGND VGND VPWR VPWR _2221_ sky130_fd_sc_hd__o31a_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1019 gpio_configure\[7\]\[5\] VGND VGND VPWR VPWR net1552 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6962_ clknet_leaf_17_csclk net1739 net512 VGND VGND VPWR VPWR gpio_configure\[15\]\[0\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_53_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5913_ _2731_ _2733_ _2735_ _2737_ VGND VGND VPWR VPWR _2738_ sky130_fd_sc_hd__or4_1
X_6893_ clknet_leaf_40_csclk net733 net516 VGND VGND VPWR VPWR gpio_configure\[6\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_21_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5844_ gpio_configure\[4\]\[7\] _2502_ _2671_ VGND VGND VPWR VPWR _2672_ sky130_fd_sc_hd__a21o_1
XFILLER_34_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5775_ gpio_configure\[5\]\[4\] net422 net420 gpio_configure\[25\]\[4\] VGND VGND
+ VPWR VPWR _2606_ sky130_fd_sc_hd__a22o_1
XFILLER_21_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4726_ _1937_ VGND VGND VPWR VPWR _1938_ sky130_fd_sc_hd__inv_2
XFILLER_175_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4657_ _1589_ net478 _1662_ VGND VGND VPWR VPWR _1869_ sky130_fd_sc_hd__and3_1
XFILLER_175_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput80 spi_sck VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_1
Xhold820 _0575_ VGND VGND VPWR VPWR net1353 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3608_ gpio_configure\[34\]\[2\] net358 _0932_ gpio_configure\[35\]\[2\] VGND VGND
+ VPWR VPWR _1197_ sky130_fd_sc_hd__a22o_1
XFILLER_174_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput91 spimemio_flash_io3_do VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_1
Xhold831 _0145_ VGND VGND VPWR VPWR net1364 sky130_fd_sc_hd__dlygate4sd3_1
X_4588_ net127 net126 net125 net128 VGND VGND VPWR VPWR _1800_ sky130_fd_sc_hd__or4bb_4
Xhold842 gpio_configure\[2\]\[6\] VGND VGND VPWR VPWR net1375 sky130_fd_sc_hd__dlygate4sd3_1
Xhold853 _0691_ VGND VGND VPWR VPWR net1386 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6327_ gpio_configure\[11\]\[12\] _2814_ _2842_ gpio_configure\[15\]\[12\] VGND VGND
+ VPWR VPWR _3137_ sky130_fd_sc_hd__a22o_1
Xhold864 gpio_configure\[18\]\[1\] VGND VGND VPWR VPWR net1397 sky130_fd_sc_hd__dlygate4sd3_1
Xhold875 _0306_ VGND VGND VPWR VPWR net1408 sky130_fd_sc_hd__dlygate4sd3_1
X_3539_ gpio_configure\[1\]\[4\] _0934_ _1129_ gpio_configure\[11\]\[12\] VGND VGND
+ VPWR VPWR _1130_ sky130_fd_sc_hd__a22o_2
XFILLER_107_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold886 gpio_configure\[25\]\[6\] VGND VGND VPWR VPWR net1419 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold897 _0731_ VGND VGND VPWR VPWR net1430 sky130_fd_sc_hd__dlygate4sd3_1
X_6258_ gpio_configure\[37\]\[9\] _2806_ net416 gpio_configure\[32\]\[9\] _3059_ VGND
+ VGND VPWR VPWR _3071_ sky130_fd_sc_hd__a221o_1
XFILLER_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5209_ net818 net451 _2394_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__mux2_1
XFILLER_103_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6189_ gpio_configure\[30\]\[6\] _2799_ _2841_ gpio_configure\[34\]\[6\] _3004_ VGND
+ VGND VPWR VPWR _3005_ sky130_fd_sc_hd__a221o_1
XFILLER_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1520 hkspi.odata\[2\] VGND VGND VPWR VPWR net2053 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1531 wbbd_addr\[4\] VGND VGND VPWR VPWR net2064 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1542 net346 VGND VGND VPWR VPWR net2075 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1553 wbbd_state\[0\] VGND VGND VPWR VPWR net2086 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1564 hkspi.state\[4\] VGND VGND VPWR VPWR net2097 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1575 serial_data_staging_2\[9\] VGND VGND VPWR VPWR net2108 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1586 hkspi.readmode VGND VGND VPWR VPWR net2119 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1597 xfer_state\[2\] VGND VGND VPWR VPWR net2130 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_189_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3890_ _1385_ _1386_ VGND VGND VPWR VPWR _1441_ sky130_fd_sc_hd__nor2_1
XFILLER_188_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5560_ net438 net1399 _2438_ VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__mux2_1
XFILLER_157_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4511_ _1643_ _1655_ _1720_ _1722_ VGND VGND VPWR VPWR _1723_ sky130_fd_sc_hd__o211a_1
XFILLER_144_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5491_ net437 net1423 _2430_ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__mux2_1
XFILLER_129_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold105 _0850_ VGND VGND VPWR VPWR net638 sky130_fd_sc_hd__dlygate4sd3_1
X_4442_ _1623_ _1647_ VGND VGND VPWR VPWR _1654_ sky130_fd_sc_hd__nor2_2
Xhold116 _0728_ VGND VGND VPWR VPWR net649 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 net442 VGND VGND VPWR VPWR net660 sky130_fd_sc_hd__clkbuf_16
Xhold138 _1513_ VGND VGND VPWR VPWR net671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 _0317_ VGND VGND VPWR VPWR net682 sky130_fd_sc_hd__dlygate4sd3_1
X_7161_ clknet_3_3_0_wb_clk_i _0763_ net499 VGND VGND VPWR VPWR serial_load_pre sky130_fd_sc_hd__dfrtp_1
XFILLER_144_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4373_ net124 _1583_ VGND VGND VPWR VPWR _1585_ sky130_fd_sc_hd__or2_2
XFILLER_98_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6112_ gpio_configure\[30\]\[3\] _2799_ _2823_ gpio_configure\[2\]\[3\] _2930_ VGND
+ VGND VPWR VPWR _2931_ sky130_fd_sc_hd__a221o_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3324_ _0873_ net381 VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__nor2_8
X_7092_ clknet_leaf_77_csclk net1671 net485 VGND VGND VPWR VPWR gpio_configure\[31\]\[10\]
+ sky130_fd_sc_hd__dfstp_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6043_ gpio_configure\[14\]\[0\] net411 _2859_ _2864_ VGND VGND VPWR VPWR _2865_
+ sky130_fd_sc_hd__a211o_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ net638 net581 net551 VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__or3b_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3186_ hkspi.pre_pass_thru_mgmt VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__inv_2
XFILLER_27_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6945_ clknet_leaf_41_csclk net1042 net517 VGND VGND VPWR VPWR gpio_configure\[12\]\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_53_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_2_0_wb_clk_i clknet_1_1_1_wb_clk_i VGND VGND VPWR VPWR clknet_2_2_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6876_ clknet_leaf_24_csclk net1659 net518 VGND VGND VPWR VPWR gpio_configure\[4\]\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_5827_ gpio_configure\[19\]\[6\] _2491_ _2531_ gpio_configure\[24\]\[6\] _2655_ VGND
+ VGND VPWR VPWR _2656_ sky130_fd_sc_hd__a221o_1
XFILLER_22_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5758_ gpio_configure\[6\]\[3\] _2490_ _2588_ _2589_ VGND VGND VPWR VPWR _2590_ sky130_fd_sc_hd__a211o_1
XFILLER_182_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4709_ _1579_ _1798_ _1889_ _1920_ VGND VGND VPWR VPWR _1921_ sky130_fd_sc_hd__o211a_1
X_5689_ _2459_ _2466_ VGND VGND VPWR VPWR _2524_ sky130_fd_sc_hd__and2_4
XFILLER_108_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold650 _0609_ VGND VGND VPWR VPWR net1183 sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 gpio_configure\[2\]\[4\] VGND VGND VPWR VPWR net1194 sky130_fd_sc_hd__dlygate4sd3_1
Xhold672 _0157_ VGND VGND VPWR VPWR net1205 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap391 _2860_ VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__buf_12
Xhold683 gpio_configure\[32\]\[10\] VGND VGND VPWR VPWR net1216 sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 _0250_ VGND VGND VPWR VPWR net1227 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1350 net1883 VGND VGND VPWR VPWR wb_dat_o[28] sky130_fd_sc_hd__buf_12
XFILLER_85_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1361 net1955 VGND VGND VPWR VPWR net1894 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1372 mgmt_gpio_data_buf\[22\] VGND VGND VPWR VPWR net1905 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1383 gpio_configure\[35\]\[6\] VGND VGND VPWR VPWR net1916 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1394 net264 VGND VGND VPWR VPWR net1927 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4991_ _2174_ _2200_ VGND VGND VPWR VPWR _2201_ sky130_fd_sc_hd__nor2_1
XFILLER_91_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6730_ clknet_leaf_18_csclk net1163 net512 VGND VGND VPWR VPWR gpio_configure\[36\]\[12\]
+ sky130_fd_sc_hd__dfstp_1
X_3942_ net474 clknet_1_1__leaf_wbbd_sck net483 _1457_ VGND VGND VPWR VPWR csclk sky130_fd_sc_hd__a22o_2
XFILLER_189_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6661_ clknet_leaf_78_csclk net1626 net485 VGND VGND VPWR VPWR gpio_configure\[8\]\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_32_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3873_ net512 net483 VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__and2_1
XFILLER_176_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5612_ pad_count_1\[1\] pad_count_1\[0\] VGND VGND VPWR VPWR _2459_ sky130_fd_sc_hd__nor2_4
X_6592_ clknet_leaf_56_csclk net743 net504 VGND VGND VPWR VPWR mgmt_gpio_data_buf\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_191_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5543_ net1262 net434 _2436_ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__mux2_1
XFILLER_129_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5474_ net1266 net434 _2428_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__mux2_1
XFILLER_117_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7213_ net87 VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__clkbuf_2
XFILLER_105_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4425_ _1612_ _1635_ VGND VGND VPWR VPWR _1637_ sky130_fd_sc_hd__nand2_1
XFILLER_144_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7144_ clknet_3_3_0_wb_clk_i _0747_ net502 VGND VGND VPWR VPWR xfer_count\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_113_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4356_ _1558_ _1565_ _1567_ _1559_ VGND VGND VPWR VPWR _1568_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout426 net427 VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__buf_8
XFILLER_86_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout437 net439 VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__buf_6
XFILLER_113_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3307_ net600 _0884_ VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__nand2_8
Xfanout448 net617 VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__buf_6
X_7075_ clknet_leaf_23_csclk net1337 net515 VGND VGND VPWR VPWR gpio_configure\[29\]\[1\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout459 net577 VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__buf_4
X_4287_ net443 net988 _1539_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__mux2_1
XFILLER_58_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6026_ _2844_ _2845_ _2846_ _2847_ VGND VGND VPWR VPWR _2848_ sky130_fd_sc_hd__or4_1
XFILLER_100_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3238_ net530 VGND VGND VPWR VPWR _0834_ sky130_fd_sc_hd__clkinv_8
XFILLER_67_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6928_ clknet_leaf_53_csclk net1347 net507 VGND VGND VPWR VPWR gpio_configure\[10\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_23_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6859_ clknet_leaf_49_csclk net887 net505 VGND VGND VPWR VPWR gpio_configure\[2\]\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_168_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold480 gpio_configure\[19\]\[12\] VGND VGND VPWR VPWR net1013 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold491 _0123_ VGND VGND VPWR VPWR net1024 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1180 gpio_configure\[32\]\[0\] VGND VGND VPWR VPWR net1713 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1191 gpio_configure\[19\]\[0\] VGND VGND VPWR VPWR net1724 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4210_ _1057_ net426 VGND VGND VPWR VPWR _1523_ sky130_fd_sc_hd__and2_2
X_5190_ net455 net1682 _2390_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__mux2_1
XFILLER_141_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4141_ _1110_ net429 VGND VGND VPWR VPWR _1513_ sky130_fd_sc_hd__nand2_2
X_4072_ net1709 _1491_ _1490_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__mux2_1
XFILLER_83_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4974_ _1599_ net432 _1772_ _1592_ VGND VGND VPWR VPWR _2184_ sky130_fd_sc_hd__a211oi_1
X_3925_ mgmt_gpio_data\[35\] net81 net79 VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__mux2_8
XFILLER_51_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6713_ clknet_leaf_8_csclk net767 net509 VGND VGND VPWR VPWR gpio_configure\[16\]\[10\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_149_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6644_ clknet_3_4_0_wb_clk_i _0257_ VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__dfxtp_1
X_3856_ hkspi.fixed\[1\] _1416_ VGND VGND VPWR VPWR _1422_ sky130_fd_sc_hd__nor2_1
XFILLER_137_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6575_ clknet_leaf_0_csclk net1731 net486 VGND VGND VPWR VPWR mgmt_gpio_data\[33\]
+ sky130_fd_sc_hd__dfrtp_1
X_3787_ gpio_configure\[21\]\[0\] _0911_ _1314_ net172 _1320_ VGND VGND VPWR VPWR
+ _1373_ sky130_fd_sc_hd__a221o_1
XFILLER_164_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5526_ net441 net952 _2434_ VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__mux2_1
X_5457_ net372 net427 VGND VGND VPWR VPWR _2427_ sky130_fd_sc_hd__nand2_8
XFILLER_160_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4408_ net125 _1610_ net126 VGND VGND VPWR VPWR _1620_ sky130_fd_sc_hd__a21oi_1
XFILLER_182_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5388_ net459 net1348 _2419_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__mux2_1
XFILLER_160_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7127_ clknet_leaf_27_csclk net1605 net521 VGND VGND VPWR VPWR gpio_configure\[36\]\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_4339_ net130 net129 net101 net100 VGND VGND VPWR VPWR _1551_ sky130_fd_sc_hd__and4_1
XFILLER_101_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7058_ clknet_leaf_26_csclk net1987 net521 VGND VGND VPWR VPWR gpio_configure\[27\]\[0\]
+ sky130_fd_sc_hd__dfstp_4
X_6009_ _2478_ _2793_ _2800_ VGND VGND VPWR VPWR _2831_ sky130_fd_sc_hd__and3_4
XFILLER_39_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_150 net297 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_161 net392 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_172 net463 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_183 clknet_2_0__leaf_mgmt_gpio_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_194 _1085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3710_ _1291_ _1293_ _1295_ _1297_ VGND VGND VPWR VPWR _1298_ sky130_fd_sc_hd__or4_1
XFILLER_147_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4690_ _1803_ _1886_ VGND VGND VPWR VPWR _1902_ sky130_fd_sc_hd__or2_1
XFILLER_186_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3641_ net26 _0900_ _1046_ gpio_configure\[28\]\[10\] _1229_ VGND VGND VPWR VPWR
+ _1230_ sky130_fd_sc_hd__a221o_1
XFILLER_146_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6360_ net170 net165 wbbd_state\[5\] VGND VGND VPWR VPWR _3160_ sky130_fd_sc_hd__a21bo_1
X_3572_ gpio_configure\[2\]\[3\] _0908_ _1095_ gpio_configure\[3\]\[11\] _1161_ VGND
+ VGND VPWR VPWR _1162_ sky130_fd_sc_hd__a221o_1
X_5311_ net438 net1379 _2410_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__mux2_1
XFILLER_127_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6291_ _3096_ _3098_ _3100_ _3102_ VGND VGND VPWR VPWR _3103_ sky130_fd_sc_hd__or4_2
XFILLER_142_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5242_ net471 net1451 net547 VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__mux2_1
XFILLER_102_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_30_csclk clknet_3_7_0_csclk VGND VGND VPWR VPWR clknet_leaf_30_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_68_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5173_ _1599_ _1655_ _2203_ _1651_ _1721_ VGND VGND VPWR VPWR _2379_ sky130_fd_sc_hd__o221a_1
X_4124_ net451 net828 _1510_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__mux2_1
XFILLER_68_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput1 debug_mode VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_2
X_4055_ net1722 _1482_ _1481_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_45_csclk clknet_3_6_0_csclk VGND VGND VPWR VPWR clknet_leaf_45_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4957_ _1574_ _2146_ VGND VGND VPWR VPWR _2167_ sky130_fd_sc_hd__nand2_1
XFILLER_52_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3908_ net475 _1445_ VGND VGND VPWR VPWR _1453_ sky130_fd_sc_hd__nand2_1
X_4888_ _1645_ _2082_ _1966_ _1698_ VGND VGND VPWR VPWR _2099_ sky130_fd_sc_hd__a211o_1
XFILLER_138_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3839_ hkspi.count\[0\] _1410_ VGND VGND VPWR VPWR _1411_ sky130_fd_sc_hd__nor2_1
X_6627_ clknet_3_5_0_wb_clk_i _0240_ VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__dfxtp_1
XFILLER_192_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6558_ clknet_leaf_56_csclk net951 net504 VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__dfrtp_1
XFILLER_192_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5509_ net437 net1367 _2432_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__mux2_1
XFILLER_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6489_ clknet_leaf_71_csclk net1004 net498 VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__dfstp_4
XFILLER_106_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire476 net544 VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__buf_4
XFILLER_171_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5860_ net2123 _2687_ net366 VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__mux2_1
XFILLER_61_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4811_ _1782_ _1801_ _1971_ _1997_ _2021_ VGND VGND VPWR VPWR _2022_ sky130_fd_sc_hd__o2111a_1
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5791_ gpio_configure\[11\]\[4\] _2505_ _2521_ gpio_configure\[21\]\[4\] _2621_ VGND
+ VGND VPWR VPWR _2622_ sky130_fd_sc_hd__a221o_1
XFILLER_61_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4742_ _1612_ _1617_ _1936_ VGND VGND VPWR VPWR _1954_ sky130_fd_sc_hd__and3_1
X_4673_ _1801_ _1872_ VGND VGND VPWR VPWR _1885_ sky130_fd_sc_hd__nor2_1
X_6412_ net492 net481 VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__and2_1
X_3624_ gpio_configure\[8\]\[2\] _0939_ _1095_ gpio_configure\[3\]\[10\] _1200_ VGND
+ VGND VPWR VPWR _1213_ sky130_fd_sc_hd__a221o_1
XFILLER_174_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6343_ serial_data_staging_2\[11\] _2444_ _2485_ VGND VGND VPWR VPWR _3153_ sky130_fd_sc_hd__o21ba_1
XFILLER_127_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3555_ gpio_configure\[0\]\[3\] _0898_ _1116_ gpio_configure\[26\]\[11\] VGND VGND
+ VPWR VPWR _1145_ sky130_fd_sc_hd__a22o_1
XFILLER_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6274_ gpio_configure\[30\]\[10\] _2799_ net408 gpio_configure\[35\]\[10\] VGND VGND
+ VPWR VPWR _3086_ sky130_fd_sc_hd__a22o_1
X_3486_ gpio_configure\[17\]\[4\] net367 _1076_ gpio_configure\[27\]\[12\] VGND VGND
+ VPWR VPWR _1077_ sky130_fd_sc_hd__a22o_1
X_5225_ _1196_ net427 VGND VGND VPWR VPWR _2400_ sky130_fd_sc_hd__and2_4
XFILLER_69_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5156_ _2280_ _2284_ _2314_ VGND VGND VPWR VPWR _2363_ sky130_fd_sc_hd__nor3_1
XFILLER_29_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4107_ net577 net814 _1508_ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__mux2_1
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5087_ _2282_ _2295_ VGND VGND VPWR VPWR _2296_ sky130_fd_sc_hd__or2_1
XFILLER_84_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4038_ net1029 net449 _1477_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__mux2_1
XFILLER_84_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5989_ _1449_ _2469_ _2796_ VGND VGND VPWR VPWR _2811_ sky130_fd_sc_hd__and3_4
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_50 _1510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_61 _2499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 _2540_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_83 gpio_configure\[11\]\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_94 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput190 net190 VGND VGND VPWR VPWR mgmt_gpio_oeb[23] sky130_fd_sc_hd__buf_12
XFILLER_94_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold309 gpio_configure\[25\]\[2\] VGND VGND VPWR VPWR net842 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3340_ net390 _0895_ VGND VGND VPWR VPWR _0936_ sky130_fd_sc_hd__nor2_8
Xclkbuf_3_4_0_wb_clk_i clknet_2_2_0_wb_clk_i VGND VGND VPWR VPWR clknet_3_4_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3271_ net627 net552 VGND VGND VPWR VPWR _0867_ sky130_fd_sc_hd__or2_4
XFILLER_97_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _2211_ _2214_ _2215_ _2219_ VGND VGND VPWR VPWR _2220_ sky130_fd_sc_hd__or4_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1009 gpio_configure\[9\]\[5\] VGND VGND VPWR VPWR net1542 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6961_ clknet_leaf_56_csclk net717 net506 VGND VGND VPWR VPWR gpio_configure\[14\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_5912_ gpio_configure\[25\]\[10\] _2511_ _2538_ gpio_configure\[1\]\[10\] _2736_
+ VGND VGND VPWR VPWR _2737_ sky130_fd_sc_hd__a221o_1
X_6892_ clknet_leaf_40_csclk net1388 net516 VGND VGND VPWR VPWR gpio_configure\[6\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_5843_ gpio_configure\[22\]\[7\] _2498_ _2517_ gpio_configure\[30\]\[7\] VGND VGND
+ VPWR VPWR _2671_ sky130_fd_sc_hd__a22o_1
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5774_ net2034 _2605_ net366 VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__mux2_1
XFILLER_166_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4725_ _1615_ _1616_ _1656_ _1548_ VGND VGND VPWR VPWR _1937_ sky130_fd_sc_hd__a211oi_4
XFILLER_135_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4656_ _1592_ _1663_ VGND VGND VPWR VPWR _1868_ sky130_fd_sc_hd__nor2_1
XFILLER_190_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3607_ net383 _0903_ VGND VGND VPWR VPWR _1196_ sky130_fd_sc_hd__nor2_2
Xinput70 mgmt_gpio_in[7] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__buf_2
Xinput81 spi_sdo VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold810 _0523_ VGND VGND VPWR VPWR net1343 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_174_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold821 gpio_configure\[21\]\[6\] VGND VGND VPWR VPWR net1354 sky130_fd_sc_hd__dlygate4sd3_1
X_4587_ _1779_ _1798_ VGND VGND VPWR VPWR _1799_ sky130_fd_sc_hd__nor2_1
XFILLER_116_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold832 gpio_configure\[11\]\[6\] VGND VGND VPWR VPWR net1365 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput92 spimemio_flash_io3_oeb VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_2
Xhold843 _0467_ VGND VGND VPWR VPWR net1376 sky130_fd_sc_hd__dlygate4sd3_1
X_6326_ gpio_configure\[2\]\[12\] net398 _2855_ gpio_configure\[27\]\[12\] _3135_
+ VGND VGND VPWR VPWR _3136_ sky130_fd_sc_hd__a221o_1
X_3538_ net582 _0973_ VGND VGND VPWR VPWR _1129_ sky130_fd_sc_hd__nor2_4
Xhold854 gpio_configure\[6\]\[2\] VGND VGND VPWR VPWR net1387 sky130_fd_sc_hd__dlygate4sd3_1
Xhold865 _0590_ VGND VGND VPWR VPWR net1398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 net2114 VGND VGND VPWR VPWR net1409 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold887 _0651_ VGND VGND VPWR VPWR net1420 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_107_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold898 gpio_configure\[31\]\[1\] VGND VGND VPWR VPWR net1431 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6257_ _3064_ _3065_ _3067_ _3069_ VGND VGND VPWR VPWR _3070_ sky130_fd_sc_hd__or4_1
XFILLER_88_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3469_ gpio_configure\[0\]\[4\] _0898_ _0917_ gpio_configure\[29\]\[4\] VGND VGND
+ VPWR VPWR _1060_ sky130_fd_sc_hd__a22o_1
XFILLER_103_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5208_ net864 net457 _2394_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__mux2_1
XFILLER_190_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6188_ gpio_configure\[14\]\[6\] net411 net406 gpio_configure\[27\]\[6\] VGND VGND
+ VPWR VPWR _3004_ sky130_fd_sc_hd__a22o_1
XFILLER_130_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1510 _0782_ VGND VGND VPWR VPWR net2043 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1521 hkspi.odata\[5\] VGND VGND VPWR VPWR net2054 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5139_ _2319_ _2329_ _2337_ _2346_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__or4_1
Xhold1532 wbbd_data\[3\] VGND VGND VPWR VPWR net2065 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1543 hkspi.pre_pass_thru_mgmt VGND VGND VPWR VPWR net2076 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1554 _0009_ VGND VGND VPWR VPWR net2087 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1565 _0081_ VGND VGND VPWR VPWR net2098 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1576 mgmt_gpio_data_buf\[3\] VGND VGND VPWR VPWR net2109 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1587 mgmt_gpio_data_buf\[7\] VGND VGND VPWR VPWR net2120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1598 mgmt_gpio_data\[10\] VGND VGND VPWR VPWR net2131 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4510_ _1660_ _1682_ _1721_ VGND VGND VPWR VPWR _1722_ sky130_fd_sc_hd__and3_1
XFILLER_117_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5490_ net440 net1556 _2430_ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__mux2_1
XFILLER_156_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold106 _0877_ VGND VGND VPWR VPWR net639 sky130_fd_sc_hd__dlygate4sd3_1
X_4441_ _1634_ _1647_ VGND VGND VPWR VPWR _1653_ sky130_fd_sc_hd__or2_2
XFILLER_172_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold117 gpio_configure\[4\]\[6\] VGND VGND VPWR VPWR net650 sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 _0198_ VGND VGND VPWR VPWR net661 sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 _0222_ VGND VGND VPWR VPWR net672 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7160_ clknet_3_2_0_wb_clk_i _0762_ net499 VGND VGND VPWR VPWR serial_clock_pre sky130_fd_sc_hd__dfrtp_1
X_4372_ net124 _1583_ VGND VGND VPWR VPWR _1584_ sky130_fd_sc_hd__nor2_8
XFILLER_171_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6111_ gpio_configure\[20\]\[3\] net396 net410 gpio_configure\[8\]\[3\] VGND VGND
+ VPWR VPWR _2930_ sky130_fd_sc_hd__a22o_1
XFILLER_125_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3323_ _0889_ net385 VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__nor2_8
XFILLER_98_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7091_ clknet_leaf_5_csclk net1446 net494 VGND VGND VPWR VPWR gpio_configure\[31\]\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6042_ gpio_configure\[17\]\[0\] net391 _2861_ gpio_configure\[28\]\[0\] _2863_ VGND
+ VGND VPWR VPWR _2864_ sky130_fd_sc_hd__a221o_1
X_3254_ net637 net1965 net474 VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__mux2_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3185_ hkspi.addr\[0\] VGND VGND VPWR VPWR _0815_ sky130_fd_sc_hd__inv_2
XFILLER_54_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6944_ clknet_leaf_53_csclk net797 net517 VGND VGND VPWR VPWR gpio_configure\[12\]\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_179_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6875_ clknet_leaf_26_csclk net566 net519 VGND VGND VPWR VPWR gpio_configure\[4\]\[1\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_22_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5826_ gpio_configure\[11\]\[6\] _2505_ _2507_ gpio_configure\[10\]\[6\] VGND VGND
+ VPWR VPWR _2655_ sky130_fd_sc_hd__a22o_1
XFILLER_139_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5757_ gpio_configure\[9\]\[3\] _2512_ _2529_ gpio_configure\[29\]\[3\] _2586_ VGND
+ VGND VPWR VPWR _2589_ sky130_fd_sc_hd__a221o_1
XFILLER_148_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4708_ _1902_ _1903_ _1918_ _1919_ VGND VGND VPWR VPWR _1920_ sky130_fd_sc_hd__and4_1
XFILLER_175_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5688_ net472 _2466_ _2489_ VGND VGND VPWR VPWR _2523_ sky130_fd_sc_hd__and3_4
XFILLER_108_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4639_ _1791_ _1833_ VGND VGND VPWR VPWR _1851_ sky130_fd_sc_hd__nor2_1
XFILLER_150_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold640 _0649_ VGND VGND VPWR VPWR net1173 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold651 gpio_configure\[28\]\[1\] VGND VGND VPWR VPWR net1184 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap370 net640 VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__buf_8
Xhold662 _0465_ VGND VGND VPWR VPWR net1195 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap381 net382 VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__buf_12
Xhold673 gpio_configure\[23\]\[5\] VGND VGND VPWR VPWR net1206 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap392 _2843_ VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__buf_12
Xhold684 _0371_ VGND VGND VPWR VPWR net1217 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6309_ gpio_configure\[34\]\[11\] net393 _2852_ gpio_configure\[19\]\[11\] _3119_
+ VGND VGND VPWR VPWR _3120_ sky130_fd_sc_hd__a221o_1
XFILLER_103_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold695 gpio_configure\[31\]\[12\] VGND VGND VPWR VPWR net1228 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1340 net1873 VGND VGND VPWR VPWR wb_dat_o[31] sky130_fd_sc_hd__buf_12
Xhold1351 net1951 VGND VGND VPWR VPWR net1884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1362 net1895 VGND VGND VPWR VPWR wb_dat_o[29] sky130_fd_sc_hd__buf_12
Xhold1373 mgmt_gpio_data_buf\[9\] VGND VGND VPWR VPWR net1906 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1384 gpio_configure\[11\]\[11\] VGND VGND VPWR VPWR net1917 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1395 net296 VGND VGND VPWR VPWR net1928 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xnet499_2 clknet_2_3__leaf_mgmt_gpio_in[4] VGND VGND VPWR VPWR net533 sky130_fd_sc_hd__inv_2
X_4990_ _2189_ _2199_ VGND VGND VPWR VPWR _2200_ sky130_fd_sc_hd__and2b_1
XFILLER_90_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3941_ net474 net533 VGND VGND VPWR VPWR _1457_ sky130_fd_sc_hd__nor2_2
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6660_ clknet_leaf_78_csclk net1624 net485 VGND VGND VPWR VPWR gpio_configure\[8\]\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_3872_ hkspi_disable gpio_configure\[3\]\[3\] net67 VGND VGND VPWR VPWR _1427_ sky130_fd_sc_hd__nor3_2
XFILLER_189_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5611_ xfer_state\[2\] _2457_ net2132 VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__mux2_1
XFILLER_149_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6591_ clknet_leaf_57_csclk net829 net504 VGND VGND VPWR VPWR mgmt_gpio_data_buf\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_5542_ net1435 net437 _2436_ VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__mux2_1
XFILLER_192_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5473_ net1443 net437 _2428_ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__mux2_1
XFILLER_132_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4424_ _1617_ _1628_ _1633_ VGND VGND VPWR VPWR _1636_ sky130_fd_sc_hd__nand3_4
XFILLER_132_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7143_ clknet_3_3_0_wb_clk_i _0746_ net499 VGND VGND VPWR VPWR serial_busy sky130_fd_sc_hd__dfrtp_1
XFILLER_99_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4355_ _1554_ _1557_ net128 VGND VGND VPWR VPWR _1567_ sky130_fd_sc_hd__a21oi_1
XFILLER_113_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout427 net645 VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__buf_12
X_3306_ net378 net601 VGND VGND VPWR VPWR _0902_ sky130_fd_sc_hd__nor2_8
X_7074_ clknet_leaf_63_csclk net1599 net501 VGND VGND VPWR VPWR gpio_configure\[29\]\[0\]
+ sky130_fd_sc_hd__dfstp_1
Xfanout438 net439 VGND VGND VPWR VPWR net438 sky130_fd_sc_hd__clkbuf_4
X_4286_ net449 net1073 _1539_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__mux2_1
Xfanout449 net451 VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__buf_8
XFILLER_113_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6025_ _2823_ net395 _2841_ net407 VGND VGND VPWR VPWR _2847_ sky130_fd_sc_hd__or4_1
X_3237_ net99 VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__inv_4
XFILLER_86_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6927_ clknet_leaf_39_csclk net1121 net517 VGND VGND VPWR VPWR gpio_configure\[10\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_81_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6858_ clknet_leaf_50_csclk net1617 net506 VGND VGND VPWR VPWR gpio_configure\[2\]\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_120_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5809_ gpio_configure\[5\]\[5\] net422 net420 gpio_configure\[25\]\[5\] VGND VGND
+ VPWR VPWR _2639_ sky130_fd_sc_hd__a22o_1
X_6789_ clknet_2_0__leaf_mgmt_gpio_in[4] _0392_ _0063_ VGND VGND VPWR VPWR hkspi.ldata\[6\]
+ sky130_fd_sc_hd__dfrtn_1
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold470 _1469_ VGND VGND VPWR VPWR net1003 sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 _0348_ VGND VGND VPWR VPWR net1014 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold492 gpio_configure\[25\]\[3\] VGND VGND VPWR VPWR net1025 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1170 _0376_ VGND VGND VPWR VPWR net1703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1181 _0698_ VGND VGND VPWR VPWR net1714 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1192 _0597_ VGND VGND VPWR VPWR net1725 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_728 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4140_ net1017 net443 _1512_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__mux2_1
XFILLER_96_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4071_ net1510 net466 _0933_ VGND VGND VPWR VPWR _1491_ sky130_fd_sc_hd__mux2_1
XFILLER_49_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4973_ _2180_ _2182_ VGND VGND VPWR VPWR _2183_ sky130_fd_sc_hd__or2_1
X_6712_ clknet_leaf_9_csclk net827 net509 VGND VGND VPWR VPWR gpio_configure\[16\]\[9\]
+ sky130_fd_sc_hd__dfrtp_4
X_3924_ mgmt_gpio_data\[33\] net78 net79 VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__mux2_8
XFILLER_20_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6643_ clknet_3_4_0_wb_clk_i _0256_ VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__dfxtp_1
X_3855_ hkspi.fixed\[2\] _1416_ _1421_ net2092 VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__o22a_1
XFILLER_164_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3786_ gpio_configure\[18\]\[0\] _0894_ _1062_ gpio_configure\[21\]\[8\] _1371_ VGND
+ VGND VPWR VPWR _1372_ sky130_fd_sc_hd__a221o_1
X_6574_ clknet_leaf_0_csclk net1743 net486 VGND VGND VPWR VPWR mgmt_gpio_data\[32\]
+ sky130_fd_sc_hd__dfrtp_1
X_5525_ net446 net1158 _2434_ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__mux2_1
XFILLER_117_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5456_ net573 net652 _2426_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__mux2_1
XFILLER_132_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4407_ net125 _1610_ VGND VGND VPWR VPWR _1619_ sky130_fd_sc_hd__xnor2_2
XFILLER_160_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5387_ net465 net848 _2419_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__mux2_1
XFILLER_99_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7126_ clknet_leaf_32_csclk net927 net524 VGND VGND VPWR VPWR gpio_configure\[35\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_4338_ net103 net102 net105 net104 VGND VGND VPWR VPWR _1550_ sky130_fd_sc_hd__and4_1
XFILLER_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4269_ net1318 net443 _1536_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__mux2_1
X_7057_ clknet_leaf_58_csclk net1273 net503 VGND VGND VPWR VPWR gpio_configure\[26\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_101_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6008_ _2469_ _2796_ _2800_ VGND VGND VPWR VPWR _2830_ sky130_fd_sc_hd__and3_4
XFILLER_67_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_140 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_151 net297 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_162 net392 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_173 net467 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_184 clknet_2_0__leaf_mgmt_gpio_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_195 _1136_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3640_ gpio_configure\[21\]\[2\] _0911_ _1047_ gpio_configure\[18\]\[10\] VGND VGND
+ VPWR VPWR _1229_ sky130_fd_sc_hd__a22o_1
XFILLER_146_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3571_ gpio_configure\[3\]\[3\] _0915_ _1119_ gpio_configure\[5\]\[11\] VGND VGND
+ VPWR VPWR _1161_ sky130_fd_sc_hd__a22o_1
X_5310_ net441 net1106 _2410_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__mux2_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6290_ gpio_configure\[3\]\[10\] _2830_ _2842_ gpio_configure\[15\]\[10\] _3101_
+ VGND VGND VPWR VPWR _3102_ sky130_fd_sc_hd__a221o_1
XFILLER_154_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5241_ net379 _0881_ net483 net546 VGND VGND VPWR VPWR _2403_ sky130_fd_sc_hd__or4_4
XFILLER_130_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5172_ _2324_ _2347_ _2349_ _2377_ VGND VGND VPWR VPWR _2378_ sky130_fd_sc_hd__nor4_1
XFILLER_68_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4123_ net457 net862 _1510_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__mux2_1
XFILLER_69_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput2 debug_oeb VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
X_4054_ net1326 net471 net356 VGND VGND VPWR VPWR _1482_ sky130_fd_sc_hd__mux2_1
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_opt_1_0_csclk clknet_3_1_0_csclk VGND VGND VPWR VPWR clknet_opt_1_0_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_37_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4956_ _1668_ _1671_ _2142_ _2154_ _1890_ VGND VGND VPWR VPWR _2166_ sky130_fd_sc_hd__o221a_1
X_3907_ net473 net307 VGND VGND VPWR VPWR _1452_ sky130_fd_sc_hd__nor2_1
XFILLER_177_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4887_ _2096_ _2097_ _1697_ _2087_ VGND VGND VPWR VPWR _2098_ sky130_fd_sc_hd__nand4b_1
XFILLER_165_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6626_ clknet_3_4_0_wb_clk_i _0239_ VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__dfxtp_1
XFILLER_138_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3838_ hkspi.state\[0\] _1382_ VGND VGND VPWR VPWR _1410_ sky130_fd_sc_hd__nand2_1
XFILLER_192_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6557_ clknet_leaf_56_csclk net965 net504 VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__dfrtp_1
XFILLER_180_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3769_ net275 _0910_ _0919_ gpio_configure\[24\]\[0\] _1354_ VGND VGND VPWR VPWR
+ _1355_ sky130_fd_sc_hd__a221o_1
XFILLER_118_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5508_ net441 net1212 _2432_ VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__mux2_1
XFILLER_193_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6488_ clknet_leaf_61_csclk net791 net498 VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__dfstp_2
XFILLER_105_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5439_ _0911_ net647 VGND VGND VPWR VPWR _2425_ sky130_fd_sc_hd__nand2_8
XFILLER_161_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7109_ clknet_leaf_55_csclk net1394 net506 VGND VGND VPWR VPWR gpio_configure\[33\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4810_ _2017_ _2020_ _1947_ _2008_ VGND VGND VPWR VPWR _2021_ sky130_fd_sc_hd__and4b_1
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5790_ gpio_configure\[19\]\[4\] _2491_ _2506_ gpio_configure\[27\]\[4\] VGND VGND
+ VPWR VPWR _2621_ sky130_fd_sc_hd__a22o_1
XFILLER_178_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4741_ _1642_ _1936_ _1943_ VGND VGND VPWR VPWR _1953_ sky130_fd_sc_hd__and3_1
XFILLER_193_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4672_ _1689_ net432 VGND VGND VPWR VPWR _1884_ sky130_fd_sc_hd__or2_1
XFILLER_186_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6411_ net492 net481 VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__and2_1
X_3623_ net63 _1007_ _1057_ gpio_configure\[9\]\[10\] _1201_ VGND VGND VPWR VPWR _1212_
+ sky130_fd_sc_hd__a221o_1
XFILLER_174_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6342_ gpio_configure\[0\]\[12\] _2851_ _3142_ _3151_ _0824_ VGND VGND VPWR VPWR
+ _3152_ sky130_fd_sc_hd__o221a_2
X_3554_ gpio_configure\[19\]\[11\] _1054_ _1098_ gpio_configure\[25\]\[11\] VGND VGND
+ VPWR VPWR _1144_ sky130_fd_sc_hd__a22o_1
XFILLER_142_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6273_ gpio_configure\[14\]\[10\] net411 _2855_ gpio_configure\[27\]\[10\] VGND VGND
+ VPWR VPWR _3085_ sky130_fd_sc_hd__a22o_1
X_3485_ net639 _0973_ VGND VGND VPWR VPWR _1076_ sky130_fd_sc_hd__nor2_8
XFILLER_143_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5224_ net470 net1771 _2399_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__mux2_1
XFILLER_102_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5155_ _2234_ _2282_ _2361_ _1893_ VGND VGND VPWR VPWR _2362_ sky130_fd_sc_hd__or4b_1
XFILLER_84_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4106_ net461 net1730 _1508_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__mux2_1
XFILLER_29_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5086_ _2284_ _2287_ _2288_ _2294_ VGND VGND VPWR VPWR _2295_ sky130_fd_sc_hd__or4_1
XFILLER_110_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4037_ net1638 net455 _1477_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__mux2_1
XFILLER_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5988_ _1448_ _2478_ _2809_ VGND VGND VPWR VPWR _2810_ sky130_fd_sc_hd__and3_4
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4939_ _2144_ _2147_ _2148_ VGND VGND VPWR VPWR _2149_ sky130_fd_sc_hd__or3_1
XFILLER_178_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_40 _1170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_51 _1779_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_62 _2502_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_73 _2791_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_84 gpio_configure\[11\]\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6609_ clknet_leaf_9_csclk net672 net509 VGND VGND VPWR VPWR gpio_configure\[2\]\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_192_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_95 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput180 net180 VGND VGND VPWR VPWR mgmt_gpio_oeb[14] sky130_fd_sc_hd__buf_12
XFILLER_121_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput191 net191 VGND VGND VPWR VPWR mgmt_gpio_oeb[24] sky130_fd_sc_hd__buf_12
XFILLER_0_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_44_csclk clknet_3_6_0_csclk VGND VGND VPWR VPWR clknet_leaf_44_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_140_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3270_ net551 net638 VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__nand2_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_59_csclk clknet_3_2_0_csclk VGND VGND VPWR VPWR clknet_leaf_59_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_97_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6960_ clknet_leaf_56_csclk net1418 net504 VGND VGND VPWR VPWR gpio_configure\[14\]\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_54_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5911_ gpio_configure\[6\]\[10\] _2490_ _2491_ gpio_configure\[19\]\[10\] VGND VGND
+ VPWR VPWR _2736_ sky130_fd_sc_hd__a22o_1
XFILLER_46_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6891_ clknet_leaf_67_csclk net879 net505 VGND VGND VPWR VPWR gpio_configure\[6\]\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_5842_ gpio_configure\[2\]\[7\] _2523_ _2531_ gpio_configure\[24\]\[7\] _2669_ VGND
+ VGND VPWR VPWR _2670_ sky130_fd_sc_hd__a221o_1
XFILLER_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5773_ net475 serial_data_staging_1\[2\] _2604_ VGND VGND VPWR VPWR _2605_ sky130_fd_sc_hd__a21o_1
XFILLER_166_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4724_ _1644_ _1656_ VGND VGND VPWR VPWR _1936_ sky130_fd_sc_hd__nor2_1
XFILLER_147_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4655_ _1678_ _1807_ VGND VGND VPWR VPWR _1867_ sky130_fd_sc_hd__nor2_2
XFILLER_135_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput60 mgmt_gpio_in[31] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_1
X_3606_ gpio_configure\[6\]\[2\] net357 _0908_ gpio_configure\[2\]\[2\] VGND VGND
+ VPWR VPWR _1195_ sky130_fd_sc_hd__a22o_1
Xhold800 _0191_ VGND VGND VPWR VPWR net1333 sky130_fd_sc_hd__dlygate4sd3_1
Xinput71 mgmt_gpio_in[8] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_2
Xhold811 gpio_configure\[3\]\[2\] VGND VGND VPWR VPWR net1344 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput82 spi_sdoenb VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dlymetal6s2s_1
X_4586_ net477 _1797_ VGND VGND VPWR VPWR _1798_ sky130_fd_sc_hd__or2_4
XFILLER_190_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput93 trap VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__buf_4
Xhold822 _0619_ VGND VGND VPWR VPWR net1355 sky130_fd_sc_hd__dlygate4sd3_1
Xhold833 _0539_ VGND VGND VPWR VPWR net1366 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6325_ gpio_configure\[7\]\[12\] _2811_ _2838_ gpio_configure\[12\]\[12\] VGND VGND
+ VPWR VPWR _3135_ sky130_fd_sc_hd__a22o_1
Xhold844 gpio_configure\[25\]\[1\] VGND VGND VPWR VPWR net1377 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3537_ gpio_configure\[24\]\[4\] _0919_ _1127_ gpio_configure\[33\]\[12\] _1126_
+ VGND VGND VPWR VPWR _1128_ sky130_fd_sc_hd__a221o_2
Xhold855 _0495_ VGND VGND VPWR VPWR net1388 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold866 net2129 VGND VGND VPWR VPWR net1399 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold877 _0420_ VGND VGND VPWR VPWR net1410 sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 gpio_configure\[9\]\[1\] VGND VGND VPWR VPWR net1421 sky130_fd_sc_hd__dlygate4sd3_1
X_6256_ gpio_configure\[16\]\[9\] _2831_ _2860_ gpio_configure\[17\]\[9\] _3068_ VGND
+ VGND VPWR VPWR _3069_ sky130_fd_sc_hd__a221o_1
Xhold899 _0121_ VGND VGND VPWR VPWR net1432 sky130_fd_sc_hd__dlygate4sd3_1
X_3468_ _1044_ _1049_ _1052_ _1058_ VGND VGND VPWR VPWR _1059_ sky130_fd_sc_hd__or4_1
X_5207_ net924 net463 _2394_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__mux2_1
XFILLER_76_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6187_ gpio_configure\[21\]\[6\] _2820_ net412 gpio_configure\[9\]\[6\] _3002_ VGND
+ VGND VPWR VPWR _3003_ sky130_fd_sc_hd__a221o_1
X_3399_ gpio_configure\[32\]\[6\] _0890_ _0902_ gpio_configure\[37\]\[6\] _0992_ VGND
+ VGND VPWR VPWR _0993_ sky130_fd_sc_hd__a221o_1
Xhold1500 serial_clock_pre VGND VGND VPWR VPWR net2033 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_191_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1511 serial_data_staging_2\[6\] VGND VGND VPWR VPWR net2044 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1522 _0073_ VGND VGND VPWR VPWR net2055 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1533 hkspi.writemode VGND VGND VPWR VPWR net2066 sky130_fd_sc_hd__dlygate4sd3_1
X_5138_ _2338_ _2345_ VGND VGND VPWR VPWR _2346_ sky130_fd_sc_hd__and2b_1
Xhold1544 irq_2_inputsrc VGND VGND VPWR VPWR net2077 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1555 hkspi.count\[2\] VGND VGND VPWR VPWR net2088 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1566 mgmt_gpio_data_buf\[19\] VGND VGND VPWR VPWR net2099 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1577 mgmt_gpio_data_buf\[0\] VGND VGND VPWR VPWR net2110 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1588 mgmt_gpio_data\[0\] VGND VGND VPWR VPWR net2121 sky130_fd_sc_hd__dlygate4sd3_1
X_5069_ _2276_ _2277_ VGND VGND VPWR VPWR _2278_ sky130_fd_sc_hd__nor2_1
Xhold1599 pad_count_1\[0\] VGND VGND VPWR VPWR net2132 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_40_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4440_ _1634_ _1647_ VGND VGND VPWR VPWR _1652_ sky130_fd_sc_hd__nor2_4
XFILLER_156_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold107 _0925_ VGND VGND VPWR VPWR net640 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold118 _0483_ VGND VGND VPWR VPWR net651 sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 mgmt_gpio_data\[9\] VGND VGND VPWR VPWR net662 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4371_ net110 net99 VGND VGND VPWR VPWR _1583_ sky130_fd_sc_hd__nand2_2
XFILLER_171_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6110_ _2919_ _2928_ VGND VGND VPWR VPWR _2929_ sky130_fd_sc_hd__or2_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3322_ _0881_ net382 VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__nor2_8
XFILLER_140_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7090_ clknet_leaf_77_csclk net1823 net485 VGND VGND VPWR VPWR gpio_configure\[31\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6041_ gpio_configure\[15\]\[0\] net407 net404 gpio_configure\[25\]\[0\] VGND VGND
+ VPWR VPWR _2863_ sky130_fd_sc_hd__a22o_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ net636 net605 _0848_ VGND VGND VPWR VPWR _0849_ sky130_fd_sc_hd__a21bo_1
XFILLER_98_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3184_ hkspi.count\[1\] VGND VGND VPWR VPWR _0814_ sky130_fd_sc_hd__inv_2
XFILLER_78_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6943_ clknet_leaf_37_csclk net1547 net522 VGND VGND VPWR VPWR gpio_configure\[12\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6874_ clknet_leaf_26_csclk net1309 net519 VGND VGND VPWR VPWR gpio_configure\[4\]\[0\]
+ sky130_fd_sc_hd__dfstp_2
X_5825_ _2647_ _2649_ _2651_ _2653_ VGND VGND VPWR VPWR _2654_ sky130_fd_sc_hd__or4_1
XFILLER_50_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5756_ gpio_configure\[5\]\[3\] net422 net420 gpio_configure\[25\]\[3\] VGND VGND
+ VPWR VPWR _2588_ sky130_fd_sc_hd__a22o_1
X_4707_ _1803_ _1863_ VGND VGND VPWR VPWR _1919_ sky130_fd_sc_hd__or2_1
XFILLER_148_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5687_ gpio_configure\[8\]\[0\] _2520_ _2521_ gpio_configure\[21\]\[0\] _2519_ VGND
+ VGND VPWR VPWR _2522_ sky130_fd_sc_hd__a221o_2
XFILLER_162_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4638_ net477 _1692_ VGND VGND VPWR VPWR _1850_ sky130_fd_sc_hd__or2_4
XFILLER_116_550 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold630 _0333_ VGND VGND VPWR VPWR net1163 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4569_ net124 _1774_ VGND VGND VPWR VPWR _1781_ sky130_fd_sc_hd__nor2_1
XFILLER_150_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold641 gpio_configure\[9\]\[4\] VGND VGND VPWR VPWR net1174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold652 _0670_ VGND VGND VPWR VPWR net1185 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap371 _0924_ VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__buf_6
Xhold663 gpio_configure\[6\]\[4\] VGND VGND VPWR VPWR net1196 sky130_fd_sc_hd__dlygate4sd3_1
X_6308_ gpio_configure\[37\]\[11\] net400 net416 gpio_configure\[32\]\[11\] _3107_
+ VGND VGND VPWR VPWR _3119_ sky130_fd_sc_hd__a221o_1
Xmax_cap382 net582 VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__buf_12
Xhold674 _0634_ VGND VGND VPWR VPWR net1207 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap393 _2841_ VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__buf_8
Xhold685 gpio_configure\[10\]\[12\] VGND VGND VPWR VPWR net1218 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold696 _0697_ VGND VGND VPWR VPWR net1229 sky130_fd_sc_hd__dlygate4sd3_1
X_6239_ gpio_configure\[31\]\[8\] _2480_ _2814_ gpio_configure\[11\]\[8\] VGND VGND
+ VPWR VPWR _3053_ sky130_fd_sc_hd__a22o_1
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1330 net1863 VGND VGND VPWR VPWR wb_dat_o[13] sky130_fd_sc_hd__buf_12
Xhold1341 net1958 VGND VGND VPWR VPWR net1874 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1352 net1885 VGND VGND VPWR VPWR wb_dat_o[4] sky130_fd_sc_hd__buf_12
XFILLER_85_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1363 net1953 VGND VGND VPWR VPWR net1896 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1374 _0438_ VGND VGND VPWR VPWR net1907 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1385 gpio_configure\[2\]\[11\] VGND VGND VPWR VPWR net1918 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1396 net332 VGND VGND VPWR VPWR net1929 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3940_ serial_load_pre serial_bb_load serial_bb_enable VGND VGND VPWR VPWR net310
+ sky130_fd_sc_hd__mux2_2
XFILLER_63_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3871_ net58 _1411_ _1426_ net2067 VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__a22o_1
XFILLER_176_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5610_ xfer_state\[0\] xfer_state\[2\] VGND VGND VPWR VPWR _2458_ sky130_fd_sc_hd__or2_1
XFILLER_177_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6590_ clknet_leaf_56_csclk net863 net504 VGND VGND VPWR VPWR mgmt_gpio_data_buf\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_31_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5541_ net794 net660 _2436_ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__mux2_1
XFILLER_157_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5472_ net1142 net441 _2428_ VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__mux2_1
XFILLER_172_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7211_ clknet_leaf_75_csclk net1008 net485 VGND VGND VPWR VPWR gpio_configure\[27\]\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_160_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4423_ _1617_ _1628_ _1633_ VGND VGND VPWR VPWR _1635_ sky130_fd_sc_hd__and3_4
X_7142_ clknet_leaf_35_csclk net604 net525 VGND VGND VPWR VPWR gpio_configure\[37\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_4354_ _1558_ _1565_ VGND VGND VPWR VPWR _1566_ sky130_fd_sc_hd__nand2_1
XFILLER_99_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3305_ net600 _0880_ VGND VGND VPWR VPWR _0901_ sky130_fd_sc_hd__nand2_8
Xfanout428 net646 VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__buf_12
XFILLER_59_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7073_ clknet_leaf_33_csclk net929 net525 VGND VGND VPWR VPWR gpio_configure\[28\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
Xfanout439 net634 VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__buf_12
X_4285_ net455 net1666 _1539_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__mux2_1
XFILLER_113_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6024_ net417 net415 net410 net409 VGND VGND VPWR VPWR _2846_ sky130_fd_sc_hd__or4_1
XFILLER_100_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3236_ net110 VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__clkinv_2
XFILLER_39_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6926_ clknet_leaf_16_csclk net1285 net512 VGND VGND VPWR VPWR gpio_configure\[10\]\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_81_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6857_ clknet_leaf_41_csclk net1044 net517 VGND VGND VPWR VPWR gpio_configure\[1\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5808_ gpio_configure\[26\]\[5\] _2534_ _2537_ gpio_configure\[17\]\[5\] _2637_ VGND
+ VGND VPWR VPWR _2638_ sky130_fd_sc_hd__a221o_1
XFILLER_167_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6788_ clknet_2_2__leaf_mgmt_gpio_in[4] net2002 _0062_ VGND VGND VPWR VPWR hkspi.ldata\[5\]
+ sky130_fd_sc_hd__dfrtn_1
XFILLER_183_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5739_ gpio_configure\[6\]\[2\] _2490_ _2498_ gpio_configure\[22\]\[2\] _2571_ VGND
+ VGND VPWR VPWR _2572_ sky130_fd_sc_hd__a221o_1
XFILLER_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold460 _0377_ VGND VGND VPWR VPWR net993 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold471 _0111_ VGND VGND VPWR VPWR net1004 sky130_fd_sc_hd__dlygate4sd3_1
Xhold482 net287 VGND VGND VPWR VPWR net1015 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold493 _0648_ VGND VGND VPWR VPWR net1026 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1160 _0106_ VGND VGND VPWR VPWR net1693 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1171 net301 VGND VGND VPWR VPWR net1704 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1182 net300 VGND VGND VPWR VPWR net1715 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1193 gpio_configure\[31\]\[2\] VGND VGND VPWR VPWR net1726 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_2__f_mgmt_gpio_in[4] clknet_0_mgmt_gpio_in[4] VGND VGND VPWR VPWR clknet_2_2__leaf_mgmt_gpio_in[4]
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_154_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4070_ _0909_ net483 _1480_ net351 net426 VGND VGND VPWR VPWR _1490_ sky130_fd_sc_hd__o221a_4
XFILLER_110_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4972_ _1768_ _2004_ _2181_ _1992_ _1693_ VGND VGND VPWR VPWR _2182_ sky130_fd_sc_hd__o32ai_4
XFILLER_17_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6711_ clknet_leaf_9_csclk net1784 net509 VGND VGND VPWR VPWR gpio_configure\[16\]\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_3923_ mgmt_gpio_data\[32\] net80 net79 VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__mux2_8
XFILLER_20_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6642_ clknet_3_4_0_wb_clk_i _0255_ VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__dfxtp_1
X_3854_ _1416_ _1420_ VGND VGND VPWR VPWR _1421_ sky130_fd_sc_hd__nor2_1
XFILLER_20_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6573_ clknet_leaf_36_csclk net805 net522 VGND VGND VPWR VPWR mgmt_gpio_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_192_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3785_ net93 _0852_ _0882_ _1047_ gpio_configure\[18\]\[8\] VGND VGND VPWR VPWR _1371_
+ sky130_fd_sc_hd__a32o_1
XFILLER_164_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5524_ net452 net972 _2434_ VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__mux2_1
XFILLER_118_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5455_ net437 net1469 _2426_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__mux2_1
XFILLER_133_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4406_ _1604_ _1615_ _1616_ VGND VGND VPWR VPWR _1618_ sky130_fd_sc_hd__nand3_2
X_5386_ net470 net1738 _2419_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__mux2_1
XFILLER_120_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7125_ clknet_leaf_33_csclk net649 net524 VGND VGND VPWR VPWR gpio_configure\[35\]\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_101_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4337_ net107 net106 net109 net108 VGND VGND VPWR VPWR _1549_ sky130_fd_sc_hd__and4_1
XFILLER_101_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7056_ clknet_leaf_58_csclk net1424 net503 VGND VGND VPWR VPWR gpio_configure\[26\]\[6\]
+ sky130_fd_sc_hd__dfrtp_2
X_4268_ net1110 net449 _1536_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__mux2_1
XFILLER_86_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6007_ _1447_ _2801_ VGND VGND VPWR VPWR _2829_ sky130_fd_sc_hd__nor2_8
X_3219_ gpio_configure\[15\]\[3\] VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__inv_2
X_4199_ net1804 net468 _1521_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__mux2_1
XFILLER_55_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6909_ clknet_leaf_29_csclk net979 net520 VGND VGND VPWR VPWR gpio_configure\[8\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_23_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold290 _0220_ VGND VGND VPWR VPWR net823 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_130 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_141 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_152 net298 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_163 net405 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_174 clknet_3_6_0_wb_clk_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_185 clknet_2_0__leaf_mgmt_gpio_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_196 _1160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3570_ gpio_configure\[16\]\[3\] _0912_ net350 gpio_configure\[4\]\[3\] _1159_ VGND
+ VGND VPWR VPWR _1160_ sky130_fd_sc_hd__a221o_1
XFILLER_115_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5240_ net435 net932 _2402_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__mux2_1
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5171_ _2322_ _2376_ VGND VGND VPWR VPWR _2377_ sky130_fd_sc_hd__nor2_1
X_4122_ net462 net1455 _1510_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__mux2_1
XFILLER_68_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4053_ _0903_ net483 _1480_ _0904_ net429 VGND VGND VPWR VPWR _1481_ sky130_fd_sc_hd__o221a_4
Xinput3 debug_out VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XFILLER_110_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4955_ _1674_ _2143_ _2039_ VGND VGND VPWR VPWR _2165_ sky130_fd_sc_hd__a21oi_1
XFILLER_51_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3906_ _1447_ _1450_ VGND VGND VPWR VPWR _1451_ sky130_fd_sc_hd__or2_1
XFILLER_189_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4886_ _1636_ _2081_ _1970_ _1669_ VGND VGND VPWR VPWR _2097_ sky130_fd_sc_hd__o211a_1
X_6625_ clknet_leaf_10_csclk net1203 net511 VGND VGND VPWR VPWR gpio_configure\[5\]\[12\]
+ sky130_fd_sc_hd__dfrtp_2
X_3837_ _0821_ net2146 _1409_ hkspi.pass_thru_user VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__a31o_1
X_6556_ clknet_leaf_56_csclk net1084 net504 VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__dfrtp_1
XFILLER_20_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3768_ gpio_configure\[23\]\[8\] _1067_ _1073_ gpio_configure\[24\]\[8\] VGND VGND
+ VPWR VPWR _1354_ sky130_fd_sc_hd__a22o_1
X_5507_ net446 net1176 _2432_ VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__mux2_1
XFILLER_180_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6487_ clknet_leaf_71_csclk net674 net498 VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__dfstp_1
X_3699_ gpio_configure\[17\]\[1\] net367 _1076_ gpio_configure\[27\]\[9\] VGND VGND
+ VPWR VPWR _1287_ sky130_fd_sc_hd__a22o_1
XFILLER_118_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5438_ net434 net1312 _2424_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__mux2_1
Xoutput340 net1888 VGND VGND VPWR VPWR net1889 sky130_fd_sc_hd__buf_12
XFILLER_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5369_ net464 net1371 _2417_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__mux2_1
XFILLER_126_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7108_ clknet_leaf_31_csclk net957 net523 VGND VGND VPWR VPWR gpio_configure\[33\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7039_ clknet_leaf_39_csclk net1143 net516 VGND VGND VPWR VPWR gpio_configure\[24\]\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_28_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire412 _2835_ VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__buf_12
XFILLER_183_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4740_ _1642_ _1936_ VGND VGND VPWR VPWR _1952_ sky130_fd_sc_hd__nand2_1
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4671_ _1689_ net432 VGND VGND VPWR VPWR _1883_ sky130_fd_sc_hd__nor2_2
XFILLER_186_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6410_ net492 net482 VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__and2_1
X_3622_ gpio_configure\[36\]\[10\] _1109_ _1205_ _1209_ _1210_ VGND VGND VPWR VPWR
+ _1211_ sky130_fd_sc_hd__a2111o_1
XFILLER_147_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6341_ net364 _3144_ _3146_ _3150_ VGND VGND VPWR VPWR _3151_ sky130_fd_sc_hd__or4_1
X_3553_ gpio_configure\[20\]\[3\] _0928_ _1047_ gpio_configure\[18\]\[11\] VGND VGND
+ VPWR VPWR _1143_ sky130_fd_sc_hd__a22o_1
XFILLER_115_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6272_ gpio_configure\[28\]\[10\] _2861_ VGND VGND VPWR VPWR _3084_ sky130_fd_sc_hd__and2_1
X_3484_ _1061_ _1066_ _1071_ _1074_ VGND VGND VPWR VPWR _1075_ sky130_fd_sc_hd__or4_1
XFILLER_170_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5223_ _1313_ net429 VGND VGND VPWR VPWR _2399_ sky130_fd_sc_hd__nand2_1
XFILLER_102_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5154_ net424 net432 _1841_ VGND VGND VPWR VPWR _2361_ sky130_fd_sc_hd__a21oi_1
X_4105_ net466 net1742 _1508_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__mux2_1
XFILLER_57_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5085_ _0832_ _1695_ _2290_ _2292_ _2293_ VGND VGND VPWR VPWR _2294_ sky130_fd_sc_hd__a2111o_1
XFILLER_56_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4036_ net1654 net461 _1477_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__mux2_1
XFILLER_52_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5987_ pad_count_2\[2\] pad_count_2\[3\] VGND VGND VPWR VPWR _2809_ sky130_fd_sc_hd__and2b_2
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4938_ net126 _1571_ _2146_ _1867_ _1718_ VGND VGND VPWR VPWR _2148_ sky130_fd_sc_hd__a311o_1
XFILLER_178_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_30 _1072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_41 _1209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4869_ _2056_ _2079_ _1582_ VGND VGND VPWR VPWR _2080_ sky130_fd_sc_hd__o21ba_1
XFILLER_20_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_52 _2407_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_63 _2506_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6608_ clknet_leaf_9_csclk net775 net509 VGND VGND VPWR VPWR gpio_configure\[2\]\[10\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA_74 _2808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_85 gpio_configure\[14\]\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_96 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6539_ clknet_leaf_2_csclk net1295 net493 VGND VGND VPWR VPWR gpio_configure\[26\]\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_106_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput181 net181 VGND VGND VPWR VPWR mgmt_gpio_oeb[15] sky130_fd_sc_hd__buf_12
Xoutput192 net192 VGND VGND VPWR VPWR mgmt_gpio_oeb[25] sky130_fd_sc_hd__buf_12
XFILLER_153_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5910_ gpio_configure\[2\]\[10\] _2523_ _2734_ VGND VGND VPWR VPWR _2735_ sky130_fd_sc_hd__a21o_1
X_6890_ clknet_leaf_15_csclk net1565 net519 VGND VGND VPWR VPWR gpio_configure\[6\]\[0\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5841_ gpio_configure\[14\]\[7\] _2494_ _2540_ gpio_configure\[12\]\[7\] VGND VGND
+ VPWR VPWR _2669_ sky130_fd_sc_hd__a22o_1
XFILLER_62_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5772_ gpio_configure\[0\]\[3\] _2526_ _2602_ _2603_ net473 VGND VGND VPWR VPWR _2604_
+ sky130_fd_sc_hd__o221a_2
X_4723_ _1862_ _1934_ _1529_ _1860_ VGND VGND VPWR VPWR _1935_ sky130_fd_sc_hd__a211o_1
XFILLER_175_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4654_ net111 _1435_ net112 VGND VGND VPWR VPWR _1866_ sky130_fd_sc_hd__or3b_4
X_3605_ gpio_configure\[32\]\[2\] _0890_ _0898_ gpio_configure\[0\]\[2\] VGND VGND
+ VPWR VPWR _1194_ sky130_fd_sc_hd__a22o_1
XFILLER_174_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput50 mgmt_gpio_in[22] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__buf_2
XFILLER_190_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput61 mgmt_gpio_in[32] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold801 gpio_configure\[0\]\[6\] VGND VGND VPWR VPWR net1334 sky130_fd_sc_hd__dlygate4sd3_1
Xinput72 mgmt_gpio_in[9] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_1
XFILLER_116_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4585_ net127 net128 _1553_ VGND VGND VPWR VPWR _1797_ sky130_fd_sc_hd__or3b_4
Xhold812 _0471_ VGND VGND VPWR VPWR net1345 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_174_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold823 gpio_configure\[1\]\[6\] VGND VGND VPWR VPWR net1356 sky130_fd_sc_hd__dlygate4sd3_1
Xinput83 spimemio_flash_clk VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__buf_2
Xinput94 uart_enabled VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_1
Xhold834 gpio_configure\[28\]\[6\] VGND VGND VPWR VPWR net1367 sky130_fd_sc_hd__dlygate4sd3_1
X_6324_ gpio_configure\[29\]\[12\] _2816_ _2820_ gpio_configure\[21\]\[12\] _3133_
+ VGND VGND VPWR VPWR _3134_ sky130_fd_sc_hd__a221o_1
XFILLER_115_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3536_ net387 _0885_ VGND VGND VPWR VPWR _1127_ sky130_fd_sc_hd__nor2_2
Xhold845 _0646_ VGND VGND VPWR VPWR net1378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 gpio_configure\[9\]\[10\] VGND VGND VPWR VPWR net1389 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold867 _0720_ VGND VGND VPWR VPWR net1400 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold878 gpio_configure\[35\]\[1\] VGND VGND VPWR VPWR net1411 sky130_fd_sc_hd__dlygate4sd3_1
X_6255_ gpio_configure\[14\]\[9\] net411 _2855_ gpio_configure\[27\]\[9\] VGND VGND
+ VPWR VPWR _3068_ sky130_fd_sc_hd__a22o_1
Xhold889 _0518_ VGND VGND VPWR VPWR net1422 sky130_fd_sc_hd__dlygate4sd3_1
X_3467_ gpio_configure\[12\]\[12\] _1056_ _1057_ gpio_configure\[9\]\[12\] _1055_
+ VGND VGND VPWR VPWR _1058_ sky130_fd_sc_hd__a221o_1
X_5206_ net1704 net469 _2394_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__mux2_1
XFILLER_88_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6186_ gpio_configure\[23\]\[6\] _2822_ _2861_ gpio_configure\[28\]\[6\] VGND VGND
+ VPWR VPWR _3002_ sky130_fd_sc_hd__a22o_1
X_3398_ gpio_configure\[19\]\[6\] _0896_ _0910_ net297 VGND VGND VPWR VPWR _0992_
+ sky130_fd_sc_hd__a22o_1
Xhold1501 serial_data_staging_1\[3\] VGND VGND VPWR VPWR net2034 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1512 hkspi.odata\[1\] VGND VGND VPWR VPWR net2045 sky130_fd_sc_hd__dlygate4sd3_1
X_5137_ _1691_ _2340_ _2342_ _2344_ VGND VGND VPWR VPWR _2345_ sky130_fd_sc_hd__or4_1
Xhold1523 serial_data_staging_1\[4\] VGND VGND VPWR VPWR net2056 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1534 hkspi.pre_pass_thru_user VGND VGND VPWR VPWR net2067 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1545 hkspi.addr\[7\] VGND VGND VPWR VPWR net2078 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1556 serial_data_staging_1\[9\] VGND VGND VPWR VPWR net2089 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_123_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1567 mgmt_gpio_data_buf\[1\] VGND VGND VPWR VPWR net2100 sky130_fd_sc_hd__dlygate4sd3_1
X_5068_ _2055_ _2140_ VGND VGND VPWR VPWR _2277_ sky130_fd_sc_hd__or2_1
XFILLER_84_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1578 mgmt_gpio_data_buf\[14\] VGND VGND VPWR VPWR net2111 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1589 xfer_count\[3\] VGND VGND VPWR VPWR net2122 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4019_ net456 net1403 _1474_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__mux2_1
XFILLER_37_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold108 _2431_ VGND VGND VPWR VPWR net641 sky130_fd_sc_hd__clkbuf_8
XFILLER_156_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold119 gpio_configure\[22\]\[7\] VGND VGND VPWR VPWR net652 sky130_fd_sc_hd__dlygate4sd3_1
X_4370_ _1576_ _1581_ wbbd_state\[9\] VGND VGND VPWR VPWR _1582_ sky130_fd_sc_hd__o21ai_1
XFILLER_125_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3321_ net387 net601 VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__nor2_8
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6040_ _2471_ _2478_ _2809_ VGND VGND VPWR VPWR _2862_ sky130_fd_sc_hd__and3_4
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ hkspi.addr\[5\] _0819_ VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__nand2_1
XFILLER_140_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6942_ clknet_leaf_15_csclk net1209 net513 VGND VGND VPWR VPWR gpio_configure\[12\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6873_ clknet_leaf_41_csclk net1052 net517 VGND VGND VPWR VPWR gpio_configure\[3\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_62_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5824_ gpio_configure\[6\]\[6\] _2490_ _2506_ gpio_configure\[27\]\[6\] _2652_ VGND
+ VGND VPWR VPWR _2653_ sky130_fd_sc_hd__a221o_1
XFILLER_179_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5755_ gpio_configure\[17\]\[3\] _2537_ _2541_ gpio_configure\[31\]\[3\] VGND VGND
+ VPWR VPWR _2587_ sky130_fd_sc_hd__a22o_1
X_4706_ _1803_ _1874_ _1904_ _1917_ VGND VGND VPWR VPWR _1918_ sky130_fd_sc_hd__o211a_1
X_5686_ pad_count_1\[4\] _2488_ _2495_ VGND VGND VPWR VPWR _2521_ sky130_fd_sc_hd__and3_4
XFILLER_148_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4637_ _1693_ _1750_ net424 _1788_ _1848_ VGND VGND VPWR VPWR _1849_ sky130_fd_sc_hd__o221a_1
XFILLER_190_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold620 _0592_ VGND VGND VPWR VPWR net1153 sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 gpio_configure\[35\]\[12\] VGND VGND VPWR VPWR net1164 sky130_fd_sc_hd__dlygate4sd3_1
X_4568_ _1776_ _1779_ VGND VGND VPWR VPWR _1780_ sky130_fd_sc_hd__or2_1
XFILLER_162_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap350 net563 VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__buf_8
XFILLER_116_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold642 _0521_ VGND VGND VPWR VPWR net1175 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold653 net2134 VGND VGND VPWR VPWR net1186 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap361 net362 VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__clkbuf_2
Xmax_cap372 _0922_ VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__buf_6
X_6307_ gpio_configure\[28\]\[11\] _2861_ _3113_ _3115_ _3117_ VGND VGND VPWR VPWR
+ _3118_ sky130_fd_sc_hd__a2111o_1
X_3519_ net554 _1008_ VGND VGND VPWR VPWR _1110_ sky130_fd_sc_hd__nor2_4
Xhold664 _0497_ VGND VGND VPWR VPWR net1197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 gpio_configure\[12\]\[4\] VGND VGND VPWR VPWR net1208 sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 _0287_ VGND VGND VPWR VPWR net1219 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4499_ _0832_ net99 _1710_ _1701_ _1696_ VGND VGND VPWR VPWR _1711_ sky130_fd_sc_hd__o311a_1
Xhold697 gpio_configure\[13\]\[12\] VGND VGND VPWR VPWR net1230 sky130_fd_sc_hd__dlygate4sd3_1
X_6238_ gpio_configure\[2\]\[8\] net398 _2843_ gpio_configure\[5\]\[8\] _3051_ VGND
+ VGND VPWR VPWR _3052_ sky130_fd_sc_hd__a221o_1
XFILLER_103_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ gpio_configure\[0\]\[5\] _2851_ _2973_ _2985_ net473 VGND VGND VPWR VPWR _2986_
+ sky130_fd_sc_hd__o221a_2
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1320 net1853 VGND VGND VPWR VPWR wb_dat_o[23] sky130_fd_sc_hd__buf_12
Xhold1331 net1944 VGND VGND VPWR VPWR net1864 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1342 net1875 VGND VGND VPWR VPWR wb_dat_o[11] sky130_fd_sc_hd__buf_12
XFILLER_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1353 net1978 VGND VGND VPWR VPWR net1886 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1364 net1897 VGND VGND VPWR VPWR wb_dat_o[16] sky130_fd_sc_hd__buf_12
XFILLER_57_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1375 gpio_configure\[37\]\[7\] VGND VGND VPWR VPWR net1908 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1386 gpio_configure\[25\]\[7\] VGND VGND VPWR VPWR net1919 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1397 net324 VGND VGND VPWR VPWR net1930 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_43_csclk clknet_3_6_0_csclk VGND VGND VPWR VPWR clknet_leaf_43_csclk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_58_csclk clknet_3_2_0_csclk VGND VGND VPWR VPWR clknet_leaf_58_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_185_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3870_ hkspi.count\[0\] hkspi.pre_pass_thru_mgmt _1410_ VGND VGND VPWR VPWR _1426_
+ sky130_fd_sc_hd__a21o_1
XFILLER_177_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5540_ net792 net445 _2436_ VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__mux2_1
XFILLER_129_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5471_ net734 net445 _2428_ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__mux2_1
XFILLER_172_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7210_ clknet_leaf_75_csclk net1056 net485 VGND VGND VPWR VPWR gpio_configure\[27\]\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_4422_ _1617_ _1633_ VGND VGND VPWR VPWR _1634_ sky130_fd_sc_hd__nand2_1
X_7141_ clknet_leaf_56_csclk net1440 net504 VGND VGND VPWR VPWR gpio_configure\[37\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_132_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4353_ _1553_ _1557_ net127 VGND VGND VPWR VPWR _1565_ sky130_fd_sc_hd__a21o_1
X_3304_ net389 _0899_ VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__nor2_4
X_7072_ clknet_leaf_51_csclk net1368 net506 VGND VGND VPWR VPWR gpio_configure\[28\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_4284_ net461 net1694 _1539_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__mux2_1
XFILLER_98_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout429 net645 VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__buf_12
XFILLER_140_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6023_ _2795_ _2806_ _2830_ _2840_ VGND VGND VPWR VPWR _2845_ sky130_fd_sc_hd__or4_1
X_3235_ pad_count_1\[4\] VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__clkinv_8
XFILLER_101_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6925_ clknet_leaf_40_csclk net729 net516 VGND VGND VPWR VPWR gpio_configure\[10\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_82_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6856_ clknet_leaf_53_csclk net1357 net506 VGND VGND VPWR VPWR gpio_configure\[1\]\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_120_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5807_ gpio_configure\[4\]\[5\] _2502_ _2510_ gpio_configure\[15\]\[5\] VGND VGND
+ VPWR VPWR _2637_ sky130_fd_sc_hd__a22o_1
XFILLER_167_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3999_ net776 net439 _1471_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__mux2_1
X_6787_ clknet_2_2__leaf_mgmt_gpio_in[4] _0390_ _0061_ VGND VGND VPWR VPWR hkspi.ldata\[4\]
+ sky130_fd_sc_hd__dfrtn_1
XFILLER_183_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5738_ gpio_configure\[18\]\[2\] _2532_ _2540_ gpio_configure\[12\]\[2\] VGND VGND
+ VPWR VPWR _2571_ sky130_fd_sc_hd__a22o_1
XFILLER_129_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5669_ pad_count_1\[2\] pad_count_1\[3\] VGND VGND VPWR VPWR _2504_ sky130_fd_sc_hd__and2b_2
XFILLER_136_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold450 _0544_ VGND VGND VPWR VPWR net983 sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 gpio_configure\[8\]\[12\] VGND VGND VPWR VPWR net994 sky130_fd_sc_hd__dlygate4sd3_1
Xhold472 net2099 VGND VGND VPWR VPWR net1005 sky130_fd_sc_hd__dlygate4sd3_1
Xhold483 _0100_ VGND VGND VPWR VPWR net1016 sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 gpio_configure\[8\]\[11\] VGND VGND VPWR VPWR net1027 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1150 _0398_ VGND VGND VPWR VPWR net1683 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_161_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1161 gpio_configure\[18\]\[9\] VGND VGND VPWR VPWR net1694 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1172 _0410_ VGND VGND VPWR VPWR net1705 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1183 _0105_ VGND VGND VPWR VPWR net1716 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1194 _0122_ VGND VGND VPWR VPWR net1727 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_699 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_1_0_wb_clk_i clknet_1_0_1_wb_clk_i VGND VGND VPWR VPWR clknet_2_1_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_68_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4971_ _1744_ _1749_ VGND VGND VPWR VPWR _2181_ sky130_fd_sc_hd__nor2_1
XFILLER_64_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6710_ clknet_leaf_5_csclk net1221 net494 VGND VGND VPWR VPWR gpio_configure\[15\]\[12\]
+ sky130_fd_sc_hd__dfrtp_2
X_3922_ _0828_ net82 net79 VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__mux2_8
XFILLER_51_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3853_ hkspi.fixed\[0\] _1419_ VGND VGND VPWR VPWR _1420_ sky130_fd_sc_hd__nor2_1
X_6641_ clknet_3_4_0_wb_clk_i _0254_ VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__dfxtp_1
XFILLER_20_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3784_ gpio_configure\[25\]\[0\] _0927_ _1098_ gpio_configure\[25\]\[8\] _1369_ VGND
+ VGND VPWR VPWR _1370_ sky130_fd_sc_hd__a221o_1
X_6572_ clknet_leaf_31_csclk net883 net523 VGND VGND VPWR VPWR mgmt_gpio_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_118_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5523_ net457 net746 _2434_ VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__mux2_1
XFILLER_157_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5454_ net660 net824 _2426_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__mux2_1
X_4405_ _1604_ _1615_ _1616_ VGND VGND VPWR VPWR _1617_ sky130_fd_sc_hd__and3_4
X_5385_ _0918_ net646 VGND VGND VPWR VPWR _2419_ sky130_fd_sc_hd__nand2_8
XFILLER_99_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7124_ clknet_leaf_32_csclk net1521 net524 VGND VGND VPWR VPWR gpio_configure\[35\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_4336_ net112 net114 net113 VGND VGND VPWR VPWR _1548_ sky130_fd_sc_hd__or3_4
XFILLER_59_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7055_ clknet_leaf_38_csclk net1557 net522 VGND VGND VPWR VPWR gpio_configure\[26\]\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_4267_ net744 net457 _1536_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__mux2_1
XFILLER_59_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6006_ _2479_ _2794_ VGND VGND VPWR VPWR _2828_ sky130_fd_sc_hd__nor2_8
X_3218_ gpio_configure\[16\]\[3\] VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__inv_2
XFILLER_39_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4198_ _1094_ net429 VGND VGND VPWR VPWR _1521_ sky130_fd_sc_hd__and2_2
XFILLER_39_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_614 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6908_ clknet_leaf_15_csclk net801 net519 VGND VGND VPWR VPWR gpio_configure\[8\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_6839_ clknet_leaf_30_csclk net975 net520 VGND VGND VPWR VPWR mgmt_gpio_data_buf\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold280 _0600_ VGND VGND VPWR VPWR net813 sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 gpio_configure\[22\]\[5\] VGND VGND VPWR VPWR net824 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_120 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_131 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_142 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_153 net298 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_164 net405 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_175 clknet_3_6_0_wb_clk_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_186 net612 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_197 _1270_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5170_ _2196_ _2299_ _2352_ _2375_ VGND VGND VPWR VPWR _2376_ sky130_fd_sc_hd__or4b_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4121_ net466 net1510 _1510_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__mux2_1
XFILLER_96_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4052_ net483 _0871_ VGND VGND VPWR VPWR _1480_ sky130_fd_sc_hd__and2b_4
Xinput4 mask_rev_in[0] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4954_ _1988_ _2160_ _2162_ _2163_ VGND VGND VPWR VPWR _2164_ sky130_fd_sc_hd__or4_1
X_3905_ _1448_ _1449_ VGND VGND VPWR VPWR _1450_ sky130_fd_sc_hd__nand2_4
XFILLER_20_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4885_ _1944_ _2092_ _2094_ _2095_ VGND VGND VPWR VPWR _2096_ sky130_fd_sc_hd__or4_1
XFILLER_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6624_ clknet_leaf_10_csclk net715 net511 VGND VGND VPWR VPWR gpio_configure\[5\]\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_165_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3836_ hkspi.state\[3\] hkspi.state\[0\] hkspi.state\[4\] VGND VGND VPWR VPWR _1409_
+ sky130_fd_sc_hd__nor3_1
XFILLER_177_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3767_ gpio_configure\[32\]\[8\] _1101_ _1116_ gpio_configure\[26\]\[8\] VGND VGND
+ VPWR VPWR _1353_ sky130_fd_sc_hd__a22o_1
X_6555_ clknet_leaf_2_csclk net1573 net492 VGND VGND VPWR VPWR mgmt_gpio_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_118_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5506_ net452 net1009 _2432_ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__mux2_1
X_6486_ clknet_leaf_72_csclk net1020 net490 VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__dfrtp_1
X_3698_ gpio_configure\[31\]\[1\] net375 _0923_ gpio_configure\[22\]\[1\] _1285_ VGND
+ VGND VPWR VPWR _1286_ sky130_fd_sc_hd__a221o_1
XFILLER_106_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5437_ net437 net1471 _2424_ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__mux2_1
XFILLER_105_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput330 net1892 VGND VGND VPWR VPWR net1893 sky130_fd_sc_hd__buf_12
XFILLER_133_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput341 net1850 VGND VGND VPWR VPWR net1851 sky130_fd_sc_hd__buf_12
X_5368_ net471 net1582 _2417_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__mux2_1
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7107_ clknet_leaf_20_csclk net1187 net511 VGND VGND VPWR VPWR gpio_configure\[33\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_4319_ net1834 net466 _1545_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__mux2_1
X_5299_ net452 net998 _2409_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__mux2_1
XFILLER_59_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7038_ clknet_leaf_60_csclk net735 net498 VGND VGND VPWR VPWR gpio_configure\[24\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_28_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4670_ _1613_ _1689_ VGND VGND VPWR VPWR _1882_ sky130_fd_sc_hd__nor2_1
XFILLER_159_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3621_ gpio_configure\[13\]\[10\] _1045_ _1121_ gpio_configure\[17\]\[10\] _1204_
+ VGND VGND VPWR VPWR _1210_ sky130_fd_sc_hd__a221o_1
XFILLER_174_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3552_ gpio_configure\[32\]\[3\] _0890_ _0974_ serial_bb_load VGND VGND VPWR VPWR
+ _1142_ sky130_fd_sc_hd__a22o_1
X_6340_ gpio_configure\[10\]\[12\] net414 _3147_ _3149_ VGND VGND VPWR VPWR _3150_
+ sky130_fd_sc_hd__a211o_1
XFILLER_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6271_ gpio_configure\[36\]\[10\] net403 net402 gpio_configure\[4\]\[10\] VGND VGND
+ VPWR VPWR _3083_ sky130_fd_sc_hd__a22o_2
XFILLER_142_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3483_ gpio_configure\[28\]\[4\] _0888_ _1073_ gpio_configure\[24\]\[12\] _1072_
+ VGND VGND VPWR VPWR _1074_ sky130_fd_sc_hd__a221o_1
XFILLER_115_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5222_ net383 _0973_ net469 net1500 net427 VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__o311a_1
XFILLER_130_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5153_ _2127_ _2293_ _2359_ VGND VGND VPWR VPWR _2360_ sky130_fd_sc_hd__or3b_1
XFILLER_96_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4104_ _1007_ net429 VGND VGND VPWR VPWR _1508_ sky130_fd_sc_hd__nand2_8
X_5084_ _1805_ _2233_ _2285_ _1798_ _2120_ VGND VGND VPWR VPWR _2293_ sky130_fd_sc_hd__o221ai_2
XFILLER_84_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4035_ net1836 net466 _1477_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__mux2_1
XFILLER_56_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5986_ gpio_configure\[36\]\[0\] net403 net402 gpio_configure\[4\]\[0\] _2807_ VGND
+ VGND VPWR VPWR _2808_ sky130_fd_sc_hd__a221o_2
XFILLER_24_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4937_ _1674_ _2146_ _2074_ VGND VGND VPWR VPWR _2147_ sky130_fd_sc_hd__a21o_1
XFILLER_33_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_20 _1004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_31 _1092_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4868_ _2049_ _2055_ _2057_ _2078_ VGND VGND VPWR VPWR _2079_ sky130_fd_sc_hd__or4_1
XANTENNA_42 _1217_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_53 _2430_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_64 _2517_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6607_ clknet_leaf_9_csclk net823 net509 VGND VGND VPWR VPWR gpio_configure\[2\]\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_75 _2808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3819_ _1398_ hkspi.addr\[5\] _1388_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__mux2_1
X_4799_ _1651_ _1745_ net424 _1807_ VGND VGND VPWR VPWR _2010_ sky130_fd_sc_hd__o22a_1
XANTENNA_86 gpio_configure\[15\]\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_97 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6538_ clknet_leaf_0_csclk net1630 net487 VGND VGND VPWR VPWR gpio_configure\[26\]\[10\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_21_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6469_ clknet_2_0__leaf_mgmt_gpio_in[4] _0091_ _0047_ VGND VGND VPWR VPWR hkspi.addr\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_161_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput171 net171 VGND VGND VPWR VPWR debug_in sky130_fd_sc_hd__buf_12
XFILLER_133_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput182 net182 VGND VGND VPWR VPWR mgmt_gpio_oeb[16] sky130_fd_sc_hd__buf_12
Xoutput193 net193 VGND VGND VPWR VPWR mgmt_gpio_oeb[26] sky130_fd_sc_hd__buf_12
XFILLER_121_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5840_ gpio_configure\[10\]\[7\] _2507_ _2529_ gpio_configure\[29\]\[7\] _2667_ VGND
+ VGND VPWR VPWR _2668_ sky130_fd_sc_hd__a221o_1
XFILLER_34_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5771_ _2590_ _2592_ _2594_ VGND VGND VPWR VPWR _2603_ sky130_fd_sc_hd__or3_1
X_4722_ _1869_ _1927_ _1932_ VGND VGND VPWR VPWR _1934_ sky130_fd_sc_hd__or3_1
XFILLER_187_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4653_ net477 _1678_ _1822_ VGND VGND VPWR VPWR _1865_ sky130_fd_sc_hd__or3_1
Xinput40 mgmt_gpio_in[13] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dlymetal6s2s_1
X_3604_ gpio_configure\[37\]\[2\] _0902_ _1136_ net303 VGND VGND VPWR VPWR _1193_
+ sky130_fd_sc_hd__a22o_1
XFILLER_175_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput51 mgmt_gpio_in[23] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_2
Xhold802 _0451_ VGND VGND VPWR VPWR net1335 sky130_fd_sc_hd__dlygate4sd3_1
X_4584_ _1689_ _1750_ _1790_ _1795_ VGND VGND VPWR VPWR _1796_ sky130_fd_sc_hd__o22a_1
Xinput62 mgmt_gpio_in[33] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_2
Xinput73 pad_flash_io0_di VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_1
Xhold813 gpio_configure\[10\]\[6\] VGND VGND VPWR VPWR net1346 sky130_fd_sc_hd__dlygate4sd3_1
Xinput84 spimemio_flash_csb VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__buf_2
Xhold824 _0459_ VGND VGND VPWR VPWR net1357 sky130_fd_sc_hd__dlygate4sd3_1
X_6323_ gpio_configure\[31\]\[12\] net423 net408 gpio_configure\[35\]\[12\] VGND VGND
+ VPWR VPWR _3133_ sky130_fd_sc_hd__a22o_1
XFILLER_155_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput95 usr1_vcc_pwrgood VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__buf_2
Xhold835 _0675_ VGND VGND VPWR VPWR net1368 sky130_fd_sc_hd__dlygate4sd3_1
X_3535_ gpio_configure\[12\]\[4\] _0921_ _1125_ gpio_configure\[22\]\[12\] VGND VGND
+ VPWR VPWR _1126_ sky130_fd_sc_hd__a22o_1
XFILLER_143_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold846 gpio_configure\[6\]\[6\] VGND VGND VPWR VPWR net1379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 _0280_ VGND VGND VPWR VPWR net1390 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold868 mgmt_gpio_data_buf\[10\] VGND VGND VPWR VPWR net1401 sky130_fd_sc_hd__dlygate4sd3_1
X_6254_ gpio_configure\[22\]\[9\] _2824_ _2829_ gpio_configure\[33\]\[9\] _3066_ VGND
+ VGND VPWR VPWR _3067_ sky130_fd_sc_hd__a221o_1
X_3466_ net554 _0885_ VGND VGND VPWR VPWR _1057_ sky130_fd_sc_hd__nor2_4
XFILLER_130_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold879 _0723_ VGND VGND VPWR VPWR net1412 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5205_ _1136_ net427 VGND VGND VPWR VPWR _2394_ sky130_fd_sc_hd__and2_1
XFILLER_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3397_ gpio_configure\[34\]\[6\] _0874_ _0908_ gpio_configure\[2\]\[6\] VGND VGND
+ VPWR VPWR _0991_ sky130_fd_sc_hd__a22o_1
X_6185_ gpio_configure\[1\]\[6\] net401 _2823_ gpio_configure\[2\]\[6\] _3000_ VGND
+ VGND VPWR VPWR _3001_ sky130_fd_sc_hd__a221o_1
Xhold1502 _0767_ VGND VGND VPWR VPWR net2035 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1513 net349 VGND VGND VPWR VPWR net2046 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5136_ _2246_ _2343_ _1971_ VGND VGND VPWR VPWR _2344_ sky130_fd_sc_hd__or3b_1
Xhold1524 net347 VGND VGND VPWR VPWR net2057 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1535 serial_data_staging_2\[7\] VGND VGND VPWR VPWR net2068 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1546 net348 VGND VGND VPWR VPWR net2079 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1557 hkspi.ldata\[0\] VGND VGND VPWR VPWR net2090 sky130_fd_sc_hd__dlygate4sd3_1
X_5067_ _2262_ _2264_ _2275_ VGND VGND VPWR VPWR _2276_ sky130_fd_sc_hd__nor3_1
Xhold1568 mgmt_gpio_data_buf\[17\] VGND VGND VPWR VPWR net2101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1579 mgmt_gpio_data_buf\[16\] VGND VGND VPWR VPWR net2112 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4018_ net462 net1479 _1474_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__mux2_1
XFILLER_37_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_550 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5969_ xfer_state\[1\] serial_data_staging_1\[11\] _2791_ VGND VGND VPWR VPWR _2792_
+ sky130_fd_sc_hd__a21o_1
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold109 _0667_ VGND VGND VPWR VPWR net642 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3320_ _0870_ net381 VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__nor2_8
XFILLER_98_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ net474 net550 _0846_ VGND VGND VPWR VPWR _0847_ sky130_fd_sc_hd__o21ai_2
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6941_ clknet_leaf_29_csclk net983 net520 VGND VGND VPWR VPWR gpio_configure\[12\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_81_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6872_ clknet_leaf_40_csclk net757 net516 VGND VGND VPWR VPWR gpio_configure\[3\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_35_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5823_ gpio_configure\[15\]\[6\] _2510_ _2537_ gpio_configure\[17\]\[6\] VGND VGND
+ VPWR VPWR _2652_ sky130_fd_sc_hd__a22o_1
XFILLER_62_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5754_ gpio_configure\[7\]\[3\] _2528_ _2538_ gpio_configure\[1\]\[3\] VGND VGND
+ VPWR VPWR _2586_ sky130_fd_sc_hd__a22o_1
XFILLER_147_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4705_ _1787_ _1863_ _1915_ _1916_ VGND VGND VPWR VPWR _1917_ sky130_fd_sc_hd__o211a_1
XFILLER_148_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5685_ net472 _2459_ _2504_ VGND VGND VPWR VPWR _2520_ sky130_fd_sc_hd__and3_4
XFILLER_8_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4636_ _1788_ net432 _1836_ net424 VGND VGND VPWR VPWR _1848_ sky130_fd_sc_hd__o22a_1
XFILLER_175_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold610 _0642_ VGND VGND VPWR VPWR net1143 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold621 gpio_configure\[0\]\[5\] VGND VGND VPWR VPWR net1154 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4567_ _0834_ _1778_ VGND VGND VPWR VPWR _1779_ sky130_fd_sc_hd__or2_4
Xhold632 _0343_ VGND VGND VPWR VPWR net1165 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap351 _0933_ VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__buf_8
Xhold643 gpio_configure\[28\]\[4\] VGND VGND VPWR VPWR net1176 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6306_ gpio_configure\[16\]\[11\] _2831_ _2860_ gpio_configure\[17\]\[11\] _3116_
+ VGND VGND VPWR VPWR _3117_ sky130_fd_sc_hd__a221o_1
XFILLER_116_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold654 _0710_ VGND VGND VPWR VPWR net1187 sky130_fd_sc_hd__dlygate4sd3_1
Xhold665 gpio_configure\[26\]\[12\] VGND VGND VPWR VPWR net1198 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap373 _0916_ VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__buf_8
XFILLER_104_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3518_ net590 net629 VGND VGND VPWR VPWR _1109_ sky130_fd_sc_hd__nor2_4
Xmax_cap384 net385 VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__buf_12
Xhold676 _0545_ VGND VGND VPWR VPWR net1209 sky130_fd_sc_hd__dlygate4sd3_1
X_4498_ _1638_ _1640_ _1639_ net124 _1605_ VGND VGND VPWR VPWR _1710_ sky130_fd_sc_hd__a2111o_1
Xmax_cap395 _2829_ VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__buf_8
Xhold687 gpio_configure\[15\]\[12\] VGND VGND VPWR VPWR net1220 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold698 _0303_ VGND VGND VPWR VPWR net1231 sky130_fd_sc_hd__dlygate4sd3_1
X_6237_ gpio_configure\[13\]\[8\] _2804_ _2862_ gpio_configure\[25\]\[8\] VGND VGND
+ VPWR VPWR _3051_ sky130_fd_sc_hd__a22o_1
XFILLER_77_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3449_ _1040_ net2001 _0970_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__mux2_1
XFILLER_76_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_588 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ net362 _2975_ _2984_ VGND VGND VPWR VPWR _2985_ sky130_fd_sc_hd__or3_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1310 net1843 VGND VGND VPWR VPWR wb_dat_o[21] sky130_fd_sc_hd__buf_12
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1321 net1940 VGND VGND VPWR VPWR net1854 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1332 net1865 VGND VGND VPWR VPWR wb_dat_o[7] sky130_fd_sc_hd__buf_12
Xhold1343 net1957 VGND VGND VPWR VPWR net1876 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5119_ _1991_ _2192_ _2326_ VGND VGND VPWR VPWR _2327_ sky130_fd_sc_hd__nor3_1
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1354 net1887 VGND VGND VPWR VPWR wb_dat_o[26] sky130_fd_sc_hd__buf_12
X_6099_ gpio_configure\[33\]\[3\] net395 _2861_ gpio_configure\[28\]\[3\] _2917_ VGND
+ VGND VPWR VPWR _2918_ sky130_fd_sc_hd__a221o_1
XFILLER_84_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1365 net1962 VGND VGND VPWR VPWR net1898 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1376 net233 VGND VGND VPWR VPWR net1909 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1387 gpio_configure\[8\]\[6\] VGND VGND VPWR VPWR net1920 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1398 net331 VGND VGND VPWR VPWR net1931 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_3_0_wb_clk_i clknet_2_1_0_wb_clk_i VGND VGND VPWR VPWR clknet_3_3_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_53_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5470_ net810 net569 _2428_ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__mux2_1
XFILLER_157_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4421_ net126 _1619_ VGND VGND VPWR VPWR _1633_ sky130_fd_sc_hd__nor2_2
XFILLER_172_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7140_ clknet_leaf_36_csclk net1533 net523 VGND VGND VPWR VPWR gpio_configure\[37\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_172_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4352_ _1548_ _1563_ VGND VGND VPWR VPWR _1564_ sky130_fd_sc_hd__or2_2
XFILLER_98_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3303_ net1971 _0884_ VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__nand2_8
X_4283_ net466 net1711 _1539_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__mux2_1
X_7071_ clknet_leaf_45_csclk net1213 net526 VGND VGND VPWR VPWR gpio_configure\[28\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_98_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6022_ _2798_ _2811_ _2836_ _2839_ VGND VGND VPWR VPWR _2844_ sky130_fd_sc_hd__or4_1
XFILLER_39_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6924_ clknet_leaf_28_csclk net1587 net520 VGND VGND VPWR VPWR gpio_configure\[10\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_35_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6855_ clknet_leaf_36_csclk net1531 net522 VGND VGND VPWR VPWR gpio_configure\[1\]\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_5806_ gpio_configure\[3\]\[5\] _2518_ _2541_ gpio_configure\[31\]\[5\] _2635_ VGND
+ VGND VPWR VPWR _2636_ sky130_fd_sc_hd__a221o_1
XFILLER_50_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6786_ clknet_2_2__leaf_mgmt_gpio_in[4] net1996 _0060_ VGND VGND VPWR VPWR hkspi.ldata\[3\]
+ sky130_fd_sc_hd__dfrtn_1
X_3998_ net1928 net660 _1471_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__mux2_1
X_5737_ gpio_configure\[3\]\[2\] _2518_ _2569_ VGND VGND VPWR VPWR _2570_ sky130_fd_sc_hd__a21o_1
XFILLER_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5668_ gpio_configure\[13\]\[0\] _2501_ _2502_ gpio_configure\[4\]\[0\] _2500_ VGND
+ VGND VPWR VPWR _2503_ sky130_fd_sc_hd__a221o_1
XFILLER_135_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4619_ _1779_ _1807_ VGND VGND VPWR VPWR _1831_ sky130_fd_sc_hd__nor2_1
XFILLER_136_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5599_ _2448_ _2449_ _2450_ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__and3_1
XFILLER_151_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold440 _0688_ VGND VGND VPWR VPWR net973 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_151_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold451 net232 VGND VGND VPWR VPWR net984 sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 _0277_ VGND VGND VPWR VPWR net995 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold473 _0196_ VGND VGND VPWR VPWR net1006 sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 gpio_configure\[1\]\[12\] VGND VGND VPWR VPWR net1017 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_145_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold495 _0276_ VGND VGND VPWR VPWR net1028 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1140 _0225_ VGND VGND VPWR VPWR net1673 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1151 gpio_configure\[1\]\[9\] VGND VGND VPWR VPWR net1684 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1162 _0335_ VGND VGND VPWR VPWR net1695 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1173 net267 VGND VGND VPWR VPWR net1706 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1184 net1963 VGND VGND VPWR VPWR net1717 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1195 net1949 VGND VGND VPWR VPWR net1728 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_450 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4970_ _1598_ net380 _1691_ _1883_ VGND VGND VPWR VPWR _2180_ sky130_fd_sc_hd__a211o_1
XFILLER_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3921_ _0827_ net90 net76 VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__mux2_2
X_6640_ clknet_3_4_0_wb_clk_i _0253_ VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__dfxtp_1
X_3852_ _1417_ _1418_ _1416_ VGND VGND VPWR VPWR _1419_ sky130_fd_sc_hd__o21ba_1
XFILLER_149_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6571_ clknet_leaf_30_csclk net1374 net518 VGND VGND VPWR VPWR mgmt_gpio_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_3783_ gpio_configure\[0\]\[0\] _0898_ _1196_ trap_output_dest VGND VGND VPWR VPWR
+ _1369_ sky130_fd_sc_hd__a22o_1
XFILLER_192_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5522_ net464 net1395 _2434_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__mux2_1
XFILLER_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5453_ net447 net1304 _2426_ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__mux2_1
XFILLER_172_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4404_ _0817_ _1552_ _1614_ VGND VGND VPWR VPWR _1616_ sky130_fd_sc_hd__nand3_2
XFILLER_99_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5384_ net573 net716 _2418_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__mux2_1
XFILLER_132_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7123_ clknet_leaf_15_csclk net1189 net519 VGND VGND VPWR VPWR gpio_configure\[35\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_4335_ net443 net1063 _1547_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__mux2_1
XFILLER_59_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7054_ clknet_leaf_25_csclk net1235 net518 VGND VGND VPWR VPWR gpio_configure\[26\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_4266_ net938 net463 _1536_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__mux2_1
XFILLER_86_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_57_csclk clknet_3_2_0_csclk VGND VGND VPWR VPWR clknet_leaf_57_csclk
+ sky130_fd_sc_hd__clkbuf_16
X_6005_ gpio_configure\[23\]\[0\] _2822_ net398 gpio_configure\[2\]\[0\] _2826_ VGND
+ VGND VPWR VPWR _2827_ sky130_fd_sc_hd__a221o_1
X_3217_ gpio_configure\[17\]\[3\] VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__inv_2
XFILLER_67_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4197_ net2057 _0969_ _1520_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__mux2_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6907_ clknet_leaf_15_csclk net873 net513 VGND VGND VPWR VPWR gpio_configure\[8\]\[1\]
+ sky130_fd_sc_hd__dfstp_4
XFILLER_23_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6838_ clknet_leaf_40_csclk net686 net516 VGND VGND VPWR VPWR mgmt_gpio_data_buf\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6769_ clknet_leaf_60_csclk net769 net498 VGND VGND VPWR VPWR gpio_configure\[32\]\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_109_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold270 _0595_ VGND VGND VPWR VPWR net803 sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 net240 VGND VGND VPWR VPWR net814 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 _0626_ VGND VGND VPWR VPWR net825 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_110 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_121 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_132 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_143 net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_154 net359 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_165 net405 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_176 clknet_2_0__leaf_mgmt_gpio_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_187 net618 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_198 _1303_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4120_ net629 _0909_ net483 net546 VGND VGND VPWR VPWR _1510_ sky130_fd_sc_hd__or4_4
XFILLER_69_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4051_ net443 net1198 _1479_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__mux2_1
XFILLER_96_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput5 mask_rev_in[10] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4953_ _1596_ _1683_ _1675_ VGND VGND VPWR VPWR _2163_ sky130_fd_sc_hd__o21a_1
X_3904_ pad_count_2\[3\] pad_count_2\[2\] VGND VGND VPWR VPWR _1449_ sky130_fd_sc_hd__and2b_4
XFILLER_51_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4884_ _1642_ _1706_ _1749_ _1956_ VGND VGND VPWR VPWR _2095_ sky130_fd_sc_hd__o31a_1
X_6623_ clknet_leaf_10_csclk net807 net511 VGND VGND VPWR VPWR gpio_configure\[5\]\[10\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_138_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3835_ net2067 hkspi.pass_thru_user_delay _1408_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__mux2_1
XFILLER_192_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6554_ clknet_leaf_78_csclk net1710 net486 VGND VGND VPWR VPWR mgmt_gpio_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3766_ gpio_configure\[32\]\[0\] _0890_ _1083_ gpio_configure\[30\]\[8\] _1322_ VGND
+ VGND VPWR VPWR _1352_ sky130_fd_sc_hd__a221o_1
X_5505_ net457 net782 _2432_ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__mux2_1
XFILLER_192_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6485_ clknet_leaf_72_csclk net1125 net490 VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__dfstp_2
XFILLER_146_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3697_ net15 _0900_ _1196_ clk2_output_dest VGND VGND VPWR VPWR _1285_ sky130_fd_sc_hd__a22o_1
XFILLER_118_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5436_ net441 net1210 _2424_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__mux2_1
Xoutput320 net1874 VGND VGND VPWR VPWR net1875 sky130_fd_sc_hd__buf_12
XFILLER_160_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput331 net1842 VGND VGND VPWR VPWR net1843 sky130_fd_sc_hd__buf_12
Xoutput342 net1872 VGND VGND VPWR VPWR net1873 sky130_fd_sc_hd__buf_12
X_5367_ _0906_ net647 VGND VGND VPWR VPWR _2417_ sky130_fd_sc_hd__nand2_8
X_7106_ clknet_leaf_29_csclk net971 net525 VGND VGND VPWR VPWR gpio_configure\[33\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_4318_ net1973 net425 VGND VGND VPWR VPWR _1545_ sky130_fd_sc_hd__and2_2
XFILLER_59_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5298_ net458 net1588 _2409_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__mux2_1
XFILLER_87_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7037_ clknet_leaf_46_csclk net811 net515 VGND VGND VPWR VPWR gpio_configure\[24\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_4249_ net456 net1407 _1533_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__mux2_1
XFILLER_75_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3620_ gpio_configure\[14\]\[10\] _1069_ _1094_ gpio_configure\[7\]\[10\] _1193_
+ VGND VGND VPWR VPWR _1209_ sky130_fd_sc_hd__a221o_2
XFILLER_186_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3551_ gpio_configure\[24\]\[3\] _0919_ _1073_ gpio_configure\[24\]\[11\] VGND VGND
+ VPWR VPWR _1141_ sky130_fd_sc_hd__a22o_1
XFILLER_128_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6270_ net2108 net366 _3081_ _3082_ VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__o22a_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3482_ net384 _0909_ VGND VGND VPWR VPWR _1073_ sky130_fd_sc_hd__nor2_8
XFILLER_170_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5221_ net1499 _0974_ VGND VGND VPWR VPWR _2398_ sky130_fd_sc_hd__or2_1
XFILLER_88_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5152_ _1798_ _2233_ _2285_ _1850_ VGND VGND VPWR VPWR _2359_ sky130_fd_sc_hd__o22a_1
XFILLER_57_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4103_ net804 _1507_ _1499_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__mux2_1
XFILLER_110_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5083_ _1840_ _1892_ _2227_ _2291_ VGND VGND VPWR VPWR _2292_ sky130_fd_sc_hd__or4_1
XFILLER_56_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4034_ _1098_ net425 VGND VGND VPWR VPWR _1477_ sky130_fd_sc_hd__and2_2
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5985_ gpio_configure\[13\]\[0\] net417 net400 gpio_configure\[37\]\[0\] _2803_ VGND
+ VGND VPWR VPWR _2807_ sky130_fd_sc_hd__a221o_1
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4936_ _2145_ VGND VGND VPWR VPWR _2146_ sky130_fd_sc_hd__inv_2
XFILLER_33_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_10 _0919_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 _1004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4867_ _1677_ _1686_ _2041_ _2058_ _2077_ VGND VGND VPWR VPWR _2078_ sky130_fd_sc_hd__a2111o_1
XANTENNA_32 _1097_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_43 _1233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_54 _2433_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6606_ clknet_leaf_10_csclk net1701 net509 VGND VGND VPWR VPWR gpio_configure\[2\]\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_3818_ _0848_ _1397_ VGND VGND VPWR VPWR _1398_ sky130_fd_sc_hd__xnor2_1
XFILLER_192_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_65 _2518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_76 _2820_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4798_ net124 _1773_ _1792_ _1645_ _1744_ VGND VGND VPWR VPWR _2009_ sky130_fd_sc_hd__a32o_1
XANTENNA_87 gpio_configure\[18\]\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_98 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6537_ clknet_leaf_0_csclk net1620 net487 VGND VGND VPWR VPWR gpio_configure\[26\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_119_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3749_ _1328_ _1330_ _1332_ _1334_ VGND VGND VPWR VPWR _1335_ sky130_fd_sc_hd__or4_2
XFILLER_134_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6468_ clknet_2_2__leaf_mgmt_gpio_in[4] _0090_ _0046_ VGND VGND VPWR VPWR hkspi.addr\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_133_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5419_ net439 net802 _2422_ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__mux2_1
X_6399_ net486 net481 VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__and2_1
Xoutput172 net172 VGND VGND VPWR VPWR irq[0] sky130_fd_sc_hd__buf_12
XFILLER_161_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput183 net183 VGND VGND VPWR VPWR mgmt_gpio_oeb[17] sky130_fd_sc_hd__buf_12
Xoutput194 net194 VGND VGND VPWR VPWR mgmt_gpio_oeb[27] sky130_fd_sc_hd__buf_12
XFILLER_153_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5770_ _2596_ _2598_ _2599_ _2601_ VGND VGND VPWR VPWR _2602_ sky130_fd_sc_hd__or4_1
XFILLER_21_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4721_ _1590_ _1592_ _1779_ VGND VGND VPWR VPWR _1933_ sky130_fd_sc_hd__or3_2
X_4652_ _1678_ _1822_ VGND VGND VPWR VPWR _1864_ sky130_fd_sc_hd__or2_1
XFILLER_30_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput30 mask_rev_in[4] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
X_3603_ _1192_ net1995 _0970_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__mux2_1
Xinput41 mgmt_gpio_in[14] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput52 mgmt_gpio_in[24] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_1
X_4583_ net477 _1782_ VGND VGND VPWR VPWR _1795_ sky130_fd_sc_hd__or2_4
XFILLER_116_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput63 mgmt_gpio_in[34] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_8
Xhold803 gpio_configure\[29\]\[1\] VGND VGND VPWR VPWR net1336 sky130_fd_sc_hd__dlygate4sd3_1
Xinput74 pad_flash_io1_di VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold814 _0531_ VGND VGND VPWR VPWR net1347 sky130_fd_sc_hd__dlygate4sd3_1
X_6322_ gpio_configure\[20\]\[12\] _2828_ net393 gpio_configure\[34\]\[12\] _3131_
+ VGND VGND VPWR VPWR _3132_ sky130_fd_sc_hd__a221o_1
X_3534_ net386 _1006_ VGND VGND VPWR VPWR _1125_ sky130_fd_sc_hd__nor2_4
Xhold825 gpio_configure\[5\]\[6\] VGND VGND VPWR VPWR net1358 sky130_fd_sc_hd__dlygate4sd3_1
Xinput85 spimemio_flash_io0_do VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__buf_2
Xinput96 usr1_vdd_pwrgood VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__buf_2
Xhold836 gpio_configure\[15\]\[6\] VGND VGND VPWR VPWR net1369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 _0499_ VGND VGND VPWR VPWR net1380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold858 gpio_configure\[36\]\[6\] VGND VGND VPWR VPWR net1391 sky130_fd_sc_hd__dlygate4sd3_1
X_6253_ gpio_configure\[18\]\[9\] _2819_ _2837_ gpio_configure\[8\]\[9\] VGND VGND
+ VPWR VPWR _3066_ sky130_fd_sc_hd__a22o_1
Xhold869 _0439_ VGND VGND VPWR VPWR net1402 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3465_ net590 net382 VGND VGND VPWR VPWR _1056_ sky130_fd_sc_hd__nor2_4
XFILLER_170_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5204_ net469 net1927 _2393_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__mux2_1
XFILLER_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6184_ gpio_configure\[11\]\[6\] net415 net410 gpio_configure\[8\]\[6\] VGND VGND
+ VPWR VPWR _3000_ sky130_fd_sc_hd__a22o_1
X_3396_ gpio_configure\[11\]\[6\] _0907_ _0915_ gpio_configure\[3\]\[6\] _0989_ VGND
+ VGND VPWR VPWR _0990_ sky130_fd_sc_hd__a221o_1
XFILLER_97_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5135_ _1636_ _2203_ _1970_ _1672_ _1669_ VGND VGND VPWR VPWR _2343_ sky130_fd_sc_hd__o2111ai_1
Xhold1503 wbbd_data\[7\] VGND VGND VPWR VPWR net2036 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1514 hkspi.odata\[3\] VGND VGND VPWR VPWR net2047 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1525 wbbd_data\[2\] VGND VGND VPWR VPWR net2058 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1536 wbbd_addr\[1\] VGND VGND VPWR VPWR net2069 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1547 net319 VGND VGND VPWR VPWR net2080 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1558 serial_data_staging_2\[8\] VGND VGND VPWR VPWR net2091 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5066_ _2271_ _2273_ _2274_ VGND VGND VPWR VPWR _2275_ sky130_fd_sc_hd__or3_1
Xhold1569 hkspi.pre_pass_thru_mgmt VGND VGND VPWR VPWR net2102 sky130_fd_sc_hd__dlygate4sd3_1
X_4017_ net468 net1810 _1474_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__mux2_1
XFILLER_37_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_710 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5968_ gpio_configure\[0\]\[12\] _2526_ _2780_ _2790_ net473 VGND VGND VPWR VPWR
+ _2791_ sky130_fd_sc_hd__o221a_2
X_4919_ _1592_ _1791_ _1877_ VGND VGND VPWR VPWR _2130_ sky130_fd_sc_hd__o21ba_1
XFILLER_21_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5899_ gpio_configure\[8\]\[9\] _2520_ _2540_ gpio_configure\[12\]\[9\] VGND VGND
+ VPWR VPWR _2725_ sky130_fd_sc_hd__a22o_1
XFILLER_166_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ net2064 net474 VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__nand2b_1
XFILLER_112_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6940_ clknet_leaf_28_csclk net1579 net521 VGND VGND VPWR VPWR gpio_configure\[12\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_19_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6871_ clknet_leaf_37_csclk net1549 net522 VGND VGND VPWR VPWR gpio_configure\[3\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5822_ gpio_configure\[31\]\[6\] _2541_ _2650_ VGND VGND VPWR VPWR _2651_ sky130_fd_sc_hd__a21o_1
XFILLER_50_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5753_ net2037 _2585_ net366 VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__mux2_1
XFILLER_50_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4704_ _1787_ _1873_ VGND VGND VPWR VPWR _1916_ sky130_fd_sc_hd__or2_1
XFILLER_148_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5684_ gpio_configure\[30\]\[0\] _2517_ _2518_ gpio_configure\[3\]\[0\] VGND VGND
+ VPWR VPWR _2519_ sky130_fd_sc_hd__a22o_1
XFILLER_148_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4635_ _1788_ net432 VGND VGND VPWR VPWR _1847_ sky130_fd_sc_hd__nor2_1
XFILLER_118_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold600 _0682_ VGND VGND VPWR VPWR net1133 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4566_ net124 _1556_ VGND VGND VPWR VPWR _1778_ sky130_fd_sc_hd__or2_2
Xhold611 gpio_configure\[22\]\[1\] VGND VGND VPWR VPWR net1144 sky130_fd_sc_hd__dlygate4sd3_1
Xhold622 _0450_ VGND VGND VPWR VPWR net1155 sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 gpio_configure\[8\]\[4\] VGND VGND VPWR VPWR net1166 sky130_fd_sc_hd__dlygate4sd3_1
X_6305_ gpio_configure\[14\]\[11\] net411 _2855_ gpio_configure\[27\]\[11\] VGND VGND
+ VPWR VPWR _3116_ sky130_fd_sc_hd__a22o_1
Xmax_cap352 _0931_ VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__buf_8
Xhold644 _0673_ VGND VGND VPWR VPWR net1177 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap363 net364 VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__clkbuf_2
X_3517_ gpio_configure\[37\]\[4\] _0902_ _0907_ gpio_configure\[11\]\[4\] _1107_ VGND
+ VGND VPWR VPWR _1108_ sky130_fd_sc_hd__a221o_1
Xhold655 gpio_configure\[35\]\[4\] VGND VGND VPWR VPWR net1188 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap374 _0894_ VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__buf_6
XFILLER_1_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold666 _0162_ VGND VGND VPWR VPWR net1199 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4497_ _1581_ _1693_ VGND VGND VPWR VPWR _1709_ sky130_fd_sc_hd__or2_1
Xmax_cap385 net386 VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__buf_12
Xhold677 gpio_configure\[20\]\[5\] VGND VGND VPWR VPWR net1210 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap396 _2828_ VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__buf_8
Xhold688 _0313_ VGND VGND VPWR VPWR net1221 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6236_ gpio_configure\[10\]\[8\] net414 _2840_ gpio_configure\[6\]\[8\] _3049_ VGND
+ VGND VPWR VPWR _3050_ sky130_fd_sc_hd__a221o_1
Xhold699 net2124 VGND VGND VPWR VPWR net1232 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3448_ _1039_ hkspi.ldata\[4\] _0837_ VGND VGND VPWR VPWR _1040_ sky130_fd_sc_hd__mux2_1
XFILLER_89_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6167_ _2977_ _2979_ _2981_ _2983_ VGND VGND VPWR VPWR _2984_ sky130_fd_sc_hd__or4_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1300 _0104_ VGND VGND VPWR VPWR net1833 sky130_fd_sc_hd__dlygate4sd3_1
X_3379_ net383 _0973_ VGND VGND VPWR VPWR _0974_ sky130_fd_sc_hd__nor2_8
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1311 net1933 VGND VGND VPWR VPWR net1844 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1322 net1855 VGND VGND VPWR VPWR wb_dat_o[5] sky130_fd_sc_hd__buf_12
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ _1610_ _1690_ _1820_ _2040_ _2325_ VGND VGND VPWR VPWR _2326_ sky130_fd_sc_hd__a2111o_1
Xhold1333 net1945 VGND VGND VPWR VPWR net1866 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1344 net1877 VGND VGND VPWR VPWR wb_dat_o[3] sky130_fd_sc_hd__buf_12
X_6098_ gpio_configure\[14\]\[3\] net411 net408 gpio_configure\[35\]\[3\] VGND VGND
+ VPWR VPWR _2917_ sky130_fd_sc_hd__a22o_1
Xhold1355 net1961 VGND VGND VPWR VPWR net1888 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1366 net1899 VGND VGND VPWR VPWR wb_dat_o[25] sky130_fd_sc_hd__buf_12
Xhold1377 _0433_ VGND VGND VPWR VPWR net1910 sky130_fd_sc_hd__dlygate4sd3_1
X_5049_ _1735_ _1948_ _2088_ _2212_ VGND VGND VPWR VPWR _2258_ sky130_fd_sc_hd__or4_1
XTAP_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1388 gpio_configure\[7\]\[1\] VGND VGND VPWR VPWR net1921 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1399 gpio_configure\[11\]\[10\] VGND VGND VPWR VPWR net1932 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4420_ _0832_ net99 net124 VGND VGND VPWR VPWR _1632_ sky130_fd_sc_hd__or3_4
XFILLER_132_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4351_ _1561_ _1562_ VGND VGND VPWR VPWR _1563_ sky130_fd_sc_hd__nand2_1
XFILLER_125_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3302_ _0889_ net383 VGND VGND VPWR VPWR _0898_ sky130_fd_sc_hd__nor2_8
X_7070_ clknet_leaf_19_csclk net1177 net510 VGND VGND VPWR VPWR gpio_configure\[28\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_4282_ _1047_ net425 VGND VGND VPWR VPWR _1539_ sky130_fd_sc_hd__nand2_2
X_6021_ _2797_ _2805_ VGND VGND VPWR VPWR _2843_ sky130_fd_sc_hd__nor2_8
X_3233_ gpio_configure\[0\]\[3\] VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__inv_2
XFILLER_101_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_1_1_csclk clknet_1_1_0_csclk VGND VGND VPWR VPWR clknet_1_1_1_csclk sky130_fd_sc_hd__clkbuf_8
XFILLER_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6923_ clknet_leaf_48_csclk net1458 net514 VGND VGND VPWR VPWR gpio_configure\[10\]\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_35_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6854_ clknet_leaf_17_csclk net1265 net512 VGND VGND VPWR VPWR gpio_configure\[1\]\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_22_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5805_ gpio_configure\[22\]\[5\] _2498_ _2501_ gpio_configure\[13\]\[5\] VGND VGND
+ VPWR VPWR _2635_ sky130_fd_sc_hd__a22o_1
X_6785_ clknet_2_1__leaf_mgmt_gpio_in[4] net1998 _0059_ VGND VGND VPWR VPWR hkspi.ldata\[2\]
+ sky130_fd_sc_hd__dfrtn_1
X_3997_ net1049 net443 _1471_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__mux2_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5736_ gpio_configure\[11\]\[2\] _2505_ _2520_ gpio_configure\[8\]\[2\] VGND VGND
+ VPWR VPWR _2569_ sky130_fd_sc_hd__a22o_1
XFILLER_182_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5667_ net472 _2459_ _2488_ VGND VGND VPWR VPWR _2502_ sky130_fd_sc_hd__and3_4
XFILLER_136_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4618_ _1829_ _1826_ _1824_ _1827_ VGND VGND VPWR VPWR _1830_ sky130_fd_sc_hd__and4b_1
XFILLER_190_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5598_ xfer_count\[0\] _2446_ VGND VGND VPWR VPWR _2450_ sky130_fd_sc_hd__or2_1
XFILLER_190_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold430 _0616_ VGND VGND VPWR VPWR net963 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4549_ _1760_ VGND VGND VPWR VPWR _1761_ sky130_fd_sc_hd__inv_2
Xhold441 net2140 VGND VGND VPWR VPWR net974 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold452 _0432_ VGND VGND VPWR VPWR net985 sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 gpio_configure\[0\]\[12\] VGND VGND VPWR VPWR net996 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold474 gpio_configure\[27\]\[12\] VGND VGND VPWR VPWR net1007 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold485 _0218_ VGND VGND VPWR VPWR net1018 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold496 gpio_configure\[25\]\[11\] VGND VGND VPWR VPWR net1029 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6219_ serial_data_staging_2\[6\] _3033_ net473 VGND VGND VPWR VPWR _3034_ sky130_fd_sc_hd__mux2_1
XFILLER_104_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7199_ clknet_3_7_0_wb_clk_i _0801_ net529 VGND VGND VPWR VPWR wbbd_data\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_58_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1130 _0216_ VGND VGND VPWR VPWR net1663 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1141 gpio_configure\[24\]\[9\] VGND VGND VPWR VPWR net1674 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1152 _0215_ VGND VGND VPWR VPWR net1685 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1163 net274 VGND VGND VPWR VPWR net1696 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_161_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1174 _0397_ VGND VGND VPWR VPWR net1707 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1185 net283 VGND VGND VPWR VPWR net1718 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1196 gpio_configure\[21\]\[10\] VGND VGND VPWR VPWR net1729 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_721 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3920_ _0826_ net92 net76 VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__mux2_2
XFILLER_17_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3851_ hkspi.fixed\[2\] hkspi.fixed\[1\] _1384_ VGND VGND VPWR VPWR _1418_ sky130_fd_sc_hd__o21ai_1
XFILLER_177_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6570_ clknet_leaf_40_csclk net913 net516 VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__dfrtp_1
X_3782_ net282 _0886_ _1262_ net271 _1321_ VGND VGND VPWR VPWR _1368_ sky130_fd_sc_hd__a221o_1
X_5521_ net470 net1798 _2434_ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__mux2_1
XFILLER_8_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5452_ net452 net960 _2426_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__mux2_1
XFILLER_172_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4403_ _1552_ _1614_ _0817_ VGND VGND VPWR VPWR _1615_ sky130_fd_sc_hd__a21o_1
X_5383_ net437 net1417 _2418_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__mux2_1
X_7122_ clknet_leaf_29_csclk net977 net521 VGND VGND VPWR VPWR gpio_configure\[35\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_4334_ net449 net992 _1547_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__mux2_1
XFILLER_87_705 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7053_ clknet_leaf_30_csclk net1076 net520 VGND VGND VPWR VPWR gpio_configure\[26\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_4265_ net1818 net467 _1536_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__mux2_1
XFILLER_115_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6004_ gpio_configure\[22\]\[0\] _2824_ net414 gpio_configure\[10\]\[0\] VGND VGND
+ VPWR VPWR _2826_ sky130_fd_sc_hd__a22o_1
XFILLER_101_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3216_ gpio_configure\[18\]\[3\] VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__inv_2
X_4196_ net2075 _1004_ _1520_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__mux2_1
XFILLER_55_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6906_ clknet_leaf_15_csclk net1795 net513 VGND VGND VPWR VPWR gpio_configure\[8\]\[0\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_23_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6837_ clknet_leaf_40_csclk net731 net516 VGND VGND VPWR VPWR mgmt_gpio_data_buf\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_10_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6768_ clknet_leaf_71_csclk net1217 net490 VGND VGND VPWR VPWR gpio_configure\[32\]\[10\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_10_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5719_ _2546_ _2548_ _2550_ _2552_ VGND VGND VPWR VPWR _2553_ sky130_fd_sc_hd__or4_1
XFILLER_148_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6699_ clknet_3_7_0_wb_clk_i _0012_ net528 VGND VGND VPWR VPWR wbbd_state\[8\] sky130_fd_sc_hd__dfrtp_4
XFILLER_148_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold260 _0702_ VGND VGND VPWR VPWR net793 sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 mgmt_gpio_data\[15\] VGND VGND VPWR VPWR net804 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 _0189_ VGND VGND VPWR VPWR net815 sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 gpio_configure\[16\]\[9\] VGND VGND VPWR VPWR net826 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_93_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_100 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_111 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_122 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_133 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_144 net121 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_155 net360 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_166 net410 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_177 clknet_2_0__leaf_mgmt_gpio_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_188 net645 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_199 _1305_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4050_ net450 net1294 _1479_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__mux2_1
XFILLER_49_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput6 mask_rev_in[11] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
XFILLER_110_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4952_ _1594_ _1928_ _2161_ VGND VGND VPWR VPWR _2162_ sky130_fd_sc_hd__or3_1
X_3903_ pad_count_2\[0\] pad_count_2\[1\] VGND VGND VPWR VPWR _1448_ sky130_fd_sc_hd__and2b_4
X_4883_ _1642_ _1662_ _1706_ _1629_ VGND VGND VPWR VPWR _2094_ sky130_fd_sc_hd__o31a_1
XFILLER_177_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3834_ hkspi.state\[0\] _1384_ VGND VGND VPWR VPWR _1408_ sky130_fd_sc_hd__nand2_1
X_6622_ clknet_leaf_10_csclk net867 net511 VGND VGND VPWR VPWR gpio_configure\[5\]\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_177_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6553_ clknet_leaf_28_csclk net763 net520 VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__dfrtp_1
X_3765_ gpio_configure\[3\]\[8\] _1095_ _1346_ _1350_ _1063_ VGND VGND VPWR VPWR _1351_
+ sky130_fd_sc_hd__a2111o_1
XFILLER_158_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5504_ net464 net1184 _2432_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__mux2_1
X_6484_ clknet_leaf_72_csclk net1693 net490 VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__dfstp_2
X_3696_ net44 _0904_ net354 net72 _1283_ VGND VGND VPWR VPWR _1284_ sky130_fd_sc_hd__a221o_1
X_5435_ net446 net1182 _2424_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__mux2_1
Xoutput310 net310 VGND VGND VPWR VPWR serial_load sky130_fd_sc_hd__buf_12
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput321 net1860 VGND VGND VPWR VPWR net1861 sky130_fd_sc_hd__buf_12
XFILLER_133_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput332 net1838 VGND VGND VPWR VPWR net1839 sky130_fd_sc_hd__buf_12
XFILLER_126_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput343 net1876 VGND VGND VPWR VPWR net1877 sky130_fd_sc_hd__buf_12
X_5366_ net435 net1041 _2416_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__mux2_1
XFILLER_113_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4317_ net1021 net443 _1544_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__mux2_1
X_7105_ clknet_leaf_24_csclk net1681 net518 VGND VGND VPWR VPWR gpio_configure\[33\]\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_59_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5297_ net463 net884 _2409_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__mux2_1
XFILLER_59_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7036_ clknet_leaf_64_csclk net847 net501 VGND VGND VPWR VPWR gpio_configure\[24\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_4248_ net462 net1463 _1533_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__mux2_1
XFILLER_19_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4179_ net444 net894 _1518_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__mux2_1
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_41_csclk clknet_3_6_0_csclk VGND VGND VPWR VPWR clknet_leaf_41_csclk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_56_csclk clknet_3_2_0_csclk VGND VGND VPWR VPWR clknet_leaf_56_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_186_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3550_ gpio_configure\[28\]\[3\] _0888_ _0927_ gpio_configure\[25\]\[3\] VGND VGND
+ VPWR VPWR _1140_ sky130_fd_sc_hd__a22o_2
XFILLER_155_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3481_ net287 _0886_ _0910_ net295 VGND VGND VPWR VPWR _1072_ sky130_fd_sc_hd__a22o_2
X_5220_ net463 net888 _2397_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__mux2_1
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5151_ _2258_ _2340_ _2356_ _2357_ VGND VGND VPWR VPWR _2358_ sky130_fd_sc_hd__or4_1
XFILLER_96_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4102_ net614 net573 net354 VGND VGND VPWR VPWR _1507_ sky130_fd_sc_hd__mux2_1
XFILLER_57_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5082_ _1801_ _2285_ _1995_ VGND VGND VPWR VPWR _2291_ sky130_fd_sc_hd__o21bai_1
XFILLER_96_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4033_ net1254 net444 _1476_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__mux2_1
XFILLER_49_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5984_ _1447_ _2805_ VGND VGND VPWR VPWR _2806_ sky130_fd_sc_hd__nor2_4
XFILLER_52_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4935_ net128 _1566_ _2142_ VGND VGND VPWR VPWR _2145_ sky130_fd_sc_hd__or3_1
Xclkbuf_3_7_0_csclk clknet_2_3_0_csclk VGND VGND VPWR VPWR clknet_3_7_0_csclk sky130_fd_sc_hd__clkbuf_8
XANTENNA_11 _0920_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 _1004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4866_ _1673_ _2042_ _2054_ _2076_ VGND VGND VPWR VPWR _2077_ sky130_fd_sc_hd__or4_1
XANTENNA_33 _1115_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6605_ clknet_leaf_77_csclk net1018 net485 VGND VGND VPWR VPWR gpio_configure\[1\]\[12\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA_44 _1306_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_55 _2494_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3817_ hkspi.state\[3\] _1390_ hkspi.addr\[4\] VGND VGND VPWR VPWR _1397_ sky130_fd_sc_hd__o21a_1
XFILLER_165_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_66 _2518_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4797_ _1771_ _2007_ VGND VGND VPWR VPWR _2008_ sky130_fd_sc_hd__nand2_1
XFILLER_165_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_77 _2829_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_88 gpio_configure\[27\]\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6536_ clknet_leaf_0_csclk net1622 net487 VGND VGND VPWR VPWR gpio_configure\[26\]\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_3748_ gpio_configure\[34\]\[0\] net358 _1042_ gpio_configure\[6\]\[8\] _1333_ VGND
+ VGND VPWR VPWR _1334_ sky130_fd_sc_hd__a221o_1
XANTENNA_99 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3679_ _1259_ _1261_ _1264_ _1266_ VGND VGND VPWR VPWR _1267_ sky130_fd_sc_hd__or4_1
X_6467_ clknet_2_2__leaf_mgmt_gpio_in[4] _0089_ _0045_ VGND VGND VPWR VPWR hkspi.addr\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_106_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5418_ net441 net1146 _2422_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__mux2_1
X_6398_ net492 net482 VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__and2_1
XFILLER_0_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput173 net173 VGND VGND VPWR VPWR irq[1] sky130_fd_sc_hd__buf_12
XFILLER_0_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5349_ _0907_ net646 VGND VGND VPWR VPWR _2415_ sky130_fd_sc_hd__nand2_8
Xoutput184 net184 VGND VGND VPWR VPWR mgmt_gpio_oeb[18] sky130_fd_sc_hd__buf_12
Xoutput195 net195 VGND VGND VPWR VPWR mgmt_gpio_oeb[28] sky130_fd_sc_hd__buf_12
XFILLER_102_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7019_ clknet_leaf_28_csclk net1145 net519 VGND VGND VPWR VPWR gpio_configure\[22\]\[1\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4720_ _1928_ _1930_ _1931_ VGND VGND VPWR VPWR _1932_ sky130_fd_sc_hd__or3_1
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4651_ _1602_ _1684_ VGND VGND VPWR VPWR _1863_ sky130_fd_sc_hd__or2_4
XFILLER_174_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput20 mask_rev_in[24] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
X_3602_ _1191_ hkspi.ldata\[2\] _0837_ VGND VGND VPWR VPWR _1192_ sky130_fd_sc_hd__mux2_1
Xinput31 mask_rev_in[5] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_1
X_4582_ _1779_ _1793_ VGND VGND VPWR VPWR _1794_ sky130_fd_sc_hd__nor2_1
Xinput42 mgmt_gpio_in[15] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_4
XFILLER_174_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput53 mgmt_gpio_in[25] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_2
Xinput64 mgmt_gpio_in[35] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_2
Xinput75 porb VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_1
X_6321_ gpio_configure\[22\]\[12\] _2824_ _2852_ gpio_configure\[19\]\[12\] VGND VGND
+ VPWR VPWR _3131_ sky130_fd_sc_hd__a22o_1
X_3533_ gpio_configure\[20\]\[4\] _0928_ _0938_ gpio_configure\[33\]\[4\] _1123_ VGND
+ VGND VPWR VPWR _1124_ sky130_fd_sc_hd__a221o_1
Xhold804 _0678_ VGND VGND VPWR VPWR net1337 sky130_fd_sc_hd__dlygate4sd3_1
Xhold815 gpio_configure\[15\]\[2\] VGND VGND VPWR VPWR net1348 sky130_fd_sc_hd__dlygate4sd3_1
Xinput86 spimemio_flash_io0_oeb VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_4
Xhold826 _0491_ VGND VGND VPWR VPWR net1359 sky130_fd_sc_hd__dlygate4sd3_1
Xhold837 _0571_ VGND VGND VPWR VPWR net1370 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput97 usr2_vcc_pwrgood VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__buf_2
XFILLER_116_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold848 gpio_configure\[16\]\[1\] VGND VGND VPWR VPWR net1381 sky130_fd_sc_hd__dlygate4sd3_1
X_6252_ gpio_configure\[23\]\[9\] _2822_ _2828_ gpio_configure\[20\]\[9\] _3061_ VGND
+ VGND VPWR VPWR _3065_ sky130_fd_sc_hd__a221o_1
XFILLER_115_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold859 _0736_ VGND VGND VPWR VPWR net1392 sky130_fd_sc_hd__dlygate4sd3_1
X_3464_ gpio_configure\[20\]\[12\] _1053_ _1054_ gpio_configure\[19\]\[12\] VGND VGND
+ VPWR VPWR _1055_ sky130_fd_sc_hd__a22o_1
X_5203_ _1316_ net645 VGND VGND VPWR VPWR _2393_ sky130_fd_sc_hd__nand2_1
X_6183_ gpio_configure\[36\]\[6\] _2795_ _2798_ gpio_configure\[4\]\[6\] _2998_ VGND
+ VGND VPWR VPWR _2999_ sky130_fd_sc_hd__a221o_1
XFILLER_130_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3395_ gpio_configure\[15\]\[6\] _0918_ _0987_ _0988_ VGND VGND VPWR VPWR _0989_
+ sky130_fd_sc_hd__a211o_1
XFILLER_97_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5134_ _1954_ _2215_ _2254_ _2341_ VGND VGND VPWR VPWR _2342_ sky130_fd_sc_hd__or4_1
Xhold1504 serial_data_staging_1\[2\] VGND VGND VPWR VPWR net2037 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1515 irq_1_inputsrc VGND VGND VPWR VPWR net2048 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1526 wbbd_data\[1\] VGND VGND VPWR VPWR net2059 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1537 serial_data_staging_1\[12\] VGND VGND VPWR VPWR net2070 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5065_ _1698_ _1871_ _2051_ _2144_ VGND VGND VPWR VPWR _2274_ sky130_fd_sc_hd__or4_1
XFILLER_123_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1548 net317 VGND VGND VPWR VPWR net2081 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1559 hkspi.fixed\[1\] VGND VGND VPWR VPWR net2092 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4016_ _1083_ net426 VGND VGND VPWR VPWR _1474_ sky130_fd_sc_hd__nand2_2
XFILLER_38_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5967_ _2782_ _2785_ _2787_ _2789_ VGND VGND VPWR VPWR _2790_ sky130_fd_sc_hd__or4_1
X_4918_ _1588_ _1779_ _1593_ VGND VGND VPWR VPWR _2129_ sky130_fd_sc_hd__a21oi_2
XFILLER_33_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5898_ gpio_configure\[6\]\[9\] _2490_ _2523_ gpio_configure\[2\]\[9\] _2723_ VGND
+ VGND VPWR VPWR _2724_ sky130_fd_sc_hd__a221o_1
XFILLER_21_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4849_ _1665_ _1671_ _1902_ VGND VGND VPWR VPWR _2060_ sky130_fd_sc_hd__o21ai_1
XFILLER_193_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6519_ clknet_leaf_3_csclk net1287 net493 VGND VGND VPWR VPWR gpio_configure\[24\]\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_107_746 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6870_ clknet_leaf_16_csclk net1307 net512 VGND VGND VPWR VPWR gpio_configure\[3\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_5821_ gpio_configure\[20\]\[6\] _2499_ _2521_ gpio_configure\[21\]\[6\] VGND VGND
+ VPWR VPWR _2650_ sky130_fd_sc_hd__a22o_1
XFILLER_22_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5752_ net475 serial_data_staging_1\[1\] _2584_ VGND VGND VPWR VPWR _2585_ sky130_fd_sc_hd__a21o_1
X_4703_ _1833_ _1873_ _1913_ _1914_ VGND VGND VPWR VPWR _1915_ sky130_fd_sc_hd__o211a_1
XFILLER_175_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5683_ net472 _2461_ _2466_ VGND VGND VPWR VPWR _2518_ sky130_fd_sc_hd__and3_4
XFILLER_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4634_ _1839_ _1843_ _1844_ _1845_ VGND VGND VPWR VPWR _1846_ sky130_fd_sc_hd__nor4_1
XFILLER_163_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold601 gpio_configure\[15\]\[7\] VGND VGND VPWR VPWR net1134 sky130_fd_sc_hd__dlygate4sd3_1
X_4565_ net125 _1776_ VGND VGND VPWR VPWR _1777_ sky130_fd_sc_hd__or2_4
Xhold612 _0622_ VGND VGND VPWR VPWR net1145 sky130_fd_sc_hd__dlygate4sd3_1
Xhold623 gpio_configure\[23\]\[4\] VGND VGND VPWR VPWR net1156 sky130_fd_sc_hd__dlygate4sd3_1
X_6304_ gpio_configure\[22\]\[11\] _2824_ _2829_ gpio_configure\[33\]\[11\] _3114_
+ VGND VGND VPWR VPWR _3115_ sky130_fd_sc_hd__a221o_1
Xhold634 _0513_ VGND VGND VPWR VPWR net1167 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3516_ gpio_configure\[14\]\[4\] net373 _0918_ gpio_configure\[15\]\[4\] VGND VGND
+ VPWR VPWR _1107_ sky130_fd_sc_hd__a22o_1
Xhold645 gpio_configure\[7\]\[3\] VGND VGND VPWR VPWR net1178 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap353 _0929_ VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__buf_8
Xmax_cap364 net365 VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__clkbuf_2
X_4496_ _1576_ _1707_ VGND VGND VPWR VPWR _1708_ sky130_fd_sc_hd__or2_1
Xhold656 _0726_ VGND VGND VPWR VPWR net1189 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap375 _0883_ VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__buf_12
Xhold667 gpio_configure\[3\]\[3\] VGND VGND VPWR VPWR net1200 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmax_cap386 _0893_ VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__buf_12
Xhold678 _0610_ VGND VGND VPWR VPWR net1211 sky130_fd_sc_hd__dlygate4sd3_1
X_6235_ gpio_configure\[9\]\[8\] net412 _2838_ gpio_configure\[12\]\[8\] VGND VGND
+ VPWR VPWR _3049_ sky130_fd_sc_hd__a22o_1
Xmax_cap397 _2824_ VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__buf_8
XFILLER_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold689 gpio_configure\[10\]\[11\] VGND VGND VPWR VPWR net1222 sky130_fd_sc_hd__dlygate4sd3_1
X_3447_ _1023_ _1025_ _1027_ _1038_ VGND VGND VPWR VPWR _1039_ sky130_fd_sc_hd__or4_4
XFILLER_103_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3378_ net608 _0884_ VGND VGND VPWR VPWR _0973_ sky130_fd_sc_hd__nand2_8
XFILLER_134_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6166_ gpio_configure\[3\]\[5\] net413 net407 gpio_configure\[15\]\[5\] _2982_ VGND
+ VGND VPWR VPWR _2983_ sky130_fd_sc_hd__a221o_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1301 gpio_configure\[21\]\[8\] VGND VGND VPWR VPWR net1834 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1312 net1845 VGND VGND VPWR VPWR wb_dat_o[14] sky130_fd_sc_hd__buf_12
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1323 net1939 VGND VGND VPWR VPWR net1856 sky130_fd_sc_hd__dlygate4sd3_1
X_5117_ _1744_ _1994_ _2182_ VGND VGND VPWR VPWR _2325_ sky130_fd_sc_hd__a21o_1
X_6097_ net2027 _2916_ net366 VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__mux2_1
XFILLER_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1334 net1867 VGND VGND VPWR VPWR wb_dat_o[9] sky130_fd_sc_hd__buf_12
XFILLER_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1345 net1954 VGND VGND VPWR VPWR net1878 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1356 net1889 VGND VGND VPWR VPWR wb_dat_o[2] sky130_fd_sc_hd__buf_12
Xhold1367 net1969 VGND VGND VPWR VPWR net1900 sky130_fd_sc_hd__dlygate4sd3_1
X_5048_ _2254_ _2255_ _2256_ VGND VGND VPWR VPWR _2257_ sky130_fd_sc_hd__or3_1
Xhold1378 net236 VGND VGND VPWR VPWR net1911 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1389 gpio_configure\[4\]\[1\] VGND VGND VPWR VPWR net1922 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6999_ clknet_leaf_50_csclk net688 net507 VGND VGND VPWR VPWR gpio_configure\[19\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_159_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_101 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_624 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4350_ net111 _1559_ _1560_ VGND VGND VPWR VPWR _1562_ sky130_fd_sc_hd__nand3_1
XFILLER_125_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3301_ net581 net551 net638 VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__or3_4
XFILLER_98_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4281_ net447 net1162 _1538_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__mux2_1
XFILLER_99_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6020_ _2469_ _2473_ _2796_ VGND VGND VPWR VPWR _2842_ sky130_fd_sc_hd__and3_4
X_3232_ gpio_configure\[1\]\[3\] VGND VGND VPWR VPWR _0829_ sky130_fd_sc_hd__inv_2
XFILLER_140_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6922_ clknet_leaf_67_csclk net1645 net505 VGND VGND VPWR VPWR gpio_configure\[10\]\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_82_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6853_ clknet_leaf_30_csclk net1078 net518 VGND VGND VPWR VPWR gpio_configure\[1\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_50_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5804_ gpio_configure\[19\]\[5\] _2491_ _2629_ _2633_ VGND VGND VPWR VPWR _2634_
+ sky130_fd_sc_hd__a211o_1
X_6784_ clknet_2_0__leaf_mgmt_gpio_in[4] net2000 _0058_ VGND VGND VPWR VPWR hkspi.ldata\[1\]
+ sky130_fd_sc_hd__dfrtn_1
X_3996_ net1059 net449 _1471_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__mux2_1
XFILLER_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5735_ gpio_configure\[5\]\[2\] net422 _2501_ gpio_configure\[13\]\[2\] _2567_ VGND
+ VGND VPWR VPWR _2568_ sky130_fd_sc_hd__a221o_1
XFILLER_148_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5666_ net472 _2493_ _2495_ VGND VGND VPWR VPWR _2501_ sky130_fd_sc_hd__and3_4
XFILLER_108_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4617_ _0832_ _0833_ net124 _1792_ _1828_ VGND VGND VPWR VPWR _1829_ sky130_fd_sc_hd__a41o_1
XFILLER_163_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5597_ xfer_count\[0\] _2446_ VGND VGND VPWR VPWR _2449_ sky130_fd_sc_hd__nand2_1
Xhold420 _0690_ VGND VGND VPWR VPWR net953 sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 net244 VGND VGND VPWR VPWR net964 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_163_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4548_ _1753_ _1759_ wbbd_state\[8\] VGND VGND VPWR VPWR _1760_ sky130_fd_sc_hd__o21ai_2
XFILLER_89_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold442 _0442_ VGND VGND VPWR VPWR net975 sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 gpio_configure\[32\]\[12\] VGND VGND VPWR VPWR net986 sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 _0213_ VGND VGND VPWR VPWR net997 sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 _0813_ VGND VGND VPWR VPWR net1008 sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 net278 VGND VGND VPWR VPWR net1019 sky130_fd_sc_hd__dlygate4sd3_1
X_4479_ _1581_ _1689_ VGND VGND VPWR VPWR _1691_ sky130_fd_sc_hd__nor2_4
Xhold497 _0151_ VGND VGND VPWR VPWR net1030 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6218_ _3016_ _3022_ _3032_ _2851_ gpio_configure\[0\]\[7\] VGND VGND VPWR VPWR _3033_
+ sky130_fd_sc_hd__o32a_1
X_7198_ clknet_3_7_0_wb_clk_i _0800_ net528 VGND VGND VPWR VPWR wbbd_data\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1120 _0732_ VGND VGND VPWR VPWR net1653 sky130_fd_sc_hd__dlygate4sd3_1
X_6149_ gpio_configure\[30\]\[5\] _2799_ net408 gpio_configure\[35\]\[5\] VGND VGND
+ VPWR VPWR _2966_ sky130_fd_sc_hd__a22o_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1131 gpio_configure\[20\]\[2\] VGND VGND VPWR VPWR net1664 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1142 _0139_ VGND VGND VPWR VPWR net1675 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1153 gpio_configure\[26\]\[2\] VGND VGND VPWR VPWR net1686 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1164 _0403_ VGND VGND VPWR VPWR net1697 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1175 net1989 VGND VGND VPWR VPWR net1708 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1186 _0097_ VGND VGND VPWR VPWR net1719 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1197 mgmt_gpio_data\[33\] VGND VGND VPWR VPWR net1730 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_733 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3850_ hkspi.state\[3\] _0821_ hkspi.state\[0\] VGND VGND VPWR VPWR _1417_ sky130_fd_sc_hd__or3_4
X_3781_ _1360_ _1362_ _1364_ _1366_ VGND VGND VPWR VPWR _1367_ sky130_fd_sc_hd__or4_1
X_5520_ _0892_ net647 VGND VGND VPWR VPWR _2434_ sky130_fd_sc_hd__nand2_8
XFILLER_157_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5451_ net457 net820 _2426_ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__mux2_1
XFILLER_145_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4402_ net128 _1554_ _1610_ VGND VGND VPWR VPWR _1614_ sky130_fd_sc_hd__and3_1
X_5382_ net440 net1538 _2418_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__mux2_1
XFILLER_132_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7121_ clknet_leaf_28_csclk net1581 net520 VGND VGND VPWR VPWR gpio_configure\[35\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_4333_ net455 net1702 _1547_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__mux2_1
XFILLER_5_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4264_ _1065_ net427 VGND VGND VPWR VPWR _1536_ sky130_fd_sc_hd__and2_2
XFILLER_101_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7052_ clknet_leaf_30_csclk net1687 net526 VGND VGND VPWR VPWR gpio_configure\[26\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_115_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6003_ _1448_ _2796_ _2809_ VGND VGND VPWR VPWR _2825_ sky130_fd_sc_hd__and3_4
X_3215_ gpio_configure\[19\]\[3\] VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__inv_2
XFILLER_140_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4195_ net2031 _1039_ _1520_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__mux2_1
XFILLER_95_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6905_ clknet_leaf_39_csclk net1070 net516 VGND VGND VPWR VPWR gpio_configure\[7\]\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_23_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6836_ clknet_leaf_40_csclk net1402 net516 VGND VGND VPWR VPWR mgmt_gpio_data_buf\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_23_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6767_ clknet_leaf_61_csclk net835 net498 VGND VGND VPWR VPWR gpio_configure\[32\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_3979_ net534 net632 net1993 VGND VGND VPWR VPWR _1468_ sky130_fd_sc_hd__mux2_2
XFILLER_183_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5718_ gpio_configure\[15\]\[1\] _2510_ _2512_ gpio_configure\[9\]\[1\] _2551_ VGND
+ VGND VPWR VPWR _2552_ sky130_fd_sc_hd__a221o_1
XFILLER_148_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6698_ clknet_3_7_0_wb_clk_i _0011_ net528 VGND VGND VPWR VPWR wbbd_state\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_40_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5649_ xfer_count\[1\] _2484_ _2483_ net2074 VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_164_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold250 _0671_ VGND VGND VPWR VPWR net783 sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 gpio_configure\[32\]\[5\] VGND VGND VPWR VPWR net794 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold272 _0186_ VGND VGND VPWR VPWR net805 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 serial_bb_resetn VGND VGND VPWR VPWR net816 sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 _0315_ VGND VGND VPWR VPWR net827 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_135 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_101 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_112 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_123 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_134 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_145 net169 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_156 net371 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_167 net423 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_178 clknet_2_0__leaf_mgmt_gpio_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_189 net1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_csclk clknet_0_csclk VGND VGND VPWR VPWR clknet_1_1_0_csclk sky130_fd_sc_hd__clkbuf_8
XFILLER_167_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput7 mask_rev_in[12] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_37_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4951_ net121 _1587_ _1686_ VGND VGND VPWR VPWR _2161_ sky130_fd_sc_hd__and3_1
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3902_ pad_count_2\[4\] pad_count_2\[5\] VGND VGND VPWR VPWR _1447_ sky130_fd_sc_hd__nand2b_4
XFILLER_44_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4882_ _1709_ _1898_ VGND VGND VPWR VPWR _2093_ sky130_fd_sc_hd__nand2_1
XFILLER_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6621_ clknet_leaf_10_csclk net1788 net511 VGND VGND VPWR VPWR gpio_configure\[5\]\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_3833_ _1407_ net2137 _1388_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__mux2_1
XFILLER_32_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6552_ clknet_leaf_27_csclk net955 net520 VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__dfrtp_1
X_3764_ net291 _1299_ _1347_ _1349_ VGND VGND VPWR VPWR _1350_ sky130_fd_sc_hd__a211o_1
X_5503_ net470 net1791 _2432_ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__mux2_1
XFILLER_173_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6483_ clknet_leaf_72_csclk net1716 net490 VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__dfstp_1
X_3695_ gpio_configure\[11\]\[1\] _0907_ _1136_ net302 VGND VGND VPWR VPWR _1283_
+ sky130_fd_sc_hd__a22o_1
XFILLER_173_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput300 net300 VGND VGND VPWR VPWR pll_trim[9] sky130_fd_sc_hd__buf_12
X_5434_ net452 net1089 _2424_ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__mux2_1
XFILLER_160_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput311 net311 VGND VGND VPWR VPWR serial_resetn sky130_fd_sc_hd__buf_12
Xoutput322 net1862 VGND VGND VPWR VPWR net1863 sky130_fd_sc_hd__buf_12
Xoutput333 net1852 VGND VGND VPWR VPWR net1853 sky130_fd_sc_hd__buf_12
XFILLER_133_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput344 net1884 VGND VGND VPWR VPWR net1885 sky130_fd_sc_hd__buf_12
X_5365_ net439 net796 _2416_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__mux2_1
XFILLER_126_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_3_0_csclk clknet_2_1_0_csclk VGND VGND VPWR VPWR clknet_3_3_0_csclk sky130_fd_sc_hd__clkbuf_8
X_7104_ clknet_leaf_26_csclk net1414 net519 VGND VGND VPWR VPWR gpio_configure\[33\]\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_4316_ net1035 net449 _1544_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__mux2_1
XFILLER_59_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5296_ net471 net1775 _2409_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__mux2_1
XFILLER_113_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7035_ clknet_leaf_60_csclk net893 net498 VGND VGND VPWR VPWR gpio_configure\[24\]\[1\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_59_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4247_ net468 net1806 _1533_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__mux2_1
XFILLER_75_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4178_ net450 net1226 _1518_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__mux2_1
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_0_0_wb_clk_i clknet_1_0_1_wb_clk_i VGND VGND VPWR VPWR clknet_2_0_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_70_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6819_ clknet_leaf_61_csclk net1501 net498 VGND VGND VPWR VPWR serial_xfer sky130_fd_sc_hd__dfrtp_1
XFILLER_11_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3480_ gpio_configure\[18\]\[4\] _0894_ _1067_ gpio_configure\[23\]\[12\] _1070_
+ VGND VGND VPWR VPWR _1071_ sky130_fd_sc_hd__a221o_1
XFILLER_155_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5150_ _1629_ _2244_ _2245_ _1956_ _2248_ VGND VGND VPWR VPWR _2357_ sky130_fd_sc_hd__a221o_1
XFILLER_170_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4101_ net882 _1506_ _1499_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__mux2_1
XFILLER_69_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5081_ _1836_ _2233_ _2289_ VGND VGND VPWR VPWR _2290_ sky130_fd_sc_hd__o21ai_1
XFILLER_2_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4032_ net1276 net450 _1476_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__mux2_1
XFILLER_96_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_764 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5983_ _1449_ _2471_ VGND VGND VPWR VPWR _2805_ sky130_fd_sc_hd__nand2_4
XFILLER_18_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4934_ _1574_ _2143_ _2053_ VGND VGND VPWR VPWR _2144_ sky130_fd_sc_hd__a21o_1
XFILLER_178_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4865_ _2052_ _2059_ _2060_ _2075_ VGND VGND VPWR VPWR _2076_ sky130_fd_sc_hd__or4_1
XFILLER_20_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_12 _0921_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 _1004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_193_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6604_ clknet_leaf_77_csclk net1080 net484 VGND VGND VPWR VPWR gpio_configure\[1\]\[11\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA_34 _1118_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3816_ hkspi.state\[3\] _1390_ VGND VGND VPWR VPWR _1396_ sky130_fd_sc_hd__nor2_1
XANTENNA_45 _1337_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_192_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_56 _2494_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4796_ net424 _1777_ _2006_ _1744_ VGND VGND VPWR VPWR _2007_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_20_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_67 _2520_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_78 _2861_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_165_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6535_ clknet_leaf_6_csclk net1205 net497 VGND VGND VPWR VPWR gpio_configure\[28\]\[12\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_89 gpio_configure\[30\]\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3747_ gpio_configure\[15\]\[0\] _0918_ _1068_ gpio_configure\[10\]\[8\] VGND VGND
+ VPWR VPWR _1333_ sky130_fd_sc_hd__a22o_1
X_6466_ clknet_2_2__leaf_mgmt_gpio_in[4] _0088_ _0044_ VGND VGND VPWR VPWR hkspi.addr\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_3678_ net35 _0891_ _1057_ gpio_configure\[9\]\[9\] _1265_ VGND VGND VPWR VPWR _1266_
+ sky130_fd_sc_hd__a221o_1
XFILLER_118_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5417_ net447 net1268 _2422_ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__mux2_1
XFILLER_161_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6397_ net443 net1007 _3182_ VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__mux2_1
Xoutput174 net174 VGND VGND VPWR VPWR irq[2] sky130_fd_sc_hd__buf_12
X_5348_ net435 net1053 _2414_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__mux2_1
Xoutput185 net185 VGND VGND VPWR VPWR mgmt_gpio_oeb[19] sky130_fd_sc_hd__buf_12
Xoutput196 net196 VGND VGND VPWR VPWR mgmt_gpio_oeb[29] sky130_fd_sc_hd__buf_12
XFILLER_102_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5279_ net465 net858 _2407_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__mux2_1
XFILLER_75_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7018_ clknet_3_1_0_csclk net1793 net505 VGND VGND VPWR VPWR gpio_configure\[22\]\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_102_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_664 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4650_ _1861_ VGND VGND VPWR VPWR _1862_ sky130_fd_sc_hd__inv_2
Xinput10 mask_rev_in[15] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
X_3601_ _1173_ _1178_ _1183_ _1190_ VGND VGND VPWR VPWR _1191_ sky130_fd_sc_hd__or4_4
XFILLER_147_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput21 mask_rev_in[25] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_1
XFILLER_175_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput32 mask_rev_in[6] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_1
X_4581_ net477 _1790_ VGND VGND VPWR VPWR _1793_ sky130_fd_sc_hd__or2_4
Xinput43 mgmt_gpio_in[16] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_1
Xinput54 mgmt_gpio_in[26] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_2
X_6320_ gpio_configure\[36\]\[12\] net403 net402 gpio_configure\[4\]\[12\] VGND VGND
+ VPWR VPWR _3130_ sky130_fd_sc_hd__a22o_1
Xhold805 gpio_configure\[33\]\[9\] VGND VGND VPWR VPWR net1338 sky130_fd_sc_hd__dlygate4sd3_1
X_3532_ gpio_configure\[17\]\[12\] _1121_ _1122_ gpio_configure\[8\]\[12\] VGND VGND
+ VPWR VPWR _1123_ sky130_fd_sc_hd__a22o_1
Xinput65 mgmt_gpio_in[36] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_4
Xinput76 qspi_enabled VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_6
Xhold816 _0567_ VGND VGND VPWR VPWR net1349 sky130_fd_sc_hd__dlygate4sd3_1
Xinput87 spimemio_flash_io1_do VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__clkbuf_4
Xinput98 usr2_vdd_pwrgood VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_4
Xhold827 gpio_configure\[7\]\[10\] VGND VGND VPWR VPWR net1360 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold838 gpio_configure\[13\]\[1\] VGND VGND VPWR VPWR net1371 sky130_fd_sc_hd__dlygate4sd3_1
X_6251_ gpio_configure\[29\]\[9\] _2816_ _2820_ gpio_configure\[21\]\[9\] _3063_ VGND
+ VGND VPWR VPWR _3064_ sky130_fd_sc_hd__a221o_1
Xhold849 _0574_ VGND VGND VPWR VPWR net1382 sky130_fd_sc_hd__dlygate4sd3_1
X_3463_ net384 _0973_ VGND VGND VPWR VPWR _1054_ sky130_fd_sc_hd__nor2_8
XFILLER_115_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5202_ net463 net854 _2392_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__mux2_1
X_6182_ gpio_configure\[31\]\[6\] net423 net392 gpio_configure\[5\]\[6\] _2997_ VGND
+ VGND VPWR VPWR _2998_ sky130_fd_sc_hd__a221o_1
XFILLER_170_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3394_ net32 _0900_ _0919_ gpio_configure\[24\]\[6\] _0976_ VGND VGND VPWR VPWR _0988_
+ sky130_fd_sc_hd__a221o_1
XFILLER_97_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5133_ _1596_ _1686_ _1882_ _2085_ VGND VGND VPWR VPWR _2341_ sky130_fd_sc_hd__a211o_1
XFILLER_69_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1505 _0766_ VGND VGND VPWR VPWR net2038 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1516 serial_data_staging_1\[5\] VGND VGND VPWR VPWR net2049 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1527 serial_data_staging_2\[1\] VGND VGND VPWR VPWR net2060 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1538 wbbd_write VGND VGND VPWR VPWR net2071 sky130_fd_sc_hd__dlygate4sd3_1
X_5064_ _2037_ _2038_ _2157_ _2272_ VGND VGND VPWR VPWR _2273_ sky130_fd_sc_hd__or4_1
Xhold1549 serial_data_staging_1\[11\] VGND VGND VPWR VPWR net2082 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4015_ net902 net444 _1473_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__mux2_1
XFILLER_72_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5966_ gpio_configure\[5\]\[12\] _2496_ net418 gpio_configure\[24\]\[12\] _2788_
+ VGND VGND VPWR VPWR _2789_ sky130_fd_sc_hd__a221o_1
X_4917_ _1678_ _1788_ _1832_ VGND VGND VPWR VPWR _2128_ sky130_fd_sc_hd__o21bai_1
X_5897_ gpio_configure\[19\]\[9\] _2491_ _2505_ gpio_configure\[11\]\[9\] VGND VGND
+ VPWR VPWR _2723_ sky130_fd_sc_hd__a22o_1
XFILLER_32_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4848_ _1678_ _1798_ _1735_ VGND VGND VPWR VPWR _2059_ sky130_fd_sc_hd__o21bai_1
XFILLER_20_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4779_ _1609_ _1880_ _1772_ VGND VGND VPWR VPWR _1990_ sky130_fd_sc_hd__a21oi_1
XFILLER_181_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6518_ clknet_leaf_78_csclk net1637 net487 VGND VGND VPWR VPWR gpio_configure\[24\]\[10\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_134_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6449_ clknet_2_3__leaf_mgmt_gpio_in[4] _0071_ _0027_ VGND VGND VPWR VPWR hkspi.odata\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_40_csclk clknet_3_6_0_csclk VGND VGND VPWR VPWR clknet_leaf_40_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_164_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_2_0_0_csclk clknet_1_0_1_csclk VGND VGND VPWR VPWR clknet_2_0_0_csclk sky130_fd_sc_hd__clkbuf_8
XFILLER_87_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_55_csclk clknet_3_3_0_csclk VGND VGND VPWR VPWR clknet_leaf_55_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_189_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5820_ gpio_configure\[2\]\[6\] _2523_ _2529_ gpio_configure\[29\]\[6\] _2648_ VGND
+ VGND VPWR VPWR _2649_ sky130_fd_sc_hd__a221o_1
XFILLER_34_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5751_ gpio_configure\[0\]\[2\] _2526_ _2573_ _2583_ _0824_ VGND VGND VPWR VPWR _2584_
+ sky130_fd_sc_hd__o221a_1
XFILLER_15_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4702_ _1787_ _1874_ _1886_ _1833_ VGND VGND VPWR VPWR _1914_ sky130_fd_sc_hd__o22a_1
X_5682_ pad_count_1\[4\] _2489_ _2493_ VGND VGND VPWR VPWR _2517_ sky130_fd_sc_hd__and3_4
XFILLER_30_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4633_ _1692_ _1791_ VGND VGND VPWR VPWR _1845_ sky130_fd_sc_hd__nor2_1
XFILLER_147_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4564_ net127 net128 net126 VGND VGND VPWR VPWR _1776_ sky130_fd_sc_hd__nand3b_4
Xhold602 _0572_ VGND VGND VPWR VPWR net1135 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold613 gpio_configure\[18\]\[5\] VGND VGND VPWR VPWR net1146 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6303_ gpio_configure\[18\]\[11\] _2819_ _2837_ gpio_configure\[8\]\[11\] VGND VGND
+ VPWR VPWR _3114_ sky130_fd_sc_hd__a22o_1
Xhold624 _0633_ VGND VGND VPWR VPWR net1157 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3515_ _1092_ _1097_ _1100_ _1105_ VGND VGND VPWR VPWR _1106_ sky130_fd_sc_hd__or4_1
Xhold635 gpio_configure\[11\]\[12\] VGND VGND VPWR VPWR net1168 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap354 _0929_ VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__buf_8
X_4495_ net530 _1584_ VGND VGND VPWR VPWR _1707_ sky130_fd_sc_hd__nand2_4
Xhold646 _0504_ VGND VGND VPWR VPWR net1179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 gpio_configure\[13\]\[4\] VGND VGND VPWR VPWR net1190 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap376 net554 VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__buf_12
Xhold668 _0472_ VGND VGND VPWR VPWR net1201 sky130_fd_sc_hd__dlygate4sd3_1
X_6234_ gpio_configure\[34\]\[8\] net393 _2852_ gpio_configure\[19\]\[8\] _3047_ VGND
+ VGND VPWR VPWR _3048_ sky130_fd_sc_hd__a221o_1
Xmax_cap387 net388 VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__buf_12
Xhold679 gpio_configure\[28\]\[5\] VGND VGND VPWR VPWR net1212 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap398 _2823_ VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__buf_12
X_3446_ _1029_ _1030_ _1032_ _1037_ VGND VGND VPWR VPWR _1038_ sky130_fd_sc_hd__or4_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6165_ gpio_configure\[26\]\[5\] _2810_ _2811_ gpio_configure\[7\]\[5\] VGND VGND
+ VPWR VPWR _2982_ sky130_fd_sc_hd__a22o_1
X_3377_ net390 _0873_ VGND VGND VPWR VPWR _0972_ sky130_fd_sc_hd__nor2_8
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1302 _0364_ VGND VGND VPWR VPWR net1835 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1313 net1935 VGND VGND VPWR VPWR net1846 sky130_fd_sc_hd__dlygate4sd3_1
X_5116_ _1666_ _1941_ _2197_ _2300_ _2323_ VGND VGND VPWR VPWR _2324_ sky130_fd_sc_hd__a2111o_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6096_ net475 serial_data_staging_2\[1\] _2915_ VGND VGND VPWR VPWR _2916_ sky130_fd_sc_hd__a21o_1
Xhold1324 net1857 VGND VGND VPWR VPWR wb_dat_o[10] sky130_fd_sc_hd__buf_12
Xhold1335 net1946 VGND VGND VPWR VPWR net1868 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1346 net1879 VGND VGND VPWR VPWR wb_dat_o[0] sky130_fd_sc_hd__buf_12
XFILLER_27_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1357 net1960 VGND VGND VPWR VPWR net1890 sky130_fd_sc_hd__dlygate4sd3_1
X_5047_ _1735_ _1948_ _2088_ _2212_ VGND VGND VPWR VPWR _2256_ sky130_fd_sc_hd__or4_1
Xhold1368 net1901 VGND VGND VPWR VPWR wb_dat_o[24] sky130_fd_sc_hd__buf_12
XFILLER_26_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1379 hkspi.odata\[1\] VGND VGND VPWR VPWR net1912 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6998_ clknet_leaf_60_csclk net721 net498 VGND VGND VPWR VPWR gpio_configure\[19\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_41_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5949_ gpio_configure\[28\]\[12\] _2513_ _2521_ gpio_configure\[21\]\[12\] VGND VGND
+ VPWR VPWR _2772_ sky130_fd_sc_hd__a22o_1
XFILLER_185_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_159_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_558 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3300_ _0893_ _0895_ VGND VGND VPWR VPWR _0896_ sky130_fd_sc_hd__nor2_8
XFILLER_4_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4280_ net569 net718 _1538_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__mux2_1
XFILLER_98_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3231_ gpio_configure\[2\]\[3\] VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__inv_2
XFILLER_101_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6921_ clknet_leaf_41_csclk net1040 net517 VGND VGND VPWR VPWR gpio_configure\[9\]\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6852_ clknet_leaf_24_csclk net1661 net518 VGND VGND VPWR VPWR gpio_configure\[1\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_90_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5803_ gpio_configure\[18\]\[5\] _2532_ _2630_ _2632_ VGND VGND VPWR VPWR _2633_
+ sky130_fd_sc_hd__a211o_1
XFILLER_22_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6783_ clknet_2_0__leaf_mgmt_gpio_in[4] _0386_ _0057_ VGND VGND VPWR VPWR hkspi.ldata\[0\]
+ sky130_fd_sc_hd__dfrtn_1
X_3995_ net1708 net455 _1471_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__mux2_1
XFILLER_22_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5734_ gpio_configure\[27\]\[2\] _2506_ _2523_ gpio_configure\[2\]\[2\] VGND VGND
+ VPWR VPWR _2567_ sky130_fd_sc_hd__a22o_1
XFILLER_50_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5665_ gpio_configure\[22\]\[0\] _2498_ _2499_ gpio_configure\[20\]\[0\] VGND VGND
+ VPWR VPWR _2500_ sky130_fd_sc_hd__a22o_1
XFILLER_129_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4616_ _1778_ _1801_ VGND VGND VPWR VPWR _1828_ sky130_fd_sc_hd__nor2_1
XFILLER_190_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5596_ xfer_state\[3\] _1446_ _2443_ VGND VGND VPWR VPWR _2448_ sky130_fd_sc_hd__or3_1
XFILLER_135_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold410 _0177_ VGND VGND VPWR VPWR net943 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_191_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4547_ _1548_ _1758_ VGND VGND VPWR VPWR _1759_ sky130_fd_sc_hd__or2_2
Xhold421 net227 VGND VGND VPWR VPWR net954 sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 _0174_ VGND VGND VPWR VPWR net965 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold443 gpio_configure\[35\]\[3\] VGND VGND VPWR VPWR net976 sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 _0373_ VGND VGND VPWR VPWR net987 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold465 gpio_configure\[5\]\[3\] VGND VGND VPWR VPWR net998 sky130_fd_sc_hd__dlygate4sd3_1
X_4478_ _1689_ VGND VGND VPWR VPWR _1690_ sky130_fd_sc_hd__inv_2
XFILLER_171_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold476 gpio_configure\[28\]\[3\] VGND VGND VPWR VPWR net1009 sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 _0108_ VGND VGND VPWR VPWR net1020 sky130_fd_sc_hd__dlygate4sd3_1
Xhold498 gpio_configure\[0\]\[11\] VGND VGND VPWR VPWR net1031 sky130_fd_sc_hd__dlygate4sd3_1
X_6217_ net361 _3024_ _3026_ _3031_ VGND VGND VPWR VPWR _3032_ sky130_fd_sc_hd__or4_1
X_3429_ gpio_configure\[34\]\[5\] net358 _0938_ gpio_configure\[33\]\[5\] _1016_ VGND
+ VGND VPWR VPWR _1021_ sky130_fd_sc_hd__a221o_1
X_7197_ clknet_3_7_0_wb_clk_i _0799_ net528 VGND VGND VPWR VPWR wbbd_data\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_58_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6148_ gpio_configure\[28\]\[5\] _2861_ VGND VGND VPWR VPWR _2965_ sky130_fd_sc_hd__and2_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1110 _0445_ VGND VGND VPWR VPWR net1643 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1121 gpio_configure\[25\]\[9\] VGND VGND VPWR VPWR net1654 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1132 _0607_ VGND VGND VPWR VPWR net1665 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1143 gpio_configure\[7\]\[2\] VGND VGND VPWR VPWR net1676 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6079_ gpio_configure\[7\]\[2\] _2811_ net395 gpio_configure\[33\]\[2\] _2898_ VGND
+ VGND VPWR VPWR _2899_ sky130_fd_sc_hd__a221o_1
Xhold1154 _0655_ VGND VGND VPWR VPWR net1687 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1165 gpio_configure\[0\]\[9\] VGND VGND VPWR VPWR net1698 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1176 net2121 VGND VGND VPWR VPWR net1709 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1187 net273 VGND VGND VPWR VPWR net1720 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1198 _0188_ VGND VGND VPWR VPWR net1731 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3780_ net11 _0864_ _1054_ gpio_configure\[19\]\[8\] _1365_ VGND VGND VPWR VPWR _1366_
+ sky130_fd_sc_hd__a221o_1
XFILLER_9_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5450_ net464 net1144 _2426_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__mux2_1
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4401_ _0833_ _1610_ VGND VGND VPWR VPWR _1613_ sky130_fd_sc_hd__nand2_2
X_5381_ net447 net1296 _2418_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__mux2_1
Xclkbuf_3_2_0_wb_clk_i clknet_2_1_0_wb_clk_i VGND VGND VPWR VPWR clknet_3_2_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_7120_ clknet_leaf_26_csclk net1412 net519 VGND VGND VPWR VPWR gpio_configure\[35\]\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_4332_ net462 net1405 _1547_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__mux2_1
XFILLER_5_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7051_ clknet_leaf_23_csclk net1329 net515 VGND VGND VPWR VPWR gpio_configure\[26\]\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_87_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4263_ net1148 net446 _1535_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__mux2_1
XFILLER_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6002_ _1450_ _2479_ VGND VGND VPWR VPWR _2824_ sky130_fd_sc_hd__nor2_8
XFILLER_39_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3214_ gpio_configure\[20\]\[3\] VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__inv_2
X_4194_ net1951 clknet_1_0__leaf__1134_ _1520_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__mux2_1
XFILLER_94_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6904_ clknet_leaf_40_csclk net749 net516 VGND VGND VPWR VPWR gpio_configure\[7\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_23_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6835_ clknet_leaf_37_csclk net548 net522 VGND VGND VPWR VPWR mgmt_gpio_data_buf\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6766_ clknet_leaf_71_csclk net1817 net490 VGND VGND VPWR VPWR gpio_configure\[32\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_3978_ net677 net660 _1461_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__mux2_1
X_5717_ gpio_configure\[11\]\[1\] _2505_ _2540_ gpio_configure\[12\]\[1\] VGND VGND
+ VPWR VPWR _2551_ sky130_fd_sc_hd__a22o_1
XFILLER_183_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6697_ clknet_3_7_0_wb_clk_i net2003 net528 VGND VGND VPWR VPWR wbbd_state\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_1__f_mgmt_gpio_in[4] clknet_0_mgmt_gpio_in[4] VGND VGND VPWR VPWR clknet_2_1__leaf_mgmt_gpio_in[4]
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_40_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5648_ xfer_count\[2\] xfer_count\[3\] _0823_ xfer_count\[0\] VGND VGND VPWR VPWR
+ _2484_ sky130_fd_sc_hd__or4b_1
XFILLER_156_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5579_ net435 net934 _2440_ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__mux2_1
XFILLER_163_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold240 _0599_ VGND VGND VPWR VPWR net773 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 serial_bb_data_1 VGND VGND VPWR VPWR net784 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 _0703_ VGND VGND VPWR VPWR net795 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 gpio_configure\[5\]\[10\] VGND VGND VPWR VPWR net806 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold284 _0418_ VGND VGND VPWR VPWR net817 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold295 net2109 VGND VGND VPWR VPWR net828 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_102 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_113 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_124 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_135 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_146 net239 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_157 net371 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_168 net434 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_179 clknet_2_0__leaf_mgmt_gpio_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput8 mask_rev_in[13] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
XFILLER_64_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_272 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4950_ _2157_ _2158_ _2159_ VGND VGND VPWR VPWR _2160_ sky130_fd_sc_hd__nand3b_1
XFILLER_64_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3901_ net2130 _1446_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__or2_1
X_4881_ _1608_ _1952_ _1618_ VGND VGND VPWR VPWR _2092_ sky130_fd_sc_hd__a21oi_1
XTAP_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6620_ clknet_leaf_9_csclk net1092 net509 VGND VGND VPWR VPWR gpio_configure\[4\]\[12\]
+ sky130_fd_sc_hd__dfrtp_4
X_3832_ _0815_ net58 hkspi.state\[3\] VGND VGND VPWR VPWR _1407_ sky130_fd_sc_hd__mux2_1
XFILLER_177_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_550 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6551_ clknet_leaf_27_csclk net1490 net519 VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__dfrtp_1
X_3763_ net4 _0900_ _0928_ gpio_configure\[20\]\[0\] _1348_ VGND VGND VPWR VPWR _1349_
+ sky130_fd_sc_hd__a221o_1
XFILLER_146_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5502_ _0888_ net647 VGND VGND VPWR VPWR _2432_ sky130_fd_sc_hd__nand2_8
XFILLER_146_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6482_ clknet_leaf_72_csclk net1833 net490 VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__dfstp_1
XFILLER_145_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3694_ net53 _0871_ _0931_ gpio_configure\[36\]\[1\] _1281_ VGND VGND VPWR VPWR _1282_
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5433_ net458 net1664 _2424_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__mux2_1
Xoutput301 net301 VGND VGND VPWR VPWR pwr_ctrl_out[0] sky130_fd_sc_hd__buf_12
XFILLER_133_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput312 net312 VGND VGND VPWR VPWR spi_sdi sky130_fd_sc_hd__buf_12
XFILLER_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput323 net1844 VGND VGND VPWR VPWR net1845 sky130_fd_sc_hd__buf_12
XFILLER_160_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput334 net1900 VGND VGND VPWR VPWR net1901 sky130_fd_sc_hd__buf_12
X_5364_ net440 net1546 _2416_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__mux2_1
Xoutput345 net1854 VGND VGND VPWR VPWR net1855 sky130_fd_sc_hd__buf_12
XFILLER_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7103_ clknet_leaf_27_csclk net1603 net521 VGND VGND VPWR VPWR gpio_configure\[33\]\[0\]
+ sky130_fd_sc_hd__dfstp_2
X_4315_ net1282 net456 _1544_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__mux2_1
X_5295_ net355 net647 VGND VGND VPWR VPWR _2409_ sky130_fd_sc_hd__nand2_8
X_7034_ clknet_leaf_64_csclk net1964 net501 VGND VGND VPWR VPWR gpio_configure\[24\]\[0\]
+ sky130_fd_sc_hd__dfstp_4
X_4246_ _1069_ net426 VGND VGND VPWR VPWR _1533_ sky130_fd_sc_hd__nand2_4
XFILLER_19_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4177_ net456 net1320 _1518_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__mux2_1
XFILLER_83_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6818_ clknet_leaf_60_csclk net889 net499 VGND VGND VPWR VPWR serial_bb_enable sky130_fd_sc_hd__dfrtp_4
XFILLER_50_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6749_ clknet_leaf_8_csclk net697 net509 VGND VGND VPWR VPWR gpio_configure\[34\]\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_149_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4100_ net656 net439 net354 VGND VGND VPWR VPWR _1506_ sky130_fd_sc_hd__mux2_1
XFILLER_123_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5080_ _1788_ _2285_ _2132_ VGND VGND VPWR VPWR _2289_ sky130_fd_sc_hd__o21ba_1
XFILLER_56_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4031_ net1363 net456 _1476_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__mux2_1
XFILLER_2_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5982_ _2471_ _2473_ _2796_ VGND VGND VPWR VPWR _2804_ sky130_fd_sc_hd__and3_2
XFILLER_80_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4933_ _1639_ _2142_ VGND VGND VPWR VPWR _2143_ sky130_fd_sc_hd__nor2_1
XFILLER_33_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4864_ _2037_ _2061_ _2073_ _2074_ VGND VGND VPWR VPWR _2075_ sky130_fd_sc_hd__or4_1
XANTENNA_13 _0935_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6603_ clknet_leaf_77_csclk net1663 net484 VGND VGND VPWR VPWR gpio_configure\[1\]\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_3815_ _1395_ net2126 _1388_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__mux2_1
XANTENNA_24 _1004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_35 _1122_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_46 _1346_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4795_ _1993_ _2003_ VGND VGND VPWR VPWR _2006_ sky130_fd_sc_hd__nor2_1
XANTENNA_57 _2494_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6534_ clknet_leaf_6_csclk net1281 net497 VGND VGND VPWR VPWR gpio_configure\[28\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_68 _2528_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_79 _2866_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3746_ gpio_configure\[12\]\[0\] _0921_ _1093_ gpio_configure\[4\]\[8\] _1331_ VGND
+ VGND VPWR VPWR _1332_ sky130_fd_sc_hd__a221o_1
XFILLER_192_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6465_ clknet_2_2__leaf_mgmt_gpio_in[4] _0087_ _0043_ VGND VGND VPWR VPWR hkspi.addr\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3677_ gpio_configure\[3\]\[9\] _1095_ _1103_ gpio_configure\[1\]\[9\] VGND VGND
+ VPWR VPWR _1265_ sky130_fd_sc_hd__a22o_1
XFILLER_173_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5416_ net453 net1152 _2422_ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__mux2_1
X_6396_ net449 net1055 _3182_ VGND VGND VPWR VPWR _0812_ sky130_fd_sc_hd__mux2_1
X_5347_ net438 net1346 _2414_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__mux2_1
XFILLER_102_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput175 net175 VGND VGND VPWR VPWR mgmt_gpio_oeb[0] sky130_fd_sc_hd__buf_12
Xoutput186 net186 VGND VGND VPWR VPWR mgmt_gpio_oeb[1] sky130_fd_sc_hd__buf_12
Xoutput197 net197 VGND VGND VPWR VPWR mgmt_gpio_oeb[2] sky130_fd_sc_hd__buf_12
XFILLER_102_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5278_ net470 net1757 _2407_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__mux2_1
XFILLER_102_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7017_ clknet_leaf_32_csclk net923 net524 VGND VGND VPWR VPWR gpio_configure\[21\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_4229_ wbbd_state\[8\] wbbd_state\[7\] wbbd_state\[9\] VGND VGND VPWR VPWR _1527_
+ sky130_fd_sc_hd__or3_2
XFILLER_75_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3600_ _1184_ _1185_ _1186_ _1189_ VGND VGND VPWR VPWR _1190_ sky130_fd_sc_hd__or4_1
Xinput11 mask_rev_in[16] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput22 mask_rev_in[26] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dlymetal6s2s_1
X_4580_ net477 _1790_ VGND VGND VPWR VPWR _1792_ sky130_fd_sc_hd__nor2_2
Xinput33 mask_rev_in[7] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
XFILLER_162_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput44 mgmt_gpio_in[17] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_2
X_3531_ net553 _0909_ VGND VGND VPWR VPWR _1122_ sky130_fd_sc_hd__nor2_8
Xinput55 mgmt_gpio_in[27] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_2
XFILLER_183_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput66 mgmt_gpio_in[37] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput77 ser_tx VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_1
Xhold806 _0360_ VGND VGND VPWR VPWR net1339 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold817 gpio_configure\[27\]\[2\] VGND VGND VPWR VPWR net1350 sky130_fd_sc_hd__dlygate4sd3_1
Xhold828 _0270_ VGND VGND VPWR VPWR net1361 sky130_fd_sc_hd__dlygate4sd3_1
Xinput88 spimemio_flash_io1_oeb VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_4
X_6250_ gpio_configure\[30\]\[9\] _2799_ net408 gpio_configure\[35\]\[9\] VGND VGND
+ VPWR VPWR _3063_ sky130_fd_sc_hd__a22o_1
XFILLER_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold839 _0550_ VGND VGND VPWR VPWR net1372 sky130_fd_sc_hd__dlygate4sd3_1
Xinput99 wb_adr_i[0] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__buf_12
X_3462_ net590 net1966 VGND VGND VPWR VPWR _1053_ sky130_fd_sc_hd__nor2_8
X_5201_ net469 net1576 _2392_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__mux2_1
XFILLER_115_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6181_ gpio_configure\[33\]\[6\] net395 _2858_ gpio_configure\[24\]\[6\] VGND VGND
+ VPWR VPWR _2997_ sky130_fd_sc_hd__a22o_1
X_3393_ gpio_configure\[28\]\[6\] _0888_ _0892_ gpio_configure\[30\]\[6\] _0977_ VGND
+ VGND VPWR VPWR _0987_ sky130_fd_sc_hd__a221o_1
XFILLER_170_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5132_ _2255_ _2339_ VGND VGND VPWR VPWR _2340_ sky130_fd_sc_hd__or2_1
XFILLER_96_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1506 serial_data_staging_2\[3\] VGND VGND VPWR VPWR net2039 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1517 _0769_ VGND VGND VPWR VPWR net2050 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5063_ _1588_ _1788_ _1725_ VGND VGND VPWR VPWR _2272_ sky130_fd_sc_hd__o21ai_1
Xhold1528 wbbd_data\[5\] VGND VGND VPWR VPWR net2061 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1539 _0808_ VGND VGND VPWR VPWR net2072 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4014_ net1274 net450 _1473_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__mux2_1
XFILLER_65_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5965_ gpio_configure\[7\]\[12\] _2528_ _2535_ gpio_configure\[23\]\[12\] VGND VGND
+ VPWR VPWR _2788_ sky130_fd_sc_hd__a22o_1
X_4916_ _1826_ _1890_ VGND VGND VPWR VPWR _2127_ sky130_fd_sc_hd__nand2_1
XFILLER_178_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5896_ gpio_configure\[21\]\[9\] _2521_ _2529_ gpio_configure\[29\]\[9\] _2721_ VGND
+ VGND VPWR VPWR _2722_ sky130_fd_sc_hd__a221o_1
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4847_ _1700_ _1898_ VGND VGND VPWR VPWR _2058_ sky130_fd_sc_hd__nand2_1
XFILLER_148_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4778_ _1584_ _1770_ VGND VGND VPWR VPWR _1989_ sky130_fd_sc_hd__nand2_1
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3729_ net390 _1006_ VGND VGND VPWR VPWR _1316_ sky130_fd_sc_hd__nor2_1
X_6517_ clknet_leaf_78_csclk net1675 net486 VGND VGND VPWR VPWR gpio_configure\[24\]\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_180_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6448_ clknet_2_3__leaf_mgmt_gpio_in[4] _0070_ _0026_ VGND VGND VPWR VPWR hkspi.odata\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_134_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6379_ wbbd_state\[9\] net153 net136 wbbd_state\[8\] _3173_ VGND VGND VPWR VPWR _3174_
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5750_ _2575_ _2578_ _2580_ _2582_ VGND VGND VPWR VPWR _2583_ sky130_fd_sc_hd__or4_1
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4701_ _1579_ net477 _1833_ _1911_ _1912_ VGND VGND VPWR VPWR _1913_ sky130_fd_sc_hd__o311a_1
X_5681_ _2497_ _2503_ _2509_ _2515_ VGND VGND VPWR VPWR _2516_ sky130_fd_sc_hd__or4_1
XFILLER_30_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4632_ _1779_ _1788_ VGND VGND VPWR VPWR _1844_ sky130_fd_sc_hd__nor2_1
XFILLER_135_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4563_ net124 _1773_ VGND VGND VPWR VPWR _1775_ sky130_fd_sc_hd__nand2_2
Xhold603 gpio_configure\[17\]\[3\] VGND VGND VPWR VPWR net1136 sky130_fd_sc_hd__dlygate4sd3_1
X_6302_ gpio_configure\[23\]\[11\] _2822_ _2828_ gpio_configure\[20\]\[11\] VGND VGND
+ VPWR VPWR _3113_ sky130_fd_sc_hd__a22o_1
X_3514_ gpio_configure\[16\]\[4\] _0912_ _1101_ gpio_configure\[32\]\[12\] _1104_
+ VGND VGND VPWR VPWR _1105_ sky130_fd_sc_hd__a221o_1
Xhold614 _0594_ VGND VGND VPWR VPWR net1147 sky130_fd_sc_hd__dlygate4sd3_1
Xhold625 gpio_configure\[30\]\[4\] VGND VGND VPWR VPWR net1158 sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 _0292_ VGND VGND VPWR VPWR net1169 sky130_fd_sc_hd__dlygate4sd3_1
X_4494_ _0834_ _1585_ VGND VGND VPWR VPWR _1706_ sky130_fd_sc_hd__nor2_4
Xmax_cap355 _0914_ VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__buf_6
Xhold647 gpio_configure\[5\]\[4\] VGND VGND VPWR VPWR net1180 sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 _0553_ VGND VGND VPWR VPWR net1191 sky130_fd_sc_hd__dlygate4sd3_1
X_6233_ gpio_configure\[37\]\[8\] _2806_ net416 gpio_configure\[32\]\[8\] _3035_ VGND
+ VGND VPWR VPWR _3047_ sky130_fd_sc_hd__a221o_1
XFILLER_171_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap377 net553 VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__buf_12
X_3445_ _1013_ _1015_ _1034_ _1036_ VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__or4_1
XFILLER_116_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold669 gpio_configure\[5\]\[12\] VGND VGND VPWR VPWR net1202 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_170_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap388 net639 VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__buf_12
Xmax_cap399 _2819_ VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__buf_8
XFILLER_170_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6164_ gpio_configure\[1\]\[5\] net401 net405 gpio_configure\[24\]\[5\] _2980_ VGND
+ VGND VPWR VPWR _2981_ sky130_fd_sc_hd__a221o_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ _0971_ net2008 _0970_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__mux2_1
XFILLER_97_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5115_ _1789_ _1832_ VGND VGND VPWR VPWR _2323_ sky130_fd_sc_hd__or2_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1303 gpio_configure\[25\]\[8\] VGND VGND VPWR VPWR net1836 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6095_ gpio_configure\[0\]\[2\] _2851_ _2905_ _2914_ _0824_ VGND VGND VPWR VPWR _2915_
+ sky130_fd_sc_hd__o221a_1
Xhold1314 net1847 VGND VGND VPWR VPWR wb_dat_o[17] sky130_fd_sc_hd__buf_12
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1325 net1941 VGND VGND VPWR VPWR net1858 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1336 net1869 VGND VGND VPWR VPWR wb_dat_o[8] sky130_fd_sc_hd__buf_12
Xhold1347 net1952 VGND VGND VPWR VPWR net1880 sky130_fd_sc_hd__dlygate4sd3_1
X_5046_ _1652_ _1670_ _1958_ _2091_ _2213_ VGND VGND VPWR VPWR _2255_ sky130_fd_sc_hd__a2111o_1
XFILLER_27_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1358 net1891 VGND VGND VPWR VPWR wb_dat_o[18] sky130_fd_sc_hd__buf_12
XFILLER_84_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1369 net2081 VGND VGND VPWR VPWR net1902 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6997_ clknet_leaf_57_csclk net813 net503 VGND VGND VPWR VPWR gpio_configure\[19\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_25_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5948_ net2082 _2771_ net366 VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__mux2_1
XFILLER_178_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5879_ _2698_ _2701_ _2703_ _2705_ VGND VGND VPWR VPWR _2706_ sky130_fd_sc_hd__or4_1
XFILLER_139_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3230_ gpio_configure\[4\]\[3\] VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__inv_2
XFILLER_100_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6920_ clknet_leaf_53_csclk net1343 net507 VGND VGND VPWR VPWR gpio_configure\[9\]\[6\]
+ sky130_fd_sc_hd__dfrtp_2
X_6851_ clknet_leaf_48_csclk net1462 net514 VGND VGND VPWR VPWR gpio_configure\[1\]\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_23_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5802_ gpio_configure\[14\]\[5\] _2494_ _2520_ gpio_configure\[8\]\[5\] _2631_ VGND
+ VGND VPWR VPWR _2632_ sky130_fd_sc_hd__a221o_1
XFILLER_90_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3994_ net1728 net461 _1471_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__mux2_1
XFILLER_62_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6782_ clknet_3_7_0_wb_clk_i _0385_ net529 VGND VGND VPWR VPWR wbbd_addr\[6\] sky130_fd_sc_hd__dfrtp_1
X_5733_ gpio_configure\[28\]\[2\] _2513_ _2535_ gpio_configure\[23\]\[2\] _2565_ VGND
+ VGND VPWR VPWR _2566_ sky130_fd_sc_hd__a221o_1
XFILLER_176_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5664_ pad_count_1\[4\] _2459_ _2488_ VGND VGND VPWR VPWR _2499_ sky130_fd_sc_hd__and3_4
XFILLER_176_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_54_csclk clknet_3_3_0_csclk VGND VGND VPWR VPWR clknet_leaf_54_csclk
+ sky130_fd_sc_hd__clkbuf_16
X_4615_ _1795_ _1803_ net432 _1798_ VGND VGND VPWR VPWR _1827_ sky130_fd_sc_hd__o22a_1
XFILLER_135_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5595_ _2446_ VGND VGND VPWR VPWR _2447_ sky130_fd_sc_hd__inv_2
XFILLER_163_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold400 _0436_ VGND VGND VPWR VPWR net933 sky130_fd_sc_hd__dlygate4sd3_1
X_4546_ _0817_ _1754_ VGND VGND VPWR VPWR _1758_ sky130_fd_sc_hd__xnor2_2
Xhold411 net234 VGND VGND VPWR VPWR net944 sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 _0169_ VGND VGND VPWR VPWR net955 sky130_fd_sc_hd__dlygate4sd3_1
Xhold433 gpio_configure\[34\]\[7\] VGND VGND VPWR VPWR net966 sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 _0725_ VGND VGND VPWR VPWR net977 sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 gpio_configure\[18\]\[12\] VGND VGND VPWR VPWR net988 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold466 _0488_ VGND VGND VPWR VPWR net999 sky130_fd_sc_hd__dlygate4sd3_1
X_4477_ _1590_ _1688_ VGND VGND VPWR VPWR _1689_ sky130_fd_sc_hd__or2_4
Xhold477 _0672_ VGND VGND VPWR VPWR net1010 sky130_fd_sc_hd__dlygate4sd3_1
Xhold488 gpio_configure\[33\]\[12\] VGND VGND VPWR VPWR net1021 sky130_fd_sc_hd__dlygate4sd3_1
Xhold499 _0212_ VGND VGND VPWR VPWR net1032 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_69_csclk clknet_3_1_0_csclk VGND VGND VPWR VPWR clknet_leaf_69_csclk
+ sky130_fd_sc_hd__clkbuf_16
X_6216_ _3014_ _3015_ _3028_ _3030_ VGND VGND VPWR VPWR _3031_ sky130_fd_sc_hd__or4_1
X_3428_ gpio_configure\[21\]\[5\] _0911_ _0917_ gpio_configure\[29\]\[5\] _1011_ VGND
+ VGND VPWR VPWR _1020_ sky130_fd_sc_hd__a221o_1
X_7196_ clknet_3_5_0_wb_clk_i _0798_ VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__dfxtp_1
XFILLER_38_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6147_ gpio_configure\[36\]\[5\] net403 net402 gpio_configure\[4\]\[5\] VGND VGND
+ VPWR VPWR _2964_ sky130_fd_sc_hd__a22o_1
X_3359_ gpio_configure\[20\]\[7\] _0928_ net351 net70 _0954_ VGND VGND VPWR VPWR _0955_
+ sky130_fd_sc_hd__a221o_1
Xhold1100 _0346_ VGND VGND VPWR VPWR net1633 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1111 gpio_configure\[10\]\[0\] VGND VGND VPWR VPWR net1644 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1122 _0149_ VGND VGND VPWR VPWR net1655 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_161_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1133 gpio_configure\[18\]\[10\] VGND VGND VPWR VPWR net1666 sky130_fd_sc_hd__dlygate4sd3_1
X_6078_ gpio_configure\[15\]\[2\] net407 net404 gpio_configure\[25\]\[2\] VGND VGND
+ VPWR VPWR _2898_ sky130_fd_sc_hd__a22o_1
Xhold1144 _0503_ VGND VGND VPWR VPWR net1677 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1155 gpio_configure\[26\]\[0\] VGND VGND VPWR VPWR net1688 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1166 _0210_ VGND VGND VPWR VPWR net1699 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1177 _0171_ VGND VGND VPWR VPWR net1710 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_638 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5029_ _2237_ _2238_ _2235_ _2236_ VGND VGND VPWR VPWR _2239_ sky130_fd_sc_hd__and4b_1
Xhold1188 _0402_ VGND VGND VPWR VPWR net1721 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1199 net2138 VGND VGND VPWR VPWR net1732 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4400_ net99 _1611_ VGND VGND VPWR VPWR _1612_ sky130_fd_sc_hd__nor2_4
X_5380_ net453 net1160 _2418_ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__mux2_1
XFILLER_126_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4331_ net467 net1769 _1547_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__mux2_1
XFILLER_5_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7050_ clknet_leaf_60_csclk net1689 net498 VGND VGND VPWR VPWR gpio_configure\[26\]\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_4262_ net681 net569 _1535_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__mux2_1
XFILLER_99_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6001_ _2797_ _2818_ VGND VGND VPWR VPWR _2823_ sky130_fd_sc_hd__nor2_8
X_3213_ gpio_configure\[21\]\[3\] VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__inv_2
X_4193_ net1957 _1191_ _1520_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__mux2_1
XFILLER_79_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6903_ clknet_leaf_38_csclk net1553 net522 VGND VGND VPWR VPWR gpio_configure\[7\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6834_ clknet_leaf_40_csclk net1452 net522 VGND VGND VPWR VPWR mgmt_gpio_data_buf\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_6765_ clknet_leaf_69_csclk net1247 net491 VGND VGND VPWR VPWR gpio_configure\[21\]\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3977_ net658 net664 wbbd_busy VGND VGND VPWR VPWR _1467_ sky130_fd_sc_hd__mux2_1
XFILLER_50_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5716_ gpio_configure\[20\]\[1\] _2499_ _2549_ VGND VGND VPWR VPWR _2550_ sky130_fd_sc_hd__a21o_1
XFILLER_148_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6696_ clknet_3_7_0_wb_clk_i _0010_ net528 VGND VGND VPWR VPWR wbbd_state\[5\] sky130_fd_sc_hd__dfrtp_4
XFILLER_109_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5647_ _1452_ net2033 _2483_ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__mux2_1
XFILLER_40_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5578_ net438 net1391 _2440_ VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__mux2_1
XFILLER_151_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold230 _0170_ VGND VGND VPWR VPWR net763 sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 gpio_configure\[2\]\[10\] VGND VGND VPWR VPWR net774 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold252 _0419_ VGND VGND VPWR VPWR net785 sky130_fd_sc_hd__dlygate4sd3_1
X_4529_ net380 _1683_ _1691_ VGND VGND VPWR VPWR _1741_ sky130_fd_sc_hd__a21oi_1
XFILLER_6_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold263 gpio_configure\[12\]\[6\] VGND VGND VPWR VPWR net796 sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 _0236_ VGND VGND VPWR VPWR net807 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold285 net304 VGND VGND VPWR VPWR net818 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold296 _0204_ VGND VGND VPWR VPWR net829 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7179_ clknet_3_3_0_wb_clk_i _0781_ net506 VGND VGND VPWR VPWR serial_data_staging_2\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_103 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_114 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_125 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_136 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_147 net261 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_158 net371 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_169 net445 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput9 mask_rev_in[14] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_76_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3900_ net473 _1445_ VGND VGND VPWR VPWR _1446_ sky130_fd_sc_hd__nor2_1
XFILLER_32_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4880_ _1652_ _1662_ _1959_ VGND VGND VPWR VPWR _2091_ sky130_fd_sc_hd__a21o_1
XTAP_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3831_ _1405_ _1406_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__xnor2_1
XFILLER_32_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3762_ gpio_configure\[19\]\[0\] _0896_ _1125_ gpio_configure\[22\]\[8\] VGND VGND
+ VPWR VPWR _1348_ sky130_fd_sc_hd__a22o_1
X_6550_ clknet_leaf_27_csclk net915 net519 VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__dfrtp_1
XFILLER_158_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5501_ net435 net1095 net641 VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__mux2_1
X_6481_ clknet_leaf_60_csclk net1259 net498 VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__dfstp_2
X_3693_ gpio_configure\[28\]\[1\] _0888_ _1056_ gpio_configure\[12\]\[9\] VGND VGND
+ VPWR VPWR _1281_ sky130_fd_sc_hd__a22o_1
XFILLER_145_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5432_ net463 net890 _2424_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__mux2_1
Xoutput302 net302 VGND VGND VPWR VPWR pwr_ctrl_out[1] sky130_fd_sc_hd__buf_12
XFILLER_133_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput313 net313 VGND VGND VPWR VPWR spimemio_flash_io0_di sky130_fd_sc_hd__buf_12
Xoutput324 net1840 VGND VGND VPWR VPWR net1841 sky130_fd_sc_hd__buf_12
X_5363_ net447 net1208 _2416_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__mux2_1
Xoutput335 net1898 VGND VGND VPWR VPWR net1899 sky130_fd_sc_hd__buf_12
Xoutput346 net1858 VGND VGND VPWR VPWR net1859 sky130_fd_sc_hd__buf_12
X_7102_ clknet_leaf_58_csclk net1263 net503 VGND VGND VPWR VPWR gpio_configure\[32\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_4314_ net1338 net462 _1544_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__mux2_1
XFILLER_87_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5294_ net435 net930 net565 VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__mux2_1
XFILLER_113_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7033_ clknet_leaf_57_csclk net1279 net504 VGND VGND VPWR VPWR gpio_configure\[23\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_4245_ net1230 net444 _1532_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__mux2_1
XFILLER_101_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4176_ net462 net1483 _1518_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__mux2_1
XFILLER_142_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6817_ clknet_leaf_60_csclk net1410 net499 VGND VGND VPWR VPWR serial_bb_data_2 sky130_fd_sc_hd__dfrtp_1
XFILLER_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6748_ clknet_leaf_8_csclk net759 net509 VGND VGND VPWR VPWR gpio_configure\[34\]\[10\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_167_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6679_ clknet_leaf_10_csclk net1169 net511 VGND VGND VPWR VPWR gpio_configure\[11\]\[12\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_109_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4030_ net1473 net462 _1476_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__mux2_1
XFILLER_111_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5981_ gpio_configure\[30\]\[0\] _2799_ net401 gpio_configure\[1\]\[0\] VGND VGND
+ VPWR VPWR _2803_ sky130_fd_sc_hd__a22o_1
XFILLER_18_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4932_ _1605_ _2141_ VGND VGND VPWR VPWR _2142_ sky130_fd_sc_hd__or2_1
XFILLER_17_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4863_ _1726_ _1904_ VGND VGND VPWR VPWR _2074_ sky130_fd_sc_hd__nand2_1
XFILLER_33_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_14 _0948_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6602_ clknet_leaf_77_csclk net1685 net484 VGND VGND VPWR VPWR gpio_configure\[1\]\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_25 _1004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3814_ _0819_ _1391_ _1394_ _0840_ VGND VGND VPWR VPWR _1395_ sky130_fd_sc_hd__a31o_1
XFILLER_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_36 _1122_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4794_ _1772_ _2003_ _2004_ VGND VGND VPWR VPWR _2005_ sky130_fd_sc_hd__or3_1
XANTENNA_47 _1365_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_58 _2496_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6533_ clknet_leaf_69_csclk net1747 net491 VGND VGND VPWR VPWR gpio_configure\[28\]\[10\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_69 _2532_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3745_ gpio_configure\[13\]\[8\] _1045_ _1069_ gpio_configure\[14\]\[8\] VGND VGND
+ VPWR VPWR _1331_ sky130_fd_sc_hd__a22o_1
XFILLER_146_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6464_ clknet_2_2__leaf_mgmt_gpio_in[4] _0086_ _0042_ VGND VGND VPWR VPWR hkspi.addr\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3676_ gpio_configure\[14\]\[9\] _1069_ _1081_ gpio_configure\[34\]\[9\] _1263_ VGND
+ VGND VPWR VPWR _1264_ sky130_fd_sc_hd__a221o_1
XFILLER_134_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5415_ net457 net850 _2422_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__mux2_1
X_6395_ net455 net1514 _3182_ VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__mux2_1
XFILLER_133_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5346_ net441 net1120 _2414_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__mux2_1
XFILLER_0_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput176 net176 VGND VGND VPWR VPWR mgmt_gpio_oeb[10] sky130_fd_sc_hd__buf_12
Xoutput187 net187 VGND VGND VPWR VPWR mgmt_gpio_oeb[20] sky130_fd_sc_hd__buf_12
XFILLER_99_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput198 net198 VGND VGND VPWR VPWR mgmt_gpio_oeb[30] sky130_fd_sc_hd__buf_12
XFILLER_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5277_ _0915_ net647 VGND VGND VPWR VPWR _2407_ sky130_fd_sc_hd__nand2_8
XFILLER_87_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7016_ clknet_leaf_51_csclk net1355 net506 VGND VGND VPWR VPWR gpio_configure\[21\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_102_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4228_ wbbd_state\[8\] wbbd_state\[7\] wbbd_state\[9\] VGND VGND VPWR VPWR _1526_
+ sky130_fd_sc_hd__nor3_1
XFILLER_28_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4159_ _1119_ net429 VGND VGND VPWR VPWR _1516_ sky130_fd_sc_hd__and2_2
XFILLER_83_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput12 mask_rev_in[17] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
Xinput23 mask_rev_in[27] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_2
Xinput34 mask_rev_in[8] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_1
XFILLER_128_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput45 mgmt_gpio_in[18] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_2
X_3530_ _0885_ net382 VGND VGND VPWR VPWR _1121_ sky130_fd_sc_hd__nor2_2
Xinput56 mgmt_gpio_in[28] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_2
Xinput67 mgmt_gpio_in[3] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__buf_6
Xhold807 gpio_configure\[3\]\[10\] VGND VGND VPWR VPWR net1340 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput78 spi_csb VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_1
XFILLER_128_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold818 _0663_ VGND VGND VPWR VPWR net1351 sky130_fd_sc_hd__dlygate4sd3_1
Xinput89 spimemio_flash_io2_do VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold829 net1981 VGND VGND VPWR VPWR net1362 sky130_fd_sc_hd__dlygate4sd3_1
X_3461_ net48 _0904_ _1051_ gpio_configure\[35\]\[12\] _1050_ VGND VGND VPWR VPWR
+ _1052_ sky130_fd_sc_hd__a221o_1
X_5200_ _1299_ net425 VGND VGND VPWR VPWR _2392_ sky130_fd_sc_hd__nand2_1
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6180_ _2989_ _2991_ _2993_ _2995_ VGND VGND VPWR VPWR _2996_ sky130_fd_sc_hd__or4_1
X_3392_ _0980_ _0982_ _0984_ _0985_ VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__or4_1
X_5131_ _1666_ _1670_ _1942_ _2089_ _2204_ VGND VGND VPWR VPWR _2339_ sky130_fd_sc_hd__a2111o_1
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1507 serial_data_staging_2\[0\] VGND VGND VPWR VPWR net2040 sky130_fd_sc_hd__dlygate4sd3_1
X_5062_ _2168_ _2266_ _2268_ _2270_ VGND VGND VPWR VPWR _2271_ sky130_fd_sc_hd__nand4_1
Xhold1518 serial_data_staging_2\[4\] VGND VGND VPWR VPWR net2051 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1529 wbbd_data\[6\] VGND VGND VPWR VPWR net2062 sky130_fd_sc_hd__dlygate4sd3_1
X_4013_ net1646 net455 _1473_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__mux2_1
XFILLER_37_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5964_ gpio_configure\[8\]\[12\] _2520_ _2529_ gpio_configure\[29\]\[12\] _2786_
+ VGND VGND VPWR VPWR _2787_ sky130_fd_sc_hd__a221o_1
XFILLER_52_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4915_ _1843_ _2118_ _2119_ _2125_ VGND VGND VPWR VPWR _2126_ sky130_fd_sc_hd__or4b_1
XFILLER_178_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5895_ gpio_configure\[20\]\[9\] _2499_ _2524_ _2720_ VGND VGND VPWR VPWR _2721_
+ sky130_fd_sc_hd__a22o_1
XFILLER_178_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4846_ net110 net124 _0834_ _1675_ VGND VGND VPWR VPWR _2057_ sky130_fd_sc_hd__and4_1
XFILLER_193_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4777_ _1707_ net424 _1576_ VGND VGND VPWR VPWR _1988_ sky130_fd_sc_hd__a21oi_2
XFILLER_165_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6516_ clknet_leaf_78_csclk net1829 net486 VGND VGND VPWR VPWR gpio_configure\[24\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_3728_ gpio_configure\[3\]\[0\] _0915_ _1110_ gpio_configure\[2\]\[8\] VGND VGND
+ VPWR VPWR _1315_ sky130_fd_sc_hd__a22o_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6447_ clknet_2_3__leaf_mgmt_gpio_in[4] _0069_ _0025_ VGND VGND VPWR VPWR hkspi.odata\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3659_ _1240_ _1242_ _1243_ _1247_ VGND VGND VPWR VPWR _1248_ sky130_fd_sc_hd__or4_1
XFILLER_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6378_ wbbd_state\[7\] net145 net159 net433 VGND VGND VPWR VPWR _3173_ sky130_fd_sc_hd__a22o_1
XFILLER_87_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5329_ net1920 net535 _2412_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__mux2_1
XFILLER_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_660 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4700_ _1863_ _1873_ _1886_ _1757_ VGND VGND VPWR VPWR _1912_ sky130_fd_sc_hd__a31o_1
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5680_ gpio_configure\[15\]\[0\] _2510_ _2511_ gpio_configure\[25\]\[0\] _2514_ VGND
+ VGND VPWR VPWR _2515_ sky130_fd_sc_hd__a221o_1
XFILLER_187_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4631_ _1840_ _1842_ VGND VGND VPWR VPWR _1843_ sky130_fd_sc_hd__nand2b_1
XFILLER_147_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4562_ net530 _1556_ VGND VGND VPWR VPWR _1774_ sky130_fd_sc_hd__or2_2
XFILLER_116_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6301_ gpio_configure\[29\]\[11\] _2816_ _2820_ gpio_configure\[21\]\[11\] _3110_
+ VGND VGND VPWR VPWR _3112_ sky130_fd_sc_hd__a221o_1
XFILLER_156_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold604 _0584_ VGND VGND VPWR VPWR net1137 sky130_fd_sc_hd__dlygate4sd3_1
X_3513_ gpio_configure\[15\]\[12\] _1102_ _1103_ gpio_configure\[1\]\[12\] VGND VGND
+ VPWR VPWR _1104_ sky130_fd_sc_hd__a22o_1
Xhold615 gpio_configure\[16\]\[12\] VGND VGND VPWR VPWR net1148 sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 _0689_ VGND VGND VPWR VPWR net1159 sky130_fd_sc_hd__dlygate4sd3_1
X_4493_ _1576_ _1678_ VGND VGND VPWR VPWR _1705_ sky130_fd_sc_hd__or2_1
Xhold637 gpio_configure\[17\]\[4\] VGND VGND VPWR VPWR net1170 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap356 _0904_ VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__buf_8
Xhold648 _0489_ VGND VGND VPWR VPWR net1181 sky130_fd_sc_hd__dlygate4sd3_1
X_6232_ _3040_ _3041_ _3043_ _3045_ VGND VGND VPWR VPWR _3046_ sky130_fd_sc_hd__or4_1
Xmax_cap367 _0937_ VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__buf_8
XFILLER_131_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold659 gpio_configure\[16\]\[3\] VGND VGND VPWR VPWR net1192 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap378 net628 VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__buf_12
XFILLER_131_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3444_ net49 net356 _0932_ gpio_configure\[35\]\[5\] _1035_ VGND VGND VPWR VPWR _1036_
+ sky130_fd_sc_hd__a221o_1
Xmax_cap389 net390 VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__buf_12
XFILLER_131_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3375_ _0969_ net2004 _0837_ VGND VGND VPWR VPWR _0971_ sky130_fd_sc_hd__mux2_1
X_6163_ gpio_configure\[31\]\[5\] net423 net415 gpio_configure\[11\]\[5\] VGND VGND
+ VPWR VPWR _2980_ sky130_fd_sc_hd__a22o_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5114_ _2001_ _2179_ _2302_ _2321_ VGND VGND VPWR VPWR _2322_ sky130_fd_sc_hd__or4_1
Xhold1304 _0148_ VGND VGND VPWR VPWR net1837 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ net365 _2907_ _2909_ _2913_ VGND VGND VPWR VPWR _2914_ sky130_fd_sc_hd__or4_1
XFILLER_111_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1315 net1934 VGND VGND VPWR VPWR net1848 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1326 net1859 VGND VGND VPWR VPWR wb_dat_o[6] sky130_fd_sc_hd__buf_12
Xhold1337 net1947 VGND VGND VPWR VPWR net1870 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1348 net1881 VGND VGND VPWR VPWR wb_dat_o[1] sky130_fd_sc_hd__buf_12
X_5045_ _2106_ _2208_ VGND VGND VPWR VPWR _2254_ sky130_fd_sc_hd__or2_1
Xhold1359 net1959 VGND VGND VPWR VPWR net1892 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6996_ clknet_leaf_65_csclk net773 net505 VGND VGND VPWR VPWR gpio_configure\[19\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5947_ xfer_state\[1\] serial_data_staging_1\[10\] _2770_ VGND VGND VPWR VPWR _2771_
+ sky130_fd_sc_hd__a21o_1
XFILLER_43_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5878_ gpio_configure\[4\]\[8\] _2502_ _2529_ gpio_configure\[29\]\[8\] _2704_ VGND
+ VGND VPWR VPWR _2705_ sky130_fd_sc_hd__a221o_1
X_4829_ _1556_ _1694_ _1700_ VGND VGND VPWR VPWR _2040_ sky130_fd_sc_hd__o21ai_1
XFILLER_138_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1 hkspi.odata\[6\] VGND VGND VPWR VPWR net534 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6850_ clknet_leaf_17_csclk net1764 net512 VGND VGND VPWR VPWR gpio_configure\[1\]\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5801_ gpio_configure\[10\]\[5\] _2507_ _2540_ gpio_configure\[12\]\[5\] VGND VGND
+ VPWR VPWR _2631_ sky130_fd_sc_hd__a22o_1
X_6781_ clknet_3_6_0_wb_clk_i _0384_ net529 VGND VGND VPWR VPWR wbbd_addr\[5\] sky130_fd_sc_hd__dfrtp_1
X_3993_ net1826 net466 _1471_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__mux2_1
X_5732_ gpio_configure\[20\]\[2\] _2499_ _2541_ gpio_configure\[31\]\[2\] VGND VGND
+ VPWR VPWR _2565_ sky130_fd_sc_hd__a22o_1
X_5663_ pad_count_1\[4\] _2488_ _2489_ VGND VGND VPWR VPWR _2498_ sky130_fd_sc_hd__and3_4
XFILLER_148_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4614_ _1692_ _1825_ VGND VGND VPWR VPWR _1826_ sky130_fd_sc_hd__or2_1
X_5594_ xfer_state\[3\] net475 xfer_state\[2\] _2444_ VGND VGND VPWR VPWR _2446_ sky130_fd_sc_hd__o31a_1
XFILLER_128_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold401 gpio_configure\[36\]\[7\] VGND VGND VPWR VPWR net934 sky130_fd_sc_hd__dlygate4sd3_1
X_4545_ _0835_ _0836_ _1755_ VGND VGND VPWR VPWR _1757_ sky130_fd_sc_hd__or3_4
XFILLER_144_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold412 _0434_ VGND VGND VPWR VPWR net945 sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 gpio_configure\[33\]\[5\] VGND VGND VPWR VPWR net956 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold434 _0721_ VGND VGND VPWR VPWR net967 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold445 gpio_configure\[8\]\[3\] VGND VGND VPWR VPWR net978 sky130_fd_sc_hd__dlygate4sd3_1
Xhold456 _0338_ VGND VGND VPWR VPWR net989 sky130_fd_sc_hd__dlygate4sd3_1
X_4476_ net127 net128 net126 net125 VGND VGND VPWR VPWR _1688_ sky130_fd_sc_hd__or4b_1
Xhold467 gpio_configure\[25\]\[12\] VGND VGND VPWR VPWR net1000 sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 net270 VGND VGND VPWR VPWR net1011 sky130_fd_sc_hd__dlygate4sd3_1
Xhold489 _0363_ VGND VGND VPWR VPWR net1022 sky130_fd_sc_hd__dlygate4sd3_1
X_6215_ gpio_configure\[1\]\[7\] net401 net405 gpio_configure\[24\]\[7\] _3029_ VGND
+ VGND VPWR VPWR _3030_ sky130_fd_sc_hd__a221o_1
X_3427_ gpio_configure\[1\]\[5\] _0934_ _1007_ net66 _1018_ VGND VGND VPWR VPWR _1019_
+ sky130_fd_sc_hd__a221o_1
X_7195_ clknet_3_5_0_wb_clk_i _0797_ VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__dfxtp_1
XFILLER_131_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6146_ net2051 _2963_ net366 VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__mux2_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3358_ net51 _0904_ net367 gpio_configure\[17\]\[7\] VGND VGND VPWR VPWR _0954_ sky130_fd_sc_hd__a22o_2
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1101 gpio_configure\[0\]\[10\] VGND VGND VPWR VPWR net1634 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1112 _0525_ VGND VGND VPWR VPWR net1645 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1123 gpio_configure\[14\]\[2\] VGND VGND VPWR VPWR net1656 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1134 _0336_ VGND VGND VPWR VPWR net1667 sky130_fd_sc_hd__dlygate4sd3_1
X_6077_ gpio_configure\[2\]\[2\] _2823_ net394 gpio_configure\[6\]\[2\] _2896_ VGND
+ VGND VPWR VPWR _2897_ sky130_fd_sc_hd__a221o_1
XFILLER_161_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1145 gpio_configure\[3\]\[8\] VGND VGND VPWR VPWR net1678 sky130_fd_sc_hd__dlygate4sd3_1
X_3289_ _0879_ _0884_ VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__nand2_8
Xhold1156 _0653_ VGND VGND VPWR VPWR net1689 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1167 gpio_configure\[2\]\[8\] VGND VGND VPWR VPWR net1700 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1178 gpio_configure\[18\]\[8\] VGND VGND VPWR VPWR net1711 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5028_ _1808_ _1992_ _1689_ VGND VGND VPWR VPWR _2238_ sky130_fd_sc_hd__a21o_1
XTAP_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1189 net220 VGND VGND VPWR VPWR net1722 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_110_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6979_ clknet_leaf_20_csclk net869 net514 VGND VGND VPWR VPWR gpio_configure\[17\]\[1\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_110_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_107 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold990 _0538_ VGND VGND VPWR VPWR net1523 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_663 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4330_ _1125_ net426 VGND VGND VPWR VPWR _1547_ sky130_fd_sc_hd__nand2_2
XFILLER_5_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4261_ net766 net577 _1535_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__mux2_1
XFILLER_5_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6000_ _1449_ _2469_ _2478_ VGND VGND VPWR VPWR _2822_ sky130_fd_sc_hd__and3_4
XFILLER_140_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3212_ gpio_configure\[22\]\[3\] VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__inv_2
XFILLER_86_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4192_ net1961 _1249_ _1520_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__mux2_1
XFILLER_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6902_ clknet_leaf_16_csclk net1303 net512 VGND VGND VPWR VPWR gpio_configure\[7\]\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_54_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6833_ clknet_leaf_33_csclk net933 net524 VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__dfrtp_1
XFILLER_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6764_ clknet_leaf_0_csclk net1245 net486 VGND VGND VPWR VPWR gpio_configure\[21\]\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_3976_ net1015 net443 _1461_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__mux2_1
X_5715_ gpio_configure\[27\]\[1\] _2506_ _2529_ gpio_configure\[29\]\[1\] VGND VGND
+ VPWR VPWR _2549_ sky130_fd_sc_hd__a22o_1
XFILLER_148_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6695_ clknet_3_7_0_wb_clk_i _0003_ net528 VGND VGND VPWR VPWR wbbd_state\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_136_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5646_ _2445_ _2457_ _2482_ xfer_state\[3\] VGND VGND VPWR VPWR _2483_ sky130_fd_sc_hd__a22o_1
XFILLER_163_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5577_ net440 net1560 _2440_ VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__mux2_1
Xhold220 _0231_ VGND VGND VPWR VPWR net753 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold231 serial_bb_load VGND VGND VPWR VPWR net764 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4528_ _1673_ _1700_ _1709_ _1739_ VGND VGND VPWR VPWR _1740_ sky130_fd_sc_hd__and4b_1
XFILLER_191_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold242 _0221_ VGND VGND VPWR VPWR net775 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 gpio_configure\[35\]\[10\] VGND VGND VPWR VPWR net786 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 _0547_ VGND VGND VPWR VPWR net797 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold275 gpio_configure\[23\]\[3\] VGND VGND VPWR VPWR net808 sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 _0413_ VGND VGND VPWR VPWR net819 sky130_fd_sc_hd__dlygate4sd3_1
X_4459_ net530 _1631_ VGND VGND VPWR VPWR _1671_ sky130_fd_sc_hd__nand2_8
XFILLER_131_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold297 gpio_configure\[17\]\[9\] VGND VGND VPWR VPWR net830 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7178_ clknet_3_3_0_wb_clk_i _0780_ net505 VGND VGND VPWR VPWR serial_data_staging_2\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_105_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6129_ gpio_configure\[18\]\[4\] _2819_ net410 gpio_configure\[8\]\[4\] VGND VGND
+ VPWR VPWR _2947_ sky130_fd_sc_hd__a22o_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_104 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_115 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_126 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_137 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_148 net263 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_159 net375 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_466 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_53_csclk clknet_3_3_0_csclk VGND VGND VPWR VPWR clknet_leaf_53_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_189_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3830_ _0815_ _1388_ VGND VGND VPWR VPWR _1406_ sky130_fd_sc_hd__nor2_1
XFILLER_32_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3761_ gpio_configure\[20\]\[8\] _1053_ _1302_ irq_1_inputsrc VGND VGND VPWR VPWR
+ _1347_ sky130_fd_sc_hd__a22o_1
XFILLER_158_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5500_ net439 net1923 net641 VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__mux2_1
XFILLER_158_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6480_ clknet_leaf_60_csclk net1450 net498 VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__dfstp_2
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3692_ gpio_configure\[2\]\[9\] _1110_ _1279_ _0972_ VGND VGND VPWR VPWR _1280_ sky130_fd_sc_hd__a211o_1
XFILLER_185_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5431_ net469 net1568 _2424_ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__mux2_1
Xoutput303 net303 VGND VGND VPWR VPWR pwr_ctrl_out[2] sky130_fd_sc_hd__buf_12
XFILLER_145_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput314 net314 VGND VGND VPWR VPWR spimemio_flash_io1_di sky130_fd_sc_hd__buf_12
XFILLER_114_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5362_ net452 net982 _2416_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__mux2_1
Xoutput325 net1896 VGND VGND VPWR VPWR net1897 sky130_fd_sc_hd__buf_12
XFILLER_160_227 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput336 net1886 VGND VGND VPWR VPWR net1887 sky130_fd_sc_hd__buf_12
X_7101_ clknet_leaf_56_csclk net1436 net504 VGND VGND VPWR VPWR gpio_configure\[32\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xoutput347 net1864 VGND VGND VPWR VPWR net1865 sky130_fd_sc_hd__buf_12
X_4313_ net1824 net467 _1544_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__mux2_1
XFILLER_99_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5293_ net439 net650 net565 VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__mux2_1
XFILLER_87_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7032_ clknet_leaf_56_csclk net1416 net504 VGND VGND VPWR VPWR gpio_configure\[23\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_4244_ net1236 net450 _1532_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__mux2_1
XFILLER_101_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4175_ net468 net1751 _1518_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__mux2_1
XFILLER_95_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6816_ clknet_leaf_60_csclk net785 net499 VGND VGND VPWR VPWR serial_bb_data_1 sky130_fd_sc_hd__dfrtp_1
XFILLER_168_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6747_ clknet_leaf_8_csclk net833 net509 VGND VGND VPWR VPWR gpio_configure\[34\]\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_149_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3959_ net36 net1 VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__and2_1
XFILLER_109_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6678_ clknet_leaf_11_csclk net570 net511 VGND VGND VPWR VPWR gpio_configure\[11\]\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_137_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5629_ pad_count_2\[1\] pad_count_2\[0\] VGND VGND VPWR VPWR _2471_ sky130_fd_sc_hd__and2b_4
XFILLER_137_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout530 net121 VGND VGND VPWR VPWR net530 sky130_fd_sc_hd__buf_12
XFILLER_116_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5980_ _2797_ _2801_ VGND VGND VPWR VPWR _2802_ sky130_fd_sc_hd__nor2_8
XFILLER_18_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4931_ _1580_ _1642_ VGND VGND VPWR VPWR _2141_ sky130_fd_sc_hd__nor2_1
XFILLER_32_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4862_ _2062_ _2063_ _2071_ _2072_ VGND VGND VPWR VPWR _2073_ sky130_fd_sc_hd__or4_1
XFILLER_177_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6601_ clknet_leaf_77_csclk net1801 net484 VGND VGND VPWR VPWR gpio_configure\[1\]\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_3813_ hkspi.addr\[5\] hkspi.addr\[4\] _1390_ hkspi.addr\[6\] VGND VGND VPWR VPWR
+ _1394_ sky130_fd_sc_hd__a31o_1
XANTENNA_15 _0950_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 _1004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4793_ _0835_ _1762_ VGND VGND VPWR VPWR _2004_ sky130_fd_sc_hd__or2_1
XFILLER_193_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_37 _1122_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 _1367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6532_ clknet_leaf_69_csclk net1492 net497 VGND VGND VPWR VPWR gpio_configure\[28\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_59 _2498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3744_ gpio_configure\[14\]\[0\] net373 _1080_ gpio_configure\[16\]\[8\] _1329_ VGND
+ VGND VPWR VPWR _1330_ sky130_fd_sc_hd__a221o_1
XFILLER_186_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6463_ clknet_2_2__leaf_mgmt_gpio_in[4] _0085_ _0041_ VGND VGND VPWR VPWR hkspi.addr\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3675_ net273 _1009_ _1262_ net265 VGND VGND VPWR VPWR _1263_ sky130_fd_sc_hd__a22o_1
X_5414_ net464 net1397 _2422_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__mux2_1
XFILLER_161_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6394_ net461 net1516 _3182_ VGND VGND VPWR VPWR _0810_ sky130_fd_sc_hd__mux2_1
X_5345_ net446 net1284 _2414_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__mux2_1
XFILLER_87_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput177 net177 VGND VGND VPWR VPWR mgmt_gpio_oeb[11] sky130_fd_sc_hd__buf_12
Xoutput188 net188 VGND VGND VPWR VPWR mgmt_gpio_oeb[21] sky130_fd_sc_hd__buf_12
XFILLER_102_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5276_ net434 net1100 _2406_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__mux2_1
Xoutput199 net199 VGND VGND VPWR VPWR mgmt_gpio_oeb[31] sky130_fd_sc_hd__buf_12
XFILLER_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7015_ clknet_leaf_32_csclk net1519 net524 VGND VGND VPWR VPWR gpio_configure\[21\]\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_4227_ net446 net1168 net584 VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__mux2_1
XFILLER_56_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4158_ net446 net1091 _1515_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__mux2_1
XFILLER_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4089_ net1759 _1500_ _1499_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__mux2_1
XFILLER_83_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput13 mask_rev_in[18] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
XFILLER_128_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput24 mask_rev_in[28] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_2
XFILLER_168_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput35 mask_rev_in[9] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_2
XFILLER_155_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput46 mgmt_gpio_in[19] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_2
Xinput57 mgmt_gpio_in[29] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_1
Xinput68 mgmt_gpio_in[5] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_4
XFILLER_143_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold808 _0226_ VGND VGND VPWR VPWR net1341 sky130_fd_sc_hd__dlygate4sd3_1
Xinput79 spi_enabled VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_4
XFILLER_6_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold819 gpio_configure\[16\]\[2\] VGND VGND VPWR VPWR net1352 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3460_ net629 _0973_ VGND VGND VPWR VPWR _1051_ sky130_fd_sc_hd__nor2_4
XFILLER_143_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3391_ net9 _0891_ _0923_ gpio_configure\[22\]\[6\] _0979_ VGND VGND VPWR VPWR _0985_
+ sky130_fd_sc_hd__a221o_2
XFILLER_170_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5130_ _1869_ _2110_ _2251_ _2259_ VGND VGND VPWR VPWR _2338_ sky130_fd_sc_hd__or4b_1
XFILLER_35_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1508 serial_data_staging_2\[11\] VGND VGND VPWR VPWR net2041 sky130_fd_sc_hd__dlygate4sd3_1
X_5061_ _2163_ _2269_ VGND VGND VPWR VPWR _2270_ sky130_fd_sc_hd__nor2_1
XFILLER_38_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1519 wbbd_data\[0\] VGND VGND VPWR VPWR net2052 sky130_fd_sc_hd__dlygate4sd3_1
X_4012_ net1467 net462 _1473_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__mux2_1
XFILLER_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5963_ gpio_configure\[19\]\[12\] _2491_ _2517_ gpio_configure\[30\]\[12\] VGND VGND
+ VPWR VPWR _2786_ sky130_fd_sc_hd__a22o_1
X_4914_ _1800_ _1886_ _2123_ _2124_ _1870_ VGND VGND VPWR VPWR _2125_ sky130_fd_sc_hd__o2111a_1
X_5894_ gpio_configure\[16\]\[9\] net472 VGND VGND VPWR VPWR _2720_ sky130_fd_sc_hd__or2_1
XFILLER_80_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4845_ _1643_ _1678_ _1576_ VGND VGND VPWR VPWR _2056_ sky130_fd_sc_hd__a21oi_1
XFILLER_178_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4776_ _1748_ _1935_ _1987_ _1530_ net2005 VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__o32a_1
XFILLER_165_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6515_ clknet_leaf_5_csclk net1094 net494 VGND VGND VPWR VPWR gpio_configure\[30\]\[12\]
+ sky130_fd_sc_hd__dfrtp_2
X_3727_ net390 _0870_ VGND VGND VPWR VPWR _1314_ sky130_fd_sc_hd__nor2_1
XFILLER_174_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6446_ clknet_2_3__leaf_mgmt_gpio_in[4] _0068_ _0024_ VGND VGND VPWR VPWR hkspi.odata\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3658_ _0972_ _1206_ _1245_ _1246_ VGND VGND VPWR VPWR _1247_ sky130_fd_sc_hd__or4_1
XFILLER_161_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6377_ _3172_ net1988 _3162_ VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__mux2_1
X_3589_ net277 _0940_ _1053_ gpio_configure\[20\]\[11\] _1141_ VGND VGND VPWR VPWR
+ _1179_ sky130_fd_sc_hd__a221o_1
XFILLER_88_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5328_ net1528 net440 _2412_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__mux2_1
XFILLER_88_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5259_ _0934_ net647 VGND VGND VPWR VPWR _2405_ sky130_fd_sc_hd__nand2_8
XFILLER_87_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4630_ net432 _1841_ VGND VGND VPWR VPWR _1842_ sky130_fd_sc_hd__or2_2
XFILLER_147_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4561_ net530 _1556_ VGND VGND VPWR VPWR _1773_ sky130_fd_sc_hd__nor2_2
XFILLER_190_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6300_ gpio_configure\[26\]\[11\] _2810_ _2811_ gpio_configure\[7\]\[11\] _3108_
+ VGND VGND VPWR VPWR _3111_ sky130_fd_sc_hd__a221o_1
X_3512_ _0885_ net383 VGND VGND VPWR VPWR _1103_ sky130_fd_sc_hd__nor2_4
XFILLER_116_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold605 gpio_configure\[9\]\[3\] VGND VGND VPWR VPWR net1138 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold616 _0318_ VGND VGND VPWR VPWR net1149 sky130_fd_sc_hd__dlygate4sd3_1
X_4492_ _1588_ _1590_ _1592_ VGND VGND VPWR VPWR _1704_ sky130_fd_sc_hd__or3_1
Xhold627 gpio_configure\[14\]\[3\] VGND VGND VPWR VPWR net1160 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold638 _0585_ VGND VGND VPWR VPWR net1171 sky130_fd_sc_hd__dlygate4sd3_1
X_6231_ gpio_configure\[16\]\[8\] _2831_ _2860_ gpio_configure\[17\]\[8\] _3044_ VGND
+ VGND VPWR VPWR _3045_ sky130_fd_sc_hd__a221o_1
Xhold649 gpio_configure\[20\]\[4\] VGND VGND VPWR VPWR net1182 sky130_fd_sc_hd__dlygate4sd3_1
X_3443_ gpio_configure\[24\]\[5\] _0919_ net350 gpio_configure\[4\]\[5\] VGND VGND
+ VPWR VPWR _1035_ sky130_fd_sc_hd__a22o_1
XFILLER_170_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap368 _0930_ VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__buf_8
Xmax_cap379 net628 VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__buf_12
XFILLER_131_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ gpio_configure\[2\]\[5\] _2823_ net392 gpio_configure\[5\]\[5\] _2978_ VGND
+ VGND VPWR VPWR _2979_ sky130_fd_sc_hd__a221o_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ hkspi.readmode hkspi.state\[2\] VGND VGND VPWR VPWR _0970_ sky130_fd_sc_hd__nand2_4
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5113_ _1646_ _1707_ _1858_ VGND VGND VPWR VPWR _2321_ sky130_fd_sc_hd__o21ai_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ gpio_configure\[23\]\[2\] _2822_ _2910_ _2912_ VGND VGND VPWR VPWR _2913_
+ sky130_fd_sc_hd__a211o_1
XFILLER_112_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1305 net1929 VGND VGND VPWR VPWR net1838 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1316 net1849 VGND VGND VPWR VPWR wb_dat_o[19] sky130_fd_sc_hd__buf_12
Xhold1327 net1943 VGND VGND VPWR VPWR net1860 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _2246_ _2250_ _2251_ _2252_ VGND VGND VPWR VPWR _2253_ sky130_fd_sc_hd__or4_1
Xhold1338 net1871 VGND VGND VPWR VPWR wb_dat_o[27] sky130_fd_sc_hd__buf_12
Xhold1349 net1983 VGND VGND VPWR VPWR net1882 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6995_ clknet_leaf_62_csclk net941 net498 VGND VGND VPWR VPWR gpio_configure\[19\]\[1\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_25_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5946_ gpio_configure\[0\]\[11\] _2526_ _2759_ _2769_ net473 VGND VGND VPWR VPWR
+ _2770_ sky130_fd_sc_hd__o221a_1
XFILLER_40_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5877_ gpio_configure\[21\]\[8\] _2521_ _2534_ gpio_configure\[26\]\[8\] VGND VGND
+ VPWR VPWR _2704_ sky130_fd_sc_hd__a22o_1
XFILLER_139_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4828_ net530 _1631_ _1635_ _1887_ VGND VGND VPWR VPWR _2039_ sky130_fd_sc_hd__a31o_1
XFILLER_193_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4759_ _1598_ _1645_ VGND VGND VPWR VPWR _1971_ sky130_fd_sc_hd__nand2_1
XFILLER_107_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6429_ net493 net481 VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__and2_1
XFILLER_134_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_715 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_707 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold2 net633 VGND VGND VPWR VPWR net535 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_67_659 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5800_ gpio_configure\[24\]\[5\] _2531_ _2535_ gpio_configure\[23\]\[5\] _2626_ VGND
+ VGND VPWR VPWR _2630_ sky130_fd_sc_hd__a221o_1
XFILLER_23_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6780_ clknet_3_6_0_wb_clk_i _0383_ net529 VGND VGND VPWR VPWR wbbd_addr\[4\] sky130_fd_sc_hd__dfrtp_1
X_3992_ _0910_ net425 VGND VGND VPWR VPWR _1471_ sky130_fd_sc_hd__and2_2
X_5731_ net2029 _2564_ net366 VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__mux2_1
XFILLER_176_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5662_ gpio_configure\[14\]\[0\] _2494_ net422 gpio_configure\[5\]\[0\] _2492_ VGND
+ VGND VPWR VPWR _2497_ sky130_fd_sc_hd__a221o_2
XFILLER_175_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4613_ net477 net432 VGND VGND VPWR VPWR _1825_ sky130_fd_sc_hd__or2_2
XFILLER_148_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5593_ xfer_state\[3\] net475 VGND VGND VPWR VPWR _2445_ sky130_fd_sc_hd__nor2_1
XFILLER_129_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4544_ net128 _1554_ VGND VGND VPWR VPWR _1756_ sky130_fd_sc_hd__and2b_4
Xhold402 _0737_ VGND VGND VPWR VPWR net935 sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 net215 VGND VGND VPWR VPWR net946 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold424 _0711_ VGND VGND VPWR VPWR net957 sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 gpio_configure\[27\]\[3\] VGND VGND VPWR VPWR net968 sky130_fd_sc_hd__dlygate4sd3_1
X_4475_ _1683_ _1686_ VGND VGND VPWR VPWR _1687_ sky130_fd_sc_hd__nand2_1
Xhold446 _0512_ VGND VGND VPWR VPWR net979 sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 gpio_configure\[4\]\[3\] VGND VGND VPWR VPWR net990 sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 _0152_ VGND VGND VPWR VPWR net1001 sky130_fd_sc_hd__dlygate4sd3_1
X_6214_ gpio_configure\[31\]\[7\] net423 net415 gpio_configure\[11\]\[7\] VGND VGND
+ VPWR VPWR _3029_ sky130_fd_sc_hd__a22o_1
Xhold479 _0400_ VGND VGND VPWR VPWR net1012 sky130_fd_sc_hd__dlygate4sd3_1
X_3426_ gpio_configure\[0\]\[5\] _0898_ net371 gpio_configure\[26\]\[5\] VGND VGND
+ VPWR VPWR _1018_ sky130_fd_sc_hd__a22o_1
X_7194_ clknet_3_6_0_wb_clk_i _0796_ VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__dfxtp_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6145_ net2039 _2962_ net473 VGND VGND VPWR VPWR _2963_ sky130_fd_sc_hd__mux2_1
X_3357_ gpio_configure\[14\]\[7\] _0916_ _0918_ gpio_configure\[15\]\[7\] _0952_ VGND
+ VGND VPWR VPWR _0953_ sky130_fd_sc_hd__a221o_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1102 _0211_ VGND VGND VPWR VPWR net1635 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1113 gpio_configure\[23\]\[10\] VGND VGND VPWR VPWR net1646 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ gpio_configure\[30\]\[2\] _2799_ net405 gpio_configure\[24\]\[2\] VGND VGND
+ VPWR VPWR _2896_ sky130_fd_sc_hd__a22o_1
Xhold1124 _0559_ VGND VGND VPWR VPWR net1657 sky130_fd_sc_hd__dlygate4sd3_1
X_3288_ net588 net560 VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__and2_4
Xhold1135 gpio_configure\[11\]\[1\] VGND VGND VPWR VPWR net1668 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 _0224_ VGND VGND VPWR VPWR net1679 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5027_ _1788_ _2233_ VGND VGND VPWR VPWR _2237_ sky130_fd_sc_hd__nor2_1
Xhold1157 gpio_configure\[35\]\[8\] VGND VGND VPWR VPWR net1690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1168 _0219_ VGND VGND VPWR VPWR net1701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1179 _0334_ VGND VGND VPWR VPWR net1712 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6978_ clknet_leaf_17_csclk net1609 net512 VGND VGND VPWR VPWR gpio_configure\[17\]\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_186_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_740 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5929_ gpio_configure\[21\]\[11\] _2521_ _2523_ gpio_configure\[2\]\[11\] VGND VGND
+ VPWR VPWR _2753_ sky130_fd_sc_hd__a22o_1
XFILLER_179_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold980 _0426_ VGND VGND VPWR VPWR net1513 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold991 gpio_configure\[4\]\[5\] VGND VGND VPWR VPWR net1524 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_675 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4260_ net826 net465 _1535_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__mux2_1
XFILLER_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3211_ gpio_configure\[23\]\[3\] VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__inv_2
XFILLER_141_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4191_ net1952 _1311_ _1520_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__mux2_1
XFILLER_95_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6901_ clknet_leaf_31_csclk net1179 net523 VGND VGND VPWR VPWR gpio_configure\[7\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_47_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6832_ clknet_leaf_33_csclk net635 net524 VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__dfrtp_1
XFILLER_35_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6763_ clknet_leaf_0_csclk net1974 net487 VGND VGND VPWR VPWR gpio_configure\[21\]\[10\]
+ sky130_fd_sc_hd__dfstp_4
X_3975_ net616 net1925 net668 VGND VGND VPWR VPWR _1466_ sky130_fd_sc_hd__mux2_4
X_5714_ gpio_configure\[30\]\[1\] _2517_ _2518_ gpio_configure\[3\]\[1\] _2547_ VGND
+ VGND VPWR VPWR _2548_ sky130_fd_sc_hd__a221o_1
X_6694_ clknet_3_7_0_wb_clk_i _0002_ net528 VGND VGND VPWR VPWR wbbd_state\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_148_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5645_ xfer_count\[2\] xfer_count\[3\] _2451_ VGND VGND VPWR VPWR _2482_ sky130_fd_sc_hd__or3b_1
XFILLER_148_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5576_ net618 net704 _2440_ VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__mux2_1
XFILLER_156_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold210 _0205_ VGND VGND VPWR VPWR net743 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold221 gpio_configure\[17\]\[10\] VGND VGND VPWR VPWR net754 sky130_fd_sc_hd__dlygate4sd3_1
X_4527_ _1632_ _1657_ _1678_ _1680_ _1737_ VGND VGND VPWR VPWR _1739_ sky130_fd_sc_hd__o221a_1
Xhold232 _0417_ VGND VGND VPWR VPWR net765 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold243 net297 VGND VGND VPWR VPWR net776 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold254 _0341_ VGND VGND VPWR VPWR net787 sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 net2118 VGND VGND VPWR VPWR net798 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold276 _0632_ VGND VGND VPWR VPWR net809 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4458_ _0834_ _1632_ VGND VGND VPWR VPWR _1670_ sky130_fd_sc_hd__nor2_4
Xhold287 gpio_configure\[22\]\[2\] VGND VGND VPWR VPWR net820 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold298 _0325_ VGND VGND VPWR VPWR net831 sky130_fd_sc_hd__dlygate4sd3_1
X_3409_ _0972_ _0990_ _0994_ _1002_ VGND VGND VPWR VPWR _1003_ sky130_fd_sc_hd__or4_1
XFILLER_131_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7177_ clknet_3_3_0_wb_clk_i net2028 net505 VGND VGND VPWR VPWR serial_data_staging_2\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4389_ net111 _1548_ VGND VGND VPWR VPWR _1601_ sky130_fd_sc_hd__nor2_8
XFILLER_131_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6128_ gpio_configure\[23\]\[4\] _2822_ net396 gpio_configure\[20\]\[4\] VGND VGND
+ VPWR VPWR _2946_ sky130_fd_sc_hd__a22o_1
XFILLER_100_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6059_ gpio_configure\[36\]\[1\] net403 net402 gpio_configure\[4\]\[1\] _2871_ VGND
+ VGND VPWR VPWR _2880_ sky130_fd_sc_hd__a221o_1
XFILLER_100_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_105 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_116 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_127 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_149 net269 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_14_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_592 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3760_ _1342_ _1343_ _1344_ _1345_ VGND VGND VPWR VPWR _1346_ sky130_fd_sc_hd__or4_4
XFILLER_158_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3691_ gpio_configure\[7\]\[1\] _0913_ net350 gpio_configure\[4\]\[1\] _1278_ VGND
+ VGND VPWR VPWR _1279_ sky130_fd_sc_hd__a221o_1
XFILLER_185_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5430_ _0928_ net427 VGND VGND VPWR VPWR _2424_ sky130_fd_sc_hd__nand2_8
XFILLER_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput304 net304 VGND VGND VPWR VPWR pwr_ctrl_out[3] sky130_fd_sc_hd__buf_12
XFILLER_161_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5361_ net458 net1578 _2416_ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__mux2_1
XFILLER_114_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput315 net315 VGND VGND VPWR VPWR spimemio_flash_io2_di sky130_fd_sc_hd__buf_12
XFILLER_99_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput326 net1846 VGND VGND VPWR VPWR net1847 sky130_fd_sc_hd__buf_12
XFILLER_114_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput337 net1870 VGND VGND VPWR VPWR net1871 sky130_fd_sc_hd__buf_12
X_4312_ _1127_ net426 VGND VGND VPWR VPWR _1544_ sky130_fd_sc_hd__and2_2
X_7100_ clknet_leaf_58_csclk net795 net503 VGND VGND VPWR VPWR gpio_configure\[32\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_160_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput348 net1868 VGND VGND VPWR VPWR net1869 sky130_fd_sc_hd__buf_12
XFILLER_113_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5292_ net440 net1524 net565 VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__mux2_1
X_7031_ clknet_leaf_44_csclk net1207 net526 VGND VGND VPWR VPWR gpio_configure\[23\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_4243_ net1322 net456 _1532_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__mux2_1
XFILLER_87_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4174_ _1042_ net426 VGND VGND VPWR VPWR _1518_ sky130_fd_sc_hd__nand2_2
XFILLER_28_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6815_ clknet_leaf_60_csclk net817 net499 VGND VGND VPWR VPWR serial_bb_resetn sky130_fd_sc_hd__dfrtp_1
XFILLER_51_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6746_ clknet_leaf_19_csclk net1649 net510 VGND VGND VPWR VPWR gpio_configure\[34\]\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_3958_ net63 net79 VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__and2_1
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6677_ clknet_leaf_11_csclk net585 net511 VGND VGND VPWR VPWR gpio_configure\[11\]\[10\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_137_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3889_ wbbd_state\[5\] _1428_ net431 net2139 VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__a22o_1
XFILLER_149_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5628_ xfer_state\[2\] pad_count_2\[1\] pad_count_2\[0\] VGND VGND VPWR VPWR _2470_
+ sky130_fd_sc_hd__and3_1
XFILLER_164_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5559_ net440 net1526 _2438_ VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__mux2_1
XFILLER_191_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout520 net521 VGND VGND VPWR VPWR net520 sky130_fd_sc_hd__buf_8
XFILLER_59_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_1_0_wb_clk_i clknet_2_0_0_wb_clk_i VGND VGND VPWR VPWR clknet_3_1_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XFILLER_27_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4930_ _1582_ _1746_ _2056_ VGND VGND VPWR VPWR _2140_ sky130_fd_sc_hd__or3_1
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4861_ _1833_ _1863_ _1660_ VGND VGND VPWR VPWR _2072_ sky130_fd_sc_hd__o21ai_1
XTAP_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6600_ clknet_leaf_73_csclk net997 net489 VGND VGND VPWR VPWR gpio_configure\[0\]\[12\]
+ sky130_fd_sc_hd__dfstp_2
X_3812_ _1388_ _1393_ _1392_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__o21ai_1
XANTENNA_16 _0950_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4792_ _1752_ _1764_ _1765_ VGND VGND VPWR VPWR _2003_ sky130_fd_sc_hd__or3_1
XFILLER_193_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_27 _1039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_38 _1130_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6531_ clknet_leaf_69_csclk net1786 net497 VGND VGND VPWR VPWR gpio_configure\[28\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_49 _1510_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3743_ gpio_configure\[12\]\[8\] _1056_ _1129_ gpio_configure\[11\]\[8\] VGND VGND
+ VPWR VPWR _1329_ sky130_fd_sc_hd__a22o_1
XFILLER_118_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3674_ net389 net601 VGND VGND VPWR VPWR _1262_ sky130_fd_sc_hd__nor2_2
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6462_ clknet_2_0__leaf_mgmt_gpio_in[4] _0084_ _0040_ VGND VGND VPWR VPWR hkspi.pass_thru_user_delay
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_146_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5413_ net467 net1781 _2422_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__mux2_1
XFILLER_146_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6393_ net466 net1502 _3182_ VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__mux2_1
X_5344_ net569 net728 _2414_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__mux2_1
XFILLER_161_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput178 net178 VGND VGND VPWR VPWR mgmt_gpio_oeb[12] sky130_fd_sc_hd__buf_12
Xoutput189 net189 VGND VGND VPWR VPWR mgmt_gpio_oeb[22] sky130_fd_sc_hd__buf_12
X_5275_ net437 net1375 _2406_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__mux2_1
XFILLER_87_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4226_ net569 net1917 net584 VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__mux2_1
X_7014_ clknet_leaf_27_csclk net1241 net519 VGND VGND VPWR VPWR gpio_configure\[21\]\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4157_ net569 net702 _1515_ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__mux2_1
XFILLER_46_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4088_ net1451 net471 net354 VGND VGND VPWR VPWR _1500_ sky130_fd_sc_hd__mux2_1
XFILLER_43_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6729_ clknet_leaf_18_csclk net719 net512 VGND VGND VPWR VPWR gpio_configure\[36\]\[11\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_177_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_52_csclk clknet_3_3_0_csclk VGND VGND VPWR VPWR clknet_leaf_52_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_124_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_67_csclk clknet_3_3_0_csclk VGND VGND VPWR VPWR clknet_leaf_67_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_132_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput14 mask_rev_in[19] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_1
Xinput25 mask_rev_in[29] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_1
Xinput36 mgmt_gpio_in[0] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_4
Xinput47 mgmt_gpio_in[1] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_2
XFILLER_6_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput58 mgmt_gpio_in[2] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_12
Xinput69 mgmt_gpio_in[6] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_1
XFILLER_182_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold809 gpio_configure\[9\]\[6\] VGND VGND VPWR VPWR net1342 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3390_ gpio_configure\[7\]\[6\] _0913_ net354 net41 _0983_ VGND VGND VPWR VPWR _0984_
+ sky130_fd_sc_hd__a221o_1
XFILLER_123_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5060_ _1686_ _2152_ VGND VGND VPWR VPWR _2269_ sky130_fd_sc_hd__and2_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1509 serial_data_staging_2\[5\] VGND VGND VPWR VPWR net2042 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4011_ net1830 net467 _1473_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__mux2_1
XFILLER_77_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5962_ gpio_configure\[13\]\[12\] _2501_ _2510_ gpio_configure\[15\]\[12\] _2784_
+ VGND VGND VPWR VPWR _2785_ sky130_fd_sc_hd__a221o_1
XFILLER_18_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4913_ _1611_ _1693_ _1805_ _1684_ VGND VGND VPWR VPWR _2124_ sky130_fd_sc_hd__o22a_1
X_5893_ gpio_configure\[9\]\[9\] _2512_ _2538_ gpio_configure\[1\]\[9\] _2718_ VGND
+ VGND VPWR VPWR _2719_ sky130_fd_sc_hd__a221o_1
X_4844_ _1704_ _1929_ VGND VGND VPWR VPWR _2055_ sky130_fd_sc_hd__nand2_1
XFILLER_178_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4775_ _1930_ _1957_ _1985_ _1986_ _1939_ VGND VGND VPWR VPWR _1987_ sky130_fd_sc_hd__o41a_1
XFILLER_193_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6514_ clknet_leaf_5_csclk net1151 net494 VGND VGND VPWR VPWR gpio_configure\[30\]\[11\]
+ sky130_fd_sc_hd__dfrtp_2
X_3726_ net629 _0885_ VGND VGND VPWR VPWR _1313_ sky130_fd_sc_hd__nor2_1
XFILLER_119_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6445_ clknet_2_1__leaf_mgmt_gpio_in[4] _0067_ _0023_ VGND VGND VPWR VPWR hkspi.pre_pass_thru_mgmt
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_161_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3657_ net389 _1008_ _1103_ gpio_configure\[1\]\[10\] VGND VGND VPWR VPWR _1246_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_174_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3588_ _1174_ _1175_ _1176_ _1177_ VGND VGND VPWR VPWR _1178_ sky130_fd_sc_hd__or4_1
X_6376_ wbbd_state\[9\] net152 net135 wbbd_state\[8\] _3171_ VGND VGND VPWR VPWR _3172_
+ sky130_fd_sc_hd__a221o_1
XFILLER_88_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5327_ net1166 net446 _2412_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__mux2_1
XFILLER_142_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5258_ net1128 net434 _2404_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__mux2_1
XFILLER_75_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4209_ net994 net443 _1522_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__mux2_1
X_5189_ net461 net1706 _2390_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__mux2_1
XFILLER_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4560_ _1604_ _1758_ VGND VGND VPWR VPWR _1772_ sky130_fd_sc_hd__nand2_2
XFILLER_128_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3511_ _0903_ net382 VGND VGND VPWR VPWR _1102_ sky130_fd_sc_hd__nor2_8
X_4491_ _1613_ _1643_ VGND VGND VPWR VPWR _1703_ sky130_fd_sc_hd__nand2_1
Xhold606 _0520_ VGND VGND VPWR VPWR net1139 sky130_fd_sc_hd__dlygate4sd3_1
Xhold617 gpio_configure\[30\]\[11\] VGND VGND VPWR VPWR net1150 sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 _0560_ VGND VGND VPWR VPWR net1161 sky130_fd_sc_hd__dlygate4sd3_1
X_6230_ gpio_configure\[14\]\[8\] net411 _2855_ gpio_configure\[27\]\[8\] VGND VGND
+ VPWR VPWR _3044_ sky130_fd_sc_hd__a22o_1
X_3442_ gpio_configure\[9\]\[5\] net368 _1009_ net263 _1033_ VGND VGND VPWR VPWR _1034_
+ sky130_fd_sc_hd__a221o_1
Xhold639 gpio_configure\[25\]\[4\] VGND VGND VPWR VPWR net1172 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap358 _0874_ VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__buf_6
XFILLER_171_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap369 net610 VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__buf_12
XFILLER_170_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3373_ _0951_ _0957_ _0968_ VGND VGND VPWR VPWR _0969_ sky130_fd_sc_hd__or3_4
XFILLER_69_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6161_ gpio_configure\[13\]\[5\] net417 net404 gpio_configure\[25\]\[5\] VGND VGND
+ VPWR VPWR _2978_ sky130_fd_sc_hd__a22o_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_170_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5112_ _1586_ _2173_ _2222_ _2306_ VGND VGND VPWR VPWR _2320_ sky130_fd_sc_hd__or4_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6092_ gpio_configure\[37\]\[2\] net400 net416 gpio_configure\[32\]\[2\] _2911_ VGND
+ VGND VPWR VPWR _2912_ sky130_fd_sc_hd__a221o_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1306 net1839 VGND VGND VPWR VPWR wb_dat_o[22] sky130_fd_sc_hd__buf_12
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1317 net1937 VGND VGND VPWR VPWR net1850 sky130_fd_sc_hd__dlygate4sd3_1
X_5043_ _1596_ _1650_ _1718_ _1966_ _2205_ VGND VGND VPWR VPWR _2252_ sky130_fd_sc_hd__a2111o_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1328 net1861 VGND VGND VPWR VPWR wb_dat_o[12] sky130_fd_sc_hd__buf_12
XFILLER_84_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1339 net1948 VGND VGND VPWR VPWR net1872 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_wbbd_sck wbbd_sck VGND VGND VPWR VPWR clknet_0_wbbd_sck sky130_fd_sc_hd__clkbuf_16
X_6994_ clknet_leaf_62_csclk net1725 net498 VGND VGND VPWR VPWR gpio_configure\[19\]\[0\]
+ sky130_fd_sc_hd__dfstp_4
XFILLER_80_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_41_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5945_ _2761_ _2764_ _2766_ _2768_ VGND VGND VPWR VPWR _2769_ sky130_fd_sc_hd__or4_1
XFILLER_43_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5876_ gpio_configure\[5\]\[8\] _2496_ _2513_ gpio_configure\[28\]\[8\] _2702_ VGND
+ VGND VPWR VPWR _2703_ sky130_fd_sc_hd__a221o_1
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4827_ _1678_ _1836_ _1721_ VGND VGND VPWR VPWR _2038_ sky130_fd_sc_hd__o21ai_1
XFILLER_178_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4758_ _1617_ _1628_ _1633_ _1749_ VGND VGND VPWR VPWR _1970_ sky130_fd_sc_hd__nand4_2
XFILLER_193_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3709_ gpio_configure\[9\]\[1\] net368 net351 net47 _1296_ VGND VGND VPWR VPWR _1297_
+ sky130_fd_sc_hd__a221o_1
X_4689_ _1588_ _1850_ VGND VGND VPWR VPWR _1901_ sky130_fd_sc_hd__or2_1
XFILLER_162_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6428_ net492 net481 VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__and2_1
XFILLER_162_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6359_ wbbd_state\[9\] _3157_ _3158_ wbbd_state\[7\] VGND VGND VPWR VPWR _3159_ sky130_fd_sc_hd__a22o_1
XFILLER_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold3 _0515_ VGND VGND VPWR VPWR net536 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_35_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3991_ net1968 net434 _1470_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__mux2_1
X_5730_ net475 serial_data_staging_1\[0\] _2563_ VGND VGND VPWR VPWR _2564_ sky130_fd_sc_hd__a21o_1
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5661_ net472 _2488_ _2495_ VGND VGND VPWR VPWR _2496_ sky130_fd_sc_hd__and3_4
XFILLER_176_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4612_ _1795_ _1797_ VGND VGND VPWR VPWR _1824_ sky130_fd_sc_hd__or2_1
XFILLER_176_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5592_ net475 net307 VGND VGND VPWR VPWR _2444_ sky130_fd_sc_hd__nand2_2
XFILLER_191_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4543_ net128 net127 VGND VGND VPWR VPWR _1755_ sky130_fd_sc_hd__nand2b_1
XFILLER_7_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold403 net246 VGND VGND VPWR VPWR net936 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold414 _0182_ VGND VGND VPWR VPWR net947 sky130_fd_sc_hd__dlygate4sd3_1
Xhold425 net221 VGND VGND VPWR VPWR net958 sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 _0664_ VGND VGND VPWR VPWR net969 sky130_fd_sc_hd__dlygate4sd3_1
X_4474_ _1564_ _1685_ VGND VGND VPWR VPWR _1686_ sky130_fd_sc_hd__nor2_4
Xhold447 gpio_configure\[37\]\[3\] VGND VGND VPWR VPWR net980 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold458 _0480_ VGND VGND VPWR VPWR net991 sky130_fd_sc_hd__dlygate4sd3_1
X_6213_ gpio_configure\[2\]\[7\] _2823_ net392 gpio_configure\[5\]\[7\] _3027_ VGND
+ VGND VPWR VPWR _3028_ sky130_fd_sc_hd__a221o_1
XFILLER_143_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold469 wbbd_data\[7\] VGND VGND VPWR VPWR net1002 sky130_fd_sc_hd__dlygate4sd3_1
X_3425_ net17 _0864_ _0910_ net296 VGND VGND VPWR VPWR _1017_ sky130_fd_sc_hd__a22o_2
X_7193_ clknet_3_4_0_wb_clk_i _0795_ VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__dfxtp_2
XFILLER_131_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3356_ gpio_configure\[23\]\[7\] net372 _0936_ net28 VGND VGND VPWR VPWR _0952_ sky130_fd_sc_hd__a22o_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6144_ _2945_ _2951_ _2961_ _2851_ gpio_configure\[0\]\[4\] VGND VGND VPWR VPWR _2962_
+ sky130_fd_sc_hd__o32a_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1103 gpio_configure\[24\]\[10\] VGND VGND VPWR VPWR net1636 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1114 _0130_ VGND VGND VPWR VPWR net1647 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3287_ net387 _0881_ VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__nor2_4
X_6075_ gpio_configure\[36\]\[2\] net403 net402 gpio_configure\[4\]\[2\] _2894_ VGND
+ VGND VPWR VPWR _2895_ sky130_fd_sc_hd__a221o_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1125 gpio_configure\[4\]\[2\] VGND VGND VPWR VPWR net1658 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1136 _0534_ VGND VGND VPWR VPWR net1669 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1147 gpio_configure\[33\]\[2\] VGND VGND VPWR VPWR net1680 sky130_fd_sc_hd__dlygate4sd3_1
X_5026_ _1798_ _1807_ _1836_ _2233_ VGND VGND VPWR VPWR _2236_ sky130_fd_sc_hd__a31o_1
Xhold1158 _0339_ VGND VGND VPWR VPWR net1691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1169 gpio_configure\[22\]\[10\] VGND VGND VPWR VPWR net1702 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6977_ clknet_leaf_53_csclk net1072 net507 VGND VGND VPWR VPWR gpio_configure\[16\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_53_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5928_ gpio_configure\[19\]\[11\] _2491_ _2513_ gpio_configure\[28\]\[11\] _2751_
+ VGND VGND VPWR VPWR _2752_ sky130_fd_sc_hd__a221o_1
XFILLER_22_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5859_ net475 serial_data_staging_1\[6\] _2686_ VGND VGND VPWR VPWR _2687_ sky130_fd_sc_hd__a21o_1
XFILLER_186_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold970 _0809_ VGND VGND VPWR VPWR net1503 sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 gpio_configure\[27\]\[10\] VGND VGND VPWR VPWR net1514 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_134_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold992 _0482_ VGND VGND VPWR VPWR net1525 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3210_ gpio_configure\[24\]\[3\] VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__inv_2
XFILLER_141_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4190_ net1954 _1376_ _1520_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__mux2_1
XFILLER_140_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_671 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6900_ clknet_leaf_24_csclk net1677 net518 VGND VGND VPWR VPWR gpio_configure\[7\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_63_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6831_ clknet_leaf_33_csclk net945 net524 VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__dfrtp_1
XFILLER_23_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6762_ clknet_leaf_0_csclk net1735 net486 VGND VGND VPWR VPWR gpio_configure\[21\]\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3974_ net1061 net449 _1461_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__mux2_1
XFILLER_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5713_ gpio_configure\[18\]\[1\] _2532_ _2537_ gpio_configure\[17\]\[1\] VGND VGND
+ VPWR VPWR _2547_ sky130_fd_sc_hd__a22o_1
XFILLER_176_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6693_ clknet_3_7_0_wb_clk_i _0001_ net528 VGND VGND VPWR VPWR wbbd_state\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_148_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5644_ xfer_state\[2\] _2480_ _2481_ pad_count_2\[5\] VGND VGND VPWR VPWR _0761_
+ sky130_fd_sc_hd__a22o_1
XFILLER_164_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5575_ net452 net1224 _2440_ VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__mux2_1
Xhold200 _0496_ VGND VGND VPWR VPWR net733 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_191_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold211 gpio_configure\[37\]\[10\] VGND VGND VPWR VPWR net744 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4526_ _1657_ _1671_ VGND VGND VPWR VPWR _1738_ sky130_fd_sc_hd__nor2_1
XFILLER_191_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold222 _0326_ VGND VGND VPWR VPWR net755 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold233 gpio_configure\[16\]\[10\] VGND VGND VPWR VPWR net766 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 _0118_ VGND VGND VPWR VPWR net777 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 gpio_configure\[34\]\[4\] VGND VGND VPWR VPWR net788 sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 _0700_ VGND VGND VPWR VPWR net799 sky130_fd_sc_hd__dlygate4sd3_1
X_4457_ _1645_ _1662_ VGND VGND VPWR VPWR _1669_ sky130_fd_sc_hd__nand2_1
XFILLER_171_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold277 gpio_configure\[24\]\[3\] VGND VGND VPWR VPWR net810 sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 _0623_ VGND VGND VPWR VPWR net821 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_132_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold299 gpio_configure\[34\]\[9\] VGND VGND VPWR VPWR net832 sky130_fd_sc_hd__dlygate4sd3_1
X_3408_ _0996_ _0998_ _0999_ _1001_ VGND VGND VPWR VPWR _1002_ sky130_fd_sc_hd__or4_1
X_7176_ clknet_3_3_0_wb_clk_i _0778_ net505 VGND VGND VPWR VPWR serial_data_staging_2\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_172_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4388_ net112 net111 VGND VGND VPWR VPWR _1600_ sky130_fd_sc_hd__nor2_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6127_ gpio_configure\[29\]\[4\] _2816_ _2820_ gpio_configure\[21\]\[4\] _2943_ VGND
+ VGND VPWR VPWR _2945_ sky130_fd_sc_hd__a221o_2
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ net376 net562 VGND VGND VPWR VPWR _0935_ sky130_fd_sc_hd__nor2_4
XFILLER_85_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6058_ _2873_ _2874_ _2876_ _2878_ VGND VGND VPWR VPWR _2879_ sky130_fd_sc_hd__or4_1
XFILLER_39_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5009_ _2207_ _2208_ _2212_ _2218_ VGND VGND VPWR VPWR _2219_ sky130_fd_sc_hd__or4_1
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_106 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_117 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_128 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_139 net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_666 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3690_ gpio_configure\[33\]\[1\] _0938_ _1109_ gpio_configure\[36\]\[9\] VGND VGND
+ VPWR VPWR _1278_ sky130_fd_sc_hd__a22o_1
XFILLER_187_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput305 net305 VGND VGND VPWR VPWR reset sky130_fd_sc_hd__buf_12
X_5360_ net464 net1437 _2416_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__mux2_1
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput316 net316 VGND VGND VPWR VPWR spimemio_flash_io3_di sky130_fd_sc_hd__buf_12
Xoutput327 net1890 VGND VGND VPWR VPWR net1891 sky130_fd_sc_hd__buf_12
X_4311_ net444 net1300 _1543_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__mux2_1
XFILLER_99_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput338 net1882 VGND VGND VPWR VPWR net1883 sky130_fd_sc_hd__buf_12
Xoutput349 net1866 VGND VGND VPWR VPWR net1867 sky130_fd_sc_hd__buf_12
XFILLER_126_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5291_ net618 net722 net565 VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__mux2_1
XFILLER_114_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7030_ clknet_leaf_21_csclk net1157 net514 VGND VGND VPWR VPWR gpio_configure\[23\]\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_4242_ net1441 net462 _1532_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__mux2_1
XFILLER_141_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4173_ net2026 _0969_ _1517_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__mux2_1
XFILLER_95_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6814_ clknet_leaf_60_csclk net765 net499 VGND VGND VPWR VPWR serial_bb_load sky130_fd_sc_hd__dfrtp_2
XFILLER_51_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6745_ clknet_leaf_75_csclk net1014 net485 VGND VGND VPWR VPWR gpio_configure\[19\]\[12\]
+ sky130_fd_sc_hd__dfrtp_4
X_3957_ net68 net94 VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__and2_1
XFILLER_176_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6676_ clknet_leaf_11_csclk net621 net511 VGND VGND VPWR VPWR gpio_configure\[11\]\[9\]
+ sky130_fd_sc_hd__dfrtp_4
X_3888_ net2139 net431 VGND VGND VPWR VPWR _1440_ sky130_fd_sc_hd__nand2_1
XFILLER_176_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5627_ pad_count_2\[1\] pad_count_2\[0\] VGND VGND VPWR VPWR _2469_ sky130_fd_sc_hd__and2_2
XFILLER_136_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5558_ net445 net788 _2438_ VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__mux2_1
XFILLER_3_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4509_ _1654_ _1670_ VGND VGND VPWR VPWR _1721_ sky130_fd_sc_hd__nand2_1
XFILLER_132_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5489_ net446 net1234 _2430_ VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__mux2_1
XFILLER_160_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout510 net511 VGND VGND VPWR VPWR net510 sky130_fd_sc_hd__buf_6
XFILLER_104_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout521 net526 VGND VGND VPWR VPWR net521 sky130_fd_sc_hd__buf_6
X_7159_ clknet_3_2_0_wb_clk_i net531 net499 VGND VGND VPWR VPWR serial_resetn_pre
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_58_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4860_ _1672_ _1896_ _2064_ _2070_ VGND VGND VPWR VPWR _2071_ sky130_fd_sc_hd__nand4_1
XTAP_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3811_ _0838_ _0839_ _1391_ VGND VGND VPWR VPWR _1393_ sky130_fd_sc_hd__mux2_1
XFILLER_32_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4791_ _1653_ _1745_ net424 _1788_ VGND VGND VPWR VPWR _2002_ sky130_fd_sc_hd__o22ai_1
XANTENNA_17 _0969_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_28 _1054_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6530_ clknet_leaf_76_csclk net1001 net488 VGND VGND VPWR VPWR gpio_configure\[25\]\[12\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA_39 _1140_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3742_ gpio_configure\[5\]\[0\] net355 _0934_ gpio_configure\[1\]\[0\] _1327_ VGND
+ VGND VPWR VPWR _1328_ sky130_fd_sc_hd__a221o_1
XFILLER_158_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6461_ clknet_2_1__leaf_mgmt_gpio_in[4] _0083_ _0039_ VGND VGND VPWR VPWR hkspi.pass_thru_user
+ sky130_fd_sc_hd__dfrtp_4
X_3673_ gpio_configure\[14\]\[1\] net373 _1121_ gpio_configure\[17\]\[9\] _1260_ VGND
+ VGND VPWR VPWR _1261_ sky130_fd_sc_hd__a221o_1
XFILLER_173_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_568 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5412_ net374 net427 VGND VGND VPWR VPWR _2422_ sky130_fd_sc_hd__nand2_8
XFILLER_161_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6392_ _1076_ net425 VGND VGND VPWR VPWR _3182_ sky130_fd_sc_hd__nand2_2
XFILLER_173_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5343_ net458 net1586 _2414_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__mux2_1
XFILLER_142_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput179 net179 VGND VGND VPWR VPWR mgmt_gpio_oeb[13] sky130_fd_sc_hd__buf_12
X_5274_ net441 net1122 _2406_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__mux2_1
XFILLER_87_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7013_ clknet_leaf_28_csclk net963 net521 VGND VGND VPWR VPWR gpio_configure\[21\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_4225_ net577 net1932 net584 VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__mux2_1
X_4156_ net577 net752 _1515_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__mux2_1
XFILLER_56_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4087_ _0881_ net483 _1480_ _0929_ net429 VGND VGND VPWR VPWR _1499_ sky130_fd_sc_hd__o221a_4
XFILLER_24_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_655 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4989_ _2190_ _2192_ _2193_ _2198_ VGND VGND VPWR VPWR _2199_ sky130_fd_sc_hd__and4bb_1
X_6728_ clknet_leaf_17_csclk net837 net512 VGND VGND VPWR VPWR gpio_configure\[36\]\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_137_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6659_ clknet_leaf_4_csclk net899 net494 VGND VGND VPWR VPWR gpio_configure\[7\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_109_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput15 mask_rev_in[1] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput26 mask_rev_in[2] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_167_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput37 mgmt_gpio_in[10] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_2
Xinput48 mgmt_gpio_in[20] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput59 mgmt_gpio_in[30] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_2
XFILLER_128_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4010_ _1067_ net426 VGND VGND VPWR VPWR _1473_ sky130_fd_sc_hd__and2_2
XFILLER_37_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5961_ gpio_configure\[26\]\[12\] _2534_ _2783_ _2524_ VGND VGND VPWR VPWR _2784_
+ sky130_fd_sc_hd__a22o_1
X_4912_ _1776_ _1886_ _2121_ _2122_ _1858_ VGND VGND VPWR VPWR _2123_ sky130_fd_sc_hd__o2111a_1
X_5892_ gpio_configure\[10\]\[9\] net421 _2528_ gpio_configure\[7\]\[9\] VGND VGND
+ VPWR VPWR _2718_ sky130_fd_sc_hd__a22o_1
XFILLER_21_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4843_ _1738_ _2043_ VGND VGND VPWR VPWR _2054_ sky130_fd_sc_hd__or2_1
X_4774_ _1929_ _1933_ VGND VGND VPWR VPWR _1986_ sky130_fd_sc_hd__nand2_1
XFILLER_193_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6513_ clknet_leaf_1_csclk net1404 net493 VGND VGND VPWR VPWR gpio_configure\[30\]\[10\]
+ sky130_fd_sc_hd__dfstp_1
X_3725_ _1312_ net1999 _0970_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__mux2_1
XFILLER_146_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6444_ clknet_2_1__leaf_mgmt_gpio_in[4] _0066_ _0022_ VGND VGND VPWR VPWR hkspi.pre_pass_thru_user
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3656_ gpio_configure\[23\]\[10\] _1067_ _1073_ gpio_configure\[24\]\[10\] _1244_
+ VGND VGND VPWR VPWR _1245_ sky130_fd_sc_hd__a221o_1
XFILLER_146_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6375_ wbbd_state\[7\] net144 net158 net433 VGND VGND VPWR VPWR _3171_ sky130_fd_sc_hd__a22o_1
XFILLER_161_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3587_ gpio_configure\[30\]\[11\] _1083_ _1117_ net269 _1140_ VGND VGND VPWR VPWR
+ _1177_ sky130_fd_sc_hd__a221o_1
X_5326_ net978 net452 _2412_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__mux2_1
XFILLER_130_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5257_ net1334 net437 _2404_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__mux2_1
XFILLER_88_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4208_ net1027 net449 _1522_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__mux2_1
XFILLER_75_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5188_ net466 net1744 _2390_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__mux2_1
XFILLER_56_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4139_ net1079 net449 _1512_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__mux2_1
XFILLER_56_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3510_ net387 _0909_ VGND VGND VPWR VPWR _1101_ sky130_fd_sc_hd__nor2_4
XFILLER_128_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4490_ _1657_ _1663_ VGND VGND VPWR VPWR _1702_ sky130_fd_sc_hd__or2_2
Xhold607 gpio_configure\[15\]\[3\] VGND VGND VPWR VPWR net1140 sky130_fd_sc_hd__dlygate4sd3_1
Xhold618 _0136_ VGND VGND VPWR VPWR net1151 sky130_fd_sc_hd__dlygate4sd3_1
Xhold629 gpio_configure\[36\]\[12\] VGND VGND VPWR VPWR net1162 sky130_fd_sc_hd__dlygate4sd3_1
X_3441_ gpio_configure\[15\]\[5\] _0918_ _0928_ gpio_configure\[20\]\[5\] VGND VGND
+ VPWR VPWR _1033_ sky130_fd_sc_hd__a22o_1
XFILLER_143_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6160_ gpio_configure\[10\]\[5\] _2825_ net394 gpio_configure\[6\]\[5\] _2976_ VGND
+ VGND VPWR VPWR _2977_ sky130_fd_sc_hd__a221o_1
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3372_ _0960_ _0967_ VGND VGND VPWR VPWR _0968_ sky130_fd_sc_hd__or2_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5111_ wbbd_addr\[4\] _1529_ _2279_ _2318_ VGND VGND VPWR VPWR _2319_ sky130_fd_sc_hd__a22o_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ gpio_configure\[29\]\[2\] _2816_ net412 gpio_configure\[9\]\[2\] VGND VGND
+ VPWR VPWR _2911_ sky130_fd_sc_hd__a22o_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1307 net1930 VGND VGND VPWR VPWR net1840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1318 net1851 VGND VGND VPWR VPWR wb_dat_o[30] sky130_fd_sc_hd__buf_12
X_5042_ _1950_ _1951_ _2211_ VGND VGND VPWR VPWR _2251_ sky130_fd_sc_hd__or3_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1329 net1942 VGND VGND VPWR VPWR net1862 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6993_ clknet_leaf_59_csclk net1315 net502 VGND VGND VPWR VPWR gpio_configure\[18\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_51_csclk clknet_3_3_0_csclk VGND VGND VPWR VPWR clknet_leaf_51_csclk
+ sky130_fd_sc_hd__clkbuf_16
X_5944_ gpio_configure\[22\]\[11\] _2498_ _2505_ gpio_configure\[11\]\[11\] _2767_
+ VGND VGND VPWR VPWR _2768_ sky130_fd_sc_hd__a221o_1
XFILLER_80_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5875_ gpio_configure\[23\]\[8\] _2535_ _2540_ gpio_configure\[12\]\[8\] VGND VGND
+ VPWR VPWR _2702_ sky130_fd_sc_hd__a22o_1
XFILLER_61_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4826_ _1787_ _1863_ _1724_ VGND VGND VPWR VPWR _2037_ sky130_fd_sc_hd__o21ai_1
XFILLER_21_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4757_ _1599_ _1707_ _1636_ VGND VGND VPWR VPWR _1969_ sky130_fd_sc_hd__a21oi_1
XFILLER_181_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3708_ gpio_configure\[34\]\[1\] _0874_ _1068_ gpio_configure\[10\]\[9\] VGND VGND
+ VPWR VPWR _1296_ sky130_fd_sc_hd__a22o_1
XFILLER_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4688_ _1592_ _1779_ _1866_ VGND VGND VPWR VPWR _1900_ sky130_fd_sc_hd__or3_1
XFILLER_107_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6427_ net492 net481 VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__and2_1
XFILLER_146_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3639_ gpio_configure\[25\]\[2\] _0927_ _0974_ serial_bb_resetn _1227_ VGND VGND
+ VPWR VPWR _1228_ sky130_fd_sc_hd__a221o_1
XFILLER_161_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6358_ net170 net167 VGND VGND VPWR VPWR _3158_ sky130_fd_sc_hd__nand2_1
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5309_ net447 net1196 _2410_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__mux2_1
XFILLER_191_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6289_ gpio_configure\[26\]\[10\] _2810_ _2811_ gpio_configure\[7\]\[10\] VGND VGND
+ VPWR VPWR _3101_ sky130_fd_sc_hd__a22o_1
XFILLER_102_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_19_csclk clknet_3_4_0_csclk VGND VGND VPWR VPWR clknet_leaf_19_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_140_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_1__f__1134_ clknet_0__1134_ VGND VGND VPWR VPWR clknet_1_1__leaf__1134_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_138_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold4 net1912 VGND VGND VPWR VPWR net537 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_81_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3990_ net790 net439 _1470_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__mux2_1
XFILLER_62_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5660_ pad_count_1\[1\] pad_count_1\[0\] VGND VGND VPWR VPWR _2495_ sky130_fd_sc_hd__and2b_2
XFILLER_31_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4611_ net477 _1822_ VGND VGND VPWR VPWR _1823_ sky130_fd_sc_hd__or2_2
X_5591_ net475 xfer_state\[2\] VGND VGND VPWR VPWR _2443_ sky130_fd_sc_hd__nor2_1
XFILLER_129_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4542_ _1560_ _1752_ VGND VGND VPWR VPWR _1754_ sky130_fd_sc_hd__nand2_1
Xhold404 _0176_ VGND VGND VPWR VPWR net937 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire390 _0851_ VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__clkbuf_16
XFILLER_128_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold415 gpio_configure\[30\]\[7\] VGND VGND VPWR VPWR net948 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold426 _0164_ VGND VGND VPWR VPWR net959 sky130_fd_sc_hd__dlygate4sd3_1
X_4473_ _1568_ _1638_ VGND VGND VPWR VPWR _1685_ sky130_fd_sc_hd__or2_2
Xhold437 gpio_configure\[33\]\[3\] VGND VGND VPWR VPWR net970 sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 _0741_ VGND VGND VPWR VPWR net981 sky130_fd_sc_hd__dlygate4sd3_1
Xhold459 gpio_configure\[22\]\[11\] VGND VGND VPWR VPWR net992 sky130_fd_sc_hd__dlygate4sd3_1
X_6212_ gpio_configure\[13\]\[7\] net417 net404 gpio_configure\[25\]\[7\] VGND VGND
+ VPWR VPWR _3027_ sky130_fd_sc_hd__a22o_1
X_3424_ net40 net354 _0939_ gpio_configure\[8\]\[5\] VGND VGND VPWR VPWR _1016_ sky130_fd_sc_hd__a22o_1
X_7192_ clknet_3_5_0_wb_clk_i _0794_ VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__dfxtp_1
X_6143_ net359 _2953_ _2960_ VGND VGND VPWR VPWR _2961_ sky130_fd_sc_hd__or3_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3355_ _0944_ _0946_ _0948_ _0950_ VGND VGND VPWR VPWR _0951_ sky130_fd_sc_hd__or4_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1104 _0140_ VGND VGND VPWR VPWR net1637 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ gpio_configure\[22\]\[2\] net397 _2825_ gpio_configure\[10\]\[2\] _2893_ VGND
+ VGND VPWR VPWR _2894_ sky130_fd_sc_hd__a221o_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3286_ _0881_ VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__inv_2
XFILLER_97_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1115 gpio_configure\[34\]\[8\] VGND VGND VPWR VPWR net1648 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1126 _0479_ VGND VGND VPWR VPWR net1659 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 gpio_configure\[31\]\[10\] VGND VGND VPWR VPWR net1670 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5025_ _1793_ _1805_ _1823_ _2233_ VGND VGND VPWR VPWR _2235_ sky130_fd_sc_hd__a31o_1
Xhold1148 _0708_ VGND VGND VPWR VPWR net1681 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1159 net276 VGND VGND VPWR VPWR net1692 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6976_ clknet_leaf_43_csclk net845 net517 VGND VGND VPWR VPWR gpio_configure\[16\]\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_41_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5927_ gpio_configure\[4\]\[11\] _2502_ _2510_ gpio_configure\[15\]\[11\] VGND VGND
+ VPWR VPWR _2751_ sky130_fd_sc_hd__a22o_1
XFILLER_139_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5858_ gpio_configure\[0\]\[7\] _2526_ _2675_ _2685_ net473 VGND VGND VPWR VPWR _2686_
+ sky130_fd_sc_hd__o221a_2
XFILLER_179_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4809_ _1990_ _2018_ _2019_ VGND VGND VPWR VPWR _2020_ sky130_fd_sc_hd__and3b_1
XFILLER_166_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5789_ gpio_configure\[28\]\[4\] _2513_ _2517_ gpio_configure\[30\]\[4\] _2619_ VGND
+ VGND VPWR VPWR _2620_ sky130_fd_sc_hd__a221o_1
XFILLER_166_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold960 gpio_configure\[20\]\[8\] VGND VGND VPWR VPWR net1493 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold971 net229 VGND VGND VPWR VPWR net1504 sky130_fd_sc_hd__dlygate4sd3_1
Xhold982 _0811_ VGND VGND VPWR VPWR net1515 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold993 gpio_configure\[34\]\[5\] VGND VGND VPWR VPWR net1526 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_189_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6830_ clknet_leaf_29_csclk net619 net524 VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__dfrtp_1
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6761_ clknet_leaf_0_csclk net1835 net486 VGND VGND VPWR VPWR gpio_configure\[21\]\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_3973_ net567 net691 net668 VGND VGND VPWR VPWR _1465_ sky130_fd_sc_hd__mux2_4
X_5712_ gpio_configure\[14\]\[1\] _2494_ _2535_ gpio_configure\[23\]\[1\] _2545_ VGND
+ VGND VPWR VPWR _2546_ sky130_fd_sc_hd__a221o_1
X_6692_ clknet_3_7_0_wb_clk_i _0000_ net528 VGND VGND VPWR VPWR wbbd_state\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5643_ _2462_ _2476_ VGND VGND VPWR VPWR _2481_ sky130_fd_sc_hd__nor2_1
XFILLER_129_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5574_ net458 net1652 _2440_ VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__mux2_1
XFILLER_191_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold201 gpio_configure\[24\]\[4\] VGND VGND VPWR VPWR net734 sky130_fd_sc_hd__dlygate4sd3_1
X_4525_ _1632_ _1668_ _1702_ _1734_ _1736_ VGND VGND VPWR VPWR _1737_ sky130_fd_sc_hd__o2111a_1
Xhold212 _0321_ VGND VGND VPWR VPWR net745 sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 gpio_configure\[3\]\[6\] VGND VGND VPWR VPWR net756 sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 _0316_ VGND VGND VPWR VPWR net767 sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 gpio_configure\[21\]\[2\] VGND VGND VPWR VPWR net778 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold256 _0718_ VGND VGND VPWR VPWR net789 sky130_fd_sc_hd__dlygate4sd3_1
X_4456_ _1649_ _1656_ VGND VGND VPWR VPWR _1668_ sky130_fd_sc_hd__or2_4
XFILLER_131_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold267 gpio_configure\[8\]\[2\] VGND VGND VPWR VPWR net800 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold278 _0640_ VGND VGND VPWR VPWR net811 sky130_fd_sc_hd__dlygate4sd3_1
X_3407_ net18 _0864_ _0871_ net59 _1000_ VGND VGND VPWR VPWR _1001_ sky130_fd_sc_hd__a221o_1
Xhold289 gpio_configure\[2\]\[9\] VGND VGND VPWR VPWR net822 sky130_fd_sc_hd__dlygate4sd3_1
X_7175_ clknet_3_0_0_wb_clk_i _0777_ net505 VGND VGND VPWR VPWR serial_data_staging_2\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_132_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4387_ net99 _1596_ VGND VGND VPWR VPWR _1599_ sky130_fd_sc_hd__nand2_8
XFILLER_86_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6126_ gpio_configure\[7\]\[4\] _2811_ net407 gpio_configure\[15\]\[4\] _2942_ VGND
+ VGND VPWR VPWR _2944_ sky130_fd_sc_hd__a221o_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3338_ net376 net609 VGND VGND VPWR VPWR _0934_ sky130_fd_sc_hd__nor2_8
XFILLER_85_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6057_ gpio_configure\[16\]\[1\] _2831_ net391 gpio_configure\[17\]\[1\] _2877_ VGND
+ VGND VPWR VPWR _2878_ sky130_fd_sc_hd__a221o_1
X_3269_ net474 net626 net580 VGND VGND VPWR VPWR _0865_ sky130_fd_sc_hd__o21ai_1
XFILLER_45_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5008_ _2204_ _2206_ _2213_ _2217_ VGND VGND VPWR VPWR _2218_ sky130_fd_sc_hd__or4_1
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_129 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6959_ clknet_leaf_37_csclk net1539 net522 VGND VGND VPWR VPWR gpio_configure\[14\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_22_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold790 _0301_ VGND VGND VPWR VPWR net1323 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_150_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1490 net341 VGND VGND VPWR VPWR net2023 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_678 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_2_0__f_mgmt_gpio_in[4] clknet_0_mgmt_gpio_in[4] VGND VGND VPWR VPWR clknet_2_0__leaf_mgmt_gpio_in[4]
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput306 net306 VGND VGND VPWR VPWR ser_rx sky130_fd_sc_hd__buf_12
Xoutput317 net1902 VGND VGND VPWR VPWR wb_ack_o sky130_fd_sc_hd__buf_12
X_4310_ net449 net1252 _1543_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__mux2_1
Xoutput328 net1848 VGND VGND VPWR VPWR net1849 sky130_fd_sc_hd__buf_12
Xoutput339 net1894 VGND VGND VPWR VPWR net1895 sky130_fd_sc_hd__buf_12
X_5290_ net452 net990 net565 VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__mux2_1
XFILLER_113_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4241_ net1773 net468 _1532_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__mux2_1
XFILLER_114_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4172_ net2009 _1004_ _1517_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__mux2_1
XFILLER_67_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6813_ clknet_leaf_60_csclk net725 net499 VGND VGND VPWR VPWR serial_bb_clock sky130_fd_sc_hd__dfrtp_1
XFILLER_168_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6744_ clknet_leaf_75_csclk net1082 net488 VGND VGND VPWR VPWR gpio_configure\[19\]\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_3956_ wbbd_state\[8\] _1429_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__and2_1
X_6675_ clknet_leaf_11_csclk net1478 net511 VGND VGND VPWR VPWR gpio_configure\[11\]\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_167_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3887_ _1431_ _1432_ _1433_ _1438_ VGND VGND VPWR VPWR _1439_ sky130_fd_sc_hd__nor4_1
X_5626_ _2458_ _0825_ pad_count_2\[0\] VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__mux2_1
XFILLER_137_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5557_ net453 net1108 _2438_ VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__mux2_1
XFILLER_191_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4508_ _1643_ _1646_ _1659_ _1717_ _1719_ VGND VGND VPWR VPWR _1720_ sky130_fd_sc_hd__o2111a_1
XFILLER_132_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5488_ net452 net1075 _2430_ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__mux2_1
XFILLER_4_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_444 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4439_ _1647_ _1649_ VGND VGND VPWR VPWR _1651_ sky130_fd_sc_hd__or2_4
Xfanout500 net508 VGND VGND VPWR VPWR net500 sky130_fd_sc_hd__buf_4
XFILLER_116_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout511 net527 VGND VGND VPWR VPWR net511 sky130_fd_sc_hd__buf_8
XFILLER_132_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout522 net523 VGND VGND VPWR VPWR net522 sky130_fd_sc_hd__buf_8
X_7158_ clknet_3_2_0_wb_clk_i _0761_ net502 VGND VGND VPWR VPWR pad_count_2\[5\] sky130_fd_sc_hd__dfrtp_4
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6109_ _2921_ _2923_ _2925_ _2927_ VGND VGND VPWR VPWR _2928_ sky130_fd_sc_hd__or4_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7089_ clknet_leaf_31_csclk net949 net523 VGND VGND VPWR VPWR gpio_configure\[30\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_86_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3810_ net2078 _1388_ VGND VGND VPWR VPWR _1392_ sky130_fd_sc_hd__nand2_1
X_4790_ _1795_ _1800_ _1971_ VGND VGND VPWR VPWR _2001_ sky130_fd_sc_hd__o21ai_1
XFILLER_32_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_18 _0972_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_29 _1061_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3741_ gpio_configure\[11\]\[0\] _0907_ _1121_ gpio_configure\[17\]\[8\] VGND VGND
+ VPWR VPWR _1327_ sky130_fd_sc_hd__a22o_1
XFILLER_158_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6460_ clknet_2_1__leaf_mgmt_gpio_in[4] _0082_ _0038_ VGND VGND VPWR VPWR hkspi.pass_thru_mgmt_delay
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3672_ gpio_configure\[15\]\[1\] _0918_ _1045_ gpio_configure\[13\]\[9\] VGND VGND
+ VPWR VPWR _1260_ sky130_fd_sc_hd__a22o_1
XFILLER_173_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5411_ net435 net1045 _2421_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__mux2_1
XFILLER_173_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6391_ net2071 wbbd_state\[6\] _1530_ _3181_ VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__o31a_1
XFILLER_127_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5342_ net464 net1457 _2414_ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__mux2_1
XFILLER_126_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_720 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5273_ net447 net1194 _2406_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__mux2_1
XFILLER_99_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7012_ clknet_leaf_67_csclk net779 net505 VGND VGND VPWR VPWR gpio_configure\[21\]\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_4224_ net465 net620 net584 VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__mux2_1
X_4155_ net465 net900 _1515_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__mux2_1
XFILLER_95_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4086_ net1506 _1498_ _1490_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__mux2_1
XFILLER_71_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4988_ _2194_ _2195_ _2196_ _2197_ VGND VGND VPWR VPWR _2198_ sky130_fd_sc_hd__nor4_1
X_6727_ clknet_leaf_17_csclk net877 net512 VGND VGND VPWR VPWR gpio_configure\[36\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_3939_ serial_resetn_pre serial_bb_resetn serial_bb_enable VGND VGND VPWR VPWR net311
+ sky130_fd_sc_hd__mux2_2
XFILLER_176_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6658_ clknet_leaf_4_csclk net919 net495 VGND VGND VPWR VPWR gpio_configure\[7\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_5609_ xfer_state\[0\] xfer_state\[2\] VGND VGND VPWR VPWR _2457_ sky130_fd_sc_hd__nor2_1
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6589_ clknet_leaf_2_csclk net1456 net492 VGND VGND VPWR VPWR mgmt_gpio_data_buf\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput16 mask_rev_in[20] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_2
Xinput27 mask_rev_in[30] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput38 mgmt_gpio_in[11] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_4
XFILLER_167_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput49 mgmt_gpio_in[21] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_182_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5960_ gpio_configure\[16\]\[12\] _0831_ VGND VGND VPWR VPWR _2783_ sky130_fd_sc_hd__or2_1
X_4911_ net424 _1779_ _1689_ VGND VGND VPWR VPWR _2122_ sky130_fd_sc_hd__a21o_1
X_5891_ _2710_ _2712_ _2714_ _2716_ VGND VGND VPWR VPWR _2717_ sky130_fd_sc_hd__or4_1
XFILLER_61_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4842_ _1790_ _1886_ _1672_ VGND VGND VPWR VPWR _2053_ sky130_fd_sc_hd__o21ai_1
X_4773_ net530 _1950_ _1951_ _1984_ _1883_ VGND VGND VPWR VPWR _1985_ sky130_fd_sc_hd__a2111o_1
XFILLER_20_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6512_ clknet_leaf_1_csclk net1480 net493 VGND VGND VPWR VPWR gpio_configure\[30\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_3724_ _1311_ hkspi.ldata\[0\] _0837_ VGND VGND VPWR VPWR _1312_ sky130_fd_sc_hd__mux2_1
XFILLER_146_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3655_ gpio_configure\[20\]\[10\] _1053_ _1098_ gpio_configure\[25\]\[10\] VGND VGND
+ VPWR VPWR _1244_ sky130_fd_sc_hd__a22o_1
X_6443_ net532 _0018_ _0020_ VGND VGND VPWR VPWR hkspi.sdoenb sky130_fd_sc_hd__dfstp_1
XFILLER_106_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6374_ _3170_ net2065 _3162_ VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__mux2_1
X_3586_ gpio_configure\[28\]\[11\] _1046_ _1076_ gpio_configure\[27\]\[11\] _1143_
+ VGND VGND VPWR VPWR _1176_ sky130_fd_sc_hd__a221o_1
XFILLER_161_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5325_ net800 net577 _2412_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__mux2_1
XFILLER_130_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5256_ net1154 net441 _2404_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__mux2_1
XFILLER_87_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4207_ net1631 net455 _1522_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__mux2_1
XFILLER_102_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5187_ _1117_ net425 VGND VGND VPWR VPWR _2390_ sky130_fd_sc_hd__nand2_2
XFILLER_96_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4138_ net1662 net455 _1512_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__mux2_1
XFILLER_56_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4069_ net762 _1489_ _1481_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__mux2_1
XFILLER_73_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_523 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold608 _0568_ VGND VGND VPWR VPWR net1141 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3440_ gpio_configure\[19\]\[5\] _0896_ _0913_ gpio_configure\[7\]\[5\] _1031_ VGND
+ VGND VPWR VPWR _1032_ sky130_fd_sc_hd__a221o_1
Xhold619 gpio_configure\[18\]\[3\] VGND VGND VPWR VPWR net1152 sky130_fd_sc_hd__dlygate4sd3_1
X_3371_ _0962_ _0963_ _0964_ _0966_ VGND VGND VPWR VPWR _0967_ sky130_fd_sc_hd__or4_1
XFILLER_112_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5110_ _2314_ _2315_ _2317_ VGND VGND VPWR VPWR _2318_ sky130_fd_sc_hd__or3_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6090_ gpio_configure\[8\]\[2\] net410 _2861_ gpio_configure\[28\]\[2\] VGND VGND
+ VPWR VPWR _2910_ sky130_fd_sc_hd__a22o_1
XFILLER_112_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _1596_ net380 _1883_ _2248_ _2249_ VGND VGND VPWR VPWR _2250_ sky130_fd_sc_hd__a2111o_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1308 net1841 VGND VGND VPWR VPWR wb_dat_o[15] sky130_fd_sc_hd__buf_12
XFILLER_84_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1319 net1938 VGND VGND VPWR VPWR net1852 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_wb_clk_i wb_clk_i VGND VGND VPWR VPWR clknet_0_wb_clk_i sky130_fd_sc_hd__clkbuf_16
XFILLER_92_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6992_ clknet_leaf_41_csclk net803 net516 VGND VGND VPWR VPWR gpio_configure\[18\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_5943_ gpio_configure\[27\]\[11\] _2506_ _2541_ gpio_configure\[31\]\[11\] VGND VGND
+ VPWR VPWR _2767_ sky130_fd_sc_hd__a22o_1
XFILLER_179_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5874_ gpio_configure\[3\]\[8\] _2518_ _2541_ gpio_configure\[31\]\[8\] _2700_ VGND
+ VGND VPWR VPWR _2701_ sky130_fd_sc_hd__a221o_1
XFILLER_178_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4825_ _1988_ _2034_ _2035_ _1761_ VGND VGND VPWR VPWR _2036_ sky130_fd_sc_hd__o31a_1
XFILLER_166_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4756_ _1629_ _1956_ _1967_ _1749_ VGND VGND VPWR VPWR _1968_ sky130_fd_sc_hd__o22a_1
XFILLER_119_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3707_ gpio_configure\[8\]\[1\] _0939_ _1053_ gpio_configure\[20\]\[9\] _1294_ VGND
+ VGND VPWR VPWR _1295_ sky130_fd_sc_hd__a221o_1
XFILLER_146_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4687_ _1613_ _1693_ VGND VGND VPWR VPWR _1899_ sky130_fd_sc_hd__nor2_1
XFILLER_174_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6426_ net486 net481 VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__and2_1
X_3638_ gpio_configure\[32\]\[10\] _1101_ _1127_ gpio_configure\[33\]\[10\] VGND VGND
+ VPWR VPWR _1227_ sky130_fd_sc_hd__a22o_1
XFILLER_162_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3569_ gpio_configure\[37\]\[3\] _0902_ _0938_ gpio_configure\[33\]\[3\] VGND VGND
+ VPWR VPWR _1159_ sky130_fd_sc_hd__a22o_1
X_6357_ net168 net170 VGND VGND VPWR VPWR _3157_ sky130_fd_sc_hd__nand2_1
X_5308_ net569 net732 _2410_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__mux2_1
X_6288_ gpio_configure\[1\]\[10\] _2802_ _2858_ gpio_configure\[24\]\[10\] _3099_
+ VGND VGND VPWR VPWR _3100_ sky130_fd_sc_hd__a221o_1
XFILLER_48_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5239_ net439 net1911 _2402_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__mux2_1
XFILLER_102_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold5 net541 VGND VGND VPWR VPWR net538 sky130_fd_sc_hd__buf_6
XFILLER_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4610_ _0836_ _1776_ VGND VGND VPWR VPWR _1822_ sky130_fd_sc_hd__or2_2
XFILLER_175_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5590_ _0822_ serial_xfer xfer_state\[3\] _1443_ _2442_ VGND VGND VPWR VPWR _0746_
+ sky130_fd_sc_hd__o311a_1
XFILLER_128_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4541_ net128 _1751_ VGND VGND VPWR VPWR _1753_ sky130_fd_sc_hd__nand2_2
XFILLER_144_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold405 gpio_configure\[37\]\[9\] VGND VGND VPWR VPWR net938 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire380 _1675_ VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__buf_2
XFILLER_190_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold416 _0692_ VGND VGND VPWR VPWR net949 sky130_fd_sc_hd__dlygate4sd3_1
X_4472_ net110 net530 net124 net99 VGND VGND VPWR VPWR _1684_ sky130_fd_sc_hd__or4bb_4
Xhold427 gpio_configure\[22\]\[3\] VGND VGND VPWR VPWR net960 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold438 _0709_ VGND VGND VPWR VPWR net971 sky130_fd_sc_hd__dlygate4sd3_1
X_3423_ gpio_configure\[18\]\[5\] _0894_ _0922_ gpio_configure\[23\]\[5\] _1014_ VGND
+ VGND VPWR VPWR _1015_ sky130_fd_sc_hd__a221o_1
X_6211_ gpio_configure\[10\]\[7\] _2825_ net394 gpio_configure\[6\]\[7\] _3025_ VGND
+ VGND VPWR VPWR _3026_ sky130_fd_sc_hd__a221o_1
XFILLER_116_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold449 gpio_configure\[12\]\[3\] VGND VGND VPWR VPWR net982 sky130_fd_sc_hd__dlygate4sd3_1
X_7191_ clknet_3_4_0_wb_clk_i _0793_ VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__dfxtp_2
XFILLER_144_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6142_ _2944_ _2955_ _2957_ _2959_ VGND VGND VPWR VPWR _2960_ sky130_fd_sc_hd__or4_4
X_3354_ gpio_configure\[37\]\[7\] _0902_ net369 gpio_configure\[25\]\[7\] _0949_ VGND
+ VGND VPWR VPWR _0950_ sky130_fd_sc_hd__a221o_4
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ gpio_configure\[20\]\[2\] net396 net408 gpio_configure\[35\]\[2\] VGND VGND
+ VPWR VPWR _2893_ sky130_fd_sc_hd__a22o_1
Xhold1105 gpio_configure\[25\]\[10\] VGND VGND VPWR VPWR net1638 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3285_ _0879_ net2006 VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__nand2_8
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1116 _0349_ VGND VGND VPWR VPWR net1649 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _1823_ _2233_ VGND VGND VPWR VPWR _2234_ sky130_fd_sc_hd__nor2_1
Xhold1127 gpio_configure\[1\]\[2\] VGND VGND VPWR VPWR net1660 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1138 _0695_ VGND VGND VPWR VPWR net1671 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1149 net268 VGND VGND VPWR VPWR net1682 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_81_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6975_ clknet_leaf_31_csclk net1545 net523 VGND VGND VPWR VPWR gpio_configure\[16\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5926_ net2073 _2750_ net366 VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__mux2_1
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5857_ _2677_ _2680_ _2682_ _2684_ VGND VGND VPWR VPWR _2685_ sky130_fd_sc_hd__or4_1
XFILLER_139_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4808_ net477 _1777_ _1782_ _1636_ _1599_ VGND VGND VPWR VPWR _2019_ sky130_fd_sc_hd__o32a_1
XFILLER_186_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5788_ gpio_configure\[20\]\[4\] _2499_ _2523_ gpio_configure\[2\]\[4\] VGND VGND
+ VPWR VPWR _2619_ sky130_fd_sc_hd__a22o_1
X_4739_ _1613_ _1949_ VGND VGND VPWR VPWR _1951_ sky130_fd_sc_hd__nor2_1
XFILLER_181_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6409_ net492 net482 VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__and2_1
XFILLER_135_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold950 gpio_configure\[6\]\[9\] VGND VGND VPWR VPWR net1483 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold961 _0354_ VGND VGND VPWR VPWR net1494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold972 _0429_ VGND VGND VPWR VPWR net1505 sky130_fd_sc_hd__dlygate4sd3_1
Xhold983 gpio_configure\[27\]\[9\] VGND VGND VPWR VPWR net1516 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold994 _0719_ VGND VGND VPWR VPWR net1527 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_50_csclk clknet_3_3_0_csclk VGND VGND VPWR VPWR clknet_leaf_50_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_99_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_65_csclk clknet_3_3_0_csclk VGND VGND VPWR VPWR clknet_leaf_65_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_47_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6760_ clknet_leaf_72_csclk net1022 net490 VGND VGND VPWR VPWR gpio_configure\[33\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_50_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3972_ net1640 net455 _1461_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__mux2_1
XFILLER_62_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5711_ gpio_configure\[26\]\[1\] _2534_ _2541_ gpio_configure\[31\]\[1\] VGND VGND
+ VPWR VPWR _2545_ sky130_fd_sc_hd__a22o_1
XFILLER_149_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6691_ clknet_3_7_0_wb_clk_i net2087 net528 VGND VGND VPWR VPWR wbbd_state\[0\] sky130_fd_sc_hd__dfstp_1
XFILLER_149_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5642_ _2469_ _2473_ _2478_ VGND VGND VPWR VPWR _2480_ sky130_fd_sc_hd__and3_4
XFILLER_176_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5573_ net464 net1429 _2440_ VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__mux2_1
XFILLER_129_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold202 _0641_ VGND VGND VPWR VPWR net735 sky130_fd_sc_hd__dlygate4sd3_1
X_4524_ _1612_ _1667_ VGND VGND VPWR VPWR _1736_ sky130_fd_sc_hd__nand2_1
Xhold213 gpio_configure\[30\]\[2\] VGND VGND VPWR VPWR net746 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 _0475_ VGND VGND VPWR VPWR net757 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_18_csclk clknet_3_4_0_csclk VGND VGND VPWR VPWR clknet_leaf_18_csclk
+ sky130_fd_sc_hd__clkbuf_16
Xhold235 gpio_configure\[32\]\[11\] VGND VGND VPWR VPWR net768 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold246 _0615_ VGND VGND VPWR VPWR net779 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4455_ _1649_ _1656_ VGND VGND VPWR VPWR _1667_ sky130_fd_sc_hd__nor2_2
Xhold257 net280 VGND VGND VPWR VPWR net790 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold268 _0511_ VGND VGND VPWR VPWR net801 sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 gpio_configure\[19\]\[3\] VGND VGND VPWR VPWR net812 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3406_ net27 _0936_ _0938_ gpio_configure\[33\]\[6\] VGND VGND VPWR VPWR _1000_ sky130_fd_sc_hd__a22o_1
X_7174_ clknet_3_2_0_wb_clk_i _0776_ net499 VGND VGND VPWR VPWR serial_data_staging_1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_4386_ _0833_ _1597_ VGND VGND VPWR VPWR _1598_ sky130_fd_sc_hd__nor2_8
XFILLER_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3337_ net628 _0909_ VGND VGND VPWR VPWR _0933_ sky130_fd_sc_hd__nor2_8
X_6125_ gpio_configure\[30\]\[4\] _2799_ net408 gpio_configure\[35\]\[4\] VGND VGND
+ VPWR VPWR _2943_ sky130_fd_sc_hd__a22o_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3268_ net390 _0863_ VGND VGND VPWR VPWR _0864_ sky130_fd_sc_hd__nor2_8
XFILLER_86_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6056_ gpio_configure\[14\]\[1\] net411 net406 gpio_configure\[27\]\[1\] VGND VGND
+ VPWR VPWR _2877_ sky130_fd_sc_hd__a22o_1
XFILLER_65_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5007_ _1944_ _2205_ _2210_ _2216_ VGND VGND VPWR VPWR _2217_ sky130_fd_sc_hd__or4_1
XFILLER_54_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3199_ gpio_configure\[35\]\[3\] VGND VGND VPWR VPWR _0828_ sky130_fd_sc_hd__clkinv_2
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_108 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_119 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6958_ clknet_leaf_16_csclk net1297 net512 VGND VGND VPWR VPWR gpio_configure\[14\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_53_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5909_ gpio_configure\[3\]\[10\] _2518_ _2528_ gpio_configure\[7\]\[10\] VGND VGND
+ VPWR VPWR _2734_ sky130_fd_sc_hd__a22o_1
X_6889_ clknet_leaf_41_csclk net1058 net517 VGND VGND VPWR VPWR gpio_configure\[5\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_139_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_667 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_1_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold780 _0612_ VGND VGND VPWR VPWR net1313 sky130_fd_sc_hd__dlygate4sd3_1
Xhold791 gpio_configure\[31\]\[11\] VGND VGND VPWR VPWR net1324 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1480 net323 VGND VGND VPWR VPWR net2013 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1491 net322 VGND VGND VPWR VPWR net2024 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput307 net307 VGND VGND VPWR VPWR serial_clock sky130_fd_sc_hd__buf_12
Xoutput318 net1878 VGND VGND VPWR VPWR net1879 sky130_fd_sc_hd__buf_12
Xoutput329 net1880 VGND VGND VPWR VPWR net1881 sky130_fd_sc_hd__buf_12
XFILLER_141_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4240_ _1045_ net426 VGND VGND VPWR VPWR _1532_ sky130_fd_sc_hd__and2_2
XFILLER_113_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4171_ net2012 _1039_ _1517_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__mux2_1
XFILLER_122_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6812_ clknet_leaf_70_csclk net1496 net491 VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__dfrtp_4
XFILLER_51_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6743_ clknet_leaf_76_csclk net1633 net484 VGND VGND VPWR VPWR gpio_configure\[19\]\[10\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_189_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3955_ wbbd_state\[5\] _1429_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__and2_1
XFILLER_188_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6674_ clknet_leaf_5_csclk net1219 net496 VGND VGND VPWR VPWR gpio_configure\[10\]\[12\]
+ sky130_fd_sc_hd__dfrtp_2
X_3886_ _1434_ _1435_ _1436_ _1437_ VGND VGND VPWR VPWR _1438_ sky130_fd_sc_hd__or4_1
X_5625_ _2468_ _0831_ _2467_ VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__mux2_1
XFILLER_137_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5556_ net458 net1732 _2438_ VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__mux2_1
XFILLER_3_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4507_ _1632_ _1663_ _1651_ VGND VGND VPWR VPWR _1719_ sky130_fd_sc_hd__a21o_1
X_5487_ net458 net1686 _2430_ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__mux2_1
XFILLER_160_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4438_ _1647_ _1649_ VGND VGND VPWR VPWR _1650_ sky130_fd_sc_hd__nor2_1
Xfanout501 net508 VGND VGND VPWR VPWR net501 sky130_fd_sc_hd__buf_8
Xfanout512 net527 VGND VGND VPWR VPWR net512 sky130_fd_sc_hd__buf_8
XFILLER_132_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout523 net526 VGND VGND VPWR VPWR net523 sky130_fd_sc_hd__buf_6
X_7157_ clknet_3_3_0_wb_clk_i _0760_ net502 VGND VGND VPWR VPWR pad_count_2\[4\] sky130_fd_sc_hd__dfstp_2
XFILLER_116_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4369_ _1555_ _1577_ VGND VGND VPWR VPWR _1581_ sky130_fd_sc_hd__or2_4
XFILLER_112_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6108_ gpio_configure\[21\]\[3\] _2820_ _2822_ gpio_configure\[23\]\[3\] _2926_ VGND
+ VGND VPWR VPWR _2927_ sky130_fd_sc_hd__a221o_1
XFILLER_59_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7088_ clknet_leaf_52_csclk net1386 net507 VGND VGND VPWR VPWR gpio_configure\[30\]\[6\]
+ sky130_fd_sc_hd__dfrtp_2
X_6039_ _2473_ _2478_ _2793_ VGND VGND VPWR VPWR _2861_ sky130_fd_sc_hd__and3_4
XFILLER_27_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_681 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_19 _1004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3740_ gpio_configure\[7\]\[0\] _0913_ _1109_ gpio_configure\[36\]\[8\] VGND VGND
+ VPWR VPWR _1326_ sky130_fd_sc_hd__a22o_1
XFILLER_119_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3671_ gpio_configure\[32\]\[1\] _0890_ _1116_ gpio_configure\[26\]\[9\] _1258_ VGND
+ VGND VPWR VPWR _1259_ sky130_fd_sc_hd__a221o_1
X_5410_ net437 net1433 _2421_ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__mux2_1
XFILLER_185_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6390_ _0820_ net433 _3160_ _3180_ net170 VGND VGND VPWR VPWR _3181_ sky130_fd_sc_hd__a32o_1
X_5341_ net469 net1644 _2414_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__mux2_1
XFILLER_114_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5272_ net451 net694 _2406_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__mux2_1
XFILLER_114_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7011_ clknet_leaf_23_csclk net1331 net514 VGND VGND VPWR VPWR gpio_configure\[21\]\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_4223_ net470 net1477 net584 VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__mux2_1
XFILLER_114_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4154_ net470 net1755 _1515_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__mux2_1
XFILLER_83_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4085_ net1288 net434 net351 VGND VGND VPWR VPWR _1498_ sky130_fd_sc_hd__mux2_1
XFILLER_55_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4987_ _1844_ _1963_ _2002_ VGND VGND VPWR VPWR _2197_ sky130_fd_sc_hd__or3_1
X_6726_ clknet_leaf_17_csclk net1595 net512 VGND VGND VPWR VPWR gpio_configure\[36\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_3938_ mgmt_gpio_data\[13\] net93 trap_output_dest VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__mux2_2
XFILLER_177_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6657_ clknet_leaf_3_csclk net1361 net493 VGND VGND VPWR VPWR gpio_configure\[7\]\[10\]
+ sky130_fd_sc_hd__dfstp_1
X_3869_ _0814_ net58 _1424_ _1425_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__a31o_1
XFILLER_164_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5608_ net2122 _2454_ _2456_ VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__o21a_1
XFILLER_137_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6588_ clknet_leaf_78_csclk net1511 net486 VGND VGND VPWR VPWR mgmt_gpio_data_buf\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_117_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5539_ net740 net451 _2436_ VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__mux2_1
XFILLER_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7209_ clknet_leaf_77_csclk net1515 net485 VGND VGND VPWR VPWR gpio_configure\[27\]\[10\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_160_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput17 mask_rev_in[21] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_1
XFILLER_168_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput28 mask_rev_in[31] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_1
XFILLER_10_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput39 mgmt_gpio_in[12] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_4
XFILLER_182_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4910_ _1757_ _1790_ _1863_ VGND VGND VPWR VPWR _2121_ sky130_fd_sc_hd__a21o_1
XFILLER_45_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5890_ gpio_configure\[13\]\[9\] _2501_ _2534_ gpio_configure\[26\]\[9\] _2715_ VGND
+ VGND VPWR VPWR _2716_ sky130_fd_sc_hd__a221o_1
XFILLER_61_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4841_ _1684_ _1798_ _1732_ VGND VGND VPWR VPWR _2052_ sky130_fd_sc_hd__o21ai_1
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4772_ _1662_ _1686_ _1982_ _1983_ VGND VGND VPWR VPWR _1984_ sky130_fd_sc_hd__a211o_1
XFILLER_159_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6511_ clknet_leaf_1_csclk net1811 net493 VGND VGND VPWR VPWR gpio_configure\[30\]\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_3723_ _1257_ _1277_ _1310_ VGND VGND VPWR VPWR _1311_ sky130_fd_sc_hd__or3_4
XFILLER_119_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6442_ clknet_2_1__leaf_mgmt_gpio_in[4] _0065_ _0019_ VGND VGND VPWR VPWR hkspi.wrstb
+ sky130_fd_sc_hd__dfrtn_1
XFILLER_146_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3654_ gpio_configure\[30\]\[2\] _0892_ net371 gpio_configure\[26\]\[2\] _1194_ VGND
+ VGND VPWR VPWR _1243_ sky130_fd_sc_hd__a221o_1
XFILLER_173_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6373_ wbbd_state\[9\] net151 net157 net433 _3169_ VGND VGND VPWR VPWR _3170_ sky130_fd_sc_hd__a221o_1
Xclkbuf_3_0_0_wb_clk_i clknet_2_0_0_wb_clk_i VGND VGND VPWR VPWR clknet_3_0_0_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
X_3585_ net261 _1009_ _1137_ net95 _1142_ VGND VGND VPWR VPWR _1175_ sky130_fd_sc_hd__a221o_1
XFILLER_161_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5324_ net872 net465 _2412_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__mux2_1
XFILLER_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5255_ net689 net445 _2404_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__mux2_1
XFILLER_130_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4206_ net1625 net461 _1522_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__mux2_1
X_5186_ net461 net1592 _2389_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__mux2_1
XFILLER_29_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4137_ net1684 net461 _1512_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__mux2_1
XFILLER_96_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4068_ net1904 net573 net356 VGND VGND VPWR VPWR _1489_ sky130_fd_sc_hd__mux2_1
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6709_ clknet_leaf_4_csclk net917 net496 VGND VGND VPWR VPWR gpio_configure\[15\]\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_177_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold609 gpio_configure\[24\]\[5\] VGND VGND VPWR VPWR net1142 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3370_ gpio_configure\[16\]\[7\] _0912_ _0915_ gpio_configure\[3\]\[7\] _0965_ VGND
+ VGND VPWR VPWR _0966_ sky130_fd_sc_hd__a221o_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _1596_ _1686_ _1869_ VGND VGND VPWR VPWR _2249_ sky130_fd_sc_hd__a21o_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1309 net1931 VGND VGND VPWR VPWR net1842 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6991_ clknet_leaf_43_csclk net1147 net517 VGND VGND VPWR VPWR gpio_configure\[18\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_25_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5942_ gpio_configure\[13\]\[11\] _2501_ _2517_ gpio_configure\[30\]\[11\] _2765_
+ VGND VGND VPWR VPWR _2766_ sky130_fd_sc_hd__a221o_1
XFILLER_18_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5873_ gpio_configure\[19\]\[8\] _2491_ _2524_ _2699_ VGND VGND VPWR VPWR _2700_
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4824_ _1747_ _1933_ VGND VGND VPWR VPWR _2035_ sky130_fd_sc_hd__nand2_1
XFILLER_21_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4755_ _1598_ _1617_ _1622_ _1628_ _1584_ VGND VGND VPWR VPWR _1967_ sky130_fd_sc_hd__a41o_1
XFILLER_159_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3706_ serial_bb_enable _0974_ _1083_ gpio_configure\[30\]\[9\] VGND VGND VPWR VPWR
+ _1294_ sky130_fd_sc_hd__a22o_1
XFILLER_119_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4686_ _1693_ net432 VGND VGND VPWR VPWR _1898_ sky130_fd_sc_hd__or2_1
XFILLER_174_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6425_ net495 net482 VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__and2_1
XFILLER_119_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3637_ net5 _0891_ _0910_ net293 _1225_ VGND VGND VPWR VPWR _1226_ sky130_fd_sc_hd__a221o_1
XFILLER_146_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6356_ net1948 _0969_ _3156_ VGND VGND VPWR VPWR _0798_ sky130_fd_sc_hd__mux2_1
X_3568_ gpio_configure\[13\]\[3\] _0906_ _1136_ net304 _1157_ VGND VGND VPWR VPWR
+ _1158_ sky130_fd_sc_hd__a221o_1
XFILLER_88_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5307_ net459 net1387 _2410_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__mux2_1
X_6287_ gpio_configure\[31\]\[10\] _2480_ _2814_ gpio_configure\[11\]\[10\] VGND VGND
+ VPWR VPWR _3099_ sky130_fd_sc_hd__a22o_1
XFILLER_88_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3499_ _1078_ _1082_ _1085_ _1089_ VGND VGND VPWR VPWR _1090_ sky130_fd_sc_hd__or4_2
X_5238_ net441 net944 _2402_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__mux2_1
XFILLER_75_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5169_ _1757_ _1795_ _1940_ _1655_ _1838_ VGND VGND VPWR VPWR _2375_ sky130_fd_sc_hd__o221a_1
XFILLER_56_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold6 net1913 VGND VGND VPWR VPWR net539 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_59_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4540_ net128 _1554_ _1749_ VGND VGND VPWR VPWR _1752_ sky130_fd_sc_hd__and3_1
XFILLER_129_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold406 _0320_ VGND VGND VPWR VPWR net939 sky130_fd_sc_hd__dlygate4sd3_1
X_4471_ net530 _1579_ VGND VGND VPWR VPWR _1683_ sky130_fd_sc_hd__nor2_1
XFILLER_183_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold417 net245 VGND VGND VPWR VPWR net950 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold428 _0624_ VGND VGND VPWR VPWR net961 sky130_fd_sc_hd__dlygate4sd3_1
X_6210_ gpio_configure\[9\]\[7\] net412 net409 gpio_configure\[12\]\[7\] VGND VGND
+ VPWR VPWR _3025_ sky130_fd_sc_hd__a22o_1
XFILLER_116_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold439 gpio_configure\[30\]\[3\] VGND VGND VPWR VPWR net972 sky130_fd_sc_hd__dlygate4sd3_1
X_3422_ net31 _0900_ _0940_ net279 VGND VGND VPWR VPWR _1014_ sky130_fd_sc_hd__a22o_2
X_7190_ clknet_3_4_0_wb_clk_i _0792_ VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__dfxtp_1
XFILLER_99_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6141_ gpio_configure\[1\]\[4\] net401 net405 gpio_configure\[24\]\[4\] _2958_ VGND
+ VGND VPWR VPWR _2959_ sky130_fd_sc_hd__a221o_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ gpio_configure\[28\]\[7\] _0888_ _0932_ gpio_configure\[35\]\[7\] VGND VGND
+ VPWR VPWR _0949_ sky130_fd_sc_hd__a22o_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6072_ net2060 _2892_ net366 VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__mux2_1
XFILLER_112_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ net588 net560 VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__nor2_8
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1106 _0150_ VGND VGND VPWR VPWR net1639 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1117 gpio_configure\[19\]\[9\] VGND VGND VPWR VPWR net1650 sky130_fd_sc_hd__dlygate4sd3_1
X_5023_ _1588_ _1684_ _1778_ VGND VGND VPWR VPWR _2233_ sky130_fd_sc_hd__and3_2
Xhold1128 _0455_ VGND VGND VPWR VPWR net1661 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1139 gpio_configure\[3\]\[9\] VGND VGND VPWR VPWR net1672 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6974_ clknet_leaf_25_csclk net1239 net518 VGND VGND VPWR VPWR gpio_configure\[16\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_5925_ xfer_state\[1\] serial_data_staging_1\[9\] _2749_ VGND VGND VPWR VPWR _2750_
+ sky130_fd_sc_hd__a21o_1
XFILLER_61_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5856_ gpio_configure\[9\]\[7\] _2512_ _2534_ gpio_configure\[26\]\[7\] _2683_ VGND
+ VGND VPWR VPWR _2684_ sky130_fd_sc_hd__a221o_1
X_4807_ _1772_ _1774_ _1822_ _2005_ _1745_ VGND VGND VPWR VPWR _2018_ sky130_fd_sc_hd__o32a_1
X_5787_ gpio_configure\[6\]\[4\] _2490_ _2606_ _2617_ VGND VGND VPWR VPWR _2618_ sky130_fd_sc_hd__a211o_1
XFILLER_166_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4738_ _1632_ _1949_ VGND VGND VPWR VPWR _1950_ sky130_fd_sc_hd__nor2_1
XFILLER_119_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4669_ _1875_ _1878_ _1879_ _1877_ _1601_ VGND VGND VPWR VPWR _1881_ sky130_fd_sc_hd__o32a_1
X_6408_ net492 net482 VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__and2_1
Xhold940 gpio_configure\[29\]\[9\] VGND VGND VPWR VPWR net1473 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold951 _0248_ VGND VGND VPWR VPWR net1484 sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 net172 VGND VGND VPWR VPWR net1495 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold973 net248 VGND VGND VPWR VPWR net1506 sky130_fd_sc_hd__dlygate4sd3_1
X_6339_ gpio_configure\[33\]\[12\] _2829_ _2862_ gpio_configure\[25\]\[12\] _3148_
+ VGND VGND VPWR VPWR _3149_ sky130_fd_sc_hd__a221o_2
Xhold984 _0810_ VGND VGND VPWR VPWR net1517 sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 gpio_configure\[8\]\[5\] VGND VGND VPWR VPWR net1528 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_438 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3971_ net575 net594 net474 VGND VGND VPWR VPWR _1464_ sky130_fd_sc_hd__mux2_4
X_5710_ net2019 _2487_ _2544_ VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__a21o_1
XFILLER_43_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6690_ clknet_leaf_5_csclk net1231 net496 VGND VGND VPWR VPWR gpio_configure\[13\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5641_ pad_count_2\[5\] pad_count_2\[4\] VGND VGND VPWR VPWR _2479_ sky130_fd_sc_hd__nand2b_4
XFILLER_148_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5572_ net471 net1604 _2440_ VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__mux2_1
XFILLER_163_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_1_csclk clknet_1_0_0_csclk VGND VGND VPWR VPWR clknet_1_0_1_csclk sky130_fd_sc_hd__clkbuf_8
XFILLER_163_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4523_ _1668_ _1671_ VGND VGND VPWR VPWR _1735_ sky130_fd_sc_hd__nor2_2
XFILLER_129_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold203 net230 VGND VGND VPWR VPWR net736 sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 _0687_ VGND VGND VPWR VPWR net747 sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 gpio_configure\[34\]\[10\] VGND VGND VPWR VPWR net758 sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 _0372_ VGND VGND VPWR VPWR net769 sky130_fd_sc_hd__dlygate4sd3_1
X_4454_ _1665_ VGND VGND VPWR VPWR _1666_ sky130_fd_sc_hd__inv_2
Xhold247 gpio_configure\[17\]\[2\] VGND VGND VPWR VPWR net780 sky130_fd_sc_hd__dlygate4sd3_1
Xhold258 _0110_ VGND VGND VPWR VPWR net791 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold269 gpio_configure\[18\]\[6\] VGND VGND VPWR VPWR net802 sky130_fd_sc_hd__dlygate4sd3_1
X_3405_ gpio_configure\[36\]\[6\] net352 net351 net69 _0978_ VGND VGND VPWR VPWR _0999_
+ sky130_fd_sc_hd__a221o_1
X_7173_ clknet_3_1_0_wb_clk_i _0775_ net488 VGND VGND VPWR VPWR serial_data_staging_1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_4385_ net530 _1595_ VGND VGND VPWR VPWR _1597_ sky130_fd_sc_hd__or2_4
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6124_ gpio_configure\[26\]\[4\] _2810_ net413 gpio_configure\[3\]\[4\] VGND VGND
+ VPWR VPWR _2942_ sky130_fd_sc_hd__a22o_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3336_ net628 _0895_ VGND VGND VPWR VPWR _0932_ sky130_fd_sc_hd__nor2_8
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0__1134_ _1134_ VGND VGND VPWR VPWR clknet_0__1134_ sky130_fd_sc_hd__clkbuf_16
X_6055_ gpio_configure\[22\]\[1\] net397 net395 gpio_configure\[33\]\[1\] _2875_ VGND
+ VGND VPWR VPWR _2876_ sky130_fd_sc_hd__a221o_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ _0857_ net589 VGND VGND VPWR VPWR _0863_ sky130_fd_sc_hd__nand2_8
XFILLER_100_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5006_ _1629_ _1635_ _1956_ _1703_ _1584_ VGND VGND VPWR VPWR _2216_ sky130_fd_sc_hd__o32a_1
XFILLER_38_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3198_ gpio_configure\[36\]\[3\] VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__clkinv_2
XFILLER_54_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_109 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6957_ clknet_leaf_36_csclk net1161 net522 VGND VGND VPWR VPWR gpio_configure\[14\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_81_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5908_ gpio_configure\[30\]\[10\] _2517_ _2520_ gpio_configure\[8\]\[10\] _2732_
+ VGND VGND VPWR VPWR _2733_ sky130_fd_sc_hd__a221o_1
X_6888_ clknet_leaf_53_csclk net1359 net507 VGND VGND VPWR VPWR gpio_configure\[5\]\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_139_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5839_ gpio_configure\[28\]\[7\] _2513_ _2521_ gpio_configure\[21\]\[7\] VGND VGND
+ VPWR VPWR _2667_ sky130_fd_sc_hd__a22o_1
XFILLER_10_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold770 _0505_ VGND VGND VPWR VPWR net1303 sky130_fd_sc_hd__dlygate4sd3_1
Xhold781 gpio_configure\[18\]\[7\] VGND VGND VPWR VPWR net1314 sky130_fd_sc_hd__dlygate4sd3_1
Xhold792 _0696_ VGND VGND VPWR VPWR net1325 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3234__1 clknet_2_3__leaf_mgmt_gpio_in[4] VGND VGND VPWR VPWR net532 sky130_fd_sc_hd__inv_2
XFILLER_162_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1470 wbbd_state\[1\] VGND VGND VPWR VPWR net2003 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1481 net328 VGND VGND VPWR VPWR net2014 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1492 wbbd_state\[4\] VGND VGND VPWR VPWR net2025 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput308 net308 VGND VGND VPWR VPWR serial_data_1 sky130_fd_sc_hd__buf_12
Xoutput319 net1856 VGND VGND VPWR VPWR net1857 sky130_fd_sc_hd__buf_12
XFILLER_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4170_ net1959 clknet_1_1__leaf__1134_ _1517_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__mux2_1
XFILLER_67_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6811_ clknet_leaf_77_csclk net1768 net487 VGND VGND VPWR VPWR reset_reg sky130_fd_sc_hd__dfrtp_1
XFILLER_36_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6742_ clknet_leaf_76_csclk net1651 net484 VGND VGND VPWR VPWR gpio_configure\[19\]\[9\]
+ sky130_fd_sc_hd__dfrtp_4
X_3954_ wbbd_state\[7\] _1429_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__and2_1
XFILLER_149_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6673_ clknet_leaf_5_csclk net1223 net496 VGND VGND VPWR VPWR gpio_configure\[10\]\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_3885_ net118 net119 net120 net117 VGND VGND VPWR VPWR _1437_ sky130_fd_sc_hd__or4bb_1
XFILLER_176_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5624_ _0831_ _2463_ VGND VGND VPWR VPWR _2468_ sky130_fd_sc_hd__nand2_1
XFILLER_176_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5555_ net463 net906 _2438_ VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__mux2_1
XFILLER_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4506_ _1651_ _1671_ VGND VGND VPWR VPWR _1718_ sky130_fd_sc_hd__nor2_2
X_5486_ net464 net1328 _2430_ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__mux2_1
XFILLER_104_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4437_ _1617_ _1648_ VGND VGND VPWR VPWR _1649_ sky130_fd_sc_hd__nand2_1
XFILLER_104_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout502 net504 VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__buf_8
XFILLER_132_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout513 net527 VGND VGND VPWR VPWR net513 sky130_fd_sc_hd__buf_6
X_7156_ clknet_3_2_0_wb_clk_i _0759_ net502 VGND VGND VPWR VPWR pad_count_2\[3\] sky130_fd_sc_hd__dfrtp_1
Xfanout524 net525 VGND VGND VPWR VPWR net524 sky130_fd_sc_hd__buf_8
X_4368_ _1555_ _1577_ VGND VGND VPWR VPWR _1580_ sky130_fd_sc_hd__nor2_2
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6107_ gpio_configure\[29\]\[3\] _2816_ net397 gpio_configure\[22\]\[3\] VGND VGND
+ VPWR VPWR _2926_ sky130_fd_sc_hd__a22o_1
XFILLER_59_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3319_ net376 _0895_ VGND VGND VPWR VPWR _0915_ sky130_fd_sc_hd__nor2_8
X_7087_ clknet_leaf_32_csclk net953 net524 VGND VGND VPWR VPWR gpio_configure\[30\]\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_4299_ net443 net1013 _1541_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__mux2_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6038_ _2479_ _2801_ VGND VGND VPWR VPWR _2860_ sky130_fd_sc_hd__nor2_8
XFILLER_100_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_64_csclk clknet_3_2_0_csclk VGND VGND VPWR VPWR clknet_leaf_64_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_41_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_17_csclk clknet_3_5_0_csclk VGND VGND VPWR VPWR clknet_leaf_17_csclk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_647 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_60_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3670_ gpio_configure\[0\]\[9\] _1087_ _1127_ gpio_configure\[33\]\[9\] VGND VGND
+ VPWR VPWR _1258_ sky130_fd_sc_hd__a22o_1
XFILLER_185_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5340_ _0920_ net427 VGND VGND VPWR VPWR _2414_ sky130_fd_sc_hd__nand2_8
XFILLER_127_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5271_ net458 net1570 _2406_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__mux2_1
XFILLER_181_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7010_ clknet_leaf_21_csclk net1215 net514 VGND VGND VPWR VPWR gpio_configure\[21\]\[0\]
+ sky130_fd_sc_hd__dfstp_2
X_4222_ net583 net429 VGND VGND VPWR VPWR _1525_ sky130_fd_sc_hd__nand2_2
XFILLER_68_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4153_ _1093_ net429 VGND VGND VPWR VPWR _1515_ sky130_fd_sc_hd__nand2_2
XFILLER_55_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4084_ net942 _1497_ _1490_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__mux2_1
XFILLER_55_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4986_ _1831_ _1964_ _2010_ VGND VGND VPWR VPWR _2196_ sky130_fd_sc_hd__or3b_1
X_6725_ clknet_leaf_9_csclk net1105 net510 VGND VGND VPWR VPWR gpio_configure\[17\]\[12\]
+ sky130_fd_sc_hd__dfrtp_2
X_3937_ mgmt_gpio_data\[14\] clknet_3_6_0_wb_clk_i clk1_output_dest VGND VGND VPWR
+ VPWR net218 sky130_fd_sc_hd__mux2_1
XFILLER_149_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6656_ clknet_leaf_2_csclk net1466 net493 VGND VGND VPWR VPWR gpio_configure\[7\]\[9\]
+ sky130_fd_sc_hd__dfrtp_4
X_3868_ _0816_ _1424_ VGND VGND VPWR VPWR _1425_ sky130_fd_sc_hd__nor2_1
XFILLER_137_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5607_ xfer_count\[3\] _2454_ _2448_ VGND VGND VPWR VPWR _2456_ sky130_fd_sc_hd__a21boi_1
XFILLER_191_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6587_ clknet_leaf_28_csclk net574 net520 VGND VGND VPWR VPWR mgmt_gpio_data_buf\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_191_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3799_ hkspi.count\[0\] _1379_ hkspi.count\[1\] VGND VGND VPWR VPWR _1383_ sky130_fd_sc_hd__a21oi_1
XFILLER_152_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5538_ net798 net457 _2436_ VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__mux2_1
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5469_ net846 net457 _2428_ VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__mux2_1
X_7208_ clknet_leaf_75_csclk net1517 net485 VGND VGND VPWR VPWR gpio_configure\[27\]\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_132_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7139_ clknet_leaf_25_csclk net699 net518 VGND VGND VPWR VPWR gpio_configure\[37\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_86_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput18 mask_rev_in[22] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_2
XFILLER_183_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput29 mask_rev_in[3] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_109_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4840_ _1684_ _1807_ _1659_ VGND VGND VPWR VPWR _2051_ sky130_fd_sc_hd__o21ai_1
XTAP_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4771_ _1662_ net380 _1882_ VGND VGND VPWR VPWR _1983_ sky130_fd_sc_hd__a21o_1
XFILLER_14_680 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6510_ clknet_leaf_4_csclk net903 net495 VGND VGND VPWR VPWR gpio_configure\[23\]\[12\]
+ sky130_fd_sc_hd__dfrtp_2
X_3722_ _1280_ _1289_ _1298_ _1309_ VGND VGND VPWR VPWR _1310_ sky130_fd_sc_hd__or4_1
XFILLER_119_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6441_ net495 net481 VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__and2_1
XFILLER_158_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3653_ gpio_configure\[19\]\[2\] _0896_ _0928_ gpio_configure\[20\]\[2\] _1241_ VGND
+ VGND VPWR VPWR _1242_ sky130_fd_sc_hd__a221o_1
XFILLER_173_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6372_ wbbd_state\[7\] net142 net134 wbbd_state\[8\] VGND VGND VPWR VPWR _3169_ sky130_fd_sc_hd__a22o_1
X_3584_ gpio_configure\[22\]\[3\] _0923_ _0936_ net23 _1149_ VGND VGND VPWR VPWR _1174_
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5323_ net1794 net470 _2412_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__mux2_1
X_5254_ net738 net451 _2404_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__mux2_1
X_4205_ net1623 net466 _1522_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__mux2_1
X_5185_ net466 net1600 _2389_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__mux2_1
Xclkbuf_3_6_0_csclk clknet_2_3_0_csclk VGND VGND VPWR VPWR clknet_3_6_0_csclk sky130_fd_sc_hd__clkbuf_8
XFILLER_68_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4136_ net1800 net466 _1512_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__mux2_1
XFILLER_113_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4067_ net954 _1488_ _1481_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__mux2_1
XFILLER_71_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4969_ _2176_ _2177_ VGND VGND VPWR VPWR _2179_ sky130_fd_sc_hd__nand2_1
XFILLER_149_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6708_ clknet_leaf_3_csclk net1982 net494 VGND VGND VPWR VPWR gpio_configure\[15\]\[10\]
+ sky130_fd_sc_hd__dfstp_4
XFILLER_20_661 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6639_ clknet_3_4_0_wb_clk_i _0252_ VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__dfxtp_1
XFILLER_164_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6990_ clknet_leaf_17_csclk net1269 net512 VGND VGND VPWR VPWR gpio_configure\[18\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_53_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5941_ gpio_configure\[10\]\[11\] net421 _2540_ gpio_configure\[12\]\[11\] VGND VGND
+ VPWR VPWR _2765_ sky130_fd_sc_hd__a22o_1
XFILLER_18_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5872_ gpio_configure\[16\]\[8\] net472 VGND VGND VPWR VPWR _2699_ sky130_fd_sc_hd__or2_1
XFILLER_34_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4823_ _1691_ _1883_ _2033_ _1989_ VGND VGND VPWR VPWR _2034_ sky130_fd_sc_hd__or4b_1
XFILLER_166_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4754_ _1646_ _1750_ VGND VGND VPWR VPWR _1966_ sky130_fd_sc_hd__nor2_1
XFILLER_193_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3705_ gpio_configure\[31\]\[9\] _1041_ _1051_ gpio_configure\[35\]\[9\] _1292_ VGND
+ VGND VPWR VPWR _1293_ sky130_fd_sc_hd__a221o_1
XFILLER_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4685_ _1693_ _1782_ _1884_ VGND VGND VPWR VPWR _1897_ sky130_fd_sc_hd__o21ai_1
XFILLER_134_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3636_ net22 _0936_ _1054_ gpio_configure\[19\]\[10\] VGND VGND VPWR VPWR _1225_
+ sky130_fd_sc_hd__a22o_1
X_6424_ net495 net481 VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__and2_1
XFILLER_146_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6355_ net2023 _1004_ _3156_ VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__mux2_1
X_3567_ gpio_configure\[13\]\[11\] _1045_ _1068_ gpio_configure\[10\]\[11\] VGND VGND
+ VPWR VPWR _1157_ sky130_fd_sc_hd__a22o_1
XFILLER_115_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5306_ net463 net878 _2410_ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__mux2_1
X_6286_ gpio_configure\[2\]\[10\] net398 _2843_ gpio_configure\[5\]\[10\] _3097_ VGND
+ VGND VPWR VPWR _3098_ sky130_fd_sc_hd__a221o_1
XFILLER_115_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3498_ gpio_configure\[25\]\[4\] _0927_ _1086_ gpio_configure\[29\]\[12\] _1088_
+ VGND VGND VPWR VPWR _1089_ sky130_fd_sc_hd__a221o_1
XFILLER_88_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5237_ net618 net1909 _2402_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__mux2_1
XFILLER_124_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_683 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5168_ net1965 _1529_ _2364_ _2374_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__a211o_1
XFILLER_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4119_ net573 net1904 net630 VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__mux2_1
XFILLER_83_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5099_ _1589_ _1591_ _1598_ _1819_ _2040_ VGND VGND VPWR VPWR _2308_ sky130_fd_sc_hd__a311o_1
XFILLER_56_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold7 net2059 VGND VGND VPWR VPWR net540 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_87_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_30_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire360 net361 VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__clkbuf_2
X_4470_ _1654_ _1662_ VGND VGND VPWR VPWR _1682_ sky130_fd_sc_hd__nand2_1
Xhold407 gpio_configure\[19\]\[1\] VGND VGND VPWR VPWR net940 sky130_fd_sc_hd__dlygate4sd3_1
Xhold418 _0175_ VGND VGND VPWR VPWR net951 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3421_ gpio_configure\[32\]\[5\] _0890_ net369 gpio_configure\[25\]\[5\] _1012_ VGND
+ VGND VPWR VPWR _1013_ sky130_fd_sc_hd__a221o_2
Xhold429 gpio_configure\[21\]\[3\] VGND VGND VPWR VPWR net962 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6140_ gpio_configure\[31\]\[4\] net423 net415 gpio_configure\[11\]\[4\] VGND VGND
+ VPWR VPWR _2958_ sky130_fd_sc_hd__a22o_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3352_ net60 _0871_ net352 gpio_configure\[36\]\[7\] _0947_ VGND VGND VPWR VPWR _0948_
+ sky130_fd_sc_hd__a221o_4
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ net475 net2040 _2891_ VGND VGND VPWR VPWR _2892_ sky130_fd_sc_hd__a21o_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283_ _0878_ VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__inv_6
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1107 net284 VGND VGND VPWR VPWR net1640 sky130_fd_sc_hd__dlygate4sd3_1
X_5022_ _1850_ _2226_ _2231_ VGND VGND VPWR VPWR _2232_ sky130_fd_sc_hd__o21ai_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1118 _0345_ VGND VGND VPWR VPWR net1651 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1129 gpio_configure\[1\]\[10\] VGND VGND VPWR VPWR net1662 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6973_ clknet_leaf_37_csclk net1193 net522 VGND VGND VPWR VPWR gpio_configure\[16\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_5924_ gpio_configure\[0\]\[10\] _2526_ _2738_ _2748_ net473 VGND VGND VPWR VPWR
+ _2749_ sky130_fd_sc_hd__o221a_1
XFILLER_22_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5855_ gpio_configure\[6\]\[7\] _2490_ _2541_ gpio_configure\[31\]\[7\] VGND VGND
+ VPWR VPWR _2683_ sky130_fd_sc_hd__a22o_1
XFILLER_167_706 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4806_ _1744_ _1771_ _1818_ _1786_ VGND VGND VPWR VPWR _2017_ sky130_fd_sc_hd__a31o_1
XFILLER_167_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5786_ gpio_configure\[7\]\[4\] _2528_ _2538_ gpio_configure\[1\]\[4\] _2607_ VGND
+ VGND VPWR VPWR _2617_ sky130_fd_sc_hd__a221o_1
XFILLER_166_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4737_ _1633_ _1937_ VGND VGND VPWR VPWR _1949_ sky130_fd_sc_hd__nand2_1
XFILLER_119_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4668_ _1592_ _1613_ VGND VGND VPWR VPWR _1880_ sky130_fd_sc_hd__or2_2
XFILLER_107_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3619_ net45 _0904_ _0913_ gpio_configure\[7\]\[2\] _1207_ VGND VGND VPWR VPWR _1208_
+ sky130_fd_sc_hd__a221o_1
XFILLER_162_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6407_ net513 net483 VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__and2_1
Xhold930 gpio_configure\[14\]\[9\] VGND VGND VPWR VPWR net1463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold941 _0144_ VGND VGND VPWR VPWR net1474 sky130_fd_sc_hd__dlygate4sd3_1
X_4599_ _1789_ _1810_ _1794_ _1796_ VGND VGND VPWR VPWR _1811_ sky130_fd_sc_hd__or4b_1
XFILLER_190_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold952 net223 VGND VGND VPWR VPWR net1485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold963 _0415_ VGND VGND VPWR VPWR net1496 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6338_ gpio_configure\[37\]\[12\] _2806_ net416 gpio_configure\[32\]\[12\] VGND VGND
+ VPWR VPWR _3148_ sky130_fd_sc_hd__a22o_1
Xhold974 _0178_ VGND VGND VPWR VPWR net1507 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold985 gpio_configure\[21\]\[5\] VGND VGND VPWR VPWR net1518 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold996 _0514_ VGND VGND VPWR VPWR net1529 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_135_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6269_ serial_data_staging_2\[8\] _2444_ _2485_ VGND VGND VPWR VPWR _3082_ sky130_fd_sc_hd__o21ba_1
XFILLER_135_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_2_3_0_csclk clknet_1_1_1_csclk VGND VGND VPWR VPWR clknet_2_3_0_csclk sky130_fd_sc_hd__clkbuf_8
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_712 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3970_ net1718 net461 _1461_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__mux2_1
XFILLER_50_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5640_ pad_count_2\[5\] pad_count_2\[4\] VGND VGND VPWR VPWR _2478_ sky130_fd_sc_hd__and2b_4
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5571_ net352 net647 VGND VGND VPWR VPWR _2440_ sky130_fd_sc_hd__nand2_8
X_4522_ _1632_ _1665_ _1731_ _1732_ _1733_ VGND VGND VPWR VPWR _1734_ sky130_fd_sc_hd__o2111a_1
XFILLER_172_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold204 _0430_ VGND VGND VPWR VPWR net737 sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 gpio_configure\[7\]\[6\] VGND VGND VPWR VPWR net748 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold226 _0351_ VGND VGND VPWR VPWR net759 sky130_fd_sc_hd__dlygate4sd3_1
X_4453_ _1618_ _1644_ _1647_ VGND VGND VPWR VPWR _1665_ sky130_fd_sc_hd__or3_4
XFILLER_172_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold237 net2101 VGND VGND VPWR VPWR net770 sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 _0583_ VGND VGND VPWR VPWR net781 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold259 gpio_configure\[32\]\[4\] VGND VGND VPWR VPWR net792 sky130_fd_sc_hd__dlygate4sd3_1
X_3404_ gpio_configure\[14\]\[6\] _0916_ net368 gpio_configure\[9\]\[6\] _0997_ VGND
+ VGND VPWR VPWR _0998_ sky130_fd_sc_hd__a221o_1
X_7172_ clknet_3_1_0_wb_clk_i _0774_ net488 VGND VGND VPWR VPWR serial_data_staging_1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_144_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4384_ net530 _1595_ VGND VGND VPWR VPWR _1596_ sky130_fd_sc_hd__nor2_8
XFILLER_98_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6123_ gpio_configure\[36\]\[4\] net403 net402 gpio_configure\[4\]\[4\] VGND VGND
+ VPWR VPWR _2941_ sky130_fd_sc_hd__a22o_1
X_3335_ net378 net562 VGND VGND VPWR VPWR _0931_ sky130_fd_sc_hd__nor2_2
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ gpio_configure\[18\]\[1\] net399 net410 gpio_configure\[8\]\[1\] VGND VGND
+ VPWR VPWR _2875_ sky130_fd_sc_hd__a22o_1
XFILLER_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3266_ net588 net560 VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__and2b_4
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _1642_ _1648_ _1937_ _2093_ _1899_ VGND VGND VPWR VPWR _2215_ sky130_fd_sc_hd__a311o_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3197_ gpio_configure\[37\]\[3\] VGND VGND VPWR VPWR _0826_ sky130_fd_sc_hd__inv_2
XFILLER_38_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6956_ clknet_leaf_24_csclk net1657 net526 VGND VGND VPWR VPWR gpio_configure\[14\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_5907_ gpio_configure\[24\]\[10\] net418 _2534_ gpio_configure\[26\]\[10\] VGND VGND
+ VPWR VPWR _2732_ sky130_fd_sc_hd__a22o_1
X_6887_ clknet_leaf_40_csclk net1066 net516 VGND VGND VPWR VPWR gpio_configure\[5\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_167_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5838_ net2017 _2666_ _2486_ VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__mux2_1
XFILLER_22_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5769_ gpio_configure\[4\]\[3\] _2502_ _2510_ gpio_configure\[15\]\[3\] _2600_ VGND
+ VGND VPWR VPWR _2601_ sky130_fd_sc_hd__a221o_1
XFILLER_6_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold760 _0227_ VGND VGND VPWR VPWR net1293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 gpio_configure\[22\]\[4\] VGND VGND VPWR VPWR net1304 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold782 _0596_ VGND VGND VPWR VPWR net1315 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold793 net2112 VGND VGND VPWR VPWR net1326 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1460 wbbd_busy VGND VGND VPWR VPWR net1993 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1471 hkspi.ldata\[6\] VGND VGND VPWR VPWR net2004 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1482 hkspi.wrstb VGND VGND VPWR VPWR net2015 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1493 net333 VGND VGND VPWR VPWR net2026 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput309 net309 VGND VGND VPWR VPWR serial_data_2 sky130_fd_sc_hd__buf_12
XFILLER_181_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6810_ clknet_leaf_57_csclk net819 net503 VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__dfrtp_4
XFILLER_63_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6741_ clknet_leaf_75_csclk net1754 net488 VGND VGND VPWR VPWR gpio_configure\[19\]\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_50_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3953_ hkspi.pass_thru_mgmt net74 VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__and2b_4
XFILLER_189_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6672_ clknet_leaf_11_csclk net578 net511 VGND VGND VPWR VPWR gpio_configure\[10\]\[10\]
+ sky130_fd_sc_hd__dfstp_1
X_3884_ net123 net122 net131 net169 VGND VGND VPWR VPWR _1436_ sky130_fd_sc_hd__or4bb_1
XFILLER_31_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5623_ pad_count_1\[3\] _2463_ _2464_ _2467_ VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__a31o_1
XFILLER_136_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5554_ net471 net1562 _2438_ VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__mux2_1
XFILLER_144_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4505_ _1632_ _1636_ _1715_ _1716_ VGND VGND VPWR VPWR _1717_ sky130_fd_sc_hd__o211a_1
X_5485_ net469 net1688 _2430_ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__mux2_1
XFILLER_145_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4436_ _0835_ _1619_ VGND VGND VPWR VPWR _1648_ sky130_fd_sc_hd__nor2_1
Xfanout503 net504 VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__buf_4
XFILLER_120_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7155_ clknet_3_3_0_wb_clk_i _0758_ net502 VGND VGND VPWR VPWR pad_count_2\[2\] sky130_fd_sc_hd__dfrtp_2
Xfanout514 net526 VGND VGND VPWR VPWR net514 sky130_fd_sc_hd__buf_8
X_4367_ net124 _1578_ VGND VGND VPWR VPWR _1579_ sky130_fd_sc_hd__nand2_2
XFILLER_86_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout525 net526 VGND VGND VPWR VPWR net525 sky130_fd_sc_hd__buf_6
X_3318_ net376 net601 VGND VGND VPWR VPWR _0914_ sky130_fd_sc_hd__nor2_4
X_6106_ gpio_configure\[3\]\[3\] net413 net392 gpio_configure\[5\]\[3\] _2924_ VGND
+ VGND VPWR VPWR _2925_ sky130_fd_sc_hd__a221o_1
X_7086_ clknet_leaf_20_csclk net1159 net515 VGND VGND VPWR VPWR gpio_configure\[30\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_4298_ net449 net1081 _1541_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__mux2_1
XFILLER_86_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3249_ net549 net605 _0844_ VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__a21bo_1
X_6037_ gpio_configure\[35\]\[0\] net408 net405 gpio_configure\[24\]\[0\] VGND VGND
+ VPWR VPWR _2859_ sky130_fd_sc_hd__a22o_1
XFILLER_73_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6939_ clknet_leaf_47_csclk net1438 net514 VGND VGND VPWR VPWR gpio_configure\[12\]\[1\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_csclk csclk VGND VGND VPWR VPWR clknet_0_csclk sky130_fd_sc_hd__clkbuf_16
XFILLER_136_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold590 _0466_ VGND VGND VPWR VPWR net1123 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_173_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_1_0_0_csclk clknet_0_csclk VGND VGND VPWR VPWR clknet_1_0_0_csclk sky130_fd_sc_hd__clkbuf_8
XFILLER_18_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1290 _0693_ VGND VGND VPWR VPWR net1823 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5270_ net463 net886 _2406_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__mux2_1
XFILLER_99_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4221_ net444 net1218 _1524_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__mux2_1
XFILLER_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4152_ net444 net1250 _1514_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__mux2_1
XFILLER_68_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4083_ net760 net439 _0933_ VGND VGND VPWR VPWR _1497_ sky130_fd_sc_hd__mux2_1
XFILLER_68_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4985_ _1851_ _1959_ _1999_ VGND VGND VPWR VPWR _2195_ sky130_fd_sc_hd__or3_1
XFILLER_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6724_ clknet_leaf_9_csclk net680 net510 VGND VGND VPWR VPWR gpio_configure\[17\]\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_3936_ mgmt_gpio_data\[15\] user_clock clk2_output_dest VGND VGND VPWR VPWR net219
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_3_2_0_csclk clknet_2_1_0_csclk VGND VGND VPWR VPWR clknet_3_2_0_csclk sky130_fd_sc_hd__clkbuf_8
XFILLER_149_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6655_ clknet_leaf_3_csclk net1805 net493 VGND VGND VPWR VPWR gpio_configure\[7\]\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_3867_ hkspi.count\[2\] hkspi.count\[0\] hkspi.state\[0\] VGND VGND VPWR VPWR _1424_
+ sky130_fd_sc_hd__and3_1
XFILLER_31_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5606_ _2448_ _2453_ _2455_ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__and3_1
XFILLER_137_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6586_ clknet_leaf_28_csclk net631 net520 VGND VGND VPWR VPWR mgmt_gpio_data_buf\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_3798_ net2088 _1381_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__xor2_1
XFILLER_118_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5537_ net904 net463 _2436_ VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__mux2_1
XFILLER_118_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5468_ net892 net463 _2428_ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__mux2_1
XFILLER_105_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7207_ clknet_leaf_76_csclk net1503 net485 VGND VGND VPWR VPWR gpio_configure\[27\]\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_78_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4419_ net124 net110 _0833_ VGND VGND VPWR VPWR _1631_ sky130_fd_sc_hd__and3b_4
XFILLER_99_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5399_ net1238 net447 _2420_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__mux2_1
XFILLER_160_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7138_ clknet_leaf_29_csclk net981 net520 VGND VGND VPWR VPWR gpio_configure\[37\]\[3\]
+ sky130_fd_sc_hd__dfrtp_2
Xfanout366 _2486_ VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__buf_8
XFILLER_101_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_86_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7069_ clknet_leaf_33_csclk net1010 net521 VGND VGND VPWR VPWR gpio_configure\[28\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_101_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput19 mask_rev_in[23] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_1
XFILLER_6_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_182_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_260 net660 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_33_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4770_ _1899_ _1981_ _1946_ _1898_ VGND VGND VPWR VPWR _1982_ sky130_fd_sc_hd__or4b_1
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3721_ _1301_ _1304_ _1306_ _1308_ VGND VGND VPWR VPWR _1309_ sky130_fd_sc_hd__or4_1
XFILLER_158_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6440_ net495 net482 VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__and2_1
X_3652_ gpio_configure\[17\]\[2\] net367 _1062_ gpio_configure\[21\]\[10\] VGND VGND
+ VPWR VPWR _1241_ sky130_fd_sc_hd__a22o_1
XFILLER_174_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3583_ _1148_ _1154_ _1163_ _1172_ VGND VGND VPWR VPWR _1173_ sky130_fd_sc_hd__or4_2
XFILLER_127_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6371_ _3168_ net2058 _3162_ VGND VGND VPWR VPWR _0801_ sky130_fd_sc_hd__mux2_1
XFILLER_173_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5322_ _0939_ net647 VGND VGND VPWR VPWR _2412_ sky130_fd_sc_hd__and2_4
XFILLER_173_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5253_ net750 net457 _2404_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__mux2_1
X_4204_ _1122_ net425 VGND VGND VPWR VPWR _1522_ sky130_fd_sc_hd__and2_2
X_5184_ _1262_ net425 VGND VGND VPWR VPWR _2389_ sky130_fd_sc_hd__nand2_1
X_4135_ _1103_ net425 VGND VGND VPWR VPWR _1512_ sky130_fd_sc_hd__and2_1
XFILLER_29_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_63_csclk clknet_3_0_0_csclk VGND VGND VPWR VPWR clknet_leaf_63_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_113_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4066_ net1905 net439 net356 VGND VGND VPWR VPWR _1488_ sky130_fd_sc_hd__mux2_1
XFILLER_71_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_78_csclk clknet_3_0_0_csclk VGND VGND VPWR VPWR clknet_leaf_78_csclk
+ sky130_fd_sc_hd__clkbuf_16
X_4968_ _2177_ VGND VGND VPWR VPWR _2178_ sky130_fd_sc_hd__clkinv_2
XFILLER_149_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6707_ clknet_leaf_2_csclk net1476 net496 VGND VGND VPWR VPWR gpio_configure\[15\]\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_165_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3919_ mgmt_gpio_data\[36\] net89 net76 VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__mux2_2
X_4899_ _1815_ _1930_ VGND VGND VPWR VPWR _2110_ sky130_fd_sc_hd__or2_1
XFILLER_20_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6638_ clknet_leaf_4_csclk net895 net494 VGND VGND VPWR VPWR gpio_configure\[6\]\[12\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_192_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6569_ clknet_leaf_40_csclk net947 net516 VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__dfrtp_1
XFILLER_118_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_16_csclk clknet_3_5_0_csclk VGND VGND VPWR VPWR clknet_leaf_16_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_79_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5940_ gpio_configure\[29\]\[11\] _2529_ _2538_ gpio_configure\[1\]\[11\] _2763_
+ VGND VGND VPWR VPWR _2764_ sky130_fd_sc_hd__a221o_1
XFILLER_46_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5871_ gpio_configure\[6\]\[8\] _2490_ _2501_ gpio_configure\[13\]\[8\] _2697_ VGND
+ VGND VPWR VPWR _2698_ sky130_fd_sc_hd__a221o_1
XFILLER_21_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4822_ _1899_ _2032_ _2013_ _1709_ VGND VGND VPWR VPWR _2033_ sky130_fd_sc_hd__or4b_1
X_4753_ _1599_ _1651_ VGND VGND VPWR VPWR _1965_ sky130_fd_sc_hd__nor2_1
XFILLER_147_634 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3704_ gpio_configure\[16\]\[9\] _1080_ _1119_ gpio_configure\[5\]\[9\] VGND VGND
+ VPWR VPWR _1292_ sky130_fd_sc_hd__a22o_1
X_4684_ _1677_ _1792_ VGND VGND VPWR VPWR _1896_ sky130_fd_sc_hd__nand2_2
X_6423_ net495 net482 VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__and2_1
X_3635_ gpio_configure\[28\]\[2\] _0888_ _0923_ gpio_configure\[22\]\[2\] _1223_ VGND
+ VGND VPWR VPWR _1224_ sky130_fd_sc_hd__a221o_1
XFILLER_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6354_ net1955 _1039_ _3156_ VGND VGND VPWR VPWR _0796_ sky130_fd_sc_hd__mux2_1
X_3566_ net46 _0904_ _0932_ gpio_configure\[35\]\[3\] _1155_ VGND VGND VPWR VPWR _1156_
+ sky130_fd_sc_hd__a221o_1
XFILLER_115_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5305_ net471 net1564 _2410_ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__mux2_1
XFILLER_130_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3497_ net262 _1009_ _1087_ gpio_configure\[0\]\[12\] VGND VGND VPWR VPWR _1088_
+ sky130_fd_sc_hd__a22o_1
X_6285_ gpio_configure\[13\]\[10\] net417 _2862_ gpio_configure\[25\]\[10\] VGND VGND
+ VPWR VPWR _3097_ sky130_fd_sc_hd__a22o_1
XFILLER_115_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5236_ net452 net984 _2402_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__mux2_1
XFILLER_69_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5167_ _2355_ _2358_ _2373_ _2354_ VGND VGND VPWR VPWR _2374_ sky130_fd_sc_hd__a211o_1
XFILLER_29_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_695 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4118_ net439 net1905 net630 VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__mux2_1
XFILLER_56_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5098_ _1668_ _1940_ _2193_ _1827_ VGND VGND VPWR VPWR _2307_ sky130_fd_sc_hd__o211ai_1
X_4049_ net455 net1629 _1479_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__mux2_1
XFILLER_56_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_692 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold8 _1463_ VGND VGND VPWR VPWR net541 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_87_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_128_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xwire383 _0897_ VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__buf_12
Xhold408 _0598_ VGND VGND VPWR VPWR net941 sky130_fd_sc_hd__dlygate4sd3_1
Xwire394 _2840_ VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__buf_8
Xhold419 gpio_configure\[30\]\[5\] VGND VGND VPWR VPWR net952 sky130_fd_sc_hd__dlygate4sd3_1
X_3420_ net288 _0886_ _0923_ gpio_configure\[22\]\[5\] VGND VGND VPWR VPWR _1012_
+ sky130_fd_sc_hd__a22o_1
XFILLER_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3351_ gpio_configure\[34\]\[7\] net358 _0911_ gpio_configure\[21\]\[7\] VGND VGND
+ VPWR VPWR _0947_ sky130_fd_sc_hd__a22o_1
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6070_ gpio_configure\[0\]\[1\] _2851_ _2890_ net473 VGND VGND VPWR VPWR _2891_ sky130_fd_sc_hd__o211a_1
X_3282_ net607 net599 VGND VGND VPWR VPWR _0878_ sky130_fd_sc_hd__nand2_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1108 _0098_ VGND VGND VPWR VPWR net1641 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5021_ _1592_ net432 _1866_ VGND VGND VPWR VPWR _2231_ sky130_fd_sc_hd__or3_1
XFILLER_112_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1119 gpio_configure\[36\]\[2\] VGND VGND VPWR VPWR net1652 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6972_ clknet_leaf_23_csclk net1353 net514 VGND VGND VPWR VPWR gpio_configure\[16\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_19_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5923_ _2740_ _2743_ _2745_ _2747_ VGND VGND VPWR VPWR _2748_ sky130_fd_sc_hd__or4_1
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5854_ gpio_configure\[18\]\[7\] _2532_ _2537_ gpio_configure\[17\]\[7\] _2681_ VGND
+ VGND VPWR VPWR _2682_ sky130_fd_sc_hd__a221o_1
XFILLER_110_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4805_ net477 _1757_ net424 _1651_ _1745_ VGND VGND VPWR VPWR _2016_ sky130_fd_sc_hd__o32a_1
XFILLER_167_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5785_ _2609_ _2611_ _2613_ _2615_ VGND VGND VPWR VPWR _2616_ sky130_fd_sc_hd__or4_1
XFILLER_166_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4736_ _1599_ _1668_ VGND VGND VPWR VPWR _1948_ sky130_fd_sc_hd__nor2_1
XFILLER_159_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4667_ _1555_ _1591_ _0833_ VGND VGND VPWR VPWR _1879_ sky130_fd_sc_hd__and3b_1
XFILLER_134_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6406_ net513 net483 VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__and2_1
Xhold920 gpio_configure\[31\]\[6\] VGND VGND VPWR VPWR net1453 sky130_fd_sc_hd__dlygate4sd3_1
X_3618_ gpio_configure\[36\]\[2\] net352 _1051_ gpio_configure\[35\]\[10\] VGND VGND
+ VPWR VPWR _1207_ sky130_fd_sc_hd__a22o_1
XFILLER_162_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold931 _0305_ VGND VGND VPWR VPWR net1464 sky130_fd_sc_hd__dlygate4sd3_1
X_4598_ _1799_ _1802_ _1806_ _1809_ VGND VGND VPWR VPWR _1810_ sky130_fd_sc_hd__or4_1
Xhold942 gpio_configure\[15\]\[9\] VGND VGND VPWR VPWR net1475 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold953 _0166_ VGND VGND VPWR VPWR net1486 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6337_ gpio_configure\[13\]\[12\] net417 net394 gpio_configure\[6\]\[12\] VGND VGND
+ VPWR VPWR _3147_ sky130_fd_sc_hd__a22o_1
Xhold964 gpio_configure\[12\]\[8\] VGND VGND VPWR VPWR net1497 sky130_fd_sc_hd__dlygate4sd3_1
X_3549_ net38 net353 _1081_ gpio_configure\[34\]\[11\] VGND VGND VPWR VPWR _1139_
+ sky130_fd_sc_hd__a22o_1
Xhold975 net222 VGND VGND VPWR VPWR net1508 sky130_fd_sc_hd__dlygate4sd3_1
Xhold986 _0618_ VGND VGND VPWR VPWR net1519 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold997 gpio_configure\[1\]\[5\] VGND VGND VPWR VPWR net1530 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6268_ gpio_configure\[0\]\[9\] _2851_ _3070_ _3080_ net473 VGND VGND VPWR VPWR _3081_
+ sky130_fd_sc_hd__o221a_1
XFILLER_135_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5219_ net437 net1409 _2397_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__mux2_1
XFILLER_76_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6199_ gpio_configure\[26\]\[7\] _2810_ net413 gpio_configure\[3\]\[7\] VGND VGND
+ VPWR VPWR _3014_ sky130_fd_sc_hd__a22o_1
XFILLER_130_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_180_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_75_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5570_ net435 net926 net648 VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__mux2_1
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4521_ _1662_ _1667_ VGND VGND VPWR VPWR _1733_ sky130_fd_sc_hd__nand2_1
XFILLER_144_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold205 gpio_configure\[0\]\[3\] VGND VGND VPWR VPWR net738 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_172_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold216 _0507_ VGND VGND VPWR VPWR net749 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4452_ _1617_ _1622_ _1628_ _1662_ VGND VGND VPWR VPWR _1664_ sky130_fd_sc_hd__nand4_1
Xhold227 net2115 VGND VGND VPWR VPWR net760 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold238 _0194_ VGND VGND VPWR VPWR net771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 gpio_configure\[28\]\[2\] VGND VGND VPWR VPWR net782 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_618 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3403_ gpio_configure\[5\]\[6\] _0914_ _0974_ net309 VGND VGND VPWR VPWR _0997_ sky130_fd_sc_hd__a22o_1
X_7171_ clknet_3_1_0_wb_clk_i _0773_ net488 VGND VGND VPWR VPWR serial_data_staging_1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_4383_ net110 net124 VGND VGND VPWR VPWR _1595_ sky130_fd_sc_hd__nand2_2
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6122_ net2039 _2940_ net366 VGND VGND VPWR VPWR _0780_ sky130_fd_sc_hd__mux2_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3334_ net381 net609 VGND VGND VPWR VPWR _0930_ sky130_fd_sc_hd__nor2_4
XFILLER_124_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6053_ gpio_configure\[20\]\[1\] net396 _2861_ gpio_configure\[28\]\[1\] _2870_ VGND
+ VGND VPWR VPWR _2874_ sky130_fd_sc_hd__a221o_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3265_ net559 net2005 net474 VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__mux2_4
XFILLER_105_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _1596_ net380 _1883_ VGND VGND VPWR VPWR _2214_ sky130_fd_sc_hd__a21o_1
XFILLER_38_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3196_ xfer_state\[2\] VGND VGND VPWR VPWR _0825_ sky130_fd_sc_hd__clkinv_2
XFILLER_38_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6955_ clknet_leaf_19_csclk net871 net510 VGND VGND VPWR VPWR gpio_configure\[14\]\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_41_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5906_ gpio_configure\[14\]\[10\] _2494_ _2502_ gpio_configure\[4\]\[10\] _2730_
+ VGND VGND VPWR VPWR _2731_ sky130_fd_sc_hd__a221o_1
XFILLER_22_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6886_ clknet_leaf_15_csclk net1181 net513 VGND VGND VPWR VPWR gpio_configure\[5\]\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_22_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5837_ net475 serial_data_staging_1\[5\] _2665_ VGND VGND VPWR VPWR _2666_ sky130_fd_sc_hd__a21o_1
XFILLER_10_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5768_ gpio_configure\[16\]\[3\] net419 _2534_ gpio_configure\[26\]\[3\] _2525_ VGND
+ VGND VPWR VPWR _2600_ sky130_fd_sc_hd__a221o_1
X_4719_ _1593_ _1779_ VGND VGND VPWR VPWR _1931_ sky130_fd_sc_hd__nor2_1
XFILLER_108_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5699_ pad_count_1\[4\] _2489_ _2504_ VGND VGND VPWR VPWR _2534_ sky130_fd_sc_hd__and3_4
XFILLER_107_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold750 _0361_ VGND VGND VPWR VPWR net1283 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold761 gpio_configure\[26\]\[11\] VGND VGND VPWR VPWR net1294 sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 _0625_ VGND VGND VPWR VPWR net1305 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap480 _1587_ VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__clkbuf_2
Xhold783 net2104 VGND VGND VPWR VPWR net1316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold794 _0193_ VGND VGND VPWR VPWR net1327 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1450 net338 VGND VGND VPWR VPWR net1983 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1461 _1468_ VGND VGND VPWR VPWR net1994 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1472 wbbd_addr\[0\] VGND VGND VPWR VPWR net2005 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1483 net337 VGND VGND VPWR VPWR net2016 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1494 serial_data_staging_2\[2\] VGND VGND VPWR VPWR net2027 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_51_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6740_ clknet_leaf_18_csclk net1165 net510 VGND VGND VPWR VPWR gpio_configure\[35\]\[12\]
+ sky130_fd_sc_hd__dfrtp_2
X_3952_ hkspi.pass_thru_mgmt_delay net73 VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__and2b_4
XFILLER_189_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6671_ clknet_leaf_5_csclk net1428 net494 VGND VGND VPWR VPWR gpio_configure\[10\]\[9\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_189_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3883_ net114 net113 VGND VGND VPWR VPWR _1435_ sky130_fd_sc_hd__or2_1
X_5622_ pad_count_1\[3\] _2464_ VGND VGND VPWR VPWR _2467_ sky130_fd_sc_hd__nor2_1
XFILLER_149_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5553_ net358 net647 VGND VGND VPWR VPWR _2438_ sky130_fd_sc_hd__nand2_8
XFILLER_157_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_144_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4504_ _1637_ _1669_ _1672_ VGND VGND VPWR VPWR _1716_ sky130_fd_sc_hd__and3_1
X_5484_ _0924_ net427 VGND VGND VPWR VPWR _2430_ sky130_fd_sc_hd__nand2_8
XFILLER_144_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4435_ _1624_ _1626_ VGND VGND VPWR VPWR _1647_ sky130_fd_sc_hd__nand2_2
XFILLER_160_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7154_ clknet_3_3_0_wb_clk_i _0757_ net500 VGND VGND VPWR VPWR pad_count_2\[1\] sky130_fd_sc_hd__dfstp_1
Xfanout504 net508 VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__buf_8
Xfanout515 net526 VGND VGND VPWR VPWR net515 sky130_fd_sc_hd__buf_4
X_4366_ _1577_ VGND VGND VPWR VPWR _1578_ sky130_fd_sc_hd__inv_2
Xfanout526 net527 VGND VGND VPWR VPWR net526 sky130_fd_sc_hd__buf_12
XFILLER_59_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_113_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6105_ gpio_configure\[1\]\[3\] net401 _2810_ gpio_configure\[26\]\[3\] VGND VGND
+ VPWR VPWR _2924_ sky130_fd_sc_hd__a22o_1
XFILLER_59_738 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3317_ net554 _0881_ VGND VGND VPWR VPWR _0913_ sky130_fd_sc_hd__nor2_8
X_7085_ clknet_leaf_29_csclk net973 net524 VGND VGND VPWR VPWR gpio_configure\[30\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_4297_ net455 net1632 _1541_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__mux2_1
XFILLER_86_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6036_ _2478_ _2793_ _2809_ VGND VGND VPWR VPWR _2858_ sky130_fd_sc_hd__and3_4
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3248_ net636 _0819_ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__nand2_1
XFILLER_27_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_100_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6938_ clknet_leaf_15_csclk net1980 net519 VGND VGND VPWR VPWR gpio_configure\[12\]\[0\]
+ sky130_fd_sc_hd__dfstp_4
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6869_ clknet_leaf_37_csclk net1201 net522 VGND VGND VPWR VPWR gpio_configure\[3\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_10_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_123_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold580 _0353_ VGND VGND VPWR VPWR net1113 sky130_fd_sc_hd__dlygate4sd3_1
Xhold591 net277 VGND VGND VPWR VPWR net1124 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1280 _0278_ VGND VGND VPWR VPWR net1813 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1291 gpio_configure\[33\]\[8\] VGND VGND VPWR VPWR net1824 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_146_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4220_ net450 net1222 _1524_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__mux2_1
XFILLER_68_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4151_ net450 net1292 _1514_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__mux2_1
XFILLER_68_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4082_ net936 _1496_ _1490_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__mux2_1
XFILLER_83_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4984_ _1794_ _1966_ _2009_ VGND VGND VPWR VPWR _2194_ sky130_fd_sc_hd__or3_1
XFILLER_51_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6723_ clknet_leaf_9_csclk net755 net509 VGND VGND VPWR VPWR gpio_configure\[17\]\[10\]
+ sky130_fd_sc_hd__dfstp_2
X_3935_ _0830_ net2 net1 VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__mux2_4
XFILLER_149_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6654_ clknet_3_4_0_wb_clk_i _0267_ VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__dfxtp_1
X_3866_ net58 net2045 _1417_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__mux2_1
X_5605_ _2454_ VGND VGND VPWR VPWR _2455_ sky130_fd_sc_hd__clkinv_2
X_6585_ clknet_leaf_27_csclk net661 net519 VGND VGND VPWR VPWR mgmt_gpio_data_buf\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_3797_ hkspi.count\[2\] hkspi.count\[1\] VGND VGND VPWR VPWR _1382_ sky130_fd_sc_hd__and2_1
XFILLER_176_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5536_ net1713 net469 _2436_ VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__mux2_1
XFILLER_145_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5467_ net1717 net469 _2428_ VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__mux2_1
X_7206_ clknet_3_6_0_wb_clk_i net2072 net529 VGND VGND VPWR VPWR wbbd_write sky130_fd_sc_hd__dfrtp_1
X_4418_ _1612_ _1629_ VGND VGND VPWR VPWR _1630_ sky130_fd_sc_hd__nand2_1
X_5398_ net1192 net453 _2420_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__mux2_1
XFILLER_120_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7137_ clknet_leaf_64_csclk net857 net508 VGND VGND VPWR VPWR gpio_configure\[37\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4349_ _1552_ _1559_ net111 VGND VGND VPWR VPWR _1561_ sky130_fd_sc_hd__a21o_1
XFILLER_86_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7068_ clknet_leaf_65_csclk net783 net505 VGND VGND VPWR VPWR gpio_configure\[28\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_86_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6019_ _1447_ _2818_ VGND VGND VPWR VPWR _2841_ sky130_fd_sc_hd__nor2_4
XFILLER_100_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_250 clk2_output_dest VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_261 _0933_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3720_ gpio_configure\[3\]\[1\] _0915_ _1129_ gpio_configure\[11\]\[9\] _1307_ VGND
+ VGND VPWR VPWR _1308_ sky130_fd_sc_hd__a221o_1
XFILLER_119_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_173_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3651_ _1233_ _1235_ _1237_ _1239_ VGND VGND VPWR VPWR _1240_ sky130_fd_sc_hd__or4_1
XFILLER_158_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6370_ wbbd_state\[9\] net150 net154 net433 _3167_ VGND VGND VPWR VPWR _3168_ sky130_fd_sc_hd__a221o_1
X_3582_ _1165_ _1167_ _1169_ _1171_ VGND VGND VPWR VPWR _1172_ sky130_fd_sc_hd__or4_1
XFILLER_127_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5321_ net435 net1069 net556 VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__mux2_1
XFILLER_142_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5252_ net880 net463 _2404_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__mux2_1
XFILLER_142_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4203_ net898 net444 _1521_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__mux2_1
XFILLER_68_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5183_ _2378_ _2381_ _2388_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__or3_1
XFILLER_3_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4134_ net996 net443 _1511_ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__mux2_1
XFILLER_68_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4065_ net1489 _1487_ _1481_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__mux2_1
XFILLER_83_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4967_ _1772_ _1777_ _1779_ _2008_ _2087_ VGND VGND VPWR VPWR _2177_ sky130_fd_sc_hd__o311a_1
X_6706_ clknet_leaf_3_csclk net1803 net496 VGND VGND VPWR VPWR gpio_configure\[15\]\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_3918_ mgmt_gpio_data\[37\] net91 net76 VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__mux2_4
XFILLER_20_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4898_ _1950_ _2084_ _2086_ _2108_ _1939_ VGND VGND VPWR VPWR _2109_ sky130_fd_sc_hd__o41a_1
XFILLER_177_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6637_ clknet_leaf_5_csclk net1227 net494 VGND VGND VPWR VPWR gpio_configure\[6\]\[11\]
+ sky130_fd_sc_hd__dfrtp_4
X_3849_ hkspi.count\[2\] hkspi.count\[1\] hkspi.state\[0\] _1415_ VGND VGND VPWR VPWR
+ _1416_ sky130_fd_sc_hd__o211a_1
XFILLER_192_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6568_ clknet_leaf_40_csclk net1541 net516 VGND VGND VPWR VPWR mgmt_gpio_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5519_ net434 net1290 _2433_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__mux2_1
XFILLER_118_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6499_ clknet_leaf_47_csclk net1432 net514 VGND VGND VPWR VPWR gpio_configure\[31\]\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_105_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_168_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5870_ gpio_configure\[22\]\[8\] _2498_ _2499_ gpio_configure\[20\]\[8\] VGND VGND
+ VPWR VPWR _2697_ sky130_fd_sc_hd__a22o_1
X_4821_ _1998_ _2029_ _2030_ _2031_ VGND VGND VPWR VPWR _2032_ sky130_fd_sc_hd__or4_1
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_178_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4752_ _1651_ _1750_ VGND VGND VPWR VPWR _1964_ sky130_fd_sc_hd__nor2_1
X_3703_ gpio_configure\[0\]\[1\] _0898_ _1094_ gpio_configure\[7\]\[9\] _1290_ VGND
+ VGND VPWR VPWR _1291_ sky130_fd_sc_hd__a221o_1
XFILLER_119_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_646 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4683_ _1757_ _1874_ VGND VGND VPWR VPWR _1895_ sky130_fd_sc_hd__or2_1
X_6422_ net495 net482 VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__and2_1
X_3634_ gpio_configure\[27\]\[2\] net370 _1086_ gpio_configure\[29\]\[10\] VGND VGND
+ VPWR VPWR _1223_ sky130_fd_sc_hd__a22o_1
X_6353_ net1983 clknet_1_0__leaf__1134_ _3156_ VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__mux2_1
X_3565_ gpio_configure\[35\]\[11\] _1051_ _1121_ gpio_configure\[17\]\[11\] VGND VGND
+ VPWR VPWR _1155_ sky130_fd_sc_hd__a22o_1
XFILLER_161_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5304_ net357 net429 VGND VGND VPWR VPWR _2410_ sky130_fd_sc_hd__nand2_8
X_6284_ gpio_configure\[10\]\[10\] net414 net394 gpio_configure\[6\]\[10\] _3095_
+ VGND VGND VPWR VPWR _3096_ sky130_fd_sc_hd__a221o_1
X_3496_ net383 _0909_ VGND VGND VPWR VPWR _1087_ sky130_fd_sc_hd__nor2_4
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5235_ net458 net1614 _2402_ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__mux2_1
XFILLER_69_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5166_ _2333_ _2370_ _2372_ _2367_ VGND VGND VPWR VPWR _2373_ sky130_fd_sc_hd__a31oi_2
XFILLER_68_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4117_ net660 net1903 net630 VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__mux2_1
X_5097_ _1706_ _1994_ _2305_ VGND VGND VPWR VPWR _2306_ sky130_fd_sc_hd__a21o_1
XFILLER_83_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4048_ net461 net1619 _1479_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__mux2_1
XFILLER_71_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_84_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5999_ gpio_configure\[18\]\[0\] net399 _2820_ gpio_configure\[21\]\[0\] _2817_ VGND
+ VGND VPWR VPWR _2821_ sky130_fd_sc_hd__a221o_1
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_149_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput290 net290 VGND VGND VPWR VPWR pll_trim[23] sky130_fd_sc_hd__buf_12
Xhold9 net538 VGND VGND VPWR VPWR net542 sky130_fd_sc_hd__buf_6
XFILLER_47_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_101_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_62_csclk clknet_3_2_0_csclk VGND VGND VPWR VPWR clknet_leaf_62_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_116_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire362 net363 VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__clkbuf_2
XFILLER_128_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold409 mgmt_gpio_data\[6\] VGND VGND VPWR VPWR net942 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_183_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3350_ net10 _0891_ net353 net42 _0945_ VGND VGND VPWR VPWR _0946_ sky130_fd_sc_hd__a221o_1
XFILLER_124_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_77_csclk clknet_3_0_0_csclk VGND VGND VPWR VPWR clknet_leaf_77_csclk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ net551 net638 net627 VGND VGND VPWR VPWR _0877_ sky130_fd_sc_hd__or3_4
XFILLER_97_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ net477 _1608_ _2130_ VGND VGND VPWR VPWR _2230_ sky130_fd_sc_hd__o21ai_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1109 gpio_configure\[0\]\[0\] VGND VGND VPWR VPWR net1642 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_65_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6971_ clknet_leaf_21_csclk net1382 net514 VGND VGND VPWR VPWR gpio_configure\[16\]\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_53_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5922_ gpio_configure\[5\]\[10\] _2496_ net421 gpio_configure\[10\]\[10\] _2746_
+ VGND VGND VPWR VPWR _2747_ sky130_fd_sc_hd__a221o_2
XFILLER_179_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5853_ gpio_configure\[19\]\[7\] _2491_ _2505_ gpio_configure\[11\]\[7\] VGND VGND
+ VPWR VPWR _2681_ sky130_fd_sc_hd__a22o_1
XFILLER_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_15_csclk clknet_3_5_0_csclk VGND VGND VPWR VPWR clknet_leaf_15_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_22_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4804_ _1601_ _1781_ _1834_ _1958_ VGND VGND VPWR VPWR _2015_ sky130_fd_sc_hd__a31o_1
X_5784_ gpio_configure\[4\]\[4\] _2502_ _2510_ gpio_configure\[15\]\[4\] _2614_ VGND
+ VGND VPWR VPWR _2615_ sky130_fd_sc_hd__a221o_1
XFILLER_166_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4735_ _1598_ _1629_ VGND VGND VPWR VPWR _1947_ sky130_fd_sc_hd__nand2_1
XFILLER_147_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4666_ _1588_ _1776_ VGND VGND VPWR VPWR _1878_ sky130_fd_sc_hd__nor2_1
XFILLER_119_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6405_ net513 net483 VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__and2_1
X_3617_ gpio_configure\[18\]\[2\] net374 _1125_ gpio_configure\[22\]\[10\] VGND VGND
+ VPWR VPWR _1206_ sky130_fd_sc_hd__a22o_1
Xhold910 gpio_configure\[24\]\[6\] VGND VGND VPWR VPWR net1443 sky130_fd_sc_hd__dlygate4sd3_1
Xhold921 _0126_ VGND VGND VPWR VPWR net1454 sky130_fd_sc_hd__dlygate4sd3_1
X_4597_ _1774_ net432 _1807_ VGND VGND VPWR VPWR _1809_ sky130_fd_sc_hd__a21oi_1
Xhold932 gpio_configure\[7\]\[9\] VGND VGND VPWR VPWR net1465 sky130_fd_sc_hd__dlygate4sd3_1
Xhold943 _0310_ VGND VGND VPWR VPWR net1476 sky130_fd_sc_hd__dlygate4sd3_1
X_6336_ gpio_configure\[14\]\[12\] net411 _2861_ gpio_configure\[28\]\[12\] _3145_
+ VGND VGND VPWR VPWR _3146_ sky130_fd_sc_hd__a221o_1
Xhold954 gpio_configure\[10\]\[8\] VGND VGND VPWR VPWR net1487 sky130_fd_sc_hd__dlygate4sd3_1
X_3548_ gpio_configure\[11\]\[3\] _0907_ _0921_ gpio_configure\[12\]\[3\] VGND VGND
+ VPWR VPWR _1138_ sky130_fd_sc_hd__a22o_1
Xhold965 _0294_ VGND VGND VPWR VPWR net1498 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold976 _0165_ VGND VGND VPWR VPWR net1509 sky130_fd_sc_hd__dlygate4sd3_1
Xhold987 gpio_configure\[35\]\[5\] VGND VGND VPWR VPWR net1520 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_142_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold998 _0458_ VGND VGND VPWR VPWR net1531 sky130_fd_sc_hd__dlygate4sd3_1
X_6267_ net359 _3072_ _3079_ VGND VGND VPWR VPWR _3080_ sky130_fd_sc_hd__or3_1
XFILLER_88_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3479_ gpio_configure\[10\]\[12\] _1068_ _1069_ gpio_configure\[14\]\[12\] VGND VGND
+ VPWR VPWR _1070_ sky130_fd_sc_hd__a22o_1
XFILLER_130_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5218_ net660 net784 _2397_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__mux2_1
XFILLER_57_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6198_ gpio_configure\[30\]\[7\] _2799_ net408 gpio_configure\[35\]\[7\] VGND VGND
+ VPWR VPWR _3013_ sky130_fd_sc_hd__a22o_1
Xhold1610 mgmt_gpio_data\[32\] VGND VGND VPWR VPWR net2143 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5149_ _1596_ _1658_ _1738_ _1961_ _2207_ VGND VGND VPWR VPWR _2356_ sky130_fd_sc_hd__a2111o_1
XFILLER_151_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4520_ _1613_ _1665_ VGND VGND VPWR VPWR _1732_ sky130_fd_sc_hd__or2_1
XFILLER_156_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold206 _0448_ VGND VGND VPWR VPWR net739 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4451_ _0833_ _1596_ VGND VGND VPWR VPWR _1663_ sky130_fd_sc_hd__nand2_2
Xhold217 gpio_configure\[0\]\[2\] VGND VGND VPWR VPWR net750 sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 _0207_ VGND VGND VPWR VPWR net761 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold239 gpio_configure\[19\]\[2\] VGND VGND VPWR VPWR net772 sky130_fd_sc_hd__dlygate4sd3_1
X_3402_ gpio_configure\[0\]\[6\] _0898_ _0904_ net50 _0995_ VGND VGND VPWR VPWR _0996_
+ sky130_fd_sc_hd__a221o_1
X_7170_ clknet_3_1_0_wb_clk_i _0772_ net488 VGND VGND VPWR VPWR serial_data_staging_1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_4382_ _1588_ _1593_ VGND VGND VPWR VPWR _1594_ sky130_fd_sc_hd__nor2_1
XFILLER_171_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6121_ net475 net2027 _2939_ VGND VGND VPWR VPWR _2940_ sky130_fd_sc_hd__a21o_1
XFILLER_98_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3333_ net629 _0881_ VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__nor2_2
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6052_ gpio_configure\[29\]\[1\] _2816_ _2820_ gpio_configure\[21\]\[1\] _2872_ VGND
+ VGND VPWR VPWR _2873_ sky130_fd_sc_hd__a221o_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3264_ net558 net58 hkspi.state\[3\] VGND VGND VPWR VPWR _0860_ sky130_fd_sc_hd__mux2_1
XFILLER_100_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _1655_ _2203_ VGND VGND VPWR VPWR _2213_ sky130_fd_sc_hd__nor2_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3195_ net475 VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__inv_6
XFILLER_39_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6954_ clknet_leaf_17_csclk net1766 net512 VGND VGND VPWR VPWR gpio_configure\[14\]\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_41_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5905_ gpio_configure\[9\]\[10\] _2512_ _2529_ gpio_configure\[29\]\[10\] VGND VGND
+ VPWR VPWR _2730_ sky130_fd_sc_hd__a22o_1
X_6885_ clknet_leaf_36_csclk net999 net522 VGND VGND VPWR VPWR gpio_configure\[5\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5836_ gpio_configure\[0\]\[6\] _2526_ _2654_ _2664_ net473 VGND VGND VPWR VPWR _2665_
+ sky130_fd_sc_hd__o221a_1
XFILLER_167_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5767_ gpio_configure\[22\]\[3\] _2498_ _2518_ gpio_configure\[3\]\[3\] _2587_ VGND
+ VGND VPWR VPWR _2599_ sky130_fd_sc_hd__a221o_1
X_4718_ _1576_ _1775_ VGND VGND VPWR VPWR _1930_ sky130_fd_sc_hd__nor2_1
X_5698_ gpio_configure\[24\]\[0\] net418 _2532_ gpio_configure\[18\]\[0\] VGND VGND
+ VPWR VPWR _2533_ sky130_fd_sc_hd__a22o_1
XFILLER_147_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4649_ _1593_ _1782_ _1526_ VGND VGND VPWR VPWR _1861_ sky130_fd_sc_hd__o21ai_1
XFILLER_190_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold740 _0660_ VGND VGND VPWR VPWR net1273 sky130_fd_sc_hd__dlygate4sd3_1
Xhold751 gpio_configure\[10\]\[4\] VGND VGND VPWR VPWR net1284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold762 _0161_ VGND VGND VPWR VPWR net1295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold773 gpio_configure\[3\]\[4\] VGND VGND VPWR VPWR net1306 sky130_fd_sc_hd__dlygate4sd3_1
X_6319_ net2041 _3129_ net366 VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__mux2_1
XFILLER_115_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold784 _0195_ VGND VGND VPWR VPWR net1317 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold795 gpio_configure\[26\]\[1\] VGND VGND VPWR VPWR net1328 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1440 _1062_ VGND VGND VPWR VPWR net1973 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1451 gpio_configure\[8\]\[10\] VGND VGND VPWR VPWR net1984 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1462 hkspi.ldata\[3\] VGND VGND VPWR VPWR net1995 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1473 _0880_ VGND VGND VPWR VPWR net2006 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1484 serial_data_staging_1\[6\] VGND VGND VPWR VPWR net2017 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_176_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1495 _0779_ VGND VGND VPWR VPWR net2028 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_765 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3951_ net85 net58 hkspi.pass_thru_mgmt_delay VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__mux2_2
XFILLER_50_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6670_ clknet_leaf_11_csclk net1488 net511 VGND VGND VPWR VPWR gpio_configure\[10\]\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_3882_ net112 net111 VGND VGND VPWR VPWR _1434_ sky130_fd_sc_hd__and2_1
X_5621_ pad_count_1\[3\] pad_count_1\[2\] VGND VGND VPWR VPWR _2466_ sky130_fd_sc_hd__nor2_2
X_5552_ net434 net1033 _2437_ VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__mux2_1
XFILLER_191_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4503_ _1714_ _1697_ _1630_ _1711_ VGND VGND VPWR VPWR _1715_ sky130_fd_sc_hd__and4b_1
XFILLER_172_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5483_ net573 net1919 net612 VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__mux2_1
XFILLER_144_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4434_ _1618_ _1625_ _1627_ _1644_ VGND VGND VPWR VPWR _1646_ sky130_fd_sc_hd__or4_4
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7153_ clknet_3_2_0_wb_clk_i _0756_ net500 VGND VGND VPWR VPWR pad_count_2\[0\] sky130_fd_sc_hd__dfstp_1
X_4365_ net110 net99 VGND VGND VPWR VPWR _1577_ sky130_fd_sc_hd__nand2b_2
Xfanout505 net508 VGND VGND VPWR VPWR net505 sky130_fd_sc_hd__buf_8
Xfanout516 net517 VGND VGND VPWR VPWR net516 sky130_fd_sc_hd__buf_8
Xfanout527 net75 VGND VGND VPWR VPWR net527 sky130_fd_sc_hd__buf_12
X_6104_ gpio_configure\[11\]\[3\] net415 net399 gpio_configure\[18\]\[3\] _2922_ VGND
+ VGND VPWR VPWR _2923_ sky130_fd_sc_hd__a221o_1
X_3316_ _0889_ net381 VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__nor2_8
X_7084_ clknet_leaf_50_csclk net747 net508 VGND VGND VPWR VPWR gpio_configure\[30\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_113_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4296_ net461 net1650 _1541_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__mux2_1
XFILLER_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6035_ gpio_configure\[12\]\[0\] net409 net394 gpio_configure\[6\]\[0\] _2856_ VGND
+ VGND VPWR VPWR _2857_ sky130_fd_sc_hd__a221o_1
X_3247_ net474 net626 net580 VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__o21bai_1
XFILLER_100_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_731 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6937_ clknet_leaf_53_csclk net1038 net507 VGND VGND VPWR VPWR gpio_configure\[11\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6868_ clknet_leaf_23_csclk net1345 net514 VGND VGND VPWR VPWR gpio_configure\[3\]\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_167_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5819_ gpio_configure\[14\]\[6\] _2494_ _2498_ gpio_configure\[22\]\[6\] VGND VGND
+ VPWR VPWR _2648_ sky130_fd_sc_hd__a22o_1
XFILLER_50_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6799_ clknet_leaf_76_csclk net1721 net484 VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__dfstp_1
XFILLER_41_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold570 _0554_ VGND VGND VPWR VPWR net1103 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold581 gpio_configure\[25\]\[5\] VGND VGND VPWR VPWR net1114 sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 _0107_ VGND VGND VPWR VPWR net1125 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1270 _0309_ VGND VGND VPWR VPWR net1803 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1281 gpio_configure\[25\]\[0\] VGND VGND VPWR VPWR net1814 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1292 _0359_ VGND VGND VPWR VPWR net1825 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4150_ net456 net1340 _1514_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__mux2_1
XFILLER_122_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4081_ net726 net660 net351 VGND VGND VPWR VPWR _1496_ sky130_fd_sc_hd__mux2_1
XFILLER_68_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4983_ _1806_ _1962_ _2000_ VGND VGND VPWR VPWR _2193_ sky130_fd_sc_hd__nor3_1
XFILLER_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6722_ clknet_leaf_9_csclk net831 net509 VGND VGND VPWR VPWR gpio_configure\[17\]\[9\]
+ sky130_fd_sc_hd__dfrtp_4
X_3934_ _0829_ hkspi.sdoenb net483 VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__mux2_8
XFILLER_189_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6653_ clknet_3_4_0_wb_clk_i _0266_ VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__dfxtp_1
X_3865_ net2045 net2053 _1417_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__mux2_1
X_5604_ xfer_count\[0\] xfer_count\[1\] xfer_count\[2\] _2446_ VGND VGND VPWR VPWR
+ _2454_ sky130_fd_sc_hd__and4_1
XFILLER_164_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3796_ hkspi.count\[1\] hkspi.count\[0\] _1379_ VGND VGND VPWR VPWR _1381_ sky130_fd_sc_hd__and3_1
X_6584_ clknet_leaf_27_csclk net713 net519 VGND VGND VPWR VPWR mgmt_gpio_data_buf\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_191_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5535_ _0890_ net427 VGND VGND VPWR VPWR _2436_ sky130_fd_sc_hd__and2_4
XFILLER_11_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5466_ _0919_ net427 VGND VGND VPWR VPWR _2428_ sky130_fd_sc_hd__and2_4
XFILLER_145_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7205_ clknet_3_6_0_wb_clk_i _0807_ net528 VGND VGND VPWR VPWR wbbd_sck sky130_fd_sc_hd__dfrtp_2
X_4417_ _1617_ _1622_ _1628_ VGND VGND VPWR VPWR _1629_ sky130_fd_sc_hd__and3_2
XFILLER_99_650 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5397_ net1352 net459 _2420_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__mux2_1
XFILLER_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_7136_ clknet_leaf_28_csclk net539 net519 VGND VGND VPWR VPWR gpio_configure\[37\]\[1\]
+ sky130_fd_sc_hd__dfstp_2
X_4348_ _1549_ _1550_ _1551_ VGND VGND VPWR VPWR _1560_ sky130_fd_sc_hd__and3_1
XFILLER_98_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7067_ clknet_leaf_28_csclk net1185 net521 VGND VGND VPWR VPWR gpio_configure\[28\]\[1\]
+ sky130_fd_sc_hd__dfstp_2
X_4279_ net577 net836 _1538_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__mux2_1
XFILLER_86_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6018_ _1450_ _2797_ VGND VGND VPWR VPWR _2840_ sky130_fd_sc_hd__nor2_8
XFILLER_55_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_563 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_184_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_240 net569 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_251 gpio_configure\[3\]\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_262 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3650_ gpio_configure\[29\]\[2\] _0917_ _0940_ net276 _1238_ VGND VGND VPWR VPWR
+ _1239_ sky130_fd_sc_hd__a221o_1
XFILLER_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3581_ gpio_configure\[15\]\[3\] _0918_ _1007_ net64 _1170_ VGND VGND VPWR VPWR _1171_
+ sky130_fd_sc_hd__a221o_1
XFILLER_173_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5320_ net439 net748 net556 VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__mux2_1
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5251_ net1642 net469 _2404_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__mux2_1
XFILLER_115_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4202_ net918 net450 _1521_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__mux2_1
XFILLER_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5182_ wbbd_addr\[6\] _1529_ _2363_ _2384_ _2387_ VGND VGND VPWR VPWR _2388_ sky130_fd_sc_hd__a221o_1
XFILLER_142_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4133_ net1031 net449 _1511_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__mux2_1
XFILLER_29_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_3_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4064_ net1903 net441 net356 VGND VGND VPWR VPWR _1487_ sky130_fd_sc_hd__mux2_1
XFILLER_83_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_767 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4966_ _1779_ _1801_ _1970_ _1997_ VGND VGND VPWR VPWR _2176_ sky130_fd_sc_hd__o211a_1
XFILLER_51_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6705_ clknet_leaf_6_csclk net1311 net497 VGND VGND VPWR VPWR gpio_configure\[14\]\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_189_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3917_ _0970_ _1454_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__and2_2
XFILLER_177_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4897_ _1883_ _2107_ _2085_ _1699_ VGND VGND VPWR VPWR _2108_ sky130_fd_sc_hd__or4b_1
XFILLER_22_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6636_ clknet_leaf_5_csclk net1321 net494 VGND VGND VPWR VPWR gpio_configure\[6\]\[10\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_165_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3848_ hkspi.count\[1\] hkspi.count\[0\] hkspi.count\[2\] VGND VGND VPWR VPWR _1415_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_165_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6567_ clknet_leaf_40_csclk net663 net516 VGND VGND VPWR VPWR mgmt_gpio_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_3779_ gpio_configure\[30\]\[0\] _0892_ net367 gpio_configure\[17\]\[0\] VGND VGND
+ VPWR VPWR _1365_ sky130_fd_sc_hd__a22o_2
XFILLER_164_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_714 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5518_ net437 net1459 _2433_ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__mux2_1
X_6498_ clknet_leaf_61_csclk net1575 net498 VGND VGND VPWR VPWR gpio_configure\[31\]\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_145_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5449_ net469 net1792 _2426_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__mux2_1
XFILLER_160_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7119_ clknet_leaf_15_csclk net1567 net527 VGND VGND VPWR VPWR gpio_configure\[35\]\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_1__f_wbbd_sck clknet_0_wbbd_sck VGND VGND VPWR VPWR clknet_1_1__leaf_wbbd_sck
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_179_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_506 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4820_ net128 _1554_ _1749_ _1771_ _1819_ VGND VGND VPWR VPWR _2031_ sky130_fd_sc_hd__a41o_1
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4751_ _1653_ _1750_ VGND VGND VPWR VPWR _1963_ sky130_fd_sc_hd__nor2_1
XFILLER_193_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3702_ net286 _0910_ _1046_ gpio_configure\[28\]\[9\] VGND VGND VPWR VPWR _1290_
+ sky130_fd_sc_hd__a22o_1
XFILLER_147_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4682_ _1588_ _1684_ _1793_ VGND VGND VPWR VPWR _1894_ sky130_fd_sc_hd__a21o_1
XFILLER_119_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_658 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6421_ net495 net482 VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__and2_1
X_3633_ _1208_ _1211_ _1216_ _1221_ VGND VGND VPWR VPWR _1222_ sky130_fd_sc_hd__or4_2
XFILLER_174_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6352_ net2016 _1191_ _3156_ VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__mux2_1
X_3564_ gpio_configure\[9\]\[3\] net368 _1152_ _1153_ VGND VGND VPWR VPWR _1154_ sky130_fd_sc_hd__a211o_1
XFILLER_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5303_ net435 net1057 _2409_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__mux2_1
X_6283_ gpio_configure\[9\]\[10\] net412 _2838_ gpio_configure\[12\]\[10\] VGND VGND
+ VPWR VPWR _3095_ sky130_fd_sc_hd__a22o_1
XFILLER_142_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3495_ net388 _0899_ VGND VGND VPWR VPWR _1086_ sky130_fd_sc_hd__nor2_4
X_5234_ net465 net736 _2402_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__mux2_1
X_5165_ _1661_ _2262_ _2371_ _1664_ VGND VGND VPWR VPWR _2372_ sky130_fd_sc_hd__and4bb_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4116_ net618 net712 net630 VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__mux2_1
X_5096_ _1584_ _1706_ _1749_ _1770_ VGND VGND VPWR VPWR _2305_ sky130_fd_sc_hd__o31a_1
XFILLER_84_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4047_ net466 net1621 _1479_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__mux2_1
XFILLER_37_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5998_ _2479_ _2805_ VGND VGND VPWR VPWR _2820_ sky130_fd_sc_hd__nor2_8
XFILLER_52_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4949_ _1605_ _1639_ _1640_ _2141_ _2048_ VGND VGND VPWR VPWR _2159_ sky130_fd_sc_hd__o41a_1
XFILLER_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6619_ clknet_leaf_18_csclk net703 net512 VGND VGND VPWR VPWR gpio_configure\[4\]\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_193_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput280 net280 VGND VGND VPWR VPWR pll_trim[14] sky130_fd_sc_hd__buf_12
Xoutput291 net291 VGND VGND VPWR VPWR pll_trim[24] sky130_fd_sc_hd__buf_12
XFILLER_121_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_58_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_499 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3280_ _0870_ net376 VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__nor2_2
XFILLER_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6970_ clknet_3_3_0_csclk net1778 net505 VGND VGND VPWR VPWR gpio_configure\[16\]\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5921_ gpio_configure\[21\]\[10\] _2521_ _2540_ gpio_configure\[12\]\[10\] VGND VGND
+ VPWR VPWR _2746_ sky130_fd_sc_hd__a22o_1
XFILLER_80_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5852_ gpio_configure\[27\]\[7\] _2506_ _2528_ gpio_configure\[7\]\[7\] _2679_ VGND
+ VGND VPWR VPWR _2680_ sky130_fd_sc_hd__a221o_1
XFILLER_61_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4803_ _1601_ _1781_ _1804_ _1948_ VGND VGND VPWR VPWR _2014_ sky130_fd_sc_hd__a31o_1
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5783_ gpio_configure\[16\]\[4\] net419 _2534_ gpio_configure\[26\]\[4\] _2525_ VGND
+ VGND VPWR VPWR _2614_ sky130_fd_sc_hd__a221o_1
X_4734_ _1657_ _1745_ VGND VGND VPWR VPWR _1946_ sky130_fd_sc_hd__nor2_1
XFILLER_119_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4665_ _1866_ _1876_ VGND VGND VPWR VPWR _1877_ sky130_fd_sc_hd__nor2_1
XFILLER_190_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_162_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6404_ net513 net483 VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__and2_1
Xhold900 gpio_configure\[17\]\[6\] VGND VGND VPWR VPWR net1433 sky130_fd_sc_hd__dlygate4sd3_1
X_3616_ net58 _0933_ _0938_ gpio_configure\[33\]\[2\] VGND VGND VPWR VPWR _1205_ sky130_fd_sc_hd__a22o_1
Xhold911 _0643_ VGND VGND VPWR VPWR net1444 sky130_fd_sc_hd__dlygate4sd3_1
Xhold922 net2100 VGND VGND VPWR VPWR net1455 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_134_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4596_ _1555_ _1556_ VGND VGND VPWR VPWR _1808_ sky130_fd_sc_hd__or2_2
Xhold933 _0269_ VGND VGND VPWR VPWR net1466 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6335_ gpio_configure\[26\]\[12\] _2810_ _2830_ gpio_configure\[3\]\[12\] VGND VGND
+ VPWR VPWR _3145_ sky130_fd_sc_hd__a22o_1
Xhold944 gpio_configure\[11\]\[8\] VGND VGND VPWR VPWR net1477 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_162_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3547_ _0870_ _0897_ VGND VGND VPWR VPWR _1137_ sky130_fd_sc_hd__nor2_1
Xhold955 _0283_ VGND VGND VPWR VPWR net1488 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold966 serial_xfer VGND VGND VPWR VPWR net1499 sky130_fd_sc_hd__dlygate4sd3_1
Xhold977 net2110 VGND VGND VPWR VPWR net1510 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold988 _0727_ VGND VGND VPWR VPWR net1521 sky130_fd_sc_hd__dlygate4sd3_1
X_6266_ _3074_ _3076_ _3077_ _3078_ VGND VGND VPWR VPWR _3079_ sky130_fd_sc_hd__or4_1
X_3478_ net382 _1006_ VGND VGND VPWR VPWR _1069_ sky130_fd_sc_hd__nor2_4
Xhold999 gpio_configure\[37\]\[5\] VGND VGND VPWR VPWR net1532 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5217_ net457 net816 _2397_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__mux2_1
XFILLER_69_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1600 mgmt_gpio_data\[14\] VGND VGND VPWR VPWR net2133 sky130_fd_sc_hd__dlygate4sd3_1
X_6197_ gpio_configure\[36\]\[7\] net403 net402 gpio_configure\[4\]\[7\] VGND VGND
+ VPWR VPWR _3012_ sky130_fd_sc_hd__a22o_1
Xhold1611 gpio_configure\[37\]\[8\] VGND VGND VPWR VPWR net2144 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5148_ _1691_ _2214_ _2338_ _2342_ VGND VGND VPWR VPWR _2355_ sky130_fd_sc_hd__nor4_1
X_5079_ _2117_ _2232_ VGND VGND VPWR VPWR _2288_ sky130_fd_sc_hd__or2_1
XFILLER_71_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_708 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4450_ net99 _1597_ VGND VGND VPWR VPWR _1662_ sky130_fd_sc_hd__nor2_8
Xhold207 gpio_configure\[32\]\[3\] VGND VGND VPWR VPWR net740 sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 _0447_ VGND VGND VPWR VPWR net751 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold229 net228 VGND VGND VPWR VPWR net762 sky130_fd_sc_hd__dlygate4sd3_1
X_3401_ gpio_configure\[27\]\[6\] net370 _0939_ gpio_configure\[8\]\[6\] VGND VGND
+ VPWR VPWR _0995_ sky130_fd_sc_hd__a22o_1
XFILLER_132_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4381_ _1589_ net478 VGND VGND VPWR VPWR _1593_ sky130_fd_sc_hd__nand2_1
XFILLER_98_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3332_ net562 net386 VGND VGND VPWR VPWR _0928_ sky130_fd_sc_hd__nor2_8
X_6120_ gpio_configure\[0\]\[3\] _2851_ _2929_ _2938_ _0824_ VGND VGND VPWR VPWR _2939_
+ sky130_fd_sc_hd__o221a_2
XFILLER_171_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ net587 net2069 net474 VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__mux2_4
X_6051_ gpio_configure\[30\]\[1\] _2799_ net408 gpio_configure\[35\]\[1\] VGND VGND
+ VPWR VPWR _2872_ sky130_fd_sc_hd__a22o_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _1665_ _2203_ VGND VGND VPWR VPWR _2212_ sky130_fd_sc_hd__nor2_1
XFILLER_85_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3194_ xfer_state\[3\] VGND VGND VPWR VPWR _0823_ sky130_fd_sc_hd__inv_2
XFILLER_39_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6953_ clknet_leaf_41_csclk net1048 net517 VGND VGND VPWR VPWR gpio_configure\[13\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_5904_ net2089 _2729_ net366 VGND VGND VPWR VPWR _0773_ sky130_fd_sc_hd__mux2_1
XFILLER_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6884_ clknet_leaf_28_csclk net1589 net520 VGND VGND VPWR VPWR gpio_configure\[5\]\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_62_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5835_ _2656_ _2659_ _2661_ _2663_ VGND VGND VPWR VPWR _2664_ sky130_fd_sc_hd__or4_1
XFILLER_61_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5766_ gpio_configure\[13\]\[3\] _2501_ _2520_ gpio_configure\[8\]\[3\] _2597_ VGND
+ VGND VPWR VPWR _2598_ sky130_fd_sc_hd__a221o_1
X_4717_ _1576_ _1671_ VGND VGND VPWR VPWR _1929_ sky130_fd_sc_hd__or2_1
XFILLER_148_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5697_ pad_count_1\[4\] _2466_ _2489_ VGND VGND VPWR VPWR _2532_ sky130_fd_sc_hd__and3_4
XFILLER_108_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_147_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4648_ _1760_ _1859_ VGND VGND VPWR VPWR _1860_ sky130_fd_sc_hd__nor2_1
XFILLER_107_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold730 _0705_ VGND VGND VPWR VPWR net1263 sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 gpio_configure\[23\]\[11\] VGND VGND VPWR VPWR net1274 sky130_fd_sc_hd__dlygate4sd3_1
X_4579_ net477 _1779_ VGND VGND VPWR VPWR _1791_ sky130_fd_sc_hd__or2_4
Xhold752 _0529_ VGND VGND VPWR VPWR net1285 sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 gpio_configure\[14\]\[4\] VGND VGND VPWR VPWR net1296 sky130_fd_sc_hd__dlygate4sd3_1
X_6318_ net2147 _3128_ net473 VGND VGND VPWR VPWR _3129_ sky130_fd_sc_hd__mux2_1
Xhold774 _0473_ VGND VGND VPWR VPWR net1307 sky130_fd_sc_hd__dlygate4sd3_1
Xhold785 gpio_configure\[37\]\[12\] VGND VGND VPWR VPWR net1318 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold796 _0654_ VGND VGND VPWR VPWR net1329 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6249_ gpio_configure\[26\]\[9\] _2810_ _2811_ gpio_configure\[7\]\[9\] VGND VGND
+ VPWR VPWR _3062_ sky130_fd_sc_hd__a22o_1
XFILLER_77_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1430 gpio_configure\[24\]\[0\] VGND VGND VPWR VPWR net1963 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1441 _0366_ VGND VGND VPWR VPWR net1974 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1452 _0275_ VGND VGND VPWR VPWR net1985 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1463 _0389_ VGND VGND VPWR VPWR net1996 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1474 net326 VGND VGND VPWR VPWR net2007 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1485 _0770_ VGND VGND VPWR VPWR net2018 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_61_csclk clknet_3_0_0_csclk VGND VGND VPWR VPWR clknet_leaf_61_csclk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1496 serial_data_staging_1\[1\] VGND VGND VPWR VPWR net2029 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_55_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_76_csclk clknet_3_0_0_csclk VGND VGND VPWR VPWR clknet_leaf_76_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_14_csclk clknet_3_5_0_csclk VGND VGND VPWR VPWR clknet_leaf_14_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_96_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold90 _0295_ VGND VGND VPWR VPWR net623 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_29_csclk clknet_3_7_0_csclk VGND VGND VPWR VPWR clknet_leaf_29_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_90_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3950_ net260 VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__inv_2
XFILLER_16_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3881_ net105 net104 net107 net106 VGND VGND VPWR VPWR _1433_ sky130_fd_sc_hd__or4_1
X_5620_ net2142 _2460_ _2463_ _2465_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__a31o_1
XFILLER_188_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5551_ net438 net1393 _2437_ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__mux2_1
XFILLER_145_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4502_ _1661_ _1713_ _1664_ VGND VGND VPWR VPWR _1714_ sky130_fd_sc_hd__or3b_1
X_5482_ net437 net1419 net612 VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__mux2_1
X_4433_ _1617_ _1619_ _1621_ _1628_ VGND VGND VPWR VPWR _1645_ sky130_fd_sc_hd__and4_2
XFILLER_144_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7152_ clknet_3_0_0_wb_clk_i _0755_ net500 VGND VGND VPWR VPWR pad_count_1\[4\] sky130_fd_sc_hd__dfstp_4
XFILLER_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4364_ _1564_ _1575_ VGND VGND VPWR VPWR _1576_ sky130_fd_sc_hd__or2_4
Xfanout506 net508 VGND VGND VPWR VPWR net506 sky130_fd_sc_hd__buf_8
Xfanout517 net526 VGND VGND VPWR VPWR net517 sky130_fd_sc_hd__buf_8
X_6103_ gpio_configure\[7\]\[3\] _2811_ net404 gpio_configure\[25\]\[3\] VGND VGND
+ VPWR VPWR _2922_ sky130_fd_sc_hd__a22o_1
X_3315_ net386 net601 VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__nor2_8
XFILLER_112_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout528 net529 VGND VGND VPWR VPWR net528 sky130_fd_sc_hd__buf_6
X_4295_ net466 net1753 _1541_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__mux2_1
XFILLER_59_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7083_ clknet_leaf_25_csclk net1396 net518 VGND VGND VPWR VPWR gpio_configure\[30\]\[1\]
+ sky130_fd_sc_hd__dfstp_4
XFILLER_113_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_98_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3246_ net579 net474 _0840_ _0841_ VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__o31a_1
XFILLER_100_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6034_ gpio_configure\[9\]\[0\] net412 net406 gpio_configure\[27\]\[0\] VGND VGND
+ VPWR VPWR _2856_ sky130_fd_sc_hd__a22o_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6936_ clknet_leaf_53_csclk net1366 net507 VGND VGND VPWR VPWR gpio_configure\[11\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6867_ clknet_leaf_21_csclk net859 net514 VGND VGND VPWR VPWR gpio_configure\[3\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_179_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5818_ gpio_configure\[4\]\[6\] _2502_ _2517_ gpio_configure\[30\]\[6\] _2646_ VGND
+ VGND VPWR VPWR _2647_ sky130_fd_sc_hd__a221o_1
X_6798_ clknet_leaf_76_csclk net1750 net484 VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__dfrtp_2
X_5749_ gpio_configure\[19\]\[2\] _2491_ _2529_ gpio_configure\[29\]\[2\] _2581_ VGND
+ VGND VPWR VPWR _2582_ sky130_fd_sc_hd__a221o_1
XFILLER_136_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_748 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold560 gpio_configure\[30\]\[12\] VGND VGND VPWR VPWR net1093 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold571 gpio_configure\[17\]\[12\] VGND VGND VPWR VPWR net1104 sky130_fd_sc_hd__dlygate4sd3_1
Xhold582 _0650_ VGND VGND VPWR VPWR net1115 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_173_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold593 net261 VGND VGND VPWR VPWR net1126 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_173_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1260 _0621_ VGND VGND VPWR VPWR net1793 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1271 gpio_configure\[7\]\[8\] VGND VGND VPWR VPWR net1804 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1282 _0645_ VGND VGND VPWR VPWR net1815 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1293 net275 VGND VGND VPWR VPWR net1826 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_684 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_186_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4080_ net950 _1495_ _1490_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__mux2_1
XFILLER_110_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_76_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_17_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4982_ _1845_ _1998_ _2191_ VGND VGND VPWR VPWR _2192_ sky130_fd_sc_hd__or3_1
X_6721_ clknet_leaf_9_csclk net1780 net509 VGND VGND VPWR VPWR gpio_configure\[17\]\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_3933_ mgmt_gpio_data\[0\] net3 net1 VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__mux2_4
X_6652_ clknet_3_4_0_wb_clk_i _0265_ VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__dfxtp_1
XFILLER_149_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3864_ net2053 net2047 _1417_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__mux2_1
X_5603_ xfer_count\[0\] xfer_count\[1\] _2446_ xfer_count\[2\] VGND VGND VPWR VPWR
+ _2453_ sky130_fd_sc_hd__a31o_1
XFILLER_118_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6583_ clknet_leaf_35_csclk net1006 net525 VGND VGND VPWR VPWR mgmt_gpio_data_buf\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_3795_ _1379_ VGND VGND VPWR VPWR _1380_ sky130_fd_sc_hd__inv_2
X_5534_ net1228 net444 _2435_ VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__mux2_1
XFILLER_117_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_191_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5465_ net434 net1278 _2427_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__mux2_1
XFILLER_105_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7204_ clknet_3_6_0_wb_clk_i _0806_ net529 VGND VGND VPWR VPWR wbbd_data\[7\] sky130_fd_sc_hd__dfrtp_1
X_4416_ _1625_ _1627_ VGND VGND VPWR VPWR _1628_ sky130_fd_sc_hd__nor2_4
X_5396_ net1381 net464 _2420_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__mux2_1
XFILLER_99_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7135_ clknet_leaf_26_csclk net1628 net519 VGND VGND VPWR VPWR gpio_configure\[37\]\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_160_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4347_ net128 _1554_ _1557_ VGND VGND VPWR VPWR _1559_ sky130_fd_sc_hd__and3_1
XFILLER_113_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7066_ clknet_leaf_15_csclk net1977 net513 VGND VGND VPWR VPWR gpio_configure\[28\]\[0\]
+ sky130_fd_sc_hd__dfstp_4
X_4278_ net465 net876 _1538_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__mux2_1
XFILLER_46_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6017_ _1447_ _2469_ _2800_ VGND VGND VPWR VPWR _2839_ sky130_fd_sc_hd__and3b_4
X_3229_ gpio_configure\[5\]\[3\] VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkinv_2
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_1_0__f_wbbd_sck clknet_0_wbbd_sck VGND VGND VPWR VPWR clknet_1_0__leaf_wbbd_sck
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6919_ clknet_leaf_31_csclk net1543 net523 VGND VGND VPWR VPWR gpio_configure\[9\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_23_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold390 _0620_ VGND VGND VPWR VPWR net923 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1090 gpio_configure\[8\]\[8\] VGND VGND VPWR VPWR net1623 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_230 net439 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_241 net612 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_252 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_263 net471 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3580_ gpio_configure\[4\]\[11\] _1093_ _1129_ gpio_configure\[11\]\[11\] VGND VGND
+ VPWR VPWR _1170_ sky130_fd_sc_hd__a22o_2
XFILLER_139_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5250_ _0898_ net427 VGND VGND VPWR VPWR _2404_ sky130_fd_sc_hd__and2_4
XFILLER_142_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4201_ net1360 net456 _1521_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__mux2_1
XFILLER_114_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5181_ _2331_ _2386_ _2367_ VGND VGND VPWR VPWR _2387_ sky130_fd_sc_hd__a21oi_2
X_4132_ net1634 net455 _1511_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__mux2_1
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4063_ net914 _1486_ _1481_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__mux2_1
XFILLER_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4965_ _1799_ _1961_ _2027_ VGND VGND VPWR VPWR _2175_ sky130_fd_sc_hd__or3b_1
XFILLER_51_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6704_ clknet_leaf_3_csclk net1261 net496 VGND VGND VPWR VPWR gpio_configure\[14\]\[11\]
+ sky130_fd_sc_hd__dfrtp_2
X_3916_ hkspi.state\[1\] hkspi.state\[4\] _0821_ VGND VGND VPWR VPWR _1454_ sky130_fd_sc_hd__o21ai_1
XFILLER_149_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4896_ _1954_ _2093_ _2105_ _2106_ VGND VGND VPWR VPWR _2107_ sky130_fd_sc_hd__or4_1
X_6635_ clknet_leaf_1_csclk net1484 net493 VGND VGND VPWR VPWR gpio_configure\[6\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3847_ net58 net2119 _1414_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__mux2_1
XFILLER_137_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_687 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6566_ clknet_leaf_40_csclk net1760 net516 VGND VGND VPWR VPWR mgmt_gpio_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_3778_ gpio_configure\[31\]\[0\] net375 _0924_ gpio_configure\[26\]\[0\] _1363_ VGND
+ VGND VPWR VPWR _1364_ sky130_fd_sc_hd__a221o_1
XFILLER_152_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5517_ net441 net1132 _2433_ VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__mux2_1
XFILLER_173_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6497_ clknet_leaf_72_csclk net1117 net488 VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__dfstp_2
XFILLER_106_726 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5448_ _0923_ net427 VGND VGND VPWR VPWR _2426_ sky130_fd_sc_hd__nand2_8
XFILLER_160_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5379_ net458 net1656 _2418_ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__mux2_1
X_7118_ clknet_leaf_34_csclk net967 net525 VGND VGND VPWR VPWR gpio_configure\[34\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_87_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7049_ clknet_leaf_37_csclk net613 net522 VGND VGND VPWR VPWR gpio_configure\[25\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_604 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_11_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_46_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_729 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4750_ _1665_ _1750_ VGND VGND VPWR VPWR _1962_ sky130_fd_sc_hd__nor2_1
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3701_ _1282_ _1284_ _1286_ _1288_ VGND VGND VPWR VPWR _1289_ sky130_fd_sc_hd__or4_1
XFILLER_186_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4681_ _1678_ _1823_ _1841_ _1581_ VGND VGND VPWR VPWR _1893_ sky130_fd_sc_hd__o22a_1
XFILLER_159_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6420_ net495 net482 VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__and2_1
X_3632_ _1217_ _1218_ _1219_ _1220_ VGND VGND VPWR VPWR _1221_ sky130_fd_sc_hd__or4_1
XFILLER_134_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6351_ net1978 _1249_ _3156_ VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__mux2_1
X_3563_ gpio_configure\[9\]\[11\] _1057_ _1094_ gpio_configure\[7\]\[11\] _1139_ VGND
+ VGND VPWR VPWR _1153_ sky130_fd_sc_hd__a221o_2
XFILLER_127_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5302_ net438 net1358 _2409_ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__mux2_1
X_6282_ gpio_configure\[34\]\[10\] net393 _2852_ gpio_configure\[19\]\[10\] _3093_
+ VGND VGND VPWR VPWR _3094_ sky130_fd_sc_hd__a221o_1
X_3494_ net56 _0871_ _0936_ net24 _1084_ VGND VGND VPWR VPWR _1085_ sky130_fd_sc_hd__a221o_2
XFILLER_88_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5233_ net471 net1504 _2402_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__mux2_1
XFILLER_68_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5164_ _1605_ _1777_ _1872_ _2159_ VGND VGND VPWR VPWR _2371_ sky130_fd_sc_hd__o31a_1
XFILLER_111_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4115_ net452 net1005 net630 VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__mux2_1
X_5095_ _1821_ _1990_ _2185_ _2303_ VGND VGND VPWR VPWR _2304_ sky130_fd_sc_hd__or4_1
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4046_ _1116_ net425 VGND VGND VPWR VPWR _1479_ sky130_fd_sc_hd__nand2_2
XFILLER_17_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5997_ _2479_ _2818_ VGND VGND VPWR VPWR _2819_ sky130_fd_sc_hd__nor2_8
XFILLER_52_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4948_ _1605_ _1638_ _1639_ _2141_ _2046_ VGND VGND VPWR VPWR _2158_ sky130_fd_sc_hd__o41a_1
X_4879_ _1651_ _1750_ _1682_ VGND VGND VPWR VPWR _2090_ sky130_fd_sc_hd__o21ai_1
XFILLER_138_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6618_ clknet_leaf_8_csclk net753 net509 VGND VGND VPWR VPWR gpio_configure\[4\]\[10\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_192_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6549_ clknet_leaf_35_csclk net1486 net525 VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__dfrtp_1
XFILLER_106_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput270 net270 VGND VGND VPWR VPWR pll_div[4] sky130_fd_sc_hd__buf_12
Xoutput281 net281 VGND VGND VPWR VPWR pll_trim[15] sky130_fd_sc_hd__buf_12
XFILLER_121_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput292 net292 VGND VGND VPWR VPWR pll_trim[25] sky130_fd_sc_hd__buf_12
XFILLER_121_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_188_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5920_ gpio_configure\[28\]\[10\] _2513_ _2537_ gpio_configure\[17\]\[10\] _2744_
+ VGND VGND VPWR VPWR _2745_ sky130_fd_sc_hd__a221o_1
XFILLER_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5851_ gpio_configure\[8\]\[7\] _2520_ net419 _2678_ VGND VGND VPWR VPWR _2679_ sky130_fd_sc_hd__a22o_1
XFILLER_34_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4802_ _1745_ _1759_ _1766_ _1993_ VGND VGND VPWR VPWR _2013_ sky130_fd_sc_hd__nor4_1
X_5782_ gpio_configure\[17\]\[4\] _2537_ _2541_ gpio_configure\[31\]\[4\] _2612_ VGND
+ VGND VPWR VPWR _2613_ sky130_fd_sc_hd__a221o_1
X_4733_ _1868_ _1879_ _1944_ _1617_ VGND VGND VPWR VPWR _1945_ sky130_fd_sc_hd__o22a_1
XFILLER_159_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4664_ _1688_ _1782_ VGND VGND VPWR VPWR _1876_ sky130_fd_sc_hd__or2_1
XFILLER_174_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6403_ net513 net483 VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__and2_1
X_3615_ gpio_configure\[11\]\[2\] _0907_ _0916_ gpio_configure\[14\]\[2\] VGND VGND
+ VPWR VPWR _1204_ sky130_fd_sc_hd__a22o_1
XFILLER_135_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold901 _0587_ VGND VGND VPWR VPWR net1434 sky130_fd_sc_hd__dlygate4sd3_1
X_4595_ _1601_ _1756_ VGND VGND VPWR VPWR _1807_ sky130_fd_sc_hd__nand2_8
Xhold912 gpio_configure\[31\]\[9\] VGND VGND VPWR VPWR net1445 sky130_fd_sc_hd__dlygate4sd3_1
Xhold923 _0202_ VGND VGND VPWR VPWR net1456 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold934 gpio_configure\[23\]\[9\] VGND VGND VPWR VPWR net1467 sky130_fd_sc_hd__dlygate4sd3_1
X_6334_ gpio_configure\[30\]\[12\] _2799_ _2819_ gpio_configure\[18\]\[12\] _3143_
+ VGND VGND VPWR VPWR _3144_ sky130_fd_sc_hd__a221o_1
XFILLER_162_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3546_ net378 _0889_ VGND VGND VPWR VPWR _1136_ sky130_fd_sc_hd__nor2_8
Xhold945 _0288_ VGND VGND VPWR VPWR net1478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold956 net226 VGND VGND VPWR VPWR net1489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 _2398_ VGND VGND VPWR VPWR net1500 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold978 _0201_ VGND VGND VPWR VPWR net1511 sky130_fd_sc_hd__dlygate4sd3_1
X_6265_ gpio_configure\[3\]\[9\] _2830_ _2842_ gpio_configure\[15\]\[9\] _3062_ VGND
+ VGND VPWR VPWR _3078_ sky130_fd_sc_hd__a221o_1
XFILLER_130_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold989 gpio_configure\[11\]\[5\] VGND VGND VPWR VPWR net1522 sky130_fd_sc_hd__dlygate4sd3_1
X_3477_ net582 _1008_ VGND VGND VPWR VPWR _1068_ sky130_fd_sc_hd__nor2_4
XFILLER_115_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5216_ net451 net764 _2397_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__mux2_1
X_6196_ net2044 _2487_ _3010_ _3011_ VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__a22o_1
XFILLER_130_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1601 gpio_configure\[33\]\[4\] VGND VGND VPWR VPWR net2134 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1612 gpio_configure\[32\]\[9\] VGND VGND VPWR VPWR net2145 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5147_ _2347_ _2353_ VGND VGND VPWR VPWR _2354_ sky130_fd_sc_hd__and2b_1
XFILLER_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5078_ _1807_ _2285_ _2286_ VGND VGND VPWR VPWR _2287_ sky130_fd_sc_hd__o21ai_1
XFILLER_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4029_ net1808 net468 _1476_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__mux2_1
XFILLER_44_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold208 _0701_ VGND VGND VPWR VPWR net741 sky130_fd_sc_hd__dlygate4sd3_1
Xhold219 gpio_configure\[4\]\[10\] VGND VGND VPWR VPWR net752 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_171_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3400_ gpio_configure\[6\]\[6\] net357 _0991_ _0993_ VGND VGND VPWR VPWR _0994_ sky130_fd_sc_hd__a211o_1
XFILLER_125_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4380_ net127 net128 net126 net125 VGND VGND VPWR VPWR _1592_ sky130_fd_sc_hd__or4_4
XFILLER_98_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_125_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3331_ net387 net609 VGND VGND VPWR VPWR _0927_ sky130_fd_sc_hd__nor2_8
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ gpio_configure\[37\]\[1\] net400 net416 gpio_configure\[32\]\[1\] VGND VGND
+ VPWR VPWR _2871_ sky130_fd_sc_hd__a22o_1
XFILLER_112_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ net586 net558 hkspi.state\[3\] VGND VGND VPWR VPWR _0858_ sky130_fd_sc_hd__mux2_1
XFILLER_140_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5001_ _1622_ _1670_ _1937_ VGND VGND VPWR VPWR _2211_ sky130_fd_sc_hd__and3_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3193_ net2113 VGND VGND VPWR VPWR _0822_ sky130_fd_sc_hd__inv_2
XFILLER_66_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6952_ clknet_leaf_44_csclk net853 net517 VGND VGND VPWR VPWR gpio_configure\[13\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_5903_ xfer_state\[1\] serial_data_staging_1\[8\] _2728_ VGND VGND VPWR VPWR _2729_
+ sky130_fd_sc_hd__a21o_1
XFILLER_179_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6883_ clknet_leaf_49_csclk net885 net505 VGND VGND VPWR VPWR gpio_configure\[5\]\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_5834_ gpio_configure\[18\]\[6\] _2532_ _2535_ gpio_configure\[23\]\[6\] _2662_ VGND
+ VGND VPWR VPWR _2663_ sky130_fd_sc_hd__a221o_1
XFILLER_179_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5765_ gpio_configure\[14\]\[3\] _2494_ _2540_ gpio_configure\[12\]\[3\] VGND VGND
+ VPWR VPWR _2597_ sky130_fd_sc_hd__a22o_1
XFILLER_148_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4716_ _1576_ _1671_ VGND VGND VPWR VPWR _1928_ sky130_fd_sc_hd__nor2_1
X_5696_ pad_count_1\[4\] _2459_ _2504_ VGND VGND VPWR VPWR _2531_ sky130_fd_sc_hd__and3_4
XFILLER_163_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4647_ _1814_ _1856_ VGND VGND VPWR VPWR _1859_ sky130_fd_sc_hd__nor2_1
XFILLER_162_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold720 _0357_ VGND VGND VPWR VPWR net1253 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_100_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold731 gpio_configure\[1\]\[4\] VGND VGND VPWR VPWR net1264 sky130_fd_sc_hd__dlygate4sd3_1
X_4578_ net127 net126 net125 net128 VGND VGND VPWR VPWR _1790_ sky130_fd_sc_hd__or4b_4
Xhold742 _0131_ VGND VGND VPWR VPWR net1275 sky130_fd_sc_hd__dlygate4sd3_1
Xhold753 gpio_configure\[24\]\[11\] VGND VGND VPWR VPWR net1286 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6317_ _3112_ _3118_ _3127_ _2851_ gpio_configure\[0\]\[11\] VGND VGND VPWR VPWR
+ _3128_ sky130_fd_sc_hd__o32a_1
Xhold764 _0561_ VGND VGND VPWR VPWR net1297 sky130_fd_sc_hd__dlygate4sd3_1
X_3529_ gpio_configure\[6\]\[4\] _0876_ _1119_ gpio_configure\[5\]\[12\] _1118_ VGND
+ VGND VPWR VPWR _1120_ sky130_fd_sc_hd__a221o_1
Xhold775 gpio_configure\[4\]\[0\] VGND VGND VPWR VPWR net1308 sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 _0323_ VGND VGND VPWR VPWR net1319 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold797 gpio_configure\[21\]\[1\] VGND VGND VPWR VPWR net1330 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6248_ gpio_configure\[28\]\[9\] _2861_ VGND VGND VPWR VPWR _3061_ sky130_fd_sc_hd__and2_1
XFILLER_77_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_698 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6179_ gpio_configure\[10\]\[6\] _2825_ _2840_ gpio_configure\[6\]\[6\] _2994_ VGND
+ VGND VPWR VPWR _2995_ sky130_fd_sc_hd__a221o_1
XFILLER_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1420 net325 VGND VGND VPWR VPWR net1953 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_130_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1431 _0637_ VGND VGND VPWR VPWR net1964 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1442 mgmt_gpio_data_buf\[4\] VGND VGND VPWR VPWR net1975 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1453 gpio_configure\[27\]\[0\] VGND VGND VPWR VPWR net1986 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1464 hkspi.ldata\[2\] VGND VGND VPWR VPWR net1997 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1475 hkspi.SDO VGND VGND VPWR VPWR net2008 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1486 serial_data_staging_1\[0\] VGND VGND VPWR VPWR net2019 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1497 _0765_ VGND VGND VPWR VPWR net2030 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_730 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold80 _0652_ VGND VGND VPWR VPWR net613 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 hkspi.addr\[7\] VGND VGND VPWR VPWR net624 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_36_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_90_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3880_ net109 net108 net115 net116 VGND VGND VPWR VPWR _1432_ sky130_fd_sc_hd__or4b_1
XFILLER_149_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5550_ net441 net956 _2437_ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__mux2_1
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4501_ _1575_ _1599_ _1605_ _1712_ VGND VGND VPWR VPWR _1713_ sky130_fd_sc_hd__o31ai_1
X_5481_ net441 net1114 net612 VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__mux2_1
XFILLER_129_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4432_ _1619_ _1621_ VGND VGND VPWR VPWR _1644_ sky130_fd_sc_hd__nand2_1
X_7151_ clknet_3_0_0_wb_clk_i _0754_ net500 VGND VGND VPWR VPWR pad_count_1\[3\] sky130_fd_sc_hd__dfrtp_1
X_4363_ _1568_ _1571_ _1573_ VGND VGND VPWR VPWR _1575_ sky130_fd_sc_hd__or3_1
XFILLER_98_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout507 net508 VGND VGND VPWR VPWR net507 sky130_fd_sc_hd__clkbuf_8
X_6102_ gpio_configure\[34\]\[3\] net393 net391 gpio_configure\[17\]\[3\] _2920_ VGND
+ VGND VPWR VPWR _2921_ sky130_fd_sc_hd__a221o_1
X_3314_ net389 _0909_ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__nor2_8
XFILLER_140_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout518 net526 VGND VGND VPWR VPWR net518 sky130_fd_sc_hd__buf_8
Xfanout529 net164 VGND VGND VPWR VPWR net529 sky130_fd_sc_hd__buf_6
X_7082_ clknet_leaf_16_csclk net1799 net527 VGND VGND VPWR VPWR gpio_configure\[30\]\[0\]
+ sky130_fd_sc_hd__dfstp_2
X_4294_ _1054_ net425 VGND VGND VPWR VPWR _1541_ sky130_fd_sc_hd__nand2_2
XFILLER_98_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6033_ _2469_ _2478_ _2809_ VGND VGND VPWR VPWR _2855_ sky130_fd_sc_hd__and3_4
X_3245_ wbbd_addr\[6\] net474 VGND VGND VPWR VPWR _0841_ sky130_fd_sc_hd__nand2b_1
XFILLER_67_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_132_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6935_ clknet_leaf_33_csclk net1523 net524 VGND VGND VPWR VPWR gpio_configure\[11\]\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6866_ clknet_leaf_20_csclk net1758 net511 VGND VGND VPWR VPWR gpio_configure\[3\]\[0\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5817_ gpio_configure\[7\]\[6\] _2528_ _2534_ gpio_configure\[26\]\[6\] VGND VGND
+ VPWR VPWR _2646_ sky130_fd_sc_hd__a22o_1
X_6797_ clknet_leaf_76_csclk net1012 net484 VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__dfrtp_4
XFILLER_167_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5748_ gpio_configure\[14\]\[2\] _2494_ _2517_ gpio_configure\[30\]\[2\] VGND VGND
+ VPWR VPWR _2581_ sky130_fd_sc_hd__a22o_1
XFILLER_157_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5679_ gpio_configure\[9\]\[0\] _2512_ _2513_ gpio_configure\[28\]\[0\] VGND VGND
+ VPWR VPWR _2514_ sky130_fd_sc_hd__a22o_1
XFILLER_135_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold550 net235 VGND VGND VPWR VPWR net1083 sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 _0137_ VGND VGND VPWR VPWR net1094 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold572 _0328_ VGND VGND VPWR VPWR net1105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 net298 VGND VGND VPWR VPWR net1116 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_150_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold594 _0404_ VGND VGND VPWR VPWR net1127 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1250 gpio_configure\[16\]\[8\] VGND VGND VPWR VPWR net1783 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1261 gpio_configure\[8\]\[0\] VGND VGND VPWR VPWR net1794 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1272 _0268_ VGND VGND VPWR VPWR net1805 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1283 gpio_configure\[32\]\[8\] VGND VGND VPWR VPWR net1816 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1294 _0112_ VGND VGND VPWR VPWR net1827 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_696 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput170 wb_we_i VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4981_ _1592_ _1599_ _1785_ VGND VGND VPWR VPWR _2191_ sky130_fd_sc_hd__nor3_1
XFILLER_23_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3932_ _1456_ net74 hkspi.pass_thru_mgmt VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__mux2_4
X_6720_ clknet_leaf_62_csclk net1319 net501 VGND VGND VPWR VPWR gpio_configure\[37\]\[12\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_16_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6651_ clknet_3_4_0_wb_clk_i _0264_ VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__dfxtp_1
XFILLER_189_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3863_ net2047 net1956 _1417_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__mux2_1
XFILLER_149_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5602_ xfer_count\[1\] _2447_ _2451_ _2452_ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__a22o_1
X_6582_ clknet_leaf_35_csclk net1317 net525 VGND VGND VPWR VPWR mgmt_gpio_data_buf\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_3794_ hkspi.state\[0\] _1378_ VGND VGND VPWR VPWR _1379_ sky130_fd_sc_hd__or2_2
XFILLER_176_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5533_ net1324 net450 _2435_ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__mux2_1
XFILLER_118_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5464_ net437 net1415 _2427_ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_60_csclk clknet_3_2_0_csclk VGND VGND VPWR VPWR clknet_leaf_60_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_133_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7203_ clknet_3_6_0_wb_clk_i _0805_ net529 VGND VGND VPWR VPWR wbbd_data\[6\] sky130_fd_sc_hd__dfrtp_1
X_4415_ _1614_ _1626_ VGND VGND VPWR VPWR _1627_ sky130_fd_sc_hd__or2_2
X_5395_ net1777 net469 _2420_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__mux2_1
X_7134_ clknet_leaf_33_csclk net935 net524 VGND VGND VPWR VPWR gpio_configure\[36\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_4346_ _1554_ _1557_ VGND VGND VPWR VPWR _1558_ sky130_fd_sc_hd__nand2_1
XFILLER_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_75_csclk clknet_3_0_0_csclk VGND VGND VPWR VPWR clknet_leaf_75_csclk
+ sky130_fd_sc_hd__clkbuf_16
X_7065_ clknet_leaf_43_csclk net1096 net517 VGND VGND VPWR VPWR gpio_configure\[27\]\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_4277_ net471 net1594 _1538_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__mux2_1
X_6016_ _2473_ _2793_ _2796_ VGND VGND VPWR VPWR _2838_ sky130_fd_sc_hd__and3_4
X_3228_ gpio_configure\[6\]\[3\] VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__inv_2
XFILLER_82_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6918_ clknet_leaf_15_csclk net1175 net513 VGND VGND VPWR VPWR gpio_configure\[9\]\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_70_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6849_ clknet_leaf_51_csclk net1129 net506 VGND VGND VPWR VPWR gpio_configure\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_168_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_167_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_109_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_28_csclk clknet_3_7_0_csclk VGND VGND VPWR VPWR clknet_leaf_28_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_136_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold380 _0183_ VGND VGND VPWR VPWR net913 sky130_fd_sc_hd__dlygate4sd3_1
Xhold391 net302 VGND VGND VPWR VPWR net924 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1080 _0428_ VGND VGND VPWR VPWR net1613 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1091 _0273_ VGND VGND VPWR VPWR net1624 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_220 net281 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_231 net445 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_242 net660 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_253 net58 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_264 net471 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4200_ net1465 net462 _1521_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__mux2_1
XFILLER_130_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5180_ _2148_ _2274_ _2372_ _2385_ VGND VGND VPWR VPWR _2386_ sky130_fd_sc_hd__and4bb_1
XFILLER_3_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4131_ net1698 net461 _1511_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__mux2_1
XFILLER_110_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4062_ net712 net618 net356 VGND VGND VPWR VPWR _1486_ sky130_fd_sc_hd__mux2_1
XFILLER_96_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4964_ _1746_ _2173_ VGND VGND VPWR VPWR _2174_ sky130_fd_sc_hd__or2_1
X_6703_ clknet_leaf_6_csclk net1408 net497 VGND VGND VPWR VPWR gpio_configure\[14\]\[10\]
+ sky130_fd_sc_hd__dfstp_1
X_3915_ _0821_ _1441_ _1384_ hkspi.state\[3\] VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_189_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4895_ _1612_ _1936_ _1943_ _1953_ VGND VGND VPWR VPWR _2106_ sky130_fd_sc_hd__a31o_1
X_3846_ hkspi.count\[2\] hkspi.count\[1\] hkspi.count\[0\] hkspi.state\[0\] VGND VGND
+ VPWR VPWR _1414_ sky130_fd_sc_hd__or4bb_1
X_6634_ clknet_leaf_5_csclk net1752 net494 VGND VGND VPWR VPWR gpio_configure\[6\]\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_165_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3777_ net34 _0891_ _0936_ net20 VGND VGND VPWR VPWR _1363_ sky130_fd_sc_hd__a22o_1
X_6565_ clknet_3_3_0_wb_clk_i _0017_ net499 VGND VGND VPWR VPWR xfer_state\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_192_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5516_ net618 net675 _2433_ VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__mux2_1
XFILLER_3_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6496_ clknet_leaf_73_csclk net777 net488 VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__dfstp_2
XFILLER_133_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5447_ net435 net922 _2425_ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__mux2_1
XFILLER_154_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5378_ net465 net870 _2418_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__mux2_1
X_4329_ net986 net443 _1546_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__mux2_1
X_7117_ clknet_leaf_55_csclk net1400 net506 VGND VGND VPWR VPWR gpio_configure\[34\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_113_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7048_ clknet_leaf_56_csclk net1420 net504 VGND VGND VPWR VPWR gpio_configure\[25\]\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_170_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_419 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_730 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_73_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3700_ gpio_configure\[24\]\[1\] _0919_ _1065_ gpio_configure\[37\]\[9\] _1287_ VGND
+ VGND VPWR VPWR _1288_ sky130_fd_sc_hd__a221o_1
X_4680_ _1777_ _1886_ VGND VGND VPWR VPWR _1892_ sky130_fd_sc_hd__nor2_1
XFILLER_174_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3631_ gpio_configure\[5\]\[2\] net355 _0934_ gpio_configure\[1\]\[2\] _1197_ VGND
+ VGND VPWR VPWR _1220_ sky130_fd_sc_hd__a221o_1
XFILLER_146_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6350_ net1962 _1311_ _3156_ VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__mux2_1
X_3562_ gpio_configure\[7\]\[3\] _0913_ net373 gpio_configure\[14\]\[3\] _1138_ VGND
+ VGND VPWR VPWR _1152_ sky130_fd_sc_hd__a221o_1
XFILLER_155_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5301_ net441 net1065 _2409_ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__mux2_1
X_6281_ gpio_configure\[37\]\[10\] _2806_ net416 gpio_configure\[32\]\[10\] _3083_
+ VGND VGND VPWR VPWR _3093_ sky130_fd_sc_hd__a221o_1
XFILLER_142_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3493_ gpio_configure\[3\]\[4\] _0915_ _1083_ gpio_configure\[30\]\[12\] VGND VGND
+ VPWR VPWR _1084_ sky130_fd_sc_hd__a22o_1
XFILLER_115_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5232_ _0871_ net647 VGND VGND VPWR VPWR _2402_ sky130_fd_sc_hd__nand2_4
XFILLER_142_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5163_ _2166_ _2168_ _2369_ VGND VGND VPWR VPWR _2370_ sky130_fd_sc_hd__and3_1
XFILLER_96_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4114_ net458 net1316 net630 VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__mux2_1
X_5094_ _1707_ _2005_ VGND VGND VPWR VPWR _2303_ sky130_fd_sc_hd__nor2_1
XFILLER_68_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4045_ net443 net1204 _1478_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__mux2_1
XFILLER_84_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_37_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5996_ _1448_ _2800_ VGND VGND VPWR VPWR _2818_ sky130_fd_sc_hd__nand2_4
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4947_ _1638_ _2145_ VGND VGND VPWR VPWR _2157_ sky130_fd_sc_hd__nor2_1
XFILLER_177_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4878_ _1729_ _1963_ VGND VGND VPWR VPWR _2089_ sky130_fd_sc_hd__or2_1
X_6617_ clknet_leaf_12_csclk net901 net512 VGND VGND VPWR VPWR gpio_configure\[4\]\[9\]
+ sky130_fd_sc_hd__dfrtp_4
X_3829_ _0819_ hkspi.state\[0\] hkspi.addr\[1\] VGND VGND VPWR VPWR _1405_ sky130_fd_sc_hd__o21ai_1
XFILLER_118_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6548_ clknet_leaf_35_csclk net1509 net525 VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__dfrtp_1
XFILLER_106_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6479_ clknet_leaf_61_csclk net678 net498 VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__dfstp_2
XFILLER_106_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput260 net260 VGND VGND VPWR VPWR pad_flash_io1_oeb sky130_fd_sc_hd__buf_12
Xoutput271 net271 VGND VGND VPWR VPWR pll_ena sky130_fd_sc_hd__buf_12
Xoutput282 net282 VGND VGND VPWR VPWR pll_trim[16] sky130_fd_sc_hd__buf_12
Xoutput293 net293 VGND VGND VPWR VPWR pll_trim[2] sky130_fd_sc_hd__buf_12
XFILLER_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_15_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xwire365 _2850_ VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__clkbuf_2
XFILLER_156_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_171_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5850_ gpio_configure\[16\]\[7\] _0831_ VGND VGND VPWR VPWR _2678_ sky130_fd_sc_hd__or2_1
X_4801_ _1601_ _1756_ _1781_ _1955_ VGND VGND VPWR VPWR _2012_ sky130_fd_sc_hd__a31o_1
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5781_ gpio_configure\[22\]\[4\] _2498_ _2518_ gpio_configure\[3\]\[4\] VGND VGND
+ VPWR VPWR _2612_ sky130_fd_sc_hd__a22o_1
XFILLER_9_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4732_ _1591_ _1612_ _1943_ VGND VGND VPWR VPWR _1944_ sky130_fd_sc_hd__and3_1
XFILLER_187_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4663_ _1688_ _1782_ VGND VGND VPWR VPWR _1875_ sky130_fd_sc_hd__nor2_1
XFILLER_174_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3614_ gpio_configure\[3\]\[2\] _0915_ net350 gpio_configure\[4\]\[2\] VGND VGND
+ VPWR VPWR _1203_ sky130_fd_sc_hd__a22o_1
X_6402_ net513 net483 VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__and2_1
X_4594_ _1779_ _1805_ VGND VGND VPWR VPWR _1806_ sky130_fd_sc_hd__nor2_1
Xhold902 net2125 VGND VGND VPWR VPWR net1435 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_128_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold913 _0694_ VGND VGND VPWR VPWR net1446 sky130_fd_sc_hd__dlygate4sd3_1
X_3545_ _1135_ hkspi.ldata\[4\] _0970_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__mux2_1
X_6333_ gpio_configure\[16\]\[12\] _2831_ net412 gpio_configure\[9\]\[12\] VGND VGND
+ VPWR VPWR _3143_ sky130_fd_sc_hd__a22o_1
Xhold924 gpio_configure\[10\]\[1\] VGND VGND VPWR VPWR net1457 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_155_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold935 _0129_ VGND VGND VPWR VPWR net1468 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_127_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold946 gpio_configure\[30\]\[9\] VGND VGND VPWR VPWR net1479 sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 _0168_ VGND VGND VPWR VPWR net1490 sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 net1992 VGND VGND VPWR VPWR net1501 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6264_ gpio_configure\[1\]\[9\] _2802_ _2858_ gpio_configure\[24\]\[9\] _3060_ VGND
+ VGND VPWR VPWR _3077_ sky130_fd_sc_hd__a221o_1
XFILLER_103_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3476_ net385 _0903_ VGND VGND VPWR VPWR _1067_ sky130_fd_sc_hd__nor2_4
XFILLER_142_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold979 trap_output_dest VGND VGND VPWR VPWR net1512 sky130_fd_sc_hd__dlygate4sd3_1
X_5215_ net445 net724 _2397_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__mux2_1
X_6195_ net473 net2042 _2486_ VGND VGND VPWR VPWR _3011_ sky130_fd_sc_hd__o21a_1
Xhold1602 pad_count_1\[1\] VGND VGND VPWR VPWR net2135 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5146_ _2324_ _2349_ _2352_ VGND VGND VPWR VPWR _2353_ sky130_fd_sc_hd__or3_1
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1613 hkspi.state\[1\] VGND VGND VPWR VPWR net2146 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5077_ _1807_ net432 _2233_ _1793_ _1896_ VGND VGND VPWR VPWR _2286_ sky130_fd_sc_hd__o221a_1
XFILLER_151_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4028_ _1086_ net426 VGND VGND VPWR VPWR _1476_ sky130_fd_sc_hd__and2_2
XFILLER_44_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5979_ _2471_ _2800_ VGND VGND VPWR VPWR _2801_ sky130_fd_sc_hd__nand2_8
XFILLER_40_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold209 net1975 VGND VGND VPWR VPWR net742 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_125_652 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_166_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3330_ net608 _0880_ VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__nand2_8
XFILLER_124_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_611 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ net607 net599 VGND VGND VPWR VPWR _0857_ sky130_fd_sc_hd__and2b_4
XFILLER_124_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _1952_ _2209_ _1618_ VGND VGND VPWR VPWR _2210_ sky130_fd_sc_hd__a21oi_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3192_ hkspi.state\[2\] VGND VGND VPWR VPWR _0821_ sky130_fd_sc_hd__inv_2
XFILLER_39_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6951_ clknet_leaf_39_csclk net1103 net517 VGND VGND VPWR VPWR gpio_configure\[13\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5902_ gpio_configure\[0\]\[9\] _2526_ _2717_ _2727_ net473 VGND VGND VPWR VPWR _2728_
+ sky130_fd_sc_hd__o221a_1
XFILLER_46_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6882_ clknet_3_5_0_csclk net1776 net513 VGND VGND VPWR VPWR gpio_configure\[5\]\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5833_ gpio_configure\[3\]\[6\] _2518_ _2520_ gpio_configure\[8\]\[6\] VGND VGND
+ VPWR VPWR _2662_ sky130_fd_sc_hd__a22o_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5764_ gpio_configure\[10\]\[3\] net421 _2535_ gpio_configure\[23\]\[3\] _2595_ VGND
+ VGND VPWR VPWR _2596_ sky130_fd_sc_hd__a221o_1
X_4715_ _1690_ _1773_ _1882_ _1926_ VGND VGND VPWR VPWR _1927_ sky130_fd_sc_hd__a211o_1
X_5695_ gpio_configure\[7\]\[0\] _2528_ _2529_ gpio_configure\[29\]\[0\] _2527_ VGND
+ VGND VPWR VPWR _2530_ sky130_fd_sc_hd__a221o_1
XFILLER_135_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4646_ _1790_ _1825_ VGND VGND VPWR VPWR _1858_ sky130_fd_sc_hd__or2_1
XFILLER_163_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold710 _0536_ VGND VGND VPWR VPWR net1243 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold721 gpio_configure\[29\]\[12\] VGND VGND VPWR VPWR net1254 sky130_fd_sc_hd__dlygate4sd3_1
X_4577_ _1782_ _1788_ VGND VGND VPWR VPWR _1789_ sky130_fd_sc_hd__nor2_1
XFILLER_162_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold732 _0457_ VGND VGND VPWR VPWR net1265 sky130_fd_sc_hd__dlygate4sd3_1
Xhold743 gpio_configure\[29\]\[11\] VGND VGND VPWR VPWR net1276 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold754 _0141_ VGND VGND VPWR VPWR net1287 sky130_fd_sc_hd__dlygate4sd3_1
X_6316_ net364 _3120_ _3126_ VGND VGND VPWR VPWR _3127_ sky130_fd_sc_hd__or3_1
XFILLER_116_674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3528_ net376 _0899_ VGND VGND VPWR VPWR _1119_ sky130_fd_sc_hd__nor2_2
XFILLER_143_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold765 gpio_configure\[15\]\[4\] VGND VGND VPWR VPWR net1298 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold776 _0477_ VGND VGND VPWR VPWR net1309 sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 gpio_configure\[6\]\[10\] VGND VGND VPWR VPWR net1320 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold798 _0614_ VGND VGND VPWR VPWR net1331 sky130_fd_sc_hd__dlygate4sd3_1
X_6247_ gpio_configure\[31\]\[9\] _2480_ _2814_ gpio_configure\[11\]\[9\] VGND VGND
+ VPWR VPWR _3060_ sky130_fd_sc_hd__a22o_1
X_3459_ gpio_configure\[13\]\[4\] _0906_ _0911_ gpio_configure\[21\]\[4\] VGND VGND
+ VPWR VPWR _1050_ sky130_fd_sc_hd__a22o_1
XFILLER_103_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6178_ gpio_configure\[32\]\[6\] _2813_ _2860_ gpio_configure\[17\]\[6\] VGND VGND
+ VPWR VPWR _2994_ sky130_fd_sc_hd__a22o_1
Xhold1410 net321 VGND VGND VPWR VPWR net1943 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1421 net318 VGND VGND VPWR VPWR net1954 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1432 wbbd_addr\[5\] VGND VGND VPWR VPWR net1965 sky130_fd_sc_hd__dlygate4sd3_1
X_5129_ _2331_ _2336_ _2277_ VGND VGND VPWR VPWR _2337_ sky130_fd_sc_hd__a21oi_2
Xhold1443 gpio_configure\[28\]\[0\] VGND VGND VPWR VPWR net1976 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1454 _0661_ VGND VGND VPWR VPWR net1987 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1465 _0388_ VGND VGND VPWR VPWR net1998 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1476 net332 VGND VGND VPWR VPWR net2009 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1487 wbbd_state\[3\] VGND VGND VPWR VPWR net2020 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1498 net345 VGND VGND VPWR VPWR net2031 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_138_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_742 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold70 _2441_ VGND VGND VPWR VPWR net603 sky130_fd_sc_hd__buf_6
XFILLER_48_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold81 mgmt_gpio_data_buf\[15\] VGND VGND VPWR VPWR net614 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_63_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold92 _0838_ VGND VGND VPWR VPWR net625 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4500_ _1561_ _1562_ _1581_ _1592_ _1603_ VGND VGND VPWR VPWR _1712_ sky130_fd_sc_hd__a2111o_1
XFILLER_129_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5480_ net446 net1172 net612 VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__mux2_1
XFILLER_8_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1 _0831_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4431_ _0834_ _1631_ VGND VGND VPWR VPWR _1643_ sky130_fd_sc_hd__nand2_4
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7150_ clknet_3_0_0_wb_clk_i _0753_ net499 VGND VGND VPWR VPWR pad_count_1\[2\] sky130_fd_sc_hd__dfrtp_1
X_4362_ _1571_ _1573_ VGND VGND VPWR VPWR _1574_ sky130_fd_sc_hd__nor2_1
X_3313_ net589 _0879_ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__nand2_8
X_6101_ gpio_configure\[13\]\[3\] net417 net406 gpio_configure\[27\]\[3\] VGND VGND
+ VPWR VPWR _2920_ sky130_fd_sc_hd__a22o_1
Xfanout508 net527 VGND VGND VPWR VPWR net508 sky130_fd_sc_hd__buf_8
X_7081_ clknet_leaf_58_csclk net1291 net502 VGND VGND VPWR VPWR gpio_configure\[29\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_59_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4293_ net446 net1164 _1540_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__mux2_1
Xfanout519 net521 VGND VGND VPWR VPWR net519 sky130_fd_sc_hd__buf_8
XFILLER_98_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3244_ hkspi.addr\[5\] net605 VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__and2_1
X_6032_ gpio_configure\[34\]\[0\] net393 net392 gpio_configure\[5\]\[0\] _2853_ VGND
+ VGND VPWR VPWR _2854_ sky130_fd_sc_hd__a221o_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6934_ clknet_leaf_25_csclk net711 net518 VGND VGND VPWR VPWR gpio_configure\[11\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6865_ clknet_leaf_52_csclk net1101 net507 VGND VGND VPWR VPWR gpio_configure\[2\]\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_5816_ net2049 _2645_ _2486_ VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__mux2_1
X_6796_ clknet_leaf_76_csclk net1068 net484 VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__dfrtp_4
XFILLER_167_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5747_ gpio_configure\[25\]\[2\] net420 _2512_ gpio_configure\[9\]\[2\] _2579_ VGND
+ VGND VPWR VPWR _2580_ sky130_fd_sc_hd__a221o_1
XFILLER_157_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5678_ pad_count_1\[4\] _2459_ _2493_ VGND VGND VPWR VPWR _2513_ sky130_fd_sc_hd__and3_4
XFILLER_163_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_175_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4629_ net477 _1777_ VGND VGND VPWR VPWR _1841_ sky130_fd_sc_hd__or2_1
Xhold540 gpio_configure\[18\]\[11\] VGND VGND VPWR VPWR net1073 sky130_fd_sc_hd__dlygate4sd3_1
Xhold551 _0173_ VGND VGND VPWR VPWR net1084 sky130_fd_sc_hd__dlygate4sd3_1
Xhold562 gpio_configure\[27\]\[7\] VGND VGND VPWR VPWR net1095 sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 gpio_configure\[6\]\[5\] VGND VGND VPWR VPWR net1106 sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 _0119_ VGND VGND VPWR VPWR net1117 sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 gpio_configure\[0\]\[7\] VGND VGND VPWR VPWR net1128 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_131_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1240 gpio_configure\[13\]\[8\] VGND VGND VPWR VPWR net1773 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_45_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1251 _0314_ VGND VGND VPWR VPWR net1784 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1262 _0509_ VGND VGND VPWR VPWR net1795 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1273 gpio_configure\[14\]\[8\] VGND VGND VPWR VPWR net1806 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1284 _0369_ VGND VGND VPWR VPWR net1817 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1295 gpio_configure\[24\]\[8\] VGND VGND VPWR VPWR net1828 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_163_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput160 wb_dat_i[6] VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_1
XFILLER_63_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4980_ _1815_ _1869_ _1988_ VGND VGND VPWR VPWR _2190_ sky130_fd_sc_hd__or3_1
X_3931_ _1455_ net38 hkspi.pass_thru_user VGND VGND VPWR VPWR _1456_ sky130_fd_sc_hd__mux2_1
XFILLER_32_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6650_ clknet_3_1_0_wb_clk_i _0263_ VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__dfxtp_1
XFILLER_177_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3862_ net1956 net2054 _1417_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__mux2_1
XFILLER_32_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5601_ xfer_count\[0\] xfer_count\[1\] xfer_state\[3\] net475 _2444_ VGND VGND VPWR
+ VPWR _2452_ sky130_fd_sc_hd__o221a_1
X_6581_ clknet_leaf_35_csclk net771 net525 VGND VGND VPWR VPWR mgmt_gpio_data_buf\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_3793_ hkspi.state\[3\] hkspi.state\[2\] VGND VGND VPWR VPWR _1378_ sky130_fd_sc_hd__or2_1
XFILLER_145_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5532_ net1670 net455 _2435_ VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__mux2_1
XFILLER_192_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_9_csclk clknet_3_4_0_csclk VGND VGND VPWR VPWR clknet_leaf_9_csclk sky130_fd_sc_hd__clkbuf_16
X_5463_ net441 net1206 _2427_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__mux2_1
XFILLER_172_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7202_ clknet_3_6_0_wb_clk_i _0804_ net529 VGND VGND VPWR VPWR wbbd_data\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_132_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4414_ _1554_ _1610_ net128 VGND VGND VPWR VPWR _1626_ sky130_fd_sc_hd__a21oi_1
X_5394_ _0912_ net647 VGND VGND VPWR VPWR _2420_ sky130_fd_sc_hd__and2_4
X_7133_ clknet_leaf_55_csclk net1392 net506 VGND VGND VPWR VPWR gpio_configure\[36\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_4345_ net110 net99 net124 net530 VGND VGND VPWR VPWR _1557_ sky130_fd_sc_hd__o211a_4
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4276_ _1109_ net429 VGND VGND VPWR VPWR _1538_ sky130_fd_sc_hd__nand2_2
X_7064_ clknet_leaf_32_csclk net642 net524 VGND VGND VPWR VPWR gpio_configure\[27\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_101_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6015_ _2793_ _2796_ _2809_ VGND VGND VPWR VPWR _2837_ sky130_fd_sc_hd__and3_4
X_3227_ gpio_configure\[7\]\[3\] VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__inv_2
XFILLER_39_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6917_ clknet_leaf_36_csclk net1139 net522 VGND VGND VPWR VPWR gpio_configure\[9\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_52_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6848_ clknet_leaf_50_csclk net1335 net506 VGND VGND VPWR VPWR gpio_configure\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_167_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6779_ clknet_3_6_0_wb_clk_i _0382_ net529 VGND VGND VPWR VPWR wbbd_addr\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_183_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_148_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_108_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold370 _0132_ VGND VGND VPWR VPWR net903 sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 net225 VGND VGND VPWR VPWR net914 sky130_fd_sc_hd__dlygate4sd3_1
Xhold392 _0411_ VGND VGND VPWR VPWR net925 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1070 _0706_ VGND VGND VPWR VPWR net1603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1081 net231 VGND VGND VPWR VPWR net1614 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1092 gpio_configure\[8\]\[9\] VGND VGND VPWR VPWR net1625 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_210 gpio_configure\[17\]\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_221 net351 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_232 net451 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_243 _0919_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_254 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_158_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_1_0__f__1134_ clknet_0__1134_ VGND VGND VPWR VPWR clknet_1_0__leaf__1134_
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_114_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_174_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4130_ net1796 net466 _1511_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__mux2_1
XFILLER_3_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4061_ net1485 _1485_ _1481_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__mux2_1
XFILLER_49_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_83_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_110_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_91_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_52_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4963_ _1760_ _2129_ VGND VGND VPWR VPWR _2173_ sky130_fd_sc_hd__or2_1
XFILLER_51_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6702_ clknet_leaf_2_csclk net1464 net493 VGND VGND VPWR VPWR gpio_configure\[14\]\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_3914_ net2067 net2076 _1408_ _1384_ _0819_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__o32ai_1
X_4894_ _1961_ _2104_ _2083_ _1702_ VGND VGND VPWR VPWR _2105_ sky130_fd_sc_hd__or4b_1
XFILLER_149_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6633_ clknet_3_5_0_wb_clk_i _0246_ VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__dfxtp_1
X_3845_ net58 net2066 _1413_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__mux2_1
XFILLER_20_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_192_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6564_ clknet_3_2_0_wb_clk_i _0016_ net499 VGND VGND VPWR VPWR xfer_state\[2\] sky130_fd_sc_hd__dfrtp_4
X_3776_ serial_busy _0974_ _1076_ gpio_configure\[27\]\[8\] _1361_ VGND VGND VPWR
+ VPWR _1362_ sky130_fd_sc_hd__a221o_1
XFILLER_138_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_164_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5515_ net451 net1924 _2433_ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__mux2_1
X_6495_ clknet_leaf_73_csclk net667 net488 VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__dfstp_2
XFILLER_173_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5446_ net437 net1354 _2425_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__mux2_1
XFILLER_133_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5377_ net470 net1765 _2418_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__mux2_1
XFILLER_99_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7116_ clknet_leaf_33_csclk net1527 net525 VGND VGND VPWR VPWR gpio_configure\[34\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_4328_ net768 net451 _1546_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__mux2_1
XFILLER_47_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_7047_ clknet_leaf_39_csclk net1115 net516 VGND VGND VPWR VPWR gpio_configure\[25\]\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_4259_ net1783 net470 _1535_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__mux2_1
XFILLER_28_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_103_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_124_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_534 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3630_ gpio_configure\[6\]\[10\] _1042_ _1080_ gpio_configure\[16\]\[10\] _1199_
+ VGND VGND VPWR VPWR _1219_ sky130_fd_sc_hd__a221o_1
XFILLER_186_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3561_ gpio_configure\[26\]\[3\] net371 _1086_ gpio_configure\[29\]\[11\] VGND VGND
+ VPWR VPWR _1151_ sky130_fd_sc_hd__a22o_1
XFILLER_115_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5300_ net447 net1180 _2409_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__mux2_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3492_ net387 _1006_ VGND VGND VPWR VPWR _1083_ sky130_fd_sc_hd__nor2_4
X_6280_ _3087_ _3088_ _3090_ _3091_ VGND VGND VPWR VPWR _3092_ sky130_fd_sc_hd__or4_1
XFILLER_142_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5231_ net461 net1612 _2401_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__mux2_1
XFILLER_103_709 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_102_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_130_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5162_ _2042_ _2052_ _2263_ _2368_ VGND VGND VPWR VPWR _2369_ sky130_fd_sc_hd__nor4_1
Xclkbuf_leaf_12_csclk clknet_3_5_0_csclk VGND VGND VPWR VPWR clknet_leaf_12_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_111_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4113_ net465 net770 net630 VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__mux2_1
XFILLER_68_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5093_ _1635_ _1706_ _1840_ _1996_ VGND VGND VPWR VPWR _2302_ sky130_fd_sc_hd__a211o_1
XFILLER_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4044_ net449 net1280 _1478_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__mux2_1
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_27_csclk clknet_3_5_0_csclk VGND VGND VPWR VPWR clknet_leaf_27_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_52_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5995_ gpio_configure\[31\]\[0\] _2480_ _2816_ gpio_configure\[29\]\[0\] VGND VGND
+ VPWR VPWR _2817_ sky130_fd_sc_hd__a22o_1
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4946_ _2038_ _2151_ _2153_ _2155_ VGND VGND VPWR VPWR _2156_ sky130_fd_sc_hd__or4b_1
XFILLER_193_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4877_ _1662_ _1667_ _1962_ VGND VGND VPWR VPWR _2088_ sky130_fd_sc_hd__a21o_1
X_6616_ clknet_leaf_12_csclk net1756 net512 VGND VGND VPWR VPWR gpio_configure\[4\]\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_3828_ _1404_ net2116 _1388_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__mux2_1
XFILLER_20_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6547_ clknet_leaf_35_csclk net959 net525 VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__dfrtp_1
X_3759_ gpio_configure\[35\]\[0\] _0932_ net350 gpio_configure\[4\]\[0\] _1323_ VGND
+ VGND VPWR VPWR _1345_ sky130_fd_sc_hd__a221o_1
XFILLER_192_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6478_ clknet_leaf_71_csclk net1016 net490 VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__dfstp_1
XFILLER_133_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5429_ net434 net1256 _2423_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__mux2_1
XFILLER_160_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput250 net250 VGND VGND VPWR VPWR mgmt_gpio_out[9] sky130_fd_sc_hd__clkbuf_1
Xoutput261 net261 VGND VGND VPWR VPWR pll90_sel[0] sky130_fd_sc_hd__buf_12
XFILLER_121_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput272 net272 VGND VGND VPWR VPWR pll_sel[0] sky130_fd_sc_hd__buf_12
Xoutput283 net283 VGND VGND VPWR VPWR pll_trim[17] sky130_fd_sc_hd__buf_12
XFILLER_59_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput294 net294 VGND VGND VPWR VPWR pll_trim[3] sky130_fd_sc_hd__buf_12
XFILLER_114_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_114_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_55_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_129_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_1_1_1_wb_clk_i clknet_1_1_0_wb_clk_i VGND VGND VPWR VPWR clknet_1_1_1_wb_clk_i
+ sky130_fd_sc_hd__clkbuf_8
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_151_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4800_ _1781_ _1792_ _1965_ VGND VGND VPWR VPWR _2011_ sky130_fd_sc_hd__a21o_1
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5780_ gpio_configure\[14\]\[4\] _2494_ _2540_ gpio_configure\[12\]\[4\] _2610_ VGND
+ VGND VPWR VPWR _2611_ sky130_fd_sc_hd__a221o_1
XFILLER_21_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4731_ _1679_ _1616_ _1615_ VGND VGND VPWR VPWR _1943_ sky130_fd_sc_hd__and3b_1
XFILLER_187_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4662_ _1580_ _1601_ VGND VGND VPWR VPWR _1874_ sky130_fd_sc_hd__nand2_2
X_6401_ net513 net483 VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__and2_1
X_3613_ gpio_configure\[13\]\[2\] _0906_ _0918_ gpio_configure\[15\]\[2\] VGND VGND
+ VPWR VPWR _1202_ sky130_fd_sc_hd__a22o_1
X_4593_ net477 _1803_ VGND VGND VPWR VPWR _1805_ sky130_fd_sc_hd__or2_4
Xhold903 _0704_ VGND VGND VPWR VPWR net1436 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_134_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6332_ _3130_ _3132_ _3141_ VGND VGND VPWR VPWR _3142_ sky130_fd_sc_hd__or3_1
Xhold914 gpio_configure\[9\]\[2\] VGND VGND VPWR VPWR net1447 sky130_fd_sc_hd__dlygate4sd3_1
X_3544_ clknet_1_0__leaf__1134_ net1995 _0837_ VGND VGND VPWR VPWR _1135_ sky130_fd_sc_hd__mux2_1
Xhold925 _0526_ VGND VGND VPWR VPWR net1458 sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 gpio_configure\[22\]\[6\] VGND VGND VPWR VPWR net1469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold947 _0134_ VGND VGND VPWR VPWR net1480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 gpio_configure\[28\]\[9\] VGND VGND VPWR VPWR net1491 sky130_fd_sc_hd__dlygate4sd3_1
X_6263_ gpio_configure\[2\]\[9\] net398 _2843_ gpio_configure\[5\]\[9\] _3075_ VGND
+ VGND VPWR VPWR _3076_ sky130_fd_sc_hd__a221o_1
Xhold969 gpio_configure\[27\]\[8\] VGND VGND VPWR VPWR net1502 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3475_ net16 _0864_ _1065_ gpio_configure\[37\]\[12\] _1064_ VGND VGND VPWR VPWR
+ _1066_ sky130_fd_sc_hd__a221o_2
XFILLER_103_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5214_ _0974_ net427 VGND VGND VPWR VPWR _2397_ sky130_fd_sc_hd__nand2_2
X_6194_ gpio_configure\[0\]\[6\] net365 _3009_ net475 VGND VGND VPWR VPWR _3010_ sky130_fd_sc_hd__a211o_1
XFILLER_130_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1603 gpio_configure\[37\]\[6\] VGND VGND VPWR VPWR net2136 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5145_ _2187_ _2304_ _2351_ VGND VGND VPWR VPWR _2352_ sky130_fd_sc_hd__or3b_1
Xhold1614 serial_data_staging_2\[10\] VGND VGND VPWR VPWR net2147 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5076_ _1581_ net424 VGND VGND VPWR VPWR _2285_ sky130_fd_sc_hd__and2_2
XFILLER_44_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4027_ net1248 net444 _1475_ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__mux2_1
XFILLER_84_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5978_ pad_count_2\[3\] pad_count_2\[2\] VGND VGND VPWR VPWR _2800_ sky130_fd_sc_hd__nor2_4
X_4929_ net2069 _1530_ _2036_ _2139_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__o22a_1
XFILLER_166_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_623 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_152_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ net598 net1991 net474 VGND VGND VPWR VPWR _0856_ sky130_fd_sc_hd__mux2_2
XFILLER_140_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3191_ net2103 VGND VGND VPWR VPWR _0820_ sky130_fd_sc_hd__inv_2
XFILLER_39_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_743 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_66_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_26_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6950_ clknet_leaf_22_csclk net1191 net514 VGND VGND VPWR VPWR gpio_configure\[13\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_53_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5901_ _2719_ _2722_ _2724_ _2726_ VGND VGND VPWR VPWR _2727_ sky130_fd_sc_hd__or4_1
XFILLER_34_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6881_ clknet_leaf_32_csclk net931 net523 VGND VGND VPWR VPWR gpio_configure\[4\]\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_5832_ gpio_configure\[13\]\[6\] _2501_ _2540_ gpio_configure\[12\]\[6\] _2660_ VGND
+ VGND VPWR VPWR _2661_ sky130_fd_sc_hd__a221o_1
XFILLER_34_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5763_ gpio_configure\[24\]\[3\] _2531_ _2532_ gpio_configure\[18\]\[3\] VGND VGND
+ VPWR VPWR _2595_ sky130_fd_sc_hd__a22o_1
XFILLER_148_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4714_ _1897_ _1925_ _1899_ _1898_ VGND VGND VPWR VPWR _1926_ sky130_fd_sc_hd__or4b_1
X_5694_ pad_count_1\[4\] _2493_ _2495_ VGND VGND VPWR VPWR _2529_ sky130_fd_sc_hd__and3_4
XFILLER_187_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4645_ net424 _1822_ VGND VGND VPWR VPWR _1857_ sky130_fd_sc_hd__or2_1
XFILLER_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold700 _0190_ VGND VGND VPWR VPWR net1233 sky130_fd_sc_hd__dlygate4sd3_1
Xhold711 gpio_configure\[21\]\[11\] VGND VGND VPWR VPWR net1244 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_146_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4576_ net477 _1787_ VGND VGND VPWR VPWR _1788_ sky130_fd_sc_hd__or2_4
Xhold722 _0147_ VGND VGND VPWR VPWR net1255 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap430 net645 VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__buf_12
Xhold733 gpio_configure\[24\]\[7\] VGND VGND VPWR VPWR net1266 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold744 _0146_ VGND VGND VPWR VPWR net1277 sky130_fd_sc_hd__dlygate4sd3_1
X_6315_ _3111_ _3122_ _3124_ _3125_ VGND VGND VPWR VPWR _3126_ sky130_fd_sc_hd__or4_1
Xhold755 net2120 VGND VGND VPWR VPWR net1288 sky130_fd_sc_hd__dlygate4sd3_1
X_3527_ gpio_configure\[26\]\[12\] _1116_ _1117_ net270 VGND VGND VPWR VPWR _1118_
+ sky130_fd_sc_hd__a22o_1
XFILLER_190_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold766 _0569_ VGND VGND VPWR VPWR net1299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 gpio_configure\[14\]\[12\] VGND VGND VPWR VPWR net1310 sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 _0249_ VGND VGND VPWR VPWR net1321 sky130_fd_sc_hd__dlygate4sd3_1
X_6246_ gpio_configure\[36\]\[9\] net403 net402 gpio_configure\[4\]\[9\] VGND VGND
+ VPWR VPWR _3059_ sky130_fd_sc_hd__a22o_2
Xhold799 net2105 VGND VGND VPWR VPWR net1332 sky130_fd_sc_hd__dlygate4sd3_1
X_3458_ gpio_configure\[13\]\[12\] _1045_ _1046_ gpio_configure\[28\]\[12\] _1048_
+ VGND VGND VPWR VPWR _1049_ sky130_fd_sc_hd__a221o_1
XFILLER_76_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6177_ gpio_configure\[20\]\[6\] net396 _2992_ VGND VGND VPWR VPWR _2993_ sky130_fd_sc_hd__a21o_1
XFILLER_162_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3389_ gpio_configure\[10\]\[6\] _0920_ _0921_ gpio_configure\[12\]\[6\] VGND VGND
+ VPWR VPWR _0983_ sky130_fd_sc_hd__a22o_1
Xhold1400 net323 VGND VGND VPWR VPWR net1933 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1411 net347 VGND VGND VPWR VPWR net1944 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1422 net339 VGND VGND VPWR VPWR net1955 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1433 _0893_ VGND VGND VPWR VPWR net1966 sky130_fd_sc_hd__dlygate4sd3_1
X_5128_ _2334_ _1884_ _2333_ _2335_ VGND VGND VPWR VPWR _2336_ sky130_fd_sc_hd__and4b_1
XFILLER_111_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1444 _0669_ VGND VGND VPWR VPWR net1977 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1455 wbbd_data\[4\] VGND VGND VPWR VPWR net1988 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1466 hkspi.ldata\[1\] VGND VGND VPWR VPWR net1999 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_84_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_29_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1477 mgmt_gpio_data_buf\[20\] VGND VGND VPWR VPWR net2010 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5059_ _1815_ _2161_ _2267_ VGND VGND VPWR VPWR _2268_ sky130_fd_sc_hd__nor3_1
Xhold1488 hkspi.odata\[7\] VGND VGND VPWR VPWR net2021 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1499 wbbd_state\[2\] VGND VGND VPWR VPWR net2032 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_111_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_111_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_21_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_642 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_153_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_697 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_656 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold60 _0297_ VGND VGND VPWR VPWR net593 sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 _0745_ VGND VGND VPWR VPWR net604 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_36_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold82 _0444_ VGND VGND VPWR VPWR net615 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 _0839_ VGND VGND VPWR VPWR net626 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_152_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_662 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4430_ net530 _1632_ VGND VGND VPWR VPWR _1642_ sky130_fd_sc_hd__nor2_4
XFILLER_6_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_2 _0874_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4361_ _1553_ _1557_ _1570_ net126 VGND VGND VPWR VPWR _1573_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_98_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6100_ gpio_configure\[36\]\[3\] net403 net402 gpio_configure\[4\]\[3\] _2918_ VGND
+ VGND VPWR VPWR _2919_ sky130_fd_sc_hd__a221o_1
X_3312_ _0873_ net376 VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__nor2_8
XFILLER_98_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_112_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7080_ clknet_leaf_59_csclk net1460 net502 VGND VGND VPWR VPWR gpio_configure\[29\]\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_112_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout509 net510 VGND VGND VPWR VPWR net509 sky130_fd_sc_hd__buf_8
X_4292_ net569 net683 _1540_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__mux2_1
XFILLER_152_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6031_ gpio_configure\[8\]\[0\] net410 _2852_ gpio_configure\[19\]\[0\] VGND VGND
+ VPWR VPWR _2853_ sky130_fd_sc_hd__a22o_1
X_3243_ net579 net605 net625 VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__a21oi_1
XFILLER_98_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6933_ clknet_leaf_37_csclk net1243 net522 VGND VGND VPWR VPWR gpio_configure\[11\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_35_673 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6864_ clknet_leaf_52_csclk net1376 net506 VGND VGND VPWR VPWR gpio_configure\[2\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_179_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_22_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5815_ net475 serial_data_staging_1\[4\] _2644_ VGND VGND VPWR VPWR _2645_ sky130_fd_sc_hd__a21o_1
XFILLER_179_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6795_ clknet_leaf_76_csclk net1683 net484 VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__dfstp_1
XFILLER_148_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5746_ gpio_configure\[4\]\[2\] _2502_ _2538_ gpio_configure\[1\]\[2\] VGND VGND
+ VPWR VPWR _2579_ sky130_fd_sc_hd__a22o_1
XFILLER_182_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5677_ net472 _2495_ _2504_ VGND VGND VPWR VPWR _2512_ sky130_fd_sc_hd__and3_4
XFILLER_108_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4628_ _1800_ _1825_ VGND VGND VPWR VPWR _1840_ sky130_fd_sc_hd__nor2_2
Xhold530 gpio_configure\[22\]\[12\] VGND VGND VPWR VPWR net1063 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold541 _0337_ VGND VGND VPWR VPWR net1074 sky130_fd_sc_hd__dlygate4sd3_1
X_4559_ _1604_ _1758_ VGND VGND VPWR VPWR _1771_ sky130_fd_sc_hd__and2_2
Xhold552 net262 VGND VGND VPWR VPWR net1085 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_739 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_9_8 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold563 _0668_ VGND VGND VPWR VPWR net1096 sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 _0498_ VGND VGND VPWR VPWR net1107 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold585 gpio_configure\[2\]\[12\] VGND VGND VPWR VPWR net1118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 _0452_ VGND VGND VPWR VPWR net1129 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6229_ gpio_configure\[22\]\[8\] _2824_ _2829_ gpio_configure\[33\]\[8\] _3042_ VGND
+ VGND VPWR VPWR _3043_ sky130_fd_sc_hd__a221o_1
XFILLER_77_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1230 gpio_configure\[1\]\[0\] VGND VGND VPWR VPWR net1763 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1241 _0299_ VGND VGND VPWR VPWR net1774 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1252 gpio_configure\[28\]\[8\] VGND VGND VPWR VPWR net1785 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1263 gpio_configure\[0\]\[8\] VGND VGND VPWR VPWR net1796 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1274 _0304_ VGND VGND VPWR VPWR net1807 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1285 net2144 VGND VGND VPWR VPWR net1818 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1296 _0138_ VGND VGND VPWR VPWR net1829 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_127_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_126_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_48_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput150 wb_dat_i[26] VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_1
Xinput161 wb_dat_i[7] VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3930_ mgmt_gpio_data\[1\] hkspi.SDO net482 VGND VGND VPWR VPWR _1455_ sky130_fd_sc_hd__mux2_1
XFILLER_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3861_ net2054 hkspi.odata\[6\] _1417_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__mux2_1
XFILLER_189_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5600_ xfer_count\[0\] xfer_count\[1\] VGND VGND VPWR VPWR _2451_ sky130_fd_sc_hd__nand2_1
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6580_ clknet_leaf_35_csclk net1327 net525 VGND VGND VPWR VPWR mgmt_gpio_data_buf\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_3792_ net2090 _0970_ _1376_ _1377_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__a22o_1
XFILLER_192_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5531_ net1445 net462 _2435_ VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__mux2_1
XFILLER_185_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5462_ net446 net1156 _2427_ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__mux2_1
X_7201_ clknet_3_6_0_wb_clk_i _0803_ net529 VGND VGND VPWR VPWR wbbd_data\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_133_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4413_ _1554_ _1610_ _1624_ VGND VGND VPWR VPWR _1625_ sky130_fd_sc_hd__a21boi_2
X_5393_ net434 net1134 _2419_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__mux2_1
X_7132_ clknet_leaf_34_csclk net1561 net525 VGND VGND VPWR VPWR gpio_configure\[36\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_4344_ net110 net99 VGND VGND VPWR VPWR _1556_ sky130_fd_sc_hd__or2_1
XFILLER_86_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7063_ clknet_leaf_31_csclk net1537 net523 VGND VGND VPWR VPWR gpio_configure\[27\]\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_4275_ net1104 net446 _1537_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__mux2_1
XFILLER_100_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6014_ _1448_ _2473_ _2796_ VGND VGND VPWR VPWR _2836_ sky130_fd_sc_hd__and3_1
XFILLER_140_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3226_ gpio_configure\[8\]\[3\] VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__inv_2
XFILLER_39_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_67_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6916_ clknet_leaf_47_csclk net1448 net514 VGND VGND VPWR VPWR gpio_configure\[9\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_70_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6847_ clknet_leaf_43_csclk net1155 net517 VGND VGND VPWR VPWR gpio_configure\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_168_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6778_ clknet_3_6_0_wb_clk_i _0381_ net529 VGND VGND VPWR VPWR wbbd_addr\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_139_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5729_ gpio_configure\[0\]\[1\] _2526_ _2553_ _2562_ _0824_ VGND VGND VPWR VPWR _2563_
+ sky130_fd_sc_hd__o221a_1
XFILLER_182_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_190_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold360 _0638_ VGND VGND VPWR VPWR net893 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_117_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold371 gpio_configure\[32\]\[1\] VGND VGND VPWR VPWR net904 sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 _0167_ VGND VGND VPWR VPWR net915 sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 gpio_configure\[35\]\[7\] VGND VGND VPWR VPWR net926 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_77_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1060 _0395_ VGND VGND VPWR VPWR net1593 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1071 gpio_configure\[36\]\[0\] VGND VGND VPWR VPWR net1604 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1082 _0431_ VGND VGND VPWR VPWR net1615 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1093 _0274_ VGND VGND VPWR VPWR net1626 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_200 _2421_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_211 gpio_configure\[21\]\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_716 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_222 net352 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_233 net457 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_244 _1086_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_255 net457 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_42_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_68_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4060_ net1005 net453 net356 VGND VGND VPWR VPWR _1485_ sky130_fd_sc_hd__mux2_1
XFILLER_49_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_24_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4962_ _2140_ _2171_ VGND VGND VPWR VPWR _2172_ sky130_fd_sc_hd__nor2_1
X_3913_ net2102 hkspi.state\[0\] _1384_ net2097 VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__a31o_1
X_6701_ clknet_leaf_2_csclk net1807 net493 VGND VGND VPWR VPWR gpio_configure\[14\]\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_51_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4893_ _1667_ _2082_ _2103_ VGND VGND VPWR VPWR _2104_ sky130_fd_sc_hd__a21o_1
X_6632_ clknet_3_5_0_wb_clk_i _0245_ VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__dfxtp_1
X_3844_ hkspi.count\[2\] hkspi.count\[1\] hkspi.count\[0\] hkspi.state\[0\] VGND VGND
+ VPWR VPWR _1413_ sky130_fd_sc_hd__or4b_1
XFILLER_20_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6563_ clknet_3_3_0_wb_clk_i _0015_ net502 VGND VGND VPWR VPWR xfer_state\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_158_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3775_ net272 _1009_ _1041_ gpio_configure\[31\]\[8\] VGND VGND VPWR VPWR _1361_
+ sky130_fd_sc_hd__a22o_1
XFILLER_164_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5514_ net457 net840 _2433_ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__mux2_1
XFILLER_145_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6494_ clknet_leaf_73_csclk net1050 net488 VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__dfstp_1
XFILLER_145_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_133_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5445_ net440 net1518 _2425_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__mux2_1
XFILLER_173_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5376_ net373 net429 VGND VGND VPWR VPWR _2418_ sky130_fd_sc_hd__nand2_8
XFILLER_154_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7115_ clknet_leaf_62_csclk net789 net508 VGND VGND VPWR VPWR gpio_configure\[34\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_59_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4327_ net1216 net456 _1546_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__mux2_1
XFILLER_99_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_7046_ clknet_leaf_19_csclk net1173 net510 VGND VGND VPWR VPWR gpio_configure\[25\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_4258_ _1080_ net429 VGND VGND VPWR VPWR _1535_ sky130_fd_sc_hd__and2_1
XFILLER_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3209_ gpio_configure\[25\]\[3\] VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__inv_2
XFILLER_27_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4189_ wbbd_state\[3\] net528 VGND VGND VPWR VPWR _1520_ sky130_fd_sc_hd__and2_4
XFILLER_28_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_10_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_151_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold190 _0481_ VGND VGND VPWR VPWR net723 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_144_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_104_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_120_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_679 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_65_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_8_csclk clknet_3_4_0_csclk VGND VGND VPWR VPWR clknet_leaf_8_csclk sky130_fd_sc_hd__clkbuf_16
XFILLER_160_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_61_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3560_ gpio_configure\[18\]\[3\] _0894_ _1062_ gpio_configure\[21\]\[11\] VGND VGND
+ VPWR VPWR _1150_ sky130_fd_sc_hd__a22o_1
XFILLER_10_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3491_ gpio_configure\[16\]\[12\] _1080_ _1081_ gpio_configure\[34\]\[12\] _1079_
+ VGND VGND VPWR VPWR _1082_ sky130_fd_sc_hd__a221o_1
XFILLER_5_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5230_ net467 net1610 _2401_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__mux2_1
XFILLER_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_676 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5161_ _1692_ _1873_ _1702_ VGND VGND VPWR VPWR _2368_ sky130_fd_sc_hd__o21ai_1
XFILLER_68_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4112_ net471 net1326 net630 VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__mux2_1
X_5092_ _1991_ _2192_ _2299_ _2300_ VGND VGND VPWR VPWR _2301_ sky130_fd_sc_hd__or4_1
XFILLER_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4043_ net455 net1746 _1478_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__mux2_1
XFILLER_84_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5994_ _2471_ _2473_ _2478_ VGND VGND VPWR VPWR _2816_ sky130_fd_sc_hd__and3_4
X_4945_ net110 _1694_ _2154_ _1681_ _1700_ VGND VGND VPWR VPWR _2155_ sky130_fd_sc_hd__o221a_1
XFILLER_177_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4876_ _1629_ _1749_ VGND VGND VPWR VPWR _2087_ sky130_fd_sc_hd__nand2_1
XFILLER_177_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_443 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6615_ clknet_leaf_3_csclk net1251 net494 VGND VGND VPWR VPWR gpio_configure\[3\]\[12\]
+ sky130_fd_sc_hd__dfrtp_2
X_3827_ hkspi.addr\[1\] hkspi.state\[3\] _1399_ _1403_ VGND VGND VPWR VPWR _1404_
+ sky130_fd_sc_hd__a22o_1
XFILLER_137_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6546_ clknet_leaf_36_csclk net1723 net525 VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__dfrtp_1
X_3758_ gpio_configure\[8\]\[0\] _0939_ _1081_ gpio_configure\[34\]\[8\] _1315_ VGND
+ VGND VPWR VPWR _1344_ sky130_fd_sc_hd__a221o_1
XFILLER_180_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6477_ clknet_leaf_71_csclk net1062 net490 VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__dfstp_1
XFILLER_118_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3689_ _1267_ _1276_ VGND VGND VPWR VPWR _1277_ sky130_fd_sc_hd__or2_1
XFILLER_133_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5428_ net437 net1425 _2423_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__mux2_1
XFILLER_161_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput240 net240 VGND VGND VPWR VPWR mgmt_gpio_out[34] sky130_fd_sc_hd__buf_12
Xoutput251 net251 VGND VGND VPWR VPWR pad_flash_clk sky130_fd_sc_hd__clkbuf_1
Xoutput262 net262 VGND VGND VPWR VPWR pll90_sel[1] sky130_fd_sc_hd__buf_12
Xoutput273 net273 VGND VGND VPWR VPWR pll_sel[1] sky130_fd_sc_hd__buf_12
XFILLER_121_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput284 net284 VGND VGND VPWR VPWR pll_trim[18] sky130_fd_sc_hd__buf_12
X_5359_ net470 net1748 _2416_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__mux2_1
Xoutput295 net295 VGND VGND VPWR VPWR pll_trim[4] sky130_fd_sc_hd__buf_12
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_160_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7029_ clknet_leaf_46_csclk net809 net515 VGND VGND VPWR VPWR gpio_configure\[23\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_74_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_169_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_137_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_136_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_686 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_20 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4730_ _1599_ _1665_ VGND VGND VPWR VPWR _1942_ sky130_fd_sc_hd__nor2_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4661_ _1588_ _1602_ VGND VGND VPWR VPWR _1873_ sky130_fd_sc_hd__or2_2
XFILLER_187_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6400_ net492 net481 VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__and2_1
X_3612_ gpio_configure\[12\]\[2\] _0921_ _1065_ gpio_configure\[37\]\[10\] VGND VGND
+ VPWR VPWR _1201_ sky130_fd_sc_hd__a22o_1
X_4592_ _1803_ VGND VGND VPWR VPWR _1804_ sky130_fd_sc_hd__inv_2
XFILLER_190_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6331_ _3134_ _3136_ _3138_ _3140_ VGND VGND VPWR VPWR _3141_ sky130_fd_sc_hd__or4_1
Xhold904 gpio_configure\[12\]\[1\] VGND VGND VPWR VPWR net1437 sky130_fd_sc_hd__dlygate4sd3_1
X_3543_ _1059_ _1075_ _1133_ VGND VGND VPWR VPWR _1134_ sky130_fd_sc_hd__or3_2
XFILLER_127_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold915 _0519_ VGND VGND VPWR VPWR net1448 sky130_fd_sc_hd__dlygate4sd3_1
Xhold926 gpio_configure\[29\]\[6\] VGND VGND VPWR VPWR net1459 sky130_fd_sc_hd__dlygate4sd3_1
Xhold937 _0627_ VGND VGND VPWR VPWR net1470 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold948 gpio_configure\[20\]\[9\] VGND VGND VPWR VPWR net1481 sky130_fd_sc_hd__dlygate4sd3_1
X_6262_ gpio_configure\[13\]\[9\] _2804_ _2862_ gpio_configure\[25\]\[9\] VGND VGND
+ VPWR VPWR _3075_ sky130_fd_sc_hd__a22o_1
Xhold959 _0154_ VGND VGND VPWR VPWR net1492 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3474_ net378 _0899_ VGND VGND VPWR VPWR _1065_ sky130_fd_sc_hd__nor2_4
XFILLER_115_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5213_ net1495 _1314_ net426 _2396_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__o211a_1
XFILLER_103_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6193_ _2996_ _2999_ _3008_ VGND VGND VPWR VPWR _3009_ sky130_fd_sc_hd__or3_1
XFILLER_142_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_97_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5144_ _1772_ _2350_ _1947_ _1842_ VGND VGND VPWR VPWR _2351_ sky130_fd_sc_hd__o211a_1
Xhold1604 hkspi.addr\[0\] VGND VGND VPWR VPWR net2137 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_57_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5075_ _1590_ _2283_ _2238_ _2223_ _2122_ VGND VGND VPWR VPWR _2284_ sky130_fd_sc_hd__o2111ai_4
XFILLER_151_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4026_ net1286 net450 _1475_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__mux2_1
XFILLER_37_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_25_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_64_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5977_ _1448_ _2473_ _2478_ VGND VGND VPWR VPWR _2799_ sky130_fd_sc_hd__and3_4
X_4928_ _1529_ _2080_ _2109_ _2138_ VGND VGND VPWR VPWR _2139_ sky130_fd_sc_hd__or4_1
XFILLER_21_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4859_ _1684_ _1793_ _2069_ _1637_ VGND VGND VPWR VPWR _2070_ sky130_fd_sc_hd__o211a_1
XFILLER_166_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6529_ clknet_leaf_76_csclk net1030 net484 VGND VGND VPWR VPWR gpio_configure\[25\]\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_180_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_106_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_134_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_88_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_73_csclk clknet_3_0_0_csclk VGND VGND VPWR VPWR clknet_leaf_73_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_11_csclk clknet_opt_2_0_csclk VGND VGND VPWR VPWR clknet_leaf_11_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_7_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_26_csclk clknet_3_5_0_csclk VGND VGND VPWR VPWR clknet_leaf_26_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_124_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_140_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_741 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3190_ net605 VGND VGND VPWR VPWR _0819_ sky130_fd_sc_hd__clkinv_2
XFILLER_94_711 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_94_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_81_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_47_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5900_ gpio_configure\[14\]\[9\] _2494_ _2535_ gpio_configure\[23\]\[9\] _2725_ VGND
+ VGND VPWR VPWR _2726_ sky130_fd_sc_hd__a221o_1
XFILLER_93_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6880_ clknet_leaf_32_csclk net651 net524 VGND VGND VPWR VPWR gpio_configure\[4\]\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_5831_ gpio_configure\[5\]\[6\] net422 net420 gpio_configure\[25\]\[6\] VGND VGND
+ VPWR VPWR _2660_ sky130_fd_sc_hd__a22o_1
XFILLER_34_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5762_ gpio_configure\[11\]\[3\] _2505_ _2521_ gpio_configure\[21\]\[3\] _2593_ VGND
+ VGND VPWR VPWR _2594_ sky130_fd_sc_hd__a221o_1
XFILLER_148_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4713_ _1870_ _1900_ _1923_ _1924_ VGND VGND VPWR VPWR _1925_ sky130_fd_sc_hd__nand4_1
X_5693_ net472 _2461_ _2488_ VGND VGND VPWR VPWR _2528_ sky130_fd_sc_hd__and3_4
XFILLER_147_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4644_ _1815_ _1820_ _1821_ _1855_ VGND VGND VPWR VPWR _1856_ sky130_fd_sc_hd__or4b_1
Xhold701 gpio_configure\[26\]\[4\] VGND VGND VPWR VPWR net1234 sky130_fd_sc_hd__dlygate4sd3_1
X_4575_ net126 _0836_ _1755_ VGND VGND VPWR VPWR _1787_ sky130_fd_sc_hd__or3_4
Xhold712 _0367_ VGND VGND VPWR VPWR net1245 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap420 _2511_ VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__buf_12
Xhold723 gpio_configure\[19\]\[7\] VGND VGND VPWR VPWR net1256 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_190_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3526_ _0873_ net383 VGND VGND VPWR VPWR _1117_ sky130_fd_sc_hd__nor2_8
Xhold734 _0644_ VGND VGND VPWR VPWR net1267 sky130_fd_sc_hd__dlygate4sd3_1
X_6314_ gpio_configure\[1\]\[11\] _2802_ _2858_ gpio_configure\[24\]\[11\] _3109_
+ VGND VGND VPWR VPWR _3125_ sky130_fd_sc_hd__a221o_1
Xhold745 gpio_configure\[23\]\[7\] VGND VGND VPWR VPWR net1278 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold756 _0208_ VGND VGND VPWR VPWR net1289 sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 gpio_configure\[20\]\[12\] VGND VGND VPWR VPWR net1300 sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 _0308_ VGND VGND VPWR VPWR net1311 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_116_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6245_ net2091 net366 _3057_ _3058_ VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__o22a_1
X_3457_ gpio_configure\[22\]\[4\] _0923_ _1047_ gpio_configure\[18\]\[12\] VGND VGND
+ VPWR VPWR _1048_ sky130_fd_sc_hd__a22o_1
Xhold789 gpio_configure\[13\]\[10\] VGND VGND VPWR VPWR net1322 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6176_ gpio_configure\[37\]\[6\] _2806_ net397 gpio_configure\[22\]\[6\] VGND VGND
+ VPWR VPWR _2992_ sky130_fd_sc_hd__a22o_1
XFILLER_162_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3388_ gpio_configure\[23\]\[6\] net372 _0934_ gpio_configure\[1\]\[6\] _0981_ VGND
+ VGND VPWR VPWR _0982_ sky130_fd_sc_hd__a221o_1
Xhold1401 net328 VGND VGND VPWR VPWR net1934 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1412 net349 VGND VGND VPWR VPWR net1945 sky130_fd_sc_hd__dlygate4sd3_1
X_5127_ _1691_ _2050_ _2269_ VGND VGND VPWR VPWR _2335_ sky130_fd_sc_hd__nor3_1
Xhold1423 hkspi.odata\[4\] VGND VGND VPWR VPWR net1956 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1434 _0896_ VGND VGND VPWR VPWR net1967 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1445 net336 VGND VGND VPWR VPWR net1978 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1456 net293 VGND VGND VPWR VPWR net1989 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1467 _0387_ VGND VGND VPWR VPWR net2000 sky130_fd_sc_hd__dlygate4sd3_1
X_5058_ _1580_ _1587_ _1675_ VGND VGND VPWR VPWR _2267_ sky130_fd_sc_hd__o21a_1
XFILLER_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1478 net324 VGND VGND VPWR VPWR net2011 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1489 _0074_ VGND VGND VPWR VPWR net2022 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4009_ net434 net1270 _1472_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__mux2_1
XTAP_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_654 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_122_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_668 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_121_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold50 _1129_ VGND VGND VPWR VPWR net583 sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 wbbd_data\[2\] VGND VGND VPWR VPWR net594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 hkspi.state\[3\] VGND VGND VPWR VPWR net605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 net1956 VGND VGND VPWR VPWR net616 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 _0865_ VGND VGND VPWR VPWR net627 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_35_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_674 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_3 _0886_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4360_ _1569_ _1570_ VGND VGND VPWR VPWR _1572_ sky130_fd_sc_hd__or2_1
XFILLER_125_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3311_ _0895_ net382 VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__nor2_8
XFILLER_125_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4291_ net577 net786 _1540_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__mux2_1
XFILLER_140_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6030_ _2469_ _2478_ _2800_ VGND VGND VPWR VPWR _2852_ sky130_fd_sc_hd__and3_4
X_3242_ net624 _0819_ VGND VGND VPWR VPWR _0838_ sky130_fd_sc_hd__and2_1
XFILLER_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6932_ clknet_leaf_28_csclk net1551 net521 VGND VGND VPWR VPWR gpio_configure\[11\]\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_47_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6863_ clknet_leaf_39_csclk net1123 net516 VGND VGND VPWR VPWR gpio_configure\[2\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_35_685 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_50_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5814_ gpio_configure\[0\]\[5\] _2526_ _2634_ _2643_ net473 VGND VGND VPWR VPWR _2644_
+ sky130_fd_sc_hd__o221a_2
X_6794_ clknet_leaf_77_csclk net1707 net484 VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__dfrtp_4
XFILLER_167_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5745_ gpio_configure\[10\]\[2\] net421 _2528_ gpio_configure\[7\]\[2\] _2577_ VGND
+ VGND VPWR VPWR _2578_ sky130_fd_sc_hd__a221o_1
X_5676_ pad_count_1\[4\] _2495_ _2504_ VGND VGND VPWR VPWR _2511_ sky130_fd_sc_hd__and3_4
XFILLER_148_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4627_ _1831_ _1832_ _1835_ _1837_ VGND VGND VPWR VPWR _1839_ sky130_fd_sc_hd__or4_1
XFILLER_163_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold520 gpio_configure\[10\]\[7\] VGND VGND VPWR VPWR net1053 sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 _0378_ VGND VGND VPWR VPWR net1064 sky130_fd_sc_hd__dlygate4sd3_1
X_4558_ _1759_ _1769_ VGND VGND VPWR VPWR _1770_ sky130_fd_sc_hd__nor2_2
XFILLER_190_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold542 gpio_configure\[26\]\[3\] VGND VGND VPWR VPWR net1075 sky130_fd_sc_hd__dlygate4sd3_1
Xhold553 _0405_ VGND VGND VPWR VPWR net1086 sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 wbbd_data\[0\] VGND VGND VPWR VPWR net1097 sky130_fd_sc_hd__dlygate4sd3_1
X_3509_ gpio_configure\[32\]\[4\] _0890_ net352 gpio_configure\[36\]\[4\] _1099_ VGND
+ VGND VPWR VPWR _1100_ sky130_fd_sc_hd__a221o_1
XFILLER_143_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold575 gpio_configure\[34\]\[3\] VGND VGND VPWR VPWR net1108 sky130_fd_sc_hd__dlygate4sd3_1
Xhold586 _0223_ VGND VGND VPWR VPWR net1119 sky130_fd_sc_hd__dlygate4sd3_1
X_4489_ _1575_ _1605_ _1684_ VGND VGND VPWR VPWR _1701_ sky130_fd_sc_hd__or3_1
XFILLER_104_657 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold597 gpio_configure\[13\]\[3\] VGND VGND VPWR VPWR net1130 sky130_fd_sc_hd__dlygate4sd3_1
X_6228_ gpio_configure\[18\]\[8\] _2819_ _2837_ gpio_configure\[8\]\[8\] VGND VGND
+ VPWR VPWR _3042_ sky130_fd_sc_hd__a22o_1
XFILLER_131_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6159_ gpio_configure\[9\]\[5\] net412 net409 gpio_configure\[12\]\[5\] VGND VGND
+ VPWR VPWR _2976_ sky130_fd_sc_hd__a22o_1
Xhold1220 gpio_configure\[19\]\[8\] VGND VGND VPWR VPWR net1753 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1231 _0453_ VGND VGND VPWR VPWR net1764 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1242 gpio_configure\[5\]\[0\] VGND VGND VPWR VPWR net1775 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1253 _0153_ VGND VGND VPWR VPWR net1786 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1264 _0209_ VGND VGND VPWR VPWR net1797 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1275 gpio_configure\[29\]\[8\] VGND VGND VPWR VPWR net1808 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1286 _0319_ VGND VGND VPWR VPWR net1819 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1297 gpio_configure\[23\]\[8\] VGND VGND VPWR VPWR net1830 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_181_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput140 wb_dat_i[17] VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_1
Xinput151 wb_dat_i[27] VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput162 wb_dat_i[8] VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_1
XFILLER_36_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_725 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3860_ hkspi.odata\[6\] net2021 _1417_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__mux2_1
XFILLER_31_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_677 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_72_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3791_ _0837_ _0970_ VGND VGND VPWR VPWR _1377_ sky130_fd_sc_hd__nor2_1
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5530_ net1822 net466 _2435_ VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__mux2_1
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5461_ net569 net808 _2427_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__mux2_1
X_4412_ _1553_ _1610_ net127 VGND VGND VPWR VPWR _1624_ sky130_fd_sc_hd__a21o_1
X_7200_ clknet_3_7_0_wb_clk_i _0802_ net529 VGND VGND VPWR VPWR wbbd_data\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_133_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5392_ net437 net1369 _2419_ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__mux2_1
XFILLER_99_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_172_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_7131_ clknet_leaf_25_csclk net705 net518 VGND VGND VPWR VPWR gpio_configure\[36\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_4343_ net124 net530 VGND VGND VPWR VPWR _1555_ sky130_fd_sc_hd__nand2_2
XFILLER_113_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7062_ clknet_leaf_23_csclk net655 net515 VGND VGND VPWR VPWR gpio_configure\[27\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_4274_ net679 net569 _1537_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__mux2_1
XFILLER_140_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6013_ _2471_ _2796_ _2809_ VGND VGND VPWR VPWR _2835_ sky130_fd_sc_hd__and3_1
X_3225_ gpio_configure\[9\]\[3\] VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__inv_2
XFILLER_140_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_36_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_54_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_82_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_27_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6915_ clknet_leaf_47_csclk net1422 net514 VGND VGND VPWR VPWR gpio_configure\[9\]\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_35_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_23_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6846_ clknet_leaf_65_csclk net690 net505 VGND VGND VPWR VPWR gpio_configure\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_167_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6777_ clknet_3_6_0_wb_clk_i _0380_ net529 VGND VGND VPWR VPWR wbbd_addr\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_167_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3989_ net673 net660 _1470_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__mux2_1
XFILLER_167_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5728_ _2555_ _2557_ _2559_ _2561_ VGND VGND VPWR VPWR _2562_ sky130_fd_sc_hd__or4_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5659_ net472 _2489_ _2493_ VGND VGND VPWR VPWR _2494_ sky130_fd_sc_hd__and3_4
XFILLER_163_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_117_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_527 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_89_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold350 _0185_ VGND VGND VPWR VPWR net883 sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 gpio_configure\[6\]\[12\] VGND VGND VPWR VPWR net894 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold372 _0699_ VGND VGND VPWR VPWR net905 sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 gpio_configure\[15\]\[11\] VGND VGND VPWR VPWR net916 sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 _0729_ VGND VGND VPWR VPWR net927 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_131_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1050 _0549_ VGND VGND VPWR VPWR net1583 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1061 gpio_configure\[36\]\[8\] VGND VGND VPWR VPWR net1594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1072 _0730_ VGND VGND VPWR VPWR net1605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1083 gpio_configure\[2\]\[0\] VGND VGND VPWR VPWR net1616 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1094 gpio_configure\[37\]\[0\] VGND VGND VPWR VPWR net1627 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_201 _2490_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_212 gpio_configure\[3\]\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_223 net368 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_234 net459 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_245 _2490_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_256 net471 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_682 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_154_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_96_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_49_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4961_ _2149_ _2170_ VGND VGND VPWR VPWR _2171_ sky130_fd_sc_hd__nor2_1
XFILLER_17_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6700_ clknet_3_7_0_wb_clk_i _0013_ net528 VGND VGND VPWR VPWR wbbd_state\[9\] sky130_fd_sc_hd__dfrtp_4
X_3912_ net2067 _0816_ hkspi.state\[0\] _1384_ net2083 VGND VGND VPWR VPWR _0005_
+ sky130_fd_sc_hd__a41o_1
X_4892_ _1666_ _2082_ _2088_ _2089_ _2102_ VGND VGND VPWR VPWR _2103_ sky130_fd_sc_hd__a2111o_1
XFILLER_189_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6631_ clknet_3_5_0_wb_clk_i _0244_ VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__dfxtp_1
X_3843_ _1378_ _1385_ _1412_ hkspi.state\[0\] VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__a211oi_1
XFILLER_149_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3774_ gpio_configure\[0\]\[8\] _1087_ _1127_ gpio_configure\[33\]\[8\] _1359_ VGND
+ VGND VPWR VPWR _1360_ sky130_fd_sc_hd__a221o_1
X_6562_ clknet_3_2_0_wb_clk_i _0014_ net499 VGND VGND VPWR VPWR xfer_state\[0\] sky130_fd_sc_hd__dfstp_1
XFILLER_164_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5513_ net464 net1336 _2433_ VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__mux2_1
X_6493_ clknet_leaf_73_csclk net1060 net488 VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__dfstp_1
XFILLER_145_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5444_ net447 net1240 _2425_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__mux2_1
XFILLER_133_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5375_ net435 net1047 _2417_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__mux2_1
X_7114_ clknet_leaf_33_csclk net1109 net525 VGND VGND VPWR VPWR gpio_configure\[34\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_4326_ net834 net463 _1546_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__mux2_1
XFILLER_59_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_99_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_141_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4257_ net1220 net444 _1534_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__mux2_1
X_7045_ clknet_leaf_31_csclk net1026 net523 VGND VGND VPWR VPWR gpio_configure\[25\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_101_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3208_ gpio_configure\[26\]\[3\] VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__inv_2
XFILLER_170_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4188_ net2011 _0969_ _1519_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__mux2_1
XFILLER_67_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_103_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6829_ clknet_leaf_29_csclk net985 net524 VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__dfrtp_1
XFILLER_168_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_183_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_105_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold180 _0197_ VGND VGND VPWR VPWR net713 sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 serial_bb_clock VGND VGND VPWR VPWR net724 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_93_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_19_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_747 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_92_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3490_ net628 _1008_ VGND VGND VPWR VPWR _1081_ sky130_fd_sc_hd__nor2_4
XFILLER_6_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_5_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_170_688 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5160_ _2277_ _2334_ _2366_ VGND VGND VPWR VPWR _2367_ sky130_fd_sc_hd__or3_1
XFILLER_69_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4111_ net629 _0903_ net483 net546 VGND VGND VPWR VPWR _1509_ sky130_fd_sc_hd__or4_4
X_5091_ _1652_ _1941_ _2195_ _1835_ _1847_ VGND VGND VPWR VPWR _2300_ sky130_fd_sc_hd__a2111o_1
XFILLER_96_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4042_ net462 net1491 _1478_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__mux2_1
XFILLER_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5993_ gpio_configure\[32\]\[0\] net416 _2814_ gpio_configure\[11\]\[0\] _2812_ VGND
+ VGND VPWR VPWR _2815_ sky130_fd_sc_hd__a221o_1
XFILLER_52_558 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_40_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4944_ _1568_ _1640_ VGND VGND VPWR VPWR _2154_ sky130_fd_sc_hd__or2_1
XFILLER_178_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4875_ _1746_ _1957_ VGND VGND VPWR VPWR _2086_ sky130_fd_sc_hd__or2_1
X_6614_ clknet_leaf_3_csclk net1293 net494 VGND VGND VPWR VPWR gpio_configure\[3\]\[11\]
+ sky130_fd_sc_hd__dfstp_2
X_3826_ hkspi.addr\[1\] hkspi.addr\[0\] hkspi.addr\[2\] VGND VGND VPWR VPWR _1403_
+ sky130_fd_sc_hd__a21o_1
XFILLER_20_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_193_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_165_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6545_ clknet_2_0__leaf_mgmt_gpio_in[4] _0008_ _0056_ VGND VGND VPWR VPWR hkspi.state\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_3757_ net43 net356 _1136_ net301 _1326_ VGND VGND VPWR VPWR _1343_ sky130_fd_sc_hd__a221o_2
XFILLER_173_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6476_ clknet_leaf_71_csclk net1641 net490 VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__dfstp_1
X_3688_ _1269_ _1271_ _1273_ _1275_ VGND VGND VPWR VPWR _1276_ sky130_fd_sc_hd__or4_1
X_5427_ net660 net687 _2423_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__mux2_1
Xoutput230 net230 VGND VGND VPWR VPWR mgmt_gpio_out[25] sky130_fd_sc_hd__buf_12
Xoutput241 net241 VGND VGND VPWR VPWR mgmt_gpio_out[35] sky130_fd_sc_hd__buf_12
XFILLER_133_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_161_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput252 net252 VGND VGND VPWR VPWR pad_flash_clk_oeb sky130_fd_sc_hd__buf_12
XFILLER_160_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput263 net263 VGND VGND VPWR VPWR pll90_sel[2] sky130_fd_sc_hd__buf_12
Xoutput274 net274 VGND VGND VPWR VPWR pll_sel[2] sky130_fd_sc_hd__buf_12
Xoutput285 net285 VGND VGND VPWR VPWR pll_trim[19] sky130_fd_sc_hd__buf_12
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5358_ _0921_ net429 VGND VGND VPWR VPWR _2416_ sky130_fd_sc_hd__nand2_8
Xoutput296 net296 VGND VGND VPWR VPWR pll_trim[5] sky130_fd_sc_hd__buf_12
XFILLER_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4309_ net455 net1761 _1543_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__mux2_1
XFILLER_87_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5289_ net458 net1658 net565 VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__mux2_1
XFILLER_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_7028_ clknet_leaf_64_csclk net839 net501 VGND VGND VPWR VPWR gpio_configure\[23\]\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_28_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7159__531 VGND VGND VPWR VPWR net531 _7159__531/LO sky130_fd_sc_hd__conb_1
XFILLER_75_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_31_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire357 _0876_ VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__buf_8
XFILLER_136_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_132 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_155_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_78_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout490 net491 VGND VGND VPWR VPWR net490 sky130_fd_sc_hd__buf_6
XFILLER_48_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_83 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_74_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4660_ _1588_ _1684_ VGND VGND VPWR VPWR _1872_ sky130_fd_sc_hd__and2_2
XFILLER_30_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3611_ gpio_configure\[10\]\[2\] _0920_ _1056_ gpio_configure\[12\]\[10\] VGND VGND
+ VPWR VPWR _1200_ sky130_fd_sc_hd__a22o_1
XFILLER_175_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4591_ net126 net125 _1755_ VGND VGND VPWR VPWR _1803_ sky130_fd_sc_hd__or3_4
XFILLER_190_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6330_ gpio_configure\[23\]\[12\] _2822_ _2843_ gpio_configure\[5\]\[12\] _3139_
+ VGND VGND VPWR VPWR _3140_ sky130_fd_sc_hd__a221o_1
XFILLER_162_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3542_ _1090_ _1106_ _1115_ _1132_ VGND VGND VPWR VPWR _1133_ sky130_fd_sc_hd__or4_2
Xhold905 _0542_ VGND VGND VPWR VPWR net1438 sky130_fd_sc_hd__dlygate4sd3_1
Xhold916 net289 VGND VGND VPWR VPWR net1449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold927 _0683_ VGND VGND VPWR VPWR net1460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold938 gpio_configure\[20\]\[6\] VGND VGND VPWR VPWR net1471 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_142_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3473_ gpio_configure\[21\]\[12\] _1062_ _1063_ _0972_ VGND VGND VPWR VPWR _1064_
+ sky130_fd_sc_hd__a211o_1
X_6261_ gpio_configure\[10\]\[9\] net414 _2840_ gpio_configure\[6\]\[9\] _3073_ VGND
+ VGND VPWR VPWR _3074_ sky130_fd_sc_hd__a221o_1
Xhold949 _0355_ VGND VGND VPWR VPWR net1482 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_89_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5212_ net390 _0870_ net467 VGND VGND VPWR VPWR _2396_ sky130_fd_sc_hd__or3_1
X_6192_ _3001_ _3003_ _3005_ _3007_ VGND VGND VPWR VPWR _3008_ sky130_fd_sc_hd__or4_1
XFILLER_123_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5143_ _1782_ _1822_ _2006_ _1706_ VGND VGND VPWR VPWR _2350_ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_96_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1605 gpio_configure\[34\]\[2\] VGND VGND VPWR VPWR net2138 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5074_ _1592_ _1808_ _1876_ VGND VGND VPWR VPWR _2283_ sky130_fd_sc_hd__o21a_1
XFILLER_57_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4025_ net1636 net455 _1475_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__mux2_1
XFILLER_71_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5976_ _2794_ _2797_ VGND VGND VPWR VPWR _2798_ sky130_fd_sc_hd__nor2_1
XFILLER_52_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4927_ _2110_ _2136_ _1862_ VGND VGND VPWR VPWR _2138_ sky130_fd_sc_hd__o21a_1
XFILLER_33_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4858_ _1636_ _1671_ _1906_ _2068_ VGND VGND VPWR VPWR _2069_ sky130_fd_sc_hd__o211a_1
XFILLER_21_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3809_ hkspi.addr\[6\] hkspi.addr\[5\] hkspi.addr\[4\] _1390_ VGND VGND VPWR VPWR
+ _1391_ sky130_fd_sc_hd__nand4_1
XFILLER_165_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4789_ _1665_ _1745_ net424 _1805_ VGND VGND VPWR VPWR _2000_ sky130_fd_sc_hd__o22ai_1
XFILLER_4_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6528_ clknet_leaf_76_csclk net1639 net484 VGND VGND VPWR VPWR gpio_configure\[25\]\[10\]
+ sky130_fd_sc_hd__dfstp_2
XFILLER_180_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_118_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6459_ clknet_2_1__leaf_mgmt_gpio_in[4] net2098 _0037_ VGND VGND VPWR VPWR hkspi.pass_thru_mgmt
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_106_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_85_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_18_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_43_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_71_653 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_713 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_12_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_757 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_156_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_753 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_59_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_62_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5830_ gpio_configure\[28\]\[6\] _2513_ _2538_ gpio_configure\[1\]\[6\] _2658_ VGND
+ VGND VPWR VPWR _2659_ sky130_fd_sc_hd__a221o_1
XFILLER_61_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5761_ gpio_configure\[19\]\[3\] _2491_ _2506_ gpio_configure\[27\]\[3\] VGND VGND
+ VPWR VPWR _2593_ sky130_fd_sc_hd__a22o_1
X_4712_ _1590_ _1782_ _1797_ VGND VGND VPWR VPWR _1924_ sky130_fd_sc_hd__or3_1
X_5692_ gpio_configure\[2\]\[0\] _2523_ _2524_ gpio_configure\[16\]\[0\] _2525_ VGND
+ VGND VPWR VPWR _2527_ sky130_fd_sc_hd__a221o_1
XFILLER_187_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4643_ _1774_ _1823_ _1854_ _1700_ _1699_ VGND VGND VPWR VPWR _1855_ sky130_fd_sc_hd__o2111a_1
XFILLER_162_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap410 _2837_ VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__buf_12
X_4574_ _1750_ _1769_ _1785_ VGND VGND VPWR VPWR _1786_ sky130_fd_sc_hd__nor3_1
Xhold702 _0657_ VGND VGND VPWR VPWR net1235 sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 gpio_configure\[21\]\[12\] VGND VGND VPWR VPWR net1246 sky130_fd_sc_hd__dlygate4sd3_1
Xmax_cap421 _2507_ VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__buf_12
XFILLER_162_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold724 _0604_ VGND VGND VPWR VPWR net1257 sky130_fd_sc_hd__dlygate4sd3_1
X_6313_ gpio_configure\[2\]\[11\] net398 _2843_ gpio_configure\[5\]\[11\] _3123_ VGND
+ VGND VPWR VPWR _3124_ sky130_fd_sc_hd__a221o_1
XFILLER_115_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3525_ net639 _1008_ VGND VGND VPWR VPWR _1116_ sky130_fd_sc_hd__nor2_4
Xhold735 gpio_configure\[18\]\[4\] VGND VGND VPWR VPWR net1268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 _0636_ VGND VGND VPWR VPWR net1279 sky130_fd_sc_hd__dlygate4sd3_1
Xhold757 gpio_configure\[29\]\[7\] VGND VGND VPWR VPWR net1290 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_115_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_143_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold768 _0358_ VGND VGND VPWR VPWR net1301 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold779 gpio_configure\[20\]\[7\] VGND VGND VPWR VPWR net1312 sky130_fd_sc_hd__dlygate4sd3_1
X_6244_ serial_data_staging_2\[7\] _2444_ _2485_ VGND VGND VPWR VPWR _3058_ sky130_fd_sc_hd__o21ba_1
XFILLER_89_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3456_ net384 _1008_ VGND VGND VPWR VPWR _1047_ sky130_fd_sc_hd__nor2_4
XFILLER_130_102 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_115_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3387_ gpio_configure\[18\]\[6\] net374 net369 gpio_configure\[25\]\[6\] VGND VGND
+ VPWR VPWR _0981_ sky130_fd_sc_hd__a22o_1
X_6175_ gpio_configure\[18\]\[6\] net399 _2839_ gpio_configure\[35\]\[6\] _2990_ VGND
+ VGND VPWR VPWR _2991_ sky130_fd_sc_hd__a221o_2
XFILLER_97_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_69_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1402 net326 VGND VGND VPWR VPWR net1935 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1413 net348 VGND VGND VPWR VPWR net1946 sky130_fd_sc_hd__dlygate4sd3_1
X_5126_ _1673_ _2041_ _2151_ _2155_ VGND VGND VPWR VPWR _2334_ sky130_fd_sc_hd__or4b_1
Xhold1424 net343 VGND VGND VPWR VPWR net1957 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_97_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1435 net281 VGND VGND VPWR VPWR net1968 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1446 gpio_configure\[12\]\[0\] VGND VGND VPWR VPWR net1979 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1457 _0114_ VGND VGND VPWR VPWR net1990 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1468 hkspi.ldata\[5\] VGND VGND VPWR VPWR net2001 sky130_fd_sc_hd__dlygate4sd3_1
X_5057_ _1605_ _1684_ _1800_ _2265_ _1630_ VGND VGND VPWR VPWR _2266_ sky130_fd_sc_hd__o311a_1
Xhold1479 net331 VGND VGND VPWR VPWR net2012 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_55_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4008_ net437 net1453 _1472_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__mux2_1
XTAP_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5959_ gpio_configure\[4\]\[12\] _2502_ _2518_ gpio_configure\[3\]\[12\] _2781_ VGND
+ VGND VPWR VPWR _2782_ sky130_fd_sc_hd__a221o_1
XFILLER_139_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_139_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_4_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold40 net436 VGND VGND VPWR VPWR net573 sky130_fd_sc_hd__buf_6
Xhold51 _1525_ VGND VGND VPWR VPWR net584 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold62 _1464_ VGND VGND VPWR VPWR net595 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 _0853_ VGND VGND VPWR VPWR net606 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 _1466_ VGND VGND VPWR VPWR net617 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 _0867_ VGND VGND VPWR VPWR net628 sky130_fd_sc_hd__buf_8
XFILLER_152_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_686 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_16_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_157_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_4 _0892_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3310_ net601 net381 VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__nor2_8
XFILLER_98_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4290_ net465 net860 _1540_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__mux2_1
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3241_ hkspi.count\[2\] hkspi.count\[1\] hkspi.count\[0\] VGND VGND VPWR VPWR _0837_
+ sky130_fd_sc_hd__or3_4
XFILLER_98_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_140_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_39_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6931_ clknet_3_6_0_csclk net1669 net517 VGND VGND VPWR VPWR gpio_configure\[11\]\[1\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6862_ clknet_leaf_15_csclk net1195 net513 VGND VGND VPWR VPWR gpio_configure\[2\]\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_34_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_179_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5813_ _2636_ _2638_ _2640_ _2642_ VGND VGND VPWR VPWR _2643_ sky130_fd_sc_hd__or4_1
XFILLER_179_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6793_ clknet_leaf_77_csclk net1745 net484 VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__dfrtp_4
XFILLER_50_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5744_ gpio_configure\[26\]\[2\] _2534_ _2576_ net419 VGND VGND VPWR VPWR _2577_
+ sky130_fd_sc_hd__a22o_1
XFILLER_148_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5675_ net472 _2461_ _2493_ VGND VGND VPWR VPWR _2510_ sky130_fd_sc_hd__and3_4
Xclkbuf_leaf_72_csclk clknet_3_0_0_csclk VGND VGND VPWR VPWR clknet_leaf_72_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_108_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4626_ _1837_ VGND VGND VPWR VPWR _1838_ sky130_fd_sc_hd__inv_2
XFILLER_135_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold510 gpio_configure\[1\]\[7\] VGND VGND VPWR VPWR net1043 sky130_fd_sc_hd__dlygate4sd3_1
Xhold521 _0532_ VGND VGND VPWR VPWR net1054 sky130_fd_sc_hd__dlygate4sd3_1
X_4557_ net126 _1762_ _1766_ VGND VGND VPWR VPWR _1769_ sky130_fd_sc_hd__or3_2
Xhold532 gpio_configure\[5\]\[5\] VGND VGND VPWR VPWR net1065 sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 _0656_ VGND VGND VPWR VPWR net1076 sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 gpio_configure\[6\]\[7\] VGND VGND VPWR VPWR net1087 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_116_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3508_ net278 _0940_ _1098_ gpio_configure\[25\]\[12\] VGND VGND VPWR VPWR _1099_
+ sky130_fd_sc_hd__a22o_2
XFILLER_1_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold565 _1462_ VGND VGND VPWR VPWR net1098 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_103_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4488_ _1598_ _1686_ VGND VGND VPWR VPWR _1700_ sky130_fd_sc_hd__nand2_2
Xhold576 _0717_ VGND VGND VPWR VPWR net1109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold587 gpio_configure\[10\]\[5\] VGND VGND VPWR VPWR net1120 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_143_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold598 _0552_ VGND VGND VPWR VPWR net1131 sky130_fd_sc_hd__dlygate4sd3_1
X_6227_ gpio_configure\[23\]\[8\] _2822_ _2828_ gpio_configure\[20\]\[8\] _3036_ VGND
+ VGND VPWR VPWR _3041_ sky130_fd_sc_hd__a221o_1
XFILLER_104_669 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3439_ net8 _0891_ _0936_ net25 VGND VGND VPWR VPWR _1031_ sky130_fd_sc_hd__a22o_2
XFILLER_58_701 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6158_ gpio_configure\[34\]\[5\] net393 _2852_ gpio_configure\[19\]\[5\] _2974_ VGND
+ VGND VPWR VPWR _2975_ sky130_fd_sc_hd__a221o_1
Xhold1210 _0187_ VGND VGND VPWR VPWR net1743 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1221 _0344_ VGND VGND VPWR VPWR net1754 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_10_csclk clknet_3_4_0_csclk VGND VGND VPWR VPWR clknet_leaf_10_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_85_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold1232 gpio_configure\[14\]\[0\] VGND VGND VPWR VPWR net1765 sky130_fd_sc_hd__dlygate4sd3_1
X_5109_ _2128_ _2237_ _2290_ _2316_ VGND VGND VPWR VPWR _2317_ sky130_fd_sc_hd__or4_1
Xhold1243 _0485_ VGND VGND VPWR VPWR net1776 sky130_fd_sc_hd__dlygate4sd3_1
X_6089_ gpio_configure\[21\]\[2\] _2820_ _2830_ gpio_configure\[3\]\[2\] _2908_ VGND
+ VGND VPWR VPWR _2909_ sky130_fd_sc_hd__a221o_1
Xhold1254 gpio_configure\[5\]\[8\] VGND VGND VPWR VPWR net1787 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1265 gpio_configure\[30\]\[0\] VGND VGND VPWR VPWR net1798 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1276 _0143_ VGND VGND VPWR VPWR net1809 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1287 net282 VGND VGND VPWR VPWR net1820 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1298 _0128_ VGND VGND VPWR VPWR net1831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_122_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_csclk clknet_3_5_0_csclk VGND VGND VPWR VPWR clknet_leaf_25_csclk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_53_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_13_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_107_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput130 wb_adr_i[9] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_1
Xinput141 wb_dat_i[18] VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_1
XFILLER_88_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput152 wb_dat_i[28] VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_1
Xinput163 wb_dat_i[9] VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_1
XFILLER_48_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_737 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_63_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_56_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_177_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_176_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_32_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3790_ _1335_ _1341_ _1351_ _1375_ VGND VGND VPWR VPWR _1376_ sky130_fd_sc_hd__or4_4
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_185_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5460_ net457 net838 _2427_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__mux2_1
XFILLER_8_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_145_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4411_ _1617_ _1622_ VGND VGND VPWR VPWR _1623_ sky130_fd_sc_hd__nand2_1
X_5391_ net440 net1534 _2419_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__mux2_1
XFILLER_99_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_7130_ clknet_leaf_27_csclk net1225 net521 VGND VGND VPWR VPWR gpio_configure\[36\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_4342_ net127 net126 net125 VGND VGND VPWR VPWR _1554_ sky130_fd_sc_hd__and3_2
XFILLER_98_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_7061_ clknet_leaf_29_csclk net969 net521 VGND VGND VPWR VPWR gpio_configure\[27\]\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_4273_ net754 net577 _1537_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__mux2_1
XFILLER_101_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6012_ _2815_ _2821_ _2827_ _2833_ VGND VGND VPWR VPWR _2834_ sky130_fd_sc_hd__or4_1
X_3224_ gpio_configure\[10\]\[3\] VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__inv_2
.ends

