module caravan_logo ();
endmodule
