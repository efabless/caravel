magic
tech sky130A
magscale 1 2
timestamp 1636751500
<< metal4 >>
tri 8320 10560 8640 10880 se
rect 8640 10560 8960 10880
rect 6720 8320 8000 8640
rect 6400 5760 8000 8320
tri 3200 5120 3840 5760 se
rect 3840 5440 5440 5760
tri 5440 5440 5760 5760 sw
tri 7040 5440 7360 5760 ne
rect 7360 5440 8000 5760
rect 8320 7040 8640 10560
tri 8640 10240 8960 10560 nw
rect 10880 9600 36160 10240
rect 8960 7360 9600 8640
rect 3840 5120 6720 5440
rect 3200 4800 6720 5120
tri 6720 4800 7360 5440 sw
rect 8320 5120 8960 7040
rect 10880 6720 13760 8960
rect 14080 6720 31040 8960
rect 31360 6720 36160 8960
rect 10880 5760 36160 6400
rect 13120 5440 14080 5760
tri 9600 4800 10240 5440 se
rect 10240 4800 16000 5440
rect 17600 5120 36160 5760
rect 3200 4160 16000 4800
rect 3200 3520 4160 4160
rect 7680 3840 9920 4160
rect 32000 3840 35840 5120
<< metal5 >>
tri 8000 9920 8320 10240 se
rect 8320 9920 9920 10240
tri 9920 9920 10240 10240 sw
tri 6080 9600 6400 9920 se
tri 6080 9280 6400 9600 ne
rect 6400 8640 10240 9920
tri 6080 8320 6400 8640 se
rect 6400 8320 6720 8640
tri 5760 7360 6080 7680 se
rect 6080 7360 6400 8320
tri 6400 8000 6720 8320 nw
rect 8000 7360 8960 8640
rect 9600 7360 10240 8640
tri 4480 7040 4800 7360 se
rect 4800 7040 10240 7360
tri 3200 6720 3520 7040 se
rect 3520 6720 10240 7040
rect 3200 5440 10240 6720
rect 10880 8960 36160 10240
rect 10880 6720 14400 8960
rect 15680 8640 16320 8960
rect 17600 8640 18240 8960
rect 14720 8000 16320 8640
rect 16640 8000 18240 8640
tri 18240 8320 18880 8960 nw
tri 18880 8320 19200 8640 se
tri 19200 8320 19520 8640 sw
tri 19520 8320 20160 8960 ne
rect 15680 7680 16320 8000
rect 17600 7680 18240 8000
tri 18560 8000 18880 8320 se
rect 18880 8000 19520 8320
tri 19520 8000 19840 8320 sw
rect 18560 7680 19840 8000
rect 14720 7040 16320 7680
rect 15680 6720 16320 7040
rect 16640 6720 18240 7680
rect 18560 6720 19840 7360
rect 20160 6720 20800 8960
tri 22080 8640 22400 8960 ne
rect 21120 8000 21760 8640
tri 21760 8320 22080 8640 sw
tri 21760 8000 22080 8320 nw
tri 22240 7840 22400 8000 se
tri 22240 7680 22400 7840 ne
rect 21120 7040 21760 7680
tri 21760 7360 22080 7680 sw
tri 21760 7040 22080 7360 nw
tri 22080 6720 22400 7040 se
rect 22400 6720 23040 8960
rect 23360 7040 24960 8960
rect 26240 8640 26880 8960
tri 26880 8640 27200 8960 nw
rect 28480 8640 29120 8960
tri 29120 8640 29440 8960 nw
rect 30720 8640 36160 8960
rect 25280 8000 26880 8640
tri 27200 8320 27520 8640 se
tri 27200 8000 27520 8320 ne
rect 27520 8000 29120 8640
tri 29440 8320 29760 8640 se
tri 29440 8000 29760 8320 ne
rect 29760 8000 36160 8640
rect 26240 7680 26880 8000
tri 26880 7680 27200 8000 sw
tri 28160 7680 28480 8000 ne
rect 28480 7680 29120 8000
tri 29120 7680 29440 8000 sw
tri 30400 7680 30720 8000 ne
rect 25280 7040 27840 7680
tri 27840 7360 28160 7680 sw
tri 27840 7040 28160 7360 nw
rect 28480 7040 30080 7680
tri 30080 7360 30400 7680 sw
tri 30080 7040 30400 7360 nw
rect 24320 6720 24960 7040
rect 26240 6720 26880 7040
tri 28160 6720 28480 7040 se
rect 28480 6720 29120 7040
tri 30400 6720 30720 7040 se
rect 30720 6720 36160 8000
rect 10880 5760 36160 6720
rect 13120 5440 14080 5760
tri 17280 5440 17600 5760 ne
rect 3200 5120 16320 5440
rect 17600 5149 36160 5760
rect 17600 5120 36182 5149
tri 2880 4800 3200 5120 se
rect 3200 4800 4160 5120
tri 4160 4800 4480 5120 nw
tri 6080 4800 6400 5120 ne
rect 2880 3840 4160 4800
tri 2880 3520 3200 3840 ne
rect 3200 3520 4160 3840
tri 4482 4340 4882 4740 se
rect 4882 4342 5682 4740
tri 5682 4342 6080 4740 sw
rect 4882 4340 6080 4342
rect 4482 3540 6080 4340
rect 6400 3840 11520 5120
tri 11520 4800 11840 5120 nw
tri 13440 4800 13760 5120 ne
tri 13760 4800 14080 5120 nw
tri 15360 4800 15680 5120 ne
rect 15680 4800 16320 5120
rect 17920 4800 23360 5120
rect 31230 4800 31870 5120
tri 31870 4800 32190 5120 nw
tri 33280 4800 33600 5120 ne
rect 33600 4800 33920 5120
tri 33920 4800 34240 5120 nw
tri 35390 4800 35710 5120 ne
rect 35710 4800 36182 5120
tri 11992 4340 12392 4740 se
rect 12392 4340 13192 4740
tri 13192 4340 13592 4740 sw
tri 4482 3140 4882 3540 ne
rect 4882 3538 6080 3540
rect 4882 3140 5682 3538
tri 5682 3140 6080 3538 nw
rect 11992 3540 13592 4340
tri 11992 3140 12392 3540 ne
rect 12392 3140 13192 3540
tri 13192 3140 13592 3540 nw
tri 13992 4340 14392 4740 se
rect 14392 4340 15192 4740
tri 15192 4340 15592 4740 sw
rect 13992 3540 15592 4340
rect 17920 4160 18240 4800
tri 31992 4340 32392 4740 se
rect 32392 4340 33192 4740
tri 33192 4340 33592 4740 sw
rect 17600 3840 18560 4160
tri 13992 3140 14392 3540 ne
rect 14392 3140 15192 3540
tri 15192 3140 15592 3540 nw
rect 31992 3540 33592 4340
tri 31992 3140 32392 3540 ne
rect 32392 3140 33192 3540
tri 33192 3140 33592 3540 nw
tri 33922 4340 34322 4740 se
rect 34322 4340 35122 4740
tri 35122 4340 35522 4740 sw
rect 33922 3540 35522 4340
rect 35860 4480 36182 4800
rect 35860 3840 36480 4480
tri 33922 3140 34322 3540 ne
rect 34322 3140 35122 3540
tri 35122 3140 35522 3540 nw
<< fillblock >>
rect 2240 2560 37000 11520
<< end >>
