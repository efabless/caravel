magic
tech sky130A
magscale 1 2
timestamp 1649097268
<< obsli1 >>
rect 1104 17 218868 31943
<< obsm1 >>
rect 65260 32000 106412 32008
rect 106 8 219774 32000
<< metal2 >>
rect 202 31200 258 32400
rect 570 31200 626 32400
rect 1030 31200 1086 32400
rect 1490 31200 1546 32400
rect 1950 31200 2006 32400
rect 2410 31200 2466 32400
rect 2870 31200 2926 32400
rect 3238 31200 3294 32400
rect 3698 31200 3754 32400
rect 4158 31200 4214 32400
rect 4618 31200 4674 32400
rect 5078 31200 5134 32400
rect 5538 31200 5594 32400
rect 5906 31200 5962 32400
rect 6366 31200 6422 32400
rect 6826 31200 6882 32400
rect 7286 31200 7342 32400
rect 7746 31200 7802 32400
rect 8206 31200 8262 32400
rect 8574 31200 8630 32400
rect 9034 31200 9090 32400
rect 9494 31200 9550 32400
rect 9954 31200 10010 32400
rect 10414 31200 10470 32400
rect 10874 31200 10930 32400
rect 11334 31200 11390 32400
rect 11702 31200 11758 32400
rect 12162 31200 12218 32400
rect 12622 31200 12678 32400
rect 13082 31200 13138 32400
rect 13542 31200 13598 32400
rect 14002 31200 14058 32400
rect 14370 31200 14426 32400
rect 14830 31200 14886 32400
rect 15290 31200 15346 32400
rect 15750 31200 15806 32400
rect 16210 31200 16266 32400
rect 16670 31200 16726 32400
rect 17038 31200 17094 32400
rect 17498 31200 17554 32400
rect 17958 31200 18014 32400
rect 18418 31200 18474 32400
rect 18878 31200 18934 32400
rect 19338 31200 19394 32400
rect 19706 31200 19762 32400
rect 20166 31200 20222 32400
rect 20626 31200 20682 32400
rect 21086 31200 21142 32400
rect 21546 31200 21602 32400
rect 22006 31200 22062 32400
rect 22466 31200 22522 32400
rect 22834 31200 22890 32400
rect 23294 31200 23350 32400
rect 23754 31200 23810 32400
rect 24214 31200 24270 32400
rect 24674 31200 24730 32400
rect 25134 31200 25190 32400
rect 25502 31200 25558 32400
rect 25962 31200 26018 32400
rect 26422 31200 26478 32400
rect 26882 31200 26938 32400
rect 27342 31200 27398 32400
rect 27802 31200 27858 32400
rect 28170 31200 28226 32400
rect 28630 31200 28686 32400
rect 29090 31200 29146 32400
rect 29550 31200 29606 32400
rect 30010 31200 30066 32400
rect 30470 31200 30526 32400
rect 30838 31200 30894 32400
rect 31298 31200 31354 32400
rect 31758 31200 31814 32400
rect 32218 31200 32274 32400
rect 32678 31200 32734 32400
rect 33138 31200 33194 32400
rect 33598 31200 33654 32400
rect 33966 31200 34022 32400
rect 34426 31200 34482 32400
rect 34886 31200 34942 32400
rect 35346 31200 35402 32400
rect 35806 31200 35862 32400
rect 36266 31200 36322 32400
rect 36634 31200 36690 32400
rect 37094 31200 37150 32400
rect 37554 31200 37610 32400
rect 38014 31200 38070 32400
rect 38474 31200 38530 32400
rect 38934 31200 38990 32400
rect 39302 31200 39358 32400
rect 39762 31200 39818 32400
rect 40222 31200 40278 32400
rect 40682 31200 40738 32400
rect 41142 31200 41198 32400
rect 41602 31200 41658 32400
rect 41970 31200 42026 32400
rect 42430 31200 42486 32400
rect 42890 31200 42946 32400
rect 43350 31200 43406 32400
rect 43810 31200 43866 32400
rect 44270 31200 44326 32400
rect 44730 31200 44786 32400
rect 45098 31200 45154 32400
rect 45558 31200 45614 32400
rect 46018 31200 46074 32400
rect 46478 31200 46534 32400
rect 46938 31200 46994 32400
rect 47398 31200 47454 32400
rect 47766 31200 47822 32400
rect 48226 31200 48282 32400
rect 48686 31200 48742 32400
rect 49146 31200 49202 32400
rect 49606 31200 49662 32400
rect 50066 31200 50122 32400
rect 50434 31200 50490 32400
rect 50894 31200 50950 32400
rect 51354 31200 51410 32400
rect 51814 31200 51870 32400
rect 52274 31200 52330 32400
rect 52734 31200 52790 32400
rect 53102 31200 53158 32400
rect 53562 31200 53618 32400
rect 54022 31200 54078 32400
rect 54482 31200 54538 32400
rect 54942 31200 54998 32400
rect 55402 31200 55458 32400
rect 55862 31200 55918 32400
rect 56230 31200 56286 32400
rect 56690 31200 56746 32400
rect 57150 31200 57206 32400
rect 57610 31200 57666 32400
rect 58070 31200 58126 32400
rect 58530 31200 58586 32400
rect 58898 31200 58954 32400
rect 59358 31200 59414 32400
rect 59818 31200 59874 32400
rect 60278 31200 60334 32400
rect 60738 31200 60794 32400
rect 61198 31200 61254 32400
rect 61566 31200 61622 32400
rect 62026 31200 62082 32400
rect 62486 31200 62542 32400
rect 62946 31200 63002 32400
rect 63406 31200 63462 32400
rect 63866 31200 63922 32400
rect 64234 31200 64290 32400
rect 64694 31200 64750 32400
rect 65154 31200 65210 32400
rect 65614 31200 65670 32400
rect 66074 31200 66130 32400
rect 66534 31200 66590 32400
rect 66994 31200 67050 32400
rect 67362 31200 67418 32400
rect 67822 31200 67878 32400
rect 68282 31200 68338 32400
rect 68742 31200 68798 32400
rect 69202 31200 69258 32400
rect 69662 31200 69718 32400
rect 70030 31200 70086 32400
rect 70490 31200 70546 32400
rect 70950 31200 71006 32400
rect 71410 31200 71466 32400
rect 71870 31200 71926 32400
rect 72330 31200 72386 32400
rect 72698 31200 72754 32400
rect 73158 31200 73214 32400
rect 73618 31200 73674 32400
rect 74078 31200 74134 32400
rect 74538 31200 74594 32400
rect 74998 31200 75054 32400
rect 75366 31200 75422 32400
rect 75826 31200 75882 32400
rect 76286 31200 76342 32400
rect 76746 31200 76802 32400
rect 77206 31200 77262 32400
rect 77666 31200 77722 32400
rect 78126 31200 78182 32400
rect 78494 31200 78550 32400
rect 78954 31200 79010 32400
rect 79414 31200 79470 32400
rect 79874 31200 79930 32400
rect 80334 31200 80390 32400
rect 80794 31200 80850 32400
rect 81162 31200 81218 32400
rect 81622 31200 81678 32400
rect 82082 31200 82138 32400
rect 82542 31200 82598 32400
rect 83002 31200 83058 32400
rect 83462 31200 83518 32400
rect 83830 31200 83886 32400
rect 84290 31200 84346 32400
rect 84750 31200 84806 32400
rect 85210 31200 85266 32400
rect 85670 31200 85726 32400
rect 86130 31200 86186 32400
rect 86498 31200 86554 32400
rect 86958 31200 87014 32400
rect 87418 31200 87474 32400
rect 87878 31200 87934 32400
rect 88338 31200 88394 32400
rect 88798 31200 88854 32400
rect 89258 31200 89314 32400
rect 89626 31200 89682 32400
rect 90086 31200 90142 32400
rect 90546 31200 90602 32400
rect 91006 31200 91062 32400
rect 91466 31200 91522 32400
rect 91926 31200 91982 32400
rect 92294 31200 92350 32400
rect 92754 31200 92810 32400
rect 93214 31200 93270 32400
rect 93674 31200 93730 32400
rect 94134 31200 94190 32400
rect 94594 31200 94650 32400
rect 94962 31200 95018 32400
rect 95422 31200 95478 32400
rect 95882 31200 95938 32400
rect 96342 31200 96398 32400
rect 96802 31200 96858 32400
rect 97262 31200 97318 32400
rect 97630 31200 97686 32400
rect 98090 31200 98146 32400
rect 98550 31200 98606 32400
rect 99010 31200 99066 32400
rect 99470 31200 99526 32400
rect 99930 31200 99986 32400
rect 100390 31200 100446 32400
rect 100758 31200 100814 32400
rect 101218 31200 101274 32400
rect 101678 31200 101734 32400
rect 102138 31200 102194 32400
rect 102598 31200 102654 32400
rect 103058 31200 103114 32400
rect 103426 31200 103482 32400
rect 103886 31200 103942 32400
rect 104346 31200 104402 32400
rect 104806 31200 104862 32400
rect 105266 31200 105322 32400
rect 105726 31200 105782 32400
rect 106094 31200 106150 32400
rect 106554 31200 106610 32400
rect 107014 31200 107070 32400
rect 107474 31200 107530 32400
rect 107934 31200 107990 32400
rect 108394 31200 108450 32400
rect 108762 31200 108818 32400
rect 109222 31200 109278 32400
rect 109682 31200 109738 32400
rect 110142 31200 110198 32400
rect 110602 31200 110658 32400
rect 111062 31200 111118 32400
rect 111522 31200 111578 32400
rect 111890 31200 111946 32400
rect 112350 31200 112406 32400
rect 112810 31200 112866 32400
rect 113270 31200 113326 32400
rect 113730 31200 113786 32400
rect 114190 31200 114246 32400
rect 114558 31200 114614 32400
rect 115018 31200 115074 32400
rect 115478 31200 115534 32400
rect 115938 31200 115994 32400
rect 116398 31200 116454 32400
rect 116858 31200 116914 32400
rect 117226 31200 117282 32400
rect 117686 31200 117742 32400
rect 118146 31200 118202 32400
rect 118606 31200 118662 32400
rect 119066 31200 119122 32400
rect 119526 31200 119582 32400
rect 119894 31200 119950 32400
rect 120354 31200 120410 32400
rect 120814 31200 120870 32400
rect 121274 31200 121330 32400
rect 121734 31200 121790 32400
rect 122194 31200 122250 32400
rect 122654 31200 122710 32400
rect 123022 31200 123078 32400
rect 123482 31200 123538 32400
rect 123942 31200 123998 32400
rect 124402 31200 124458 32400
rect 124862 31200 124918 32400
rect 125322 31200 125378 32400
rect 125690 31200 125746 32400
rect 126150 31200 126206 32400
rect 126610 31200 126666 32400
rect 127070 31200 127126 32400
rect 127530 31200 127586 32400
rect 127990 31200 128046 32400
rect 128358 31200 128414 32400
rect 128818 31200 128874 32400
rect 129278 31200 129334 32400
rect 129738 31200 129794 32400
rect 130198 31200 130254 32400
rect 130658 31200 130714 32400
rect 131026 31200 131082 32400
rect 131486 31200 131542 32400
rect 131946 31200 132002 32400
rect 132406 31200 132462 32400
rect 132866 31200 132922 32400
rect 133326 31200 133382 32400
rect 133786 31200 133842 32400
rect 134154 31200 134210 32400
rect 134614 31200 134670 32400
rect 135074 31200 135130 32400
rect 135534 31200 135590 32400
rect 135994 31200 136050 32400
rect 136454 31200 136510 32400
rect 136822 31200 136878 32400
rect 137282 31200 137338 32400
rect 137742 31200 137798 32400
rect 138202 31200 138258 32400
rect 138662 31200 138718 32400
rect 139122 31200 139178 32400
rect 139490 31200 139546 32400
rect 139950 31200 140006 32400
rect 140410 31200 140466 32400
rect 140870 31200 140926 32400
rect 141330 31200 141386 32400
rect 141790 31200 141846 32400
rect 142158 31200 142214 32400
rect 142618 31200 142674 32400
rect 143078 31200 143134 32400
rect 143538 31200 143594 32400
rect 143998 31200 144054 32400
rect 144458 31200 144514 32400
rect 144918 31200 144974 32400
rect 145286 31200 145342 32400
rect 145746 31200 145802 32400
rect 146206 31200 146262 32400
rect 146666 31200 146722 32400
rect 147126 31200 147182 32400
rect 147586 31200 147642 32400
rect 147954 31200 148010 32400
rect 148414 31200 148470 32400
rect 148874 31200 148930 32400
rect 149334 31200 149390 32400
rect 149794 31200 149850 32400
rect 150254 31200 150310 32400
rect 150622 31200 150678 32400
rect 151082 31200 151138 32400
rect 151542 31200 151598 32400
rect 152002 31200 152058 32400
rect 152462 31200 152518 32400
rect 152922 31200 152978 32400
rect 153290 31200 153346 32400
rect 153750 31200 153806 32400
rect 154210 31200 154266 32400
rect 154670 31200 154726 32400
rect 155130 31200 155186 32400
rect 155590 31200 155646 32400
rect 156050 31200 156106 32400
rect 156418 31200 156474 32400
rect 156878 31200 156934 32400
rect 157338 31200 157394 32400
rect 157798 31200 157854 32400
rect 158258 31200 158314 32400
rect 158718 31200 158774 32400
rect 159086 31200 159142 32400
rect 159546 31200 159602 32400
rect 160006 31200 160062 32400
rect 160466 31200 160522 32400
rect 160926 31200 160982 32400
rect 161386 31200 161442 32400
rect 161754 31200 161810 32400
rect 162214 31200 162270 32400
rect 162674 31200 162730 32400
rect 163134 31200 163190 32400
rect 163594 31200 163650 32400
rect 164054 31200 164110 32400
rect 164422 31200 164478 32400
rect 164882 31200 164938 32400
rect 165342 31200 165398 32400
rect 165802 31200 165858 32400
rect 166262 31200 166318 32400
rect 166722 31200 166778 32400
rect 167182 31200 167238 32400
rect 167550 31200 167606 32400
rect 168010 31200 168066 32400
rect 168470 31200 168526 32400
rect 168930 31200 168986 32400
rect 169390 31200 169446 32400
rect 169850 31200 169906 32400
rect 170218 31200 170274 32400
rect 170678 31200 170734 32400
rect 171138 31200 171194 32400
rect 171598 31200 171654 32400
rect 172058 31200 172114 32400
rect 172518 31200 172574 32400
rect 172886 31200 172942 32400
rect 173346 31200 173402 32400
rect 173806 31200 173862 32400
rect 174266 31200 174322 32400
rect 174726 31200 174782 32400
rect 175186 31200 175242 32400
rect 175554 31200 175610 32400
rect 176014 31200 176070 32400
rect 176474 31200 176530 32400
rect 176934 31200 176990 32400
rect 177394 31200 177450 32400
rect 177854 31200 177910 32400
rect 178314 31200 178370 32400
rect 178682 31200 178738 32400
rect 179142 31200 179198 32400
rect 179602 31200 179658 32400
rect 180062 31200 180118 32400
rect 180522 31200 180578 32400
rect 180982 31200 181038 32400
rect 181350 31200 181406 32400
rect 181810 31200 181866 32400
rect 182270 31200 182326 32400
rect 182730 31200 182786 32400
rect 183190 31200 183246 32400
rect 183650 31200 183706 32400
rect 184018 31200 184074 32400
rect 184478 31200 184534 32400
rect 184938 31200 184994 32400
rect 185398 31200 185454 32400
rect 185858 31200 185914 32400
rect 186318 31200 186374 32400
rect 186686 31200 186742 32400
rect 187146 31200 187202 32400
rect 187606 31200 187662 32400
rect 188066 31200 188122 32400
rect 188526 31200 188582 32400
rect 188986 31200 189042 32400
rect 189446 31200 189502 32400
rect 189814 31200 189870 32400
rect 190274 31200 190330 32400
rect 190734 31200 190790 32400
rect 191194 31200 191250 32400
rect 191654 31200 191710 32400
rect 192114 31200 192170 32400
rect 192482 31200 192538 32400
rect 192942 31200 192998 32400
rect 193402 31200 193458 32400
rect 193862 31200 193918 32400
rect 194322 31200 194378 32400
rect 194782 31200 194838 32400
rect 195150 31200 195206 32400
rect 195610 31200 195666 32400
rect 196070 31200 196126 32400
rect 196530 31200 196586 32400
rect 196990 31200 197046 32400
rect 197450 31200 197506 32400
rect 197818 31200 197874 32400
rect 198278 31200 198334 32400
rect 198738 31200 198794 32400
rect 199198 31200 199254 32400
rect 199658 31200 199714 32400
rect 200118 31200 200174 32400
rect 200578 31200 200634 32400
rect 200946 31200 201002 32400
rect 201406 31200 201462 32400
rect 201866 31200 201922 32400
rect 202326 31200 202382 32400
rect 202786 31200 202842 32400
rect 203246 31200 203302 32400
rect 203614 31200 203670 32400
rect 204074 31200 204130 32400
rect 204534 31200 204590 32400
rect 204994 31200 205050 32400
rect 205454 31200 205510 32400
rect 205914 31200 205970 32400
rect 206282 31200 206338 32400
rect 206742 31200 206798 32400
rect 207202 31200 207258 32400
rect 207662 31200 207718 32400
rect 208122 31200 208178 32400
rect 208582 31200 208638 32400
rect 208950 31200 209006 32400
rect 209410 31200 209466 32400
rect 209870 31200 209926 32400
rect 210330 31200 210386 32400
rect 210790 31200 210846 32400
rect 211250 31200 211306 32400
rect 211710 31200 211766 32400
rect 212078 31200 212134 32400
rect 212538 31200 212594 32400
rect 212998 31200 213054 32400
rect 213458 31200 213514 32400
rect 213918 31200 213974 32400
rect 214378 31200 214434 32400
rect 214746 31200 214802 32400
rect 215206 31200 215262 32400
rect 215666 31200 215722 32400
rect 216126 31200 216182 32400
rect 216586 31200 216642 32400
rect 217046 31200 217102 32400
rect 217414 31200 217470 32400
rect 217874 31200 217930 32400
rect 218334 31200 218390 32400
rect 218794 31200 218850 32400
rect 219254 31200 219310 32400
rect 219714 31200 219770 32400
rect 110 -400 166 800
rect 386 -400 442 800
rect 754 -400 810 800
rect 1122 -400 1178 800
rect 1490 -400 1546 800
rect 1858 -400 1914 800
rect 2226 -400 2282 800
rect 2594 -400 2650 800
rect 2962 -400 3018 800
rect 3238 -400 3294 800
rect 3606 -400 3662 800
rect 3974 -400 4030 800
rect 4342 -400 4398 800
rect 4710 -400 4766 800
rect 5078 -400 5134 800
rect 5446 -400 5502 800
rect 5814 -400 5870 800
rect 6090 -400 6146 800
rect 6458 -400 6514 800
rect 6826 -400 6882 800
rect 7194 -400 7250 800
rect 7562 -400 7618 800
rect 7930 -400 7986 800
rect 8298 -400 8354 800
rect 8666 -400 8722 800
rect 8942 -400 8998 800
rect 9310 -400 9366 800
rect 9678 -400 9734 800
rect 10046 -400 10102 800
rect 10414 -400 10470 800
rect 10782 -400 10838 800
rect 11150 -400 11206 800
rect 11518 -400 11574 800
rect 11794 -400 11850 800
rect 12162 -400 12218 800
rect 12530 -400 12586 800
rect 12898 -400 12954 800
rect 13266 -400 13322 800
rect 13634 -400 13690 800
rect 14002 -400 14058 800
rect 14370 -400 14426 800
rect 14646 -400 14702 800
rect 15014 -400 15070 800
rect 15382 -400 15438 800
rect 15750 -400 15806 800
rect 16118 -400 16174 800
rect 16486 -400 16542 800
rect 16854 -400 16910 800
rect 17222 -400 17278 800
rect 17498 -400 17554 800
rect 17866 -400 17922 800
rect 18234 -400 18290 800
rect 18602 -400 18658 800
rect 18970 -400 19026 800
rect 19338 -400 19394 800
rect 19706 -400 19762 800
rect 20074 -400 20130 800
rect 20350 -400 20406 800
rect 20718 -400 20774 800
rect 21086 -400 21142 800
rect 21454 -400 21510 800
rect 21822 -400 21878 800
rect 22190 -400 22246 800
rect 22558 -400 22614 800
rect 22926 -400 22982 800
rect 23202 -400 23258 800
rect 23570 -400 23626 800
rect 23938 -400 23994 800
rect 24306 -400 24362 800
rect 24674 -400 24730 800
rect 25042 -400 25098 800
rect 25410 -400 25466 800
rect 25778 -400 25834 800
rect 26054 -400 26110 800
rect 26422 -400 26478 800
rect 26790 -400 26846 800
rect 27158 -400 27214 800
rect 27526 -400 27582 800
rect 27894 -400 27950 800
rect 28262 -400 28318 800
rect 28630 -400 28686 800
rect 28906 -400 28962 800
rect 29274 -400 29330 800
rect 29642 -400 29698 800
rect 30010 -400 30066 800
rect 30378 -400 30434 800
rect 30746 -400 30802 800
rect 31114 -400 31170 800
rect 31482 -400 31538 800
rect 31758 -400 31814 800
rect 32126 -400 32182 800
rect 32494 -400 32550 800
rect 32862 -400 32918 800
rect 33230 -400 33286 800
rect 33598 -400 33654 800
rect 33966 -400 34022 800
rect 34334 -400 34390 800
rect 34610 -400 34666 800
rect 34978 -400 35034 800
rect 35346 -400 35402 800
rect 35714 -400 35770 800
rect 36082 -400 36138 800
rect 36450 -400 36506 800
rect 36818 -400 36874 800
rect 37186 -400 37242 800
rect 37462 -400 37518 800
rect 37830 -400 37886 800
rect 38198 -400 38254 800
rect 38566 -400 38622 800
rect 38934 -400 38990 800
rect 39302 -400 39358 800
rect 39670 -400 39726 800
rect 40038 -400 40094 800
rect 40314 -400 40370 800
rect 40682 -400 40738 800
rect 41050 -400 41106 800
rect 41418 -400 41474 800
rect 41786 -400 41842 800
rect 42154 -400 42210 800
rect 42522 -400 42578 800
rect 42890 -400 42946 800
rect 43166 -400 43222 800
rect 43534 -400 43590 800
rect 43902 -400 43958 800
rect 44270 -400 44326 800
rect 44638 -400 44694 800
rect 45006 -400 45062 800
rect 45374 -400 45430 800
rect 45742 -400 45798 800
rect 46018 -400 46074 800
rect 46386 -400 46442 800
rect 46754 -400 46810 800
rect 47122 -400 47178 800
rect 47490 -400 47546 800
rect 47858 -400 47914 800
rect 48226 -400 48282 800
rect 48594 -400 48650 800
rect 48870 -400 48926 800
rect 49238 -400 49294 800
rect 49606 -400 49662 800
rect 49974 -400 50030 800
rect 50342 -400 50398 800
rect 50710 -400 50766 800
rect 51078 -400 51134 800
rect 51446 -400 51502 800
rect 51722 -400 51778 800
rect 52090 -400 52146 800
rect 52458 -400 52514 800
rect 52826 -400 52882 800
rect 53194 -400 53250 800
rect 53562 -400 53618 800
rect 53930 -400 53986 800
rect 54298 -400 54354 800
rect 54574 -400 54630 800
rect 54942 -400 54998 800
rect 55310 -400 55366 800
rect 55678 -400 55734 800
rect 56046 -400 56102 800
rect 56414 -400 56470 800
rect 56782 -400 56838 800
rect 57150 -400 57206 800
rect 57426 -400 57482 800
rect 57794 -400 57850 800
rect 58162 -400 58218 800
rect 58530 -400 58586 800
rect 58898 -400 58954 800
rect 59266 -400 59322 800
rect 59634 -400 59690 800
rect 60002 -400 60058 800
rect 60278 -400 60334 800
rect 60646 -400 60702 800
rect 61014 -400 61070 800
rect 61382 -400 61438 800
rect 61750 -400 61806 800
rect 62118 -400 62174 800
rect 62486 -400 62542 800
rect 62854 -400 62910 800
rect 63130 -400 63186 800
rect 63498 -400 63554 800
rect 63866 -400 63922 800
rect 64234 -400 64290 800
rect 64602 -400 64658 800
rect 64970 -400 65026 800
rect 65338 -400 65394 800
rect 65706 -400 65762 800
rect 65982 -400 66038 800
rect 66350 -400 66406 800
rect 66718 -400 66774 800
rect 67086 -400 67142 800
rect 67454 -400 67510 800
rect 67822 -400 67878 800
rect 68190 -400 68246 800
rect 68558 -400 68614 800
rect 68834 -400 68890 800
rect 69202 -400 69258 800
rect 69570 -400 69626 800
rect 69938 -400 69994 800
rect 70306 -400 70362 800
rect 70674 -400 70730 800
rect 71042 -400 71098 800
rect 71410 -400 71466 800
rect 71686 -400 71742 800
rect 72054 -400 72110 800
rect 72422 -400 72478 800
rect 72790 -400 72846 800
rect 73158 -400 73214 800
rect 73526 -400 73582 800
rect 73894 -400 73950 800
rect 74262 -400 74318 800
rect 74538 -400 74594 800
rect 74906 -400 74962 800
rect 75274 -400 75330 800
rect 75642 -400 75698 800
rect 76010 -400 76066 800
rect 76378 -400 76434 800
rect 76746 -400 76802 800
rect 77114 -400 77170 800
rect 77390 -400 77446 800
rect 77758 -400 77814 800
rect 78126 -400 78182 800
rect 78494 -400 78550 800
rect 78862 -400 78918 800
rect 79230 -400 79286 800
rect 79598 -400 79654 800
rect 79966 -400 80022 800
rect 80242 -400 80298 800
rect 80610 -400 80666 800
rect 80978 -400 81034 800
rect 81346 -400 81402 800
rect 81714 -400 81770 800
rect 82082 -400 82138 800
rect 82450 -400 82506 800
rect 82818 -400 82874 800
rect 83094 -400 83150 800
rect 83462 -400 83518 800
rect 83830 -400 83886 800
rect 84198 -400 84254 800
rect 84566 -400 84622 800
rect 84934 -400 84990 800
rect 85302 -400 85358 800
rect 85670 -400 85726 800
rect 85946 -400 86002 800
rect 86314 -400 86370 800
rect 86682 -400 86738 800
rect 87050 -400 87106 800
rect 87418 -400 87474 800
rect 87786 -400 87842 800
rect 88154 -400 88210 800
rect 88522 -400 88578 800
rect 88798 -400 88854 800
rect 89166 -400 89222 800
rect 89534 -400 89590 800
rect 89902 -400 89958 800
rect 90270 -400 90326 800
rect 90638 -400 90694 800
rect 91006 -400 91062 800
rect 91374 -400 91430 800
rect 91650 -400 91706 800
rect 92018 -400 92074 800
rect 92386 -400 92442 800
rect 92754 -400 92810 800
rect 93122 -400 93178 800
rect 93490 -400 93546 800
rect 93858 -400 93914 800
rect 94226 -400 94282 800
rect 94502 -400 94558 800
rect 94870 -400 94926 800
rect 95238 -400 95294 800
rect 95606 -400 95662 800
rect 95974 -400 96030 800
rect 96342 -400 96398 800
rect 96710 -400 96766 800
rect 97078 -400 97134 800
rect 97354 -400 97410 800
rect 97722 -400 97778 800
rect 98090 -400 98146 800
rect 98458 -400 98514 800
rect 98826 -400 98882 800
rect 99194 -400 99250 800
rect 99562 -400 99618 800
rect 99930 -400 99986 800
rect 100206 -400 100262 800
rect 100574 -400 100630 800
rect 100942 -400 100998 800
rect 101310 -400 101366 800
rect 101678 -400 101734 800
rect 102046 -400 102102 800
rect 102414 -400 102470 800
rect 102782 -400 102838 800
rect 103058 -400 103114 800
rect 103426 -400 103482 800
rect 103794 -400 103850 800
rect 104162 -400 104218 800
rect 104530 -400 104586 800
rect 104898 -400 104954 800
rect 105266 -400 105322 800
rect 105634 -400 105690 800
rect 105910 -400 105966 800
rect 106278 -400 106334 800
rect 106646 -400 106702 800
rect 107014 -400 107070 800
rect 107382 -400 107438 800
rect 107750 -400 107806 800
rect 108118 -400 108174 800
rect 108486 -400 108542 800
rect 108762 -400 108818 800
rect 109130 -400 109186 800
rect 109498 -400 109554 800
rect 109866 -400 109922 800
rect 110234 -400 110290 800
rect 110602 -400 110658 800
rect 110970 -400 111026 800
rect 111338 -400 111394 800
rect 111614 -400 111670 800
rect 111982 -400 112038 800
rect 112350 -400 112406 800
rect 112718 -400 112774 800
rect 113086 -400 113142 800
rect 113454 -400 113510 800
rect 113822 -400 113878 800
rect 114190 -400 114246 800
rect 114466 -400 114522 800
rect 114834 -400 114890 800
rect 115202 -400 115258 800
rect 115570 -400 115626 800
rect 115938 -400 115994 800
rect 116306 -400 116362 800
rect 116674 -400 116730 800
rect 117042 -400 117098 800
rect 117318 -400 117374 800
rect 117686 -400 117742 800
rect 118054 -400 118110 800
rect 118422 -400 118478 800
rect 118790 -400 118846 800
rect 119158 -400 119214 800
rect 119526 -400 119582 800
rect 119894 -400 119950 800
rect 120170 -400 120226 800
rect 120538 -400 120594 800
rect 120906 -400 120962 800
rect 121274 -400 121330 800
rect 121642 -400 121698 800
rect 122010 -400 122066 800
rect 122378 -400 122434 800
rect 122746 -400 122802 800
rect 123022 -400 123078 800
rect 123390 -400 123446 800
rect 123758 -400 123814 800
rect 124126 -400 124182 800
rect 124494 -400 124550 800
rect 124862 -400 124918 800
rect 125230 -400 125286 800
rect 125598 -400 125654 800
rect 125874 -400 125930 800
rect 126242 -400 126298 800
rect 126610 -400 126666 800
rect 126978 -400 127034 800
rect 127346 -400 127402 800
rect 127714 -400 127770 800
rect 128082 -400 128138 800
rect 128450 -400 128506 800
rect 128726 -400 128782 800
rect 129094 -400 129150 800
rect 129462 -400 129518 800
rect 129830 -400 129886 800
rect 130198 -400 130254 800
rect 130566 -400 130622 800
rect 130934 -400 130990 800
rect 131302 -400 131358 800
rect 131578 -400 131634 800
rect 131946 -400 132002 800
rect 132314 -400 132370 800
rect 132682 -400 132738 800
rect 133050 -400 133106 800
rect 133418 -400 133474 800
rect 133786 -400 133842 800
rect 134154 -400 134210 800
rect 134430 -400 134486 800
rect 134798 -400 134854 800
rect 135166 -400 135222 800
rect 135534 -400 135590 800
rect 135902 -400 135958 800
rect 136270 -400 136326 800
rect 136638 -400 136694 800
rect 137006 -400 137062 800
rect 137282 -400 137338 800
rect 137650 -400 137706 800
rect 138018 -400 138074 800
rect 138386 -400 138442 800
rect 138754 -400 138810 800
rect 139122 -400 139178 800
rect 139490 -400 139546 800
rect 139858 -400 139914 800
rect 140134 -400 140190 800
rect 140502 -400 140558 800
rect 140870 -400 140926 800
rect 141238 -400 141294 800
rect 141606 -400 141662 800
rect 141974 -400 142030 800
rect 142342 -400 142398 800
rect 142710 -400 142766 800
rect 142986 -400 143042 800
rect 143354 -400 143410 800
rect 143722 -400 143778 800
rect 144090 -400 144146 800
rect 144458 -400 144514 800
rect 144826 -400 144882 800
rect 145194 -400 145250 800
rect 145562 -400 145618 800
rect 145838 -400 145894 800
rect 146206 -400 146262 800
rect 146574 -400 146630 800
rect 146942 -400 146998 800
rect 147310 -400 147366 800
rect 147678 -400 147734 800
rect 148046 -400 148102 800
rect 148414 -400 148470 800
rect 148690 -400 148746 800
rect 149058 -400 149114 800
rect 149426 -400 149482 800
rect 149794 -400 149850 800
rect 150162 -400 150218 800
rect 150530 -400 150586 800
rect 150898 -400 150954 800
rect 151266 -400 151322 800
rect 151542 -400 151598 800
rect 151910 -400 151966 800
rect 152278 -400 152334 800
rect 152646 -400 152702 800
rect 153014 -400 153070 800
rect 153382 -400 153438 800
rect 153750 -400 153806 800
rect 154118 -400 154174 800
rect 154394 -400 154450 800
rect 154762 -400 154818 800
rect 155130 -400 155186 800
rect 155498 -400 155554 800
rect 155866 -400 155922 800
rect 156234 -400 156290 800
rect 156602 -400 156658 800
rect 156970 -400 157026 800
rect 157246 -400 157302 800
rect 157614 -400 157670 800
rect 157982 -400 158038 800
rect 158350 -400 158406 800
rect 158718 -400 158774 800
rect 159086 -400 159142 800
rect 159454 -400 159510 800
rect 159822 -400 159878 800
rect 160098 -400 160154 800
rect 160466 -400 160522 800
rect 160834 -400 160890 800
rect 161202 -400 161258 800
rect 161570 -400 161626 800
rect 161938 -400 161994 800
rect 162306 -400 162362 800
rect 162674 -400 162730 800
rect 162950 -400 163006 800
rect 163318 -400 163374 800
rect 163686 -400 163742 800
rect 164054 -400 164110 800
rect 164422 -400 164478 800
rect 164790 -400 164846 800
rect 165158 -400 165214 800
rect 165526 -400 165582 800
rect 165802 -400 165858 800
rect 166170 -400 166226 800
rect 166538 -400 166594 800
rect 166906 -400 166962 800
rect 167274 -400 167330 800
rect 167642 -400 167698 800
rect 168010 -400 168066 800
rect 168378 -400 168434 800
rect 168654 -400 168710 800
rect 169022 -400 169078 800
rect 169390 -400 169446 800
rect 169758 -400 169814 800
rect 170126 -400 170182 800
rect 170494 -400 170550 800
rect 170862 -400 170918 800
rect 171230 -400 171286 800
rect 171506 -400 171562 800
rect 171874 -400 171930 800
rect 172242 -400 172298 800
rect 172610 -400 172666 800
rect 172978 -400 173034 800
rect 173346 -400 173402 800
rect 173714 -400 173770 800
rect 174082 -400 174138 800
rect 174358 -400 174414 800
rect 174726 -400 174782 800
rect 175094 -400 175150 800
rect 175462 -400 175518 800
rect 175830 -400 175886 800
rect 176198 -400 176254 800
rect 176566 -400 176622 800
rect 176934 -400 176990 800
rect 177210 -400 177266 800
rect 177578 -400 177634 800
rect 177946 -400 178002 800
rect 178314 -400 178370 800
rect 178682 -400 178738 800
rect 179050 -400 179106 800
rect 179418 -400 179474 800
rect 179786 -400 179842 800
rect 180062 -400 180118 800
rect 180430 -400 180486 800
rect 180798 -400 180854 800
rect 181166 -400 181222 800
rect 181534 -400 181590 800
rect 181902 -400 181958 800
rect 182270 -400 182326 800
rect 182638 -400 182694 800
rect 182914 -400 182970 800
rect 183282 -400 183338 800
rect 183650 -400 183706 800
rect 184018 -400 184074 800
rect 184386 -400 184442 800
rect 184754 -400 184810 800
rect 185122 -400 185178 800
rect 185490 -400 185546 800
rect 185766 -400 185822 800
rect 186134 -400 186190 800
rect 186502 -400 186558 800
rect 186870 -400 186926 800
rect 187238 -400 187294 800
rect 187606 -400 187662 800
rect 187974 -400 188030 800
rect 188342 -400 188398 800
rect 188618 -400 188674 800
rect 188986 -400 189042 800
rect 189354 -400 189410 800
rect 189722 -400 189778 800
rect 190090 -400 190146 800
rect 190458 -400 190514 800
rect 190826 -400 190882 800
rect 191194 -400 191250 800
rect 191470 -400 191526 800
rect 191838 -400 191894 800
rect 192206 -400 192262 800
rect 192574 -400 192630 800
rect 192942 -400 192998 800
rect 193310 -400 193366 800
rect 193678 -400 193734 800
rect 194046 -400 194102 800
rect 194322 -400 194378 800
rect 194690 -400 194746 800
rect 195058 -400 195114 800
rect 195426 -400 195482 800
rect 195794 -400 195850 800
rect 196162 -400 196218 800
rect 196530 -400 196586 800
rect 196898 -400 196954 800
rect 197174 -400 197230 800
rect 197542 -400 197598 800
rect 197910 -400 197966 800
rect 198278 -400 198334 800
rect 198646 -400 198702 800
rect 199014 -400 199070 800
rect 199382 -400 199438 800
rect 199750 -400 199806 800
rect 200026 -400 200082 800
rect 200394 -400 200450 800
rect 200762 -400 200818 800
rect 201130 -400 201186 800
rect 201498 -400 201554 800
rect 201866 -400 201922 800
rect 202234 -400 202290 800
rect 202602 -400 202658 800
rect 202878 -400 202934 800
rect 203246 -400 203302 800
rect 203614 -400 203670 800
rect 203982 -400 204038 800
rect 204350 -400 204406 800
rect 204718 -400 204774 800
rect 205086 -400 205142 800
rect 205454 -400 205510 800
rect 205730 -400 205786 800
rect 206098 -400 206154 800
rect 206466 -400 206522 800
rect 206834 -400 206890 800
rect 207202 -400 207258 800
rect 207570 -400 207626 800
rect 207938 -400 207994 800
rect 208306 -400 208362 800
rect 208582 -400 208638 800
rect 208950 -400 209006 800
rect 209318 -400 209374 800
rect 209686 -400 209742 800
rect 210054 -400 210110 800
rect 210422 -400 210478 800
rect 210790 -400 210846 800
rect 211158 -400 211214 800
rect 211434 -400 211490 800
rect 211802 -400 211858 800
rect 212170 -400 212226 800
rect 212538 -400 212594 800
rect 212906 -400 212962 800
rect 213274 -400 213330 800
rect 213642 -400 213698 800
rect 214010 -400 214066 800
rect 214286 -400 214342 800
rect 214654 -400 214710 800
rect 215022 -400 215078 800
rect 215390 -400 215446 800
rect 215758 -400 215814 800
rect 216126 -400 216182 800
rect 216494 -400 216550 800
rect 216862 -400 216918 800
rect 217138 -400 217194 800
rect 217506 -400 217562 800
rect 217874 -400 217930 800
rect 218242 -400 218298 800
rect 218610 -400 218666 800
rect 218978 -400 219034 800
rect 219346 -400 219402 800
rect 219714 -400 219770 800
<< obsm2 >>
rect 112 31144 146 31958
rect 314 31144 514 31958
rect 682 31144 974 31958
rect 1142 31144 1434 31958
rect 1602 31144 1894 31958
rect 2062 31144 2354 31958
rect 2522 31144 2814 31958
rect 2982 31144 3182 31958
rect 3350 31144 3642 31958
rect 3810 31144 4102 31958
rect 4270 31144 4562 31958
rect 4730 31144 5022 31958
rect 5190 31144 5482 31958
rect 5650 31144 5850 31958
rect 6018 31144 6310 31958
rect 6478 31144 6770 31958
rect 6938 31144 7230 31958
rect 7398 31144 7690 31958
rect 7858 31144 8150 31958
rect 8318 31144 8518 31958
rect 8686 31144 8978 31958
rect 9146 31144 9438 31958
rect 9606 31144 9898 31958
rect 10066 31144 10358 31958
rect 10526 31144 10818 31958
rect 10986 31144 11278 31958
rect 11446 31144 11646 31958
rect 11814 31144 12106 31958
rect 12274 31144 12566 31958
rect 12734 31144 13026 31958
rect 13194 31144 13486 31958
rect 13654 31144 13946 31958
rect 14114 31144 14314 31958
rect 14482 31144 14774 31958
rect 14942 31144 15234 31958
rect 15402 31144 15694 31958
rect 15862 31144 16154 31958
rect 16322 31144 16614 31958
rect 16782 31144 16982 31958
rect 17150 31144 17442 31958
rect 17610 31144 17902 31958
rect 18070 31144 18362 31958
rect 18530 31144 18822 31958
rect 18990 31144 19282 31958
rect 19450 31144 19650 31958
rect 19818 31144 20110 31958
rect 20278 31144 20570 31958
rect 20738 31144 21030 31958
rect 21198 31144 21490 31958
rect 21658 31144 21950 31958
rect 22118 31144 22410 31958
rect 22578 31144 22778 31958
rect 22946 31144 23238 31958
rect 23406 31144 23698 31958
rect 23866 31144 24158 31958
rect 24326 31144 24618 31958
rect 24786 31144 25078 31958
rect 25246 31144 25446 31958
rect 25614 31144 25906 31958
rect 26074 31144 26366 31958
rect 26534 31144 26826 31958
rect 26994 31144 27286 31958
rect 27454 31144 27746 31958
rect 27914 31144 28114 31958
rect 28282 31144 28574 31958
rect 28742 31144 29034 31958
rect 29202 31144 29494 31958
rect 29662 31144 29954 31958
rect 30122 31144 30414 31958
rect 30582 31144 30782 31958
rect 30950 31144 31242 31958
rect 31410 31144 31702 31958
rect 31870 31144 32162 31958
rect 32330 31144 32622 31958
rect 32790 31144 33082 31958
rect 33250 31144 33542 31958
rect 33710 31144 33910 31958
rect 34078 31144 34370 31958
rect 34538 31144 34830 31958
rect 34998 31144 35290 31958
rect 35458 31144 35750 31958
rect 35918 31144 36210 31958
rect 36378 31144 36578 31958
rect 36746 31144 37038 31958
rect 37206 31144 37498 31958
rect 37666 31144 37958 31958
rect 38126 31144 38418 31958
rect 38586 31144 38878 31958
rect 39046 31144 39246 31958
rect 39414 31144 39706 31958
rect 39874 31144 40166 31958
rect 40334 31144 40626 31958
rect 40794 31144 41086 31958
rect 41254 31144 41546 31958
rect 41714 31144 41914 31958
rect 42082 31144 42374 31958
rect 42542 31144 42834 31958
rect 43002 31144 43294 31958
rect 43462 31144 43754 31958
rect 43922 31144 44214 31958
rect 44382 31144 44674 31958
rect 44842 31144 45042 31958
rect 45210 31144 45502 31958
rect 45670 31144 45962 31958
rect 46130 31144 46422 31958
rect 46590 31144 46882 31958
rect 47050 31144 47342 31958
rect 47510 31144 47710 31958
rect 47878 31144 48170 31958
rect 48338 31144 48630 31958
rect 48798 31144 49090 31958
rect 49258 31144 49550 31958
rect 49718 31144 50010 31958
rect 50178 31144 50378 31958
rect 50546 31144 50838 31958
rect 51006 31144 51298 31958
rect 51466 31144 51758 31958
rect 51926 31144 52218 31958
rect 52386 31144 52678 31958
rect 52846 31144 53046 31958
rect 53214 31144 53506 31958
rect 53674 31144 53966 31958
rect 54134 31144 54426 31958
rect 54594 31144 54886 31958
rect 55054 31144 55346 31958
rect 55514 31144 55806 31958
rect 55974 31144 56174 31958
rect 56342 31144 56634 31958
rect 56802 31144 57094 31958
rect 57262 31144 57554 31958
rect 57722 31144 58014 31958
rect 58182 31144 58474 31958
rect 58642 31144 58842 31958
rect 59010 31144 59302 31958
rect 59470 31144 59762 31958
rect 59930 31144 60222 31958
rect 60390 31144 60682 31958
rect 60850 31144 61142 31958
rect 61310 31144 61510 31958
rect 61678 31144 61970 31958
rect 62138 31144 62430 31958
rect 62598 31144 62890 31958
rect 63058 31144 63350 31958
rect 63518 31144 63810 31958
rect 63978 31144 64178 31958
rect 64346 31144 64638 31958
rect 64806 31144 65098 31958
rect 65266 31144 65558 31958
rect 65726 31144 66018 31958
rect 66186 31144 66478 31958
rect 66646 31144 66938 31958
rect 67106 31144 67306 31958
rect 67474 31144 67766 31958
rect 67934 31144 68226 31958
rect 68394 31144 68686 31958
rect 68854 31144 69146 31958
rect 69314 31144 69606 31958
rect 69774 31144 69974 31958
rect 70142 31144 70434 31958
rect 70602 31144 70894 31958
rect 71062 31144 71354 31958
rect 71522 31144 71814 31958
rect 71982 31144 72274 31958
rect 72442 31144 72642 31958
rect 72810 31144 73102 31958
rect 73270 31144 73562 31958
rect 73730 31144 74022 31958
rect 74190 31144 74482 31958
rect 74650 31144 74942 31958
rect 75110 31144 75310 31958
rect 75478 31144 75770 31958
rect 75938 31144 76230 31958
rect 76398 31144 76690 31958
rect 76858 31144 77150 31958
rect 77318 31144 77610 31958
rect 77778 31144 78070 31958
rect 78238 31144 78438 31958
rect 78606 31144 78898 31958
rect 79066 31144 79358 31958
rect 79526 31144 79818 31958
rect 79986 31144 80278 31958
rect 80446 31144 80738 31958
rect 80906 31144 81106 31958
rect 81274 31144 81566 31958
rect 81734 31144 82026 31958
rect 82194 31144 82486 31958
rect 82654 31144 82946 31958
rect 83114 31144 83406 31958
rect 83574 31144 83774 31958
rect 83942 31144 84234 31958
rect 84402 31144 84694 31958
rect 84862 31144 85154 31958
rect 85322 31144 85614 31958
rect 85782 31144 86074 31958
rect 86242 31144 86442 31958
rect 86610 31144 86902 31958
rect 87070 31144 87362 31958
rect 87530 31144 87822 31958
rect 87990 31144 88282 31958
rect 88450 31144 88742 31958
rect 88910 31144 89202 31958
rect 89370 31144 89570 31958
rect 89738 31144 90030 31958
rect 90198 31144 90490 31958
rect 90658 31144 90950 31958
rect 91118 31144 91410 31958
rect 91578 31144 91870 31958
rect 92038 31144 92238 31958
rect 92406 31144 92698 31958
rect 92866 31144 93158 31958
rect 93326 31144 93618 31958
rect 93786 31144 94078 31958
rect 94246 31144 94538 31958
rect 94706 31144 94906 31958
rect 95074 31144 95366 31958
rect 95534 31144 95826 31958
rect 95994 31144 96286 31958
rect 96454 31144 96746 31958
rect 96914 31144 97206 31958
rect 97374 31144 97574 31958
rect 97742 31144 98034 31958
rect 98202 31144 98494 31958
rect 98662 31144 98954 31958
rect 99122 31144 99414 31958
rect 99582 31144 99874 31958
rect 100042 31144 100334 31958
rect 100502 31144 100702 31958
rect 100870 31144 101162 31958
rect 101330 31144 101622 31958
rect 101790 31144 102082 31958
rect 102250 31144 102542 31958
rect 102710 31144 103002 31958
rect 103170 31144 103370 31958
rect 103538 31144 103830 31958
rect 103998 31144 104290 31958
rect 104458 31144 104750 31958
rect 104918 31144 105210 31958
rect 105378 31144 105670 31958
rect 105838 31144 106038 31958
rect 106206 31144 106498 31958
rect 106666 31144 106958 31958
rect 107126 31144 107418 31958
rect 107586 31144 107878 31958
rect 108046 31144 108338 31958
rect 108506 31144 108706 31958
rect 108874 31144 109166 31958
rect 109334 31144 109626 31958
rect 109794 31144 110086 31958
rect 110254 31144 110546 31958
rect 110714 31144 111006 31958
rect 111174 31144 111466 31958
rect 111634 31144 111834 31958
rect 112002 31144 112294 31958
rect 112462 31144 112754 31958
rect 112922 31144 113214 31958
rect 113382 31144 113674 31958
rect 113842 31144 114134 31958
rect 114302 31144 114502 31958
rect 114670 31144 114962 31958
rect 115130 31144 115422 31958
rect 115590 31144 115882 31958
rect 116050 31144 116342 31958
rect 116510 31144 116802 31958
rect 116970 31144 117170 31958
rect 117338 31144 117630 31958
rect 117798 31144 118090 31958
rect 118258 31144 118550 31958
rect 118718 31144 119010 31958
rect 119178 31144 119470 31958
rect 119638 31144 119838 31958
rect 120006 31144 120298 31958
rect 120466 31144 120758 31958
rect 120926 31144 121218 31958
rect 121386 31144 121678 31958
rect 121846 31144 122138 31958
rect 122306 31144 122598 31958
rect 122766 31144 122966 31958
rect 123134 31144 123426 31958
rect 123594 31144 123886 31958
rect 124054 31144 124346 31958
rect 124514 31144 124806 31958
rect 124974 31144 125266 31958
rect 125434 31144 125634 31958
rect 125802 31144 126094 31958
rect 126262 31144 126554 31958
rect 126722 31144 127014 31958
rect 127182 31144 127474 31958
rect 127642 31144 127934 31958
rect 128102 31144 128302 31958
rect 128470 31144 128762 31958
rect 128930 31144 129222 31958
rect 129390 31144 129682 31958
rect 129850 31144 130142 31958
rect 130310 31144 130602 31958
rect 130770 31144 130970 31958
rect 131138 31144 131430 31958
rect 131598 31144 131890 31958
rect 132058 31144 132350 31958
rect 132518 31144 132810 31958
rect 132978 31144 133270 31958
rect 133438 31144 133730 31958
rect 133898 31144 134098 31958
rect 134266 31144 134558 31958
rect 134726 31144 135018 31958
rect 135186 31144 135478 31958
rect 135646 31144 135938 31958
rect 136106 31144 136398 31958
rect 136566 31144 136766 31958
rect 136934 31144 137226 31958
rect 137394 31144 137686 31958
rect 137854 31144 138146 31958
rect 138314 31144 138606 31958
rect 138774 31144 139066 31958
rect 139234 31144 139434 31958
rect 139602 31144 139894 31958
rect 140062 31144 140354 31958
rect 140522 31144 140814 31958
rect 140982 31144 141274 31958
rect 141442 31144 141734 31958
rect 141902 31144 142102 31958
rect 142270 31144 142562 31958
rect 142730 31144 143022 31958
rect 143190 31144 143482 31958
rect 143650 31144 143942 31958
rect 144110 31144 144402 31958
rect 144570 31144 144862 31958
rect 145030 31144 145230 31958
rect 145398 31144 145690 31958
rect 145858 31144 146150 31958
rect 146318 31144 146610 31958
rect 146778 31144 147070 31958
rect 147238 31144 147530 31958
rect 147698 31144 147898 31958
rect 148066 31144 148358 31958
rect 148526 31144 148818 31958
rect 148986 31144 149278 31958
rect 149446 31144 149738 31958
rect 149906 31144 150198 31958
rect 150366 31144 150566 31958
rect 150734 31144 151026 31958
rect 151194 31144 151486 31958
rect 151654 31144 151946 31958
rect 152114 31144 152406 31958
rect 152574 31144 152866 31958
rect 153034 31144 153234 31958
rect 153402 31144 153694 31958
rect 153862 31144 154154 31958
rect 154322 31144 154614 31958
rect 154782 31144 155074 31958
rect 155242 31144 155534 31958
rect 155702 31144 155994 31958
rect 156162 31144 156362 31958
rect 156530 31144 156822 31958
rect 156990 31144 157282 31958
rect 157450 31144 157742 31958
rect 157910 31144 158202 31958
rect 158370 31144 158662 31958
rect 158830 31144 159030 31958
rect 159198 31144 159490 31958
rect 159658 31144 159950 31958
rect 160118 31144 160410 31958
rect 160578 31144 160870 31958
rect 161038 31144 161330 31958
rect 161498 31144 161698 31958
rect 161866 31144 162158 31958
rect 162326 31144 162618 31958
rect 162786 31144 163078 31958
rect 163246 31144 163538 31958
rect 163706 31144 163998 31958
rect 164166 31144 164366 31958
rect 164534 31144 164826 31958
rect 164994 31144 165286 31958
rect 165454 31144 165746 31958
rect 165914 31144 166206 31958
rect 166374 31144 166666 31958
rect 166834 31144 167126 31958
rect 167294 31144 167494 31958
rect 167662 31144 167954 31958
rect 168122 31144 168414 31958
rect 168582 31144 168874 31958
rect 169042 31144 169334 31958
rect 169502 31144 169794 31958
rect 169962 31144 170162 31958
rect 170330 31144 170622 31958
rect 170790 31144 171082 31958
rect 171250 31144 171542 31958
rect 171710 31144 172002 31958
rect 172170 31144 172462 31958
rect 172630 31144 172830 31958
rect 172998 31144 173290 31958
rect 173458 31144 173750 31958
rect 173918 31144 174210 31958
rect 174378 31144 174670 31958
rect 174838 31144 175130 31958
rect 175298 31144 175498 31958
rect 175666 31144 175958 31958
rect 176126 31144 176418 31958
rect 176586 31144 176878 31958
rect 177046 31144 177338 31958
rect 177506 31144 177798 31958
rect 177966 31144 178258 31958
rect 178426 31144 178626 31958
rect 178794 31144 179086 31958
rect 179254 31144 179546 31958
rect 179714 31144 180006 31958
rect 180174 31144 180466 31958
rect 180634 31144 180926 31958
rect 181094 31144 181294 31958
rect 181462 31144 181754 31958
rect 181922 31144 182214 31958
rect 182382 31144 182674 31958
rect 182842 31144 183134 31958
rect 183302 31144 183594 31958
rect 183762 31144 183962 31958
rect 184130 31144 184422 31958
rect 184590 31144 184882 31958
rect 185050 31144 185342 31958
rect 185510 31144 185802 31958
rect 185970 31144 186262 31958
rect 186430 31144 186630 31958
rect 186798 31144 187090 31958
rect 187258 31144 187550 31958
rect 187718 31144 188010 31958
rect 188178 31144 188470 31958
rect 188638 31144 188930 31958
rect 189098 31144 189390 31958
rect 189558 31144 189758 31958
rect 189926 31144 190218 31958
rect 190386 31144 190678 31958
rect 190846 31144 191138 31958
rect 191306 31144 191598 31958
rect 191766 31144 192058 31958
rect 192226 31144 192426 31958
rect 192594 31144 192886 31958
rect 193054 31144 193346 31958
rect 193514 31144 193806 31958
rect 193974 31144 194266 31958
rect 194434 31144 194726 31958
rect 194894 31144 195094 31958
rect 195262 31144 195554 31958
rect 195722 31144 196014 31958
rect 196182 31144 196474 31958
rect 196642 31144 196934 31958
rect 197102 31144 197394 31958
rect 197562 31144 197762 31958
rect 197930 31144 198222 31958
rect 198390 31144 198682 31958
rect 198850 31144 199142 31958
rect 199310 31144 199602 31958
rect 199770 31144 200062 31958
rect 200230 31144 200522 31958
rect 200690 31144 200890 31958
rect 201058 31144 201350 31958
rect 201518 31144 201810 31958
rect 201978 31144 202270 31958
rect 202438 31144 202730 31958
rect 202898 31144 203190 31958
rect 203358 31144 203558 31958
rect 203726 31144 204018 31958
rect 204186 31144 204478 31958
rect 204646 31144 204938 31958
rect 205106 31144 205398 31958
rect 205566 31144 205858 31958
rect 206026 31144 206226 31958
rect 206394 31144 206686 31958
rect 206854 31144 207146 31958
rect 207314 31144 207606 31958
rect 207774 31144 208066 31958
rect 208234 31144 208526 31958
rect 208694 31144 208894 31958
rect 209062 31144 209354 31958
rect 209522 31144 209814 31958
rect 209982 31144 210274 31958
rect 210442 31144 210734 31958
rect 210902 31144 211194 31958
rect 211362 31144 211654 31958
rect 211822 31144 212022 31958
rect 212190 31144 212482 31958
rect 212650 31144 212942 31958
rect 213110 31144 213402 31958
rect 213570 31144 213862 31958
rect 214030 31144 214322 31958
rect 214490 31144 214690 31958
rect 214858 31144 215150 31958
rect 215318 31144 215610 31958
rect 215778 31144 216070 31958
rect 216238 31144 216530 31958
rect 216698 31144 216990 31958
rect 217158 31144 217358 31958
rect 217526 31144 217818 31958
rect 217986 31144 218278 31958
rect 218446 31144 218738 31958
rect 218906 31144 219198 31958
rect 219366 31144 219658 31958
rect 112 856 219768 31144
rect 222 2 330 856
rect 498 2 698 856
rect 866 2 1066 856
rect 1234 2 1434 856
rect 1602 2 1802 856
rect 1970 2 2170 856
rect 2338 2 2538 856
rect 2706 2 2906 856
rect 3074 2 3182 856
rect 3350 2 3550 856
rect 3718 2 3918 856
rect 4086 2 4286 856
rect 4454 2 4654 856
rect 4822 2 5022 856
rect 5190 2 5390 856
rect 5558 2 5758 856
rect 5926 2 6034 856
rect 6202 2 6402 856
rect 6570 2 6770 856
rect 6938 2 7138 856
rect 7306 2 7506 856
rect 7674 2 7874 856
rect 8042 2 8242 856
rect 8410 2 8610 856
rect 8778 2 8886 856
rect 9054 2 9254 856
rect 9422 2 9622 856
rect 9790 2 9990 856
rect 10158 2 10358 856
rect 10526 2 10726 856
rect 10894 2 11094 856
rect 11262 2 11462 856
rect 11630 2 11738 856
rect 11906 2 12106 856
rect 12274 2 12474 856
rect 12642 2 12842 856
rect 13010 2 13210 856
rect 13378 2 13578 856
rect 13746 2 13946 856
rect 14114 2 14314 856
rect 14482 2 14590 856
rect 14758 2 14958 856
rect 15126 2 15326 856
rect 15494 2 15694 856
rect 15862 2 16062 856
rect 16230 2 16430 856
rect 16598 2 16798 856
rect 16966 2 17166 856
rect 17334 2 17442 856
rect 17610 2 17810 856
rect 17978 2 18178 856
rect 18346 2 18546 856
rect 18714 2 18914 856
rect 19082 2 19282 856
rect 19450 2 19650 856
rect 19818 2 20018 856
rect 20186 2 20294 856
rect 20462 2 20662 856
rect 20830 2 21030 856
rect 21198 2 21398 856
rect 21566 2 21766 856
rect 21934 2 22134 856
rect 22302 2 22502 856
rect 22670 2 22870 856
rect 23038 2 23146 856
rect 23314 2 23514 856
rect 23682 2 23882 856
rect 24050 2 24250 856
rect 24418 2 24618 856
rect 24786 2 24986 856
rect 25154 2 25354 856
rect 25522 2 25722 856
rect 25890 2 25998 856
rect 26166 2 26366 856
rect 26534 2 26734 856
rect 26902 2 27102 856
rect 27270 2 27470 856
rect 27638 2 27838 856
rect 28006 2 28206 856
rect 28374 2 28574 856
rect 28742 2 28850 856
rect 29018 2 29218 856
rect 29386 2 29586 856
rect 29754 2 29954 856
rect 30122 2 30322 856
rect 30490 2 30690 856
rect 30858 2 31058 856
rect 31226 2 31426 856
rect 31594 2 31702 856
rect 31870 2 32070 856
rect 32238 2 32438 856
rect 32606 2 32806 856
rect 32974 2 33174 856
rect 33342 2 33542 856
rect 33710 2 33910 856
rect 34078 2 34278 856
rect 34446 2 34554 856
rect 34722 2 34922 856
rect 35090 2 35290 856
rect 35458 2 35658 856
rect 35826 2 36026 856
rect 36194 2 36394 856
rect 36562 2 36762 856
rect 36930 2 37130 856
rect 37298 2 37406 856
rect 37574 2 37774 856
rect 37942 2 38142 856
rect 38310 2 38510 856
rect 38678 2 38878 856
rect 39046 2 39246 856
rect 39414 2 39614 856
rect 39782 2 39982 856
rect 40150 2 40258 856
rect 40426 2 40626 856
rect 40794 2 40994 856
rect 41162 2 41362 856
rect 41530 2 41730 856
rect 41898 2 42098 856
rect 42266 2 42466 856
rect 42634 2 42834 856
rect 43002 2 43110 856
rect 43278 2 43478 856
rect 43646 2 43846 856
rect 44014 2 44214 856
rect 44382 2 44582 856
rect 44750 2 44950 856
rect 45118 2 45318 856
rect 45486 2 45686 856
rect 45854 2 45962 856
rect 46130 2 46330 856
rect 46498 2 46698 856
rect 46866 2 47066 856
rect 47234 2 47434 856
rect 47602 2 47802 856
rect 47970 2 48170 856
rect 48338 2 48538 856
rect 48706 2 48814 856
rect 48982 2 49182 856
rect 49350 2 49550 856
rect 49718 2 49918 856
rect 50086 2 50286 856
rect 50454 2 50654 856
rect 50822 2 51022 856
rect 51190 2 51390 856
rect 51558 2 51666 856
rect 51834 2 52034 856
rect 52202 2 52402 856
rect 52570 2 52770 856
rect 52938 2 53138 856
rect 53306 2 53506 856
rect 53674 2 53874 856
rect 54042 2 54242 856
rect 54410 2 54518 856
rect 54686 2 54886 856
rect 55054 2 55254 856
rect 55422 2 55622 856
rect 55790 2 55990 856
rect 56158 2 56358 856
rect 56526 2 56726 856
rect 56894 2 57094 856
rect 57262 2 57370 856
rect 57538 2 57738 856
rect 57906 2 58106 856
rect 58274 2 58474 856
rect 58642 2 58842 856
rect 59010 2 59210 856
rect 59378 2 59578 856
rect 59746 2 59946 856
rect 60114 2 60222 856
rect 60390 2 60590 856
rect 60758 2 60958 856
rect 61126 2 61326 856
rect 61494 2 61694 856
rect 61862 2 62062 856
rect 62230 2 62430 856
rect 62598 2 62798 856
rect 62966 2 63074 856
rect 63242 2 63442 856
rect 63610 2 63810 856
rect 63978 2 64178 856
rect 64346 2 64546 856
rect 64714 2 64914 856
rect 65082 2 65282 856
rect 65450 2 65650 856
rect 65818 2 65926 856
rect 66094 2 66294 856
rect 66462 2 66662 856
rect 66830 2 67030 856
rect 67198 2 67398 856
rect 67566 2 67766 856
rect 67934 2 68134 856
rect 68302 2 68502 856
rect 68670 2 68778 856
rect 68946 2 69146 856
rect 69314 2 69514 856
rect 69682 2 69882 856
rect 70050 2 70250 856
rect 70418 2 70618 856
rect 70786 2 70986 856
rect 71154 2 71354 856
rect 71522 2 71630 856
rect 71798 2 71998 856
rect 72166 2 72366 856
rect 72534 2 72734 856
rect 72902 2 73102 856
rect 73270 2 73470 856
rect 73638 2 73838 856
rect 74006 2 74206 856
rect 74374 2 74482 856
rect 74650 2 74850 856
rect 75018 2 75218 856
rect 75386 2 75586 856
rect 75754 2 75954 856
rect 76122 2 76322 856
rect 76490 2 76690 856
rect 76858 2 77058 856
rect 77226 2 77334 856
rect 77502 2 77702 856
rect 77870 2 78070 856
rect 78238 2 78438 856
rect 78606 2 78806 856
rect 78974 2 79174 856
rect 79342 2 79542 856
rect 79710 2 79910 856
rect 80078 2 80186 856
rect 80354 2 80554 856
rect 80722 2 80922 856
rect 81090 2 81290 856
rect 81458 2 81658 856
rect 81826 2 82026 856
rect 82194 2 82394 856
rect 82562 2 82762 856
rect 82930 2 83038 856
rect 83206 2 83406 856
rect 83574 2 83774 856
rect 83942 2 84142 856
rect 84310 2 84510 856
rect 84678 2 84878 856
rect 85046 2 85246 856
rect 85414 2 85614 856
rect 85782 2 85890 856
rect 86058 2 86258 856
rect 86426 2 86626 856
rect 86794 2 86994 856
rect 87162 2 87362 856
rect 87530 2 87730 856
rect 87898 2 88098 856
rect 88266 2 88466 856
rect 88634 2 88742 856
rect 88910 2 89110 856
rect 89278 2 89478 856
rect 89646 2 89846 856
rect 90014 2 90214 856
rect 90382 2 90582 856
rect 90750 2 90950 856
rect 91118 2 91318 856
rect 91486 2 91594 856
rect 91762 2 91962 856
rect 92130 2 92330 856
rect 92498 2 92698 856
rect 92866 2 93066 856
rect 93234 2 93434 856
rect 93602 2 93802 856
rect 93970 2 94170 856
rect 94338 2 94446 856
rect 94614 2 94814 856
rect 94982 2 95182 856
rect 95350 2 95550 856
rect 95718 2 95918 856
rect 96086 2 96286 856
rect 96454 2 96654 856
rect 96822 2 97022 856
rect 97190 2 97298 856
rect 97466 2 97666 856
rect 97834 2 98034 856
rect 98202 2 98402 856
rect 98570 2 98770 856
rect 98938 2 99138 856
rect 99306 2 99506 856
rect 99674 2 99874 856
rect 100042 2 100150 856
rect 100318 2 100518 856
rect 100686 2 100886 856
rect 101054 2 101254 856
rect 101422 2 101622 856
rect 101790 2 101990 856
rect 102158 2 102358 856
rect 102526 2 102726 856
rect 102894 2 103002 856
rect 103170 2 103370 856
rect 103538 2 103738 856
rect 103906 2 104106 856
rect 104274 2 104474 856
rect 104642 2 104842 856
rect 105010 2 105210 856
rect 105378 2 105578 856
rect 105746 2 105854 856
rect 106022 2 106222 856
rect 106390 2 106590 856
rect 106758 2 106958 856
rect 107126 2 107326 856
rect 107494 2 107694 856
rect 107862 2 108062 856
rect 108230 2 108430 856
rect 108598 2 108706 856
rect 108874 2 109074 856
rect 109242 2 109442 856
rect 109610 2 109810 856
rect 109978 2 110178 856
rect 110346 2 110546 856
rect 110714 2 110914 856
rect 111082 2 111282 856
rect 111450 2 111558 856
rect 111726 2 111926 856
rect 112094 2 112294 856
rect 112462 2 112662 856
rect 112830 2 113030 856
rect 113198 2 113398 856
rect 113566 2 113766 856
rect 113934 2 114134 856
rect 114302 2 114410 856
rect 114578 2 114778 856
rect 114946 2 115146 856
rect 115314 2 115514 856
rect 115682 2 115882 856
rect 116050 2 116250 856
rect 116418 2 116618 856
rect 116786 2 116986 856
rect 117154 2 117262 856
rect 117430 2 117630 856
rect 117798 2 117998 856
rect 118166 2 118366 856
rect 118534 2 118734 856
rect 118902 2 119102 856
rect 119270 2 119470 856
rect 119638 2 119838 856
rect 120006 2 120114 856
rect 120282 2 120482 856
rect 120650 2 120850 856
rect 121018 2 121218 856
rect 121386 2 121586 856
rect 121754 2 121954 856
rect 122122 2 122322 856
rect 122490 2 122690 856
rect 122858 2 122966 856
rect 123134 2 123334 856
rect 123502 2 123702 856
rect 123870 2 124070 856
rect 124238 2 124438 856
rect 124606 2 124806 856
rect 124974 2 125174 856
rect 125342 2 125542 856
rect 125710 2 125818 856
rect 125986 2 126186 856
rect 126354 2 126554 856
rect 126722 2 126922 856
rect 127090 2 127290 856
rect 127458 2 127658 856
rect 127826 2 128026 856
rect 128194 2 128394 856
rect 128562 2 128670 856
rect 128838 2 129038 856
rect 129206 2 129406 856
rect 129574 2 129774 856
rect 129942 2 130142 856
rect 130310 2 130510 856
rect 130678 2 130878 856
rect 131046 2 131246 856
rect 131414 2 131522 856
rect 131690 2 131890 856
rect 132058 2 132258 856
rect 132426 2 132626 856
rect 132794 2 132994 856
rect 133162 2 133362 856
rect 133530 2 133730 856
rect 133898 2 134098 856
rect 134266 2 134374 856
rect 134542 2 134742 856
rect 134910 2 135110 856
rect 135278 2 135478 856
rect 135646 2 135846 856
rect 136014 2 136214 856
rect 136382 2 136582 856
rect 136750 2 136950 856
rect 137118 2 137226 856
rect 137394 2 137594 856
rect 137762 2 137962 856
rect 138130 2 138330 856
rect 138498 2 138698 856
rect 138866 2 139066 856
rect 139234 2 139434 856
rect 139602 2 139802 856
rect 139970 2 140078 856
rect 140246 2 140446 856
rect 140614 2 140814 856
rect 140982 2 141182 856
rect 141350 2 141550 856
rect 141718 2 141918 856
rect 142086 2 142286 856
rect 142454 2 142654 856
rect 142822 2 142930 856
rect 143098 2 143298 856
rect 143466 2 143666 856
rect 143834 2 144034 856
rect 144202 2 144402 856
rect 144570 2 144770 856
rect 144938 2 145138 856
rect 145306 2 145506 856
rect 145674 2 145782 856
rect 145950 2 146150 856
rect 146318 2 146518 856
rect 146686 2 146886 856
rect 147054 2 147254 856
rect 147422 2 147622 856
rect 147790 2 147990 856
rect 148158 2 148358 856
rect 148526 2 148634 856
rect 148802 2 149002 856
rect 149170 2 149370 856
rect 149538 2 149738 856
rect 149906 2 150106 856
rect 150274 2 150474 856
rect 150642 2 150842 856
rect 151010 2 151210 856
rect 151378 2 151486 856
rect 151654 2 151854 856
rect 152022 2 152222 856
rect 152390 2 152590 856
rect 152758 2 152958 856
rect 153126 2 153326 856
rect 153494 2 153694 856
rect 153862 2 154062 856
rect 154230 2 154338 856
rect 154506 2 154706 856
rect 154874 2 155074 856
rect 155242 2 155442 856
rect 155610 2 155810 856
rect 155978 2 156178 856
rect 156346 2 156546 856
rect 156714 2 156914 856
rect 157082 2 157190 856
rect 157358 2 157558 856
rect 157726 2 157926 856
rect 158094 2 158294 856
rect 158462 2 158662 856
rect 158830 2 159030 856
rect 159198 2 159398 856
rect 159566 2 159766 856
rect 159934 2 160042 856
rect 160210 2 160410 856
rect 160578 2 160778 856
rect 160946 2 161146 856
rect 161314 2 161514 856
rect 161682 2 161882 856
rect 162050 2 162250 856
rect 162418 2 162618 856
rect 162786 2 162894 856
rect 163062 2 163262 856
rect 163430 2 163630 856
rect 163798 2 163998 856
rect 164166 2 164366 856
rect 164534 2 164734 856
rect 164902 2 165102 856
rect 165270 2 165470 856
rect 165638 2 165746 856
rect 165914 2 166114 856
rect 166282 2 166482 856
rect 166650 2 166850 856
rect 167018 2 167218 856
rect 167386 2 167586 856
rect 167754 2 167954 856
rect 168122 2 168322 856
rect 168490 2 168598 856
rect 168766 2 168966 856
rect 169134 2 169334 856
rect 169502 2 169702 856
rect 169870 2 170070 856
rect 170238 2 170438 856
rect 170606 2 170806 856
rect 170974 2 171174 856
rect 171342 2 171450 856
rect 171618 2 171818 856
rect 171986 2 172186 856
rect 172354 2 172554 856
rect 172722 2 172922 856
rect 173090 2 173290 856
rect 173458 2 173658 856
rect 173826 2 174026 856
rect 174194 2 174302 856
rect 174470 2 174670 856
rect 174838 2 175038 856
rect 175206 2 175406 856
rect 175574 2 175774 856
rect 175942 2 176142 856
rect 176310 2 176510 856
rect 176678 2 176878 856
rect 177046 2 177154 856
rect 177322 2 177522 856
rect 177690 2 177890 856
rect 178058 2 178258 856
rect 178426 2 178626 856
rect 178794 2 178994 856
rect 179162 2 179362 856
rect 179530 2 179730 856
rect 179898 2 180006 856
rect 180174 2 180374 856
rect 180542 2 180742 856
rect 180910 2 181110 856
rect 181278 2 181478 856
rect 181646 2 181846 856
rect 182014 2 182214 856
rect 182382 2 182582 856
rect 182750 2 182858 856
rect 183026 2 183226 856
rect 183394 2 183594 856
rect 183762 2 183962 856
rect 184130 2 184330 856
rect 184498 2 184698 856
rect 184866 2 185066 856
rect 185234 2 185434 856
rect 185602 2 185710 856
rect 185878 2 186078 856
rect 186246 2 186446 856
rect 186614 2 186814 856
rect 186982 2 187182 856
rect 187350 2 187550 856
rect 187718 2 187918 856
rect 188086 2 188286 856
rect 188454 2 188562 856
rect 188730 2 188930 856
rect 189098 2 189298 856
rect 189466 2 189666 856
rect 189834 2 190034 856
rect 190202 2 190402 856
rect 190570 2 190770 856
rect 190938 2 191138 856
rect 191306 2 191414 856
rect 191582 2 191782 856
rect 191950 2 192150 856
rect 192318 2 192518 856
rect 192686 2 192886 856
rect 193054 2 193254 856
rect 193422 2 193622 856
rect 193790 2 193990 856
rect 194158 2 194266 856
rect 194434 2 194634 856
rect 194802 2 195002 856
rect 195170 2 195370 856
rect 195538 2 195738 856
rect 195906 2 196106 856
rect 196274 2 196474 856
rect 196642 2 196842 856
rect 197010 2 197118 856
rect 197286 2 197486 856
rect 197654 2 197854 856
rect 198022 2 198222 856
rect 198390 2 198590 856
rect 198758 2 198958 856
rect 199126 2 199326 856
rect 199494 2 199694 856
rect 199862 2 199970 856
rect 200138 2 200338 856
rect 200506 2 200706 856
rect 200874 2 201074 856
rect 201242 2 201442 856
rect 201610 2 201810 856
rect 201978 2 202178 856
rect 202346 2 202546 856
rect 202714 2 202822 856
rect 202990 2 203190 856
rect 203358 2 203558 856
rect 203726 2 203926 856
rect 204094 2 204294 856
rect 204462 2 204662 856
rect 204830 2 205030 856
rect 205198 2 205398 856
rect 205566 2 205674 856
rect 205842 2 206042 856
rect 206210 2 206410 856
rect 206578 2 206778 856
rect 206946 2 207146 856
rect 207314 2 207514 856
rect 207682 2 207882 856
rect 208050 2 208250 856
rect 208418 2 208526 856
rect 208694 2 208894 856
rect 209062 2 209262 856
rect 209430 2 209630 856
rect 209798 2 209998 856
rect 210166 2 210366 856
rect 210534 2 210734 856
rect 210902 2 211102 856
rect 211270 2 211378 856
rect 211546 2 211746 856
rect 211914 2 212114 856
rect 212282 2 212482 856
rect 212650 2 212850 856
rect 213018 2 213218 856
rect 213386 2 213586 856
rect 213754 2 213954 856
rect 214122 2 214230 856
rect 214398 2 214598 856
rect 214766 2 214966 856
rect 215134 2 215334 856
rect 215502 2 215702 856
rect 215870 2 216070 856
rect 216238 2 216438 856
rect 216606 2 216806 856
rect 216974 2 217082 856
rect 217250 2 217450 856
rect 217618 2 217818 856
rect 217986 2 218186 856
rect 218354 2 218554 856
rect 218722 2 218922 856
rect 219090 2 219290 856
rect 219458 2 219658 856
<< metal3 >>
rect 219200 30200 220400 30320
rect 219200 27072 220400 27192
rect -400 26528 800 26648
rect 219200 23808 220400 23928
rect 219200 20680 220400 20800
rect 219200 17416 220400 17536
rect -400 15920 800 16040
rect 219200 14288 220400 14408
rect 219200 11024 220400 11144
rect 219200 7896 220400 8016
rect -400 5312 800 5432
rect 219200 4632 220400 4752
rect 219200 1504 220400 1624
<< obsm3 >>
rect 800 30400 219200 31109
rect 800 30120 219120 30400
rect 800 27272 219200 30120
rect 800 26992 219120 27272
rect 800 26728 219200 26992
rect 880 26448 219200 26728
rect 800 24008 219200 26448
rect 800 23728 219120 24008
rect 800 20880 219200 23728
rect 800 20600 219120 20880
rect 800 17616 219200 20600
rect 800 17336 219120 17616
rect 800 16120 219200 17336
rect 880 15840 219200 16120
rect 800 14488 219200 15840
rect 800 14208 219120 14488
rect 800 11224 219200 14208
rect 800 10944 219120 11224
rect 800 8096 219200 10944
rect 800 7816 219120 8096
rect 800 5512 219200 7816
rect 880 5232 219200 5512
rect 800 4832 219200 5232
rect 800 4552 219120 4832
rect 800 1704 219200 4552
rect 800 1424 219120 1704
rect 800 35 219200 1424
<< metal4 >>
rect 4014 1040 4194 30512
rect 4834 1088 5014 30464
rect 5654 1088 5834 30464
rect 19064 1040 19244 30512
rect 19884 1088 20064 30464
rect 20704 1088 20884 30464
rect 34114 1040 34294 30512
rect 34934 1088 35114 30464
rect 35754 1088 35934 30464
rect 49164 1040 49344 30512
rect 49984 1088 50164 30464
rect 50804 1088 50984 30464
rect 64214 1040 64394 30512
rect 65034 1088 65214 30464
rect 65854 1088 66034 30464
rect 79264 1040 79444 30512
rect 80084 1088 80264 30464
rect 80904 1088 81084 30464
rect 94314 1040 94494 30512
rect 95134 1088 95314 30464
rect 95954 1088 96134 30464
rect 109364 1040 109544 30512
rect 110184 1088 110364 30464
rect 111004 1088 111184 30464
rect 124414 1040 124594 30512
rect 125234 1088 125414 30464
rect 126054 1088 126234 30464
rect 139464 1040 139644 30512
rect 140284 1088 140464 30464
rect 141104 1088 141284 30464
rect 154514 1040 154694 30512
rect 155334 1088 155514 30464
rect 156154 1088 156334 30464
rect 169564 1040 169744 30512
rect 170384 1088 170564 30464
rect 171204 1088 171384 30464
rect 184614 1040 184794 30512
rect 185434 1088 185614 30464
rect 186254 1088 186434 30464
rect 186814 1088 186994 30464
rect 187414 1088 187594 30464
rect 199664 1040 199844 30512
rect 200484 1088 200664 30464
rect 201304 1088 201484 30464
rect 201864 1088 202044 30464
rect 202464 1088 202644 30464
rect 214714 1040 214894 30512
rect 215534 1088 215714 30464
rect 216354 1088 216534 30464
rect 216914 1088 217094 30464
rect 217514 1088 217694 30464
<< obsm4 >>
rect 67403 960 79184 29477
rect 79524 1008 80004 29477
rect 80344 1008 80824 29477
rect 81164 1008 94234 29477
rect 79524 960 94234 1008
rect 94574 1008 95054 29477
rect 95394 1008 95874 29477
rect 96214 1008 109284 29477
rect 94574 960 109284 1008
rect 109624 1008 110104 29477
rect 110444 1008 110924 29477
rect 111264 1008 124334 29477
rect 109624 960 124334 1008
rect 124674 1008 125154 29477
rect 125494 1008 125974 29477
rect 126314 1008 139384 29477
rect 124674 960 139384 1008
rect 139724 1008 140204 29477
rect 140544 1008 141024 29477
rect 141364 1008 154434 29477
rect 139724 960 154434 1008
rect 154774 1008 155254 29477
rect 155594 1008 156074 29477
rect 156414 1008 169484 29477
rect 154774 960 169484 1008
rect 169824 1008 170304 29477
rect 170644 1008 171124 29477
rect 171464 1008 184534 29477
rect 169824 960 184534 1008
rect 184874 1008 185354 29477
rect 185694 1008 186174 29477
rect 186514 1008 186734 29477
rect 187074 1008 187334 29477
rect 187674 1008 199584 29477
rect 184874 960 199584 1008
rect 199924 1008 200404 29477
rect 200744 1008 201224 29477
rect 201564 1008 201784 29477
rect 202124 1008 202384 29477
rect 202724 1008 213013 29477
rect 199924 960 213013 1008
rect 67403 35 213013 960
<< labels >>
rlabel metal3 s -400 5312 800 5432 6 caravel_clk
port 1 nsew signal input
rlabel metal3 s -400 15920 800 16040 6 caravel_clk2
port 2 nsew signal input
rlabel metal3 s -400 26528 800 26648 6 caravel_rstn
port 3 nsew signal input
rlabel metal2 s 47398 31200 47454 32400 6 la_data_in_core[0]
port 4 nsew signal output
rlabel metal2 s 180982 31200 181038 32400 6 la_data_in_core[100]
port 5 nsew signal output
rlabel metal2 s 182270 31200 182326 32400 6 la_data_in_core[101]
port 6 nsew signal output
rlabel metal2 s 183650 31200 183706 32400 6 la_data_in_core[102]
port 7 nsew signal output
rlabel metal2 s 184938 31200 184994 32400 6 la_data_in_core[103]
port 8 nsew signal output
rlabel metal2 s 186318 31200 186374 32400 6 la_data_in_core[104]
port 9 nsew signal output
rlabel metal2 s 187606 31200 187662 32400 6 la_data_in_core[105]
port 10 nsew signal output
rlabel metal2 s 188986 31200 189042 32400 6 la_data_in_core[106]
port 11 nsew signal output
rlabel metal2 s 190274 31200 190330 32400 6 la_data_in_core[107]
port 12 nsew signal output
rlabel metal2 s 191654 31200 191710 32400 6 la_data_in_core[108]
port 13 nsew signal output
rlabel metal2 s 192942 31200 192998 32400 6 la_data_in_core[109]
port 14 nsew signal output
rlabel metal2 s 60738 31200 60794 32400 6 la_data_in_core[10]
port 15 nsew signal output
rlabel metal2 s 194322 31200 194378 32400 6 la_data_in_core[110]
port 16 nsew signal output
rlabel metal2 s 195610 31200 195666 32400 6 la_data_in_core[111]
port 17 nsew signal output
rlabel metal2 s 196990 31200 197046 32400 6 la_data_in_core[112]
port 18 nsew signal output
rlabel metal2 s 198278 31200 198334 32400 6 la_data_in_core[113]
port 19 nsew signal output
rlabel metal2 s 199658 31200 199714 32400 6 la_data_in_core[114]
port 20 nsew signal output
rlabel metal2 s 200946 31200 201002 32400 6 la_data_in_core[115]
port 21 nsew signal output
rlabel metal2 s 202326 31200 202382 32400 6 la_data_in_core[116]
port 22 nsew signal output
rlabel metal2 s 203614 31200 203670 32400 6 la_data_in_core[117]
port 23 nsew signal output
rlabel metal2 s 204994 31200 205050 32400 6 la_data_in_core[118]
port 24 nsew signal output
rlabel metal2 s 206282 31200 206338 32400 6 la_data_in_core[119]
port 25 nsew signal output
rlabel metal2 s 62026 31200 62082 32400 6 la_data_in_core[11]
port 26 nsew signal output
rlabel metal2 s 207662 31200 207718 32400 6 la_data_in_core[120]
port 27 nsew signal output
rlabel metal2 s 208950 31200 209006 32400 6 la_data_in_core[121]
port 28 nsew signal output
rlabel metal2 s 210330 31200 210386 32400 6 la_data_in_core[122]
port 29 nsew signal output
rlabel metal2 s 211710 31200 211766 32400 6 la_data_in_core[123]
port 30 nsew signal output
rlabel metal2 s 212998 31200 213054 32400 6 la_data_in_core[124]
port 31 nsew signal output
rlabel metal2 s 214378 31200 214434 32400 6 la_data_in_core[125]
port 32 nsew signal output
rlabel metal2 s 215666 31200 215722 32400 6 la_data_in_core[126]
port 33 nsew signal output
rlabel metal2 s 217046 31200 217102 32400 6 la_data_in_core[127]
port 34 nsew signal output
rlabel metal2 s 63406 31200 63462 32400 6 la_data_in_core[12]
port 35 nsew signal output
rlabel metal2 s 64694 31200 64750 32400 6 la_data_in_core[13]
port 36 nsew signal output
rlabel metal2 s 66074 31200 66130 32400 6 la_data_in_core[14]
port 37 nsew signal output
rlabel metal2 s 67362 31200 67418 32400 6 la_data_in_core[15]
port 38 nsew signal output
rlabel metal2 s 68742 31200 68798 32400 6 la_data_in_core[16]
port 39 nsew signal output
rlabel metal2 s 70030 31200 70086 32400 6 la_data_in_core[17]
port 40 nsew signal output
rlabel metal2 s 71410 31200 71466 32400 6 la_data_in_core[18]
port 41 nsew signal output
rlabel metal2 s 72698 31200 72754 32400 6 la_data_in_core[19]
port 42 nsew signal output
rlabel metal2 s 48686 31200 48742 32400 6 la_data_in_core[1]
port 43 nsew signal output
rlabel metal2 s 74078 31200 74134 32400 6 la_data_in_core[20]
port 44 nsew signal output
rlabel metal2 s 75366 31200 75422 32400 6 la_data_in_core[21]
port 45 nsew signal output
rlabel metal2 s 76746 31200 76802 32400 6 la_data_in_core[22]
port 46 nsew signal output
rlabel metal2 s 78126 31200 78182 32400 6 la_data_in_core[23]
port 47 nsew signal output
rlabel metal2 s 79414 31200 79470 32400 6 la_data_in_core[24]
port 48 nsew signal output
rlabel metal2 s 80794 31200 80850 32400 6 la_data_in_core[25]
port 49 nsew signal output
rlabel metal2 s 82082 31200 82138 32400 6 la_data_in_core[26]
port 50 nsew signal output
rlabel metal2 s 83462 31200 83518 32400 6 la_data_in_core[27]
port 51 nsew signal output
rlabel metal2 s 84750 31200 84806 32400 6 la_data_in_core[28]
port 52 nsew signal output
rlabel metal2 s 86130 31200 86186 32400 6 la_data_in_core[29]
port 53 nsew signal output
rlabel metal2 s 50066 31200 50122 32400 6 la_data_in_core[2]
port 54 nsew signal output
rlabel metal2 s 87418 31200 87474 32400 6 la_data_in_core[30]
port 55 nsew signal output
rlabel metal2 s 88798 31200 88854 32400 6 la_data_in_core[31]
port 56 nsew signal output
rlabel metal2 s 90086 31200 90142 32400 6 la_data_in_core[32]
port 57 nsew signal output
rlabel metal2 s 91466 31200 91522 32400 6 la_data_in_core[33]
port 58 nsew signal output
rlabel metal2 s 92754 31200 92810 32400 6 la_data_in_core[34]
port 59 nsew signal output
rlabel metal2 s 94134 31200 94190 32400 6 la_data_in_core[35]
port 60 nsew signal output
rlabel metal2 s 95422 31200 95478 32400 6 la_data_in_core[36]
port 61 nsew signal output
rlabel metal2 s 96802 31200 96858 32400 6 la_data_in_core[37]
port 62 nsew signal output
rlabel metal2 s 98090 31200 98146 32400 6 la_data_in_core[38]
port 63 nsew signal output
rlabel metal2 s 99470 31200 99526 32400 6 la_data_in_core[39]
port 64 nsew signal output
rlabel metal2 s 51354 31200 51410 32400 6 la_data_in_core[3]
port 65 nsew signal output
rlabel metal2 s 100758 31200 100814 32400 6 la_data_in_core[40]
port 66 nsew signal output
rlabel metal2 s 102138 31200 102194 32400 6 la_data_in_core[41]
port 67 nsew signal output
rlabel metal2 s 103426 31200 103482 32400 6 la_data_in_core[42]
port 68 nsew signal output
rlabel metal2 s 104806 31200 104862 32400 6 la_data_in_core[43]
port 69 nsew signal output
rlabel metal2 s 106094 31200 106150 32400 6 la_data_in_core[44]
port 70 nsew signal output
rlabel metal2 s 107474 31200 107530 32400 6 la_data_in_core[45]
port 71 nsew signal output
rlabel metal2 s 108762 31200 108818 32400 6 la_data_in_core[46]
port 72 nsew signal output
rlabel metal2 s 110142 31200 110198 32400 6 la_data_in_core[47]
port 73 nsew signal output
rlabel metal2 s 111522 31200 111578 32400 6 la_data_in_core[48]
port 74 nsew signal output
rlabel metal2 s 112810 31200 112866 32400 6 la_data_in_core[49]
port 75 nsew signal output
rlabel metal2 s 52734 31200 52790 32400 6 la_data_in_core[4]
port 76 nsew signal output
rlabel metal2 s 114190 31200 114246 32400 6 la_data_in_core[50]
port 77 nsew signal output
rlabel metal2 s 115478 31200 115534 32400 6 la_data_in_core[51]
port 78 nsew signal output
rlabel metal2 s 116858 31200 116914 32400 6 la_data_in_core[52]
port 79 nsew signal output
rlabel metal2 s 118146 31200 118202 32400 6 la_data_in_core[53]
port 80 nsew signal output
rlabel metal2 s 119526 31200 119582 32400 6 la_data_in_core[54]
port 81 nsew signal output
rlabel metal2 s 120814 31200 120870 32400 6 la_data_in_core[55]
port 82 nsew signal output
rlabel metal2 s 122194 31200 122250 32400 6 la_data_in_core[56]
port 83 nsew signal output
rlabel metal2 s 123482 31200 123538 32400 6 la_data_in_core[57]
port 84 nsew signal output
rlabel metal2 s 124862 31200 124918 32400 6 la_data_in_core[58]
port 85 nsew signal output
rlabel metal2 s 126150 31200 126206 32400 6 la_data_in_core[59]
port 86 nsew signal output
rlabel metal2 s 54022 31200 54078 32400 6 la_data_in_core[5]
port 87 nsew signal output
rlabel metal2 s 127530 31200 127586 32400 6 la_data_in_core[60]
port 88 nsew signal output
rlabel metal2 s 128818 31200 128874 32400 6 la_data_in_core[61]
port 89 nsew signal output
rlabel metal2 s 130198 31200 130254 32400 6 la_data_in_core[62]
port 90 nsew signal output
rlabel metal2 s 131486 31200 131542 32400 6 la_data_in_core[63]
port 91 nsew signal output
rlabel metal2 s 132866 31200 132922 32400 6 la_data_in_core[64]
port 92 nsew signal output
rlabel metal2 s 134154 31200 134210 32400 6 la_data_in_core[65]
port 93 nsew signal output
rlabel metal2 s 135534 31200 135590 32400 6 la_data_in_core[66]
port 94 nsew signal output
rlabel metal2 s 136822 31200 136878 32400 6 la_data_in_core[67]
port 95 nsew signal output
rlabel metal2 s 138202 31200 138258 32400 6 la_data_in_core[68]
port 96 nsew signal output
rlabel metal2 s 139490 31200 139546 32400 6 la_data_in_core[69]
port 97 nsew signal output
rlabel metal2 s 55402 31200 55458 32400 6 la_data_in_core[6]
port 98 nsew signal output
rlabel metal2 s 140870 31200 140926 32400 6 la_data_in_core[70]
port 99 nsew signal output
rlabel metal2 s 142158 31200 142214 32400 6 la_data_in_core[71]
port 100 nsew signal output
rlabel metal2 s 143538 31200 143594 32400 6 la_data_in_core[72]
port 101 nsew signal output
rlabel metal2 s 144918 31200 144974 32400 6 la_data_in_core[73]
port 102 nsew signal output
rlabel metal2 s 146206 31200 146262 32400 6 la_data_in_core[74]
port 103 nsew signal output
rlabel metal2 s 147586 31200 147642 32400 6 la_data_in_core[75]
port 104 nsew signal output
rlabel metal2 s 148874 31200 148930 32400 6 la_data_in_core[76]
port 105 nsew signal output
rlabel metal2 s 150254 31200 150310 32400 6 la_data_in_core[77]
port 106 nsew signal output
rlabel metal2 s 151542 31200 151598 32400 6 la_data_in_core[78]
port 107 nsew signal output
rlabel metal2 s 152922 31200 152978 32400 6 la_data_in_core[79]
port 108 nsew signal output
rlabel metal2 s 56690 31200 56746 32400 6 la_data_in_core[7]
port 109 nsew signal output
rlabel metal2 s 154210 31200 154266 32400 6 la_data_in_core[80]
port 110 nsew signal output
rlabel metal2 s 155590 31200 155646 32400 6 la_data_in_core[81]
port 111 nsew signal output
rlabel metal2 s 156878 31200 156934 32400 6 la_data_in_core[82]
port 112 nsew signal output
rlabel metal2 s 158258 31200 158314 32400 6 la_data_in_core[83]
port 113 nsew signal output
rlabel metal2 s 159546 31200 159602 32400 6 la_data_in_core[84]
port 114 nsew signal output
rlabel metal2 s 160926 31200 160982 32400 6 la_data_in_core[85]
port 115 nsew signal output
rlabel metal2 s 162214 31200 162270 32400 6 la_data_in_core[86]
port 116 nsew signal output
rlabel metal2 s 163594 31200 163650 32400 6 la_data_in_core[87]
port 117 nsew signal output
rlabel metal2 s 164882 31200 164938 32400 6 la_data_in_core[88]
port 118 nsew signal output
rlabel metal2 s 166262 31200 166318 32400 6 la_data_in_core[89]
port 119 nsew signal output
rlabel metal2 s 58070 31200 58126 32400 6 la_data_in_core[8]
port 120 nsew signal output
rlabel metal2 s 167550 31200 167606 32400 6 la_data_in_core[90]
port 121 nsew signal output
rlabel metal2 s 168930 31200 168986 32400 6 la_data_in_core[91]
port 122 nsew signal output
rlabel metal2 s 170218 31200 170274 32400 6 la_data_in_core[92]
port 123 nsew signal output
rlabel metal2 s 171598 31200 171654 32400 6 la_data_in_core[93]
port 124 nsew signal output
rlabel metal2 s 172886 31200 172942 32400 6 la_data_in_core[94]
port 125 nsew signal output
rlabel metal2 s 174266 31200 174322 32400 6 la_data_in_core[95]
port 126 nsew signal output
rlabel metal2 s 175554 31200 175610 32400 6 la_data_in_core[96]
port 127 nsew signal output
rlabel metal2 s 176934 31200 176990 32400 6 la_data_in_core[97]
port 128 nsew signal output
rlabel metal2 s 178314 31200 178370 32400 6 la_data_in_core[98]
port 129 nsew signal output
rlabel metal2 s 179602 31200 179658 32400 6 la_data_in_core[99]
port 130 nsew signal output
rlabel metal2 s 59358 31200 59414 32400 6 la_data_in_core[9]
port 131 nsew signal output
rlabel metal2 s 110 -400 166 800 6 la_data_in_mprj[0]
port 132 nsew signal output
rlabel metal2 s 142710 -400 142766 800 6 la_data_in_mprj[100]
port 133 nsew signal output
rlabel metal2 s 144090 -400 144146 800 6 la_data_in_mprj[101]
port 134 nsew signal output
rlabel metal2 s 145562 -400 145618 800 6 la_data_in_mprj[102]
port 135 nsew signal output
rlabel metal2 s 146942 -400 146998 800 6 la_data_in_mprj[103]
port 136 nsew signal output
rlabel metal2 s 148414 -400 148470 800 6 la_data_in_mprj[104]
port 137 nsew signal output
rlabel metal2 s 149794 -400 149850 800 6 la_data_in_mprj[105]
port 138 nsew signal output
rlabel metal2 s 151266 -400 151322 800 6 la_data_in_mprj[106]
port 139 nsew signal output
rlabel metal2 s 152646 -400 152702 800 6 la_data_in_mprj[107]
port 140 nsew signal output
rlabel metal2 s 154118 -400 154174 800 6 la_data_in_mprj[108]
port 141 nsew signal output
rlabel metal2 s 155498 -400 155554 800 6 la_data_in_mprj[109]
port 142 nsew signal output
rlabel metal2 s 14370 -400 14426 800 6 la_data_in_mprj[10]
port 143 nsew signal output
rlabel metal2 s 156970 -400 157026 800 6 la_data_in_mprj[110]
port 144 nsew signal output
rlabel metal2 s 158350 -400 158406 800 6 la_data_in_mprj[111]
port 145 nsew signal output
rlabel metal2 s 159822 -400 159878 800 6 la_data_in_mprj[112]
port 146 nsew signal output
rlabel metal2 s 161202 -400 161258 800 6 la_data_in_mprj[113]
port 147 nsew signal output
rlabel metal2 s 162674 -400 162730 800 6 la_data_in_mprj[114]
port 148 nsew signal output
rlabel metal2 s 164054 -400 164110 800 6 la_data_in_mprj[115]
port 149 nsew signal output
rlabel metal2 s 165526 -400 165582 800 6 la_data_in_mprj[116]
port 150 nsew signal output
rlabel metal2 s 166906 -400 166962 800 6 la_data_in_mprj[117]
port 151 nsew signal output
rlabel metal2 s 168378 -400 168434 800 6 la_data_in_mprj[118]
port 152 nsew signal output
rlabel metal2 s 169758 -400 169814 800 6 la_data_in_mprj[119]
port 153 nsew signal output
rlabel metal2 s 15750 -400 15806 800 6 la_data_in_mprj[11]
port 154 nsew signal output
rlabel metal2 s 171230 -400 171286 800 6 la_data_in_mprj[120]
port 155 nsew signal output
rlabel metal2 s 172610 -400 172666 800 6 la_data_in_mprj[121]
port 156 nsew signal output
rlabel metal2 s 174082 -400 174138 800 6 la_data_in_mprj[122]
port 157 nsew signal output
rlabel metal2 s 175462 -400 175518 800 6 la_data_in_mprj[123]
port 158 nsew signal output
rlabel metal2 s 176934 -400 176990 800 6 la_data_in_mprj[124]
port 159 nsew signal output
rlabel metal2 s 178314 -400 178370 800 6 la_data_in_mprj[125]
port 160 nsew signal output
rlabel metal2 s 179786 -400 179842 800 6 la_data_in_mprj[126]
port 161 nsew signal output
rlabel metal2 s 181166 -400 181222 800 6 la_data_in_mprj[127]
port 162 nsew signal output
rlabel metal2 s 17222 -400 17278 800 6 la_data_in_mprj[12]
port 163 nsew signal output
rlabel metal2 s 18602 -400 18658 800 6 la_data_in_mprj[13]
port 164 nsew signal output
rlabel metal2 s 20074 -400 20130 800 6 la_data_in_mprj[14]
port 165 nsew signal output
rlabel metal2 s 21454 -400 21510 800 6 la_data_in_mprj[15]
port 166 nsew signal output
rlabel metal2 s 22926 -400 22982 800 6 la_data_in_mprj[16]
port 167 nsew signal output
rlabel metal2 s 24306 -400 24362 800 6 la_data_in_mprj[17]
port 168 nsew signal output
rlabel metal2 s 25778 -400 25834 800 6 la_data_in_mprj[18]
port 169 nsew signal output
rlabel metal2 s 27158 -400 27214 800 6 la_data_in_mprj[19]
port 170 nsew signal output
rlabel metal2 s 1490 -400 1546 800 6 la_data_in_mprj[1]
port 171 nsew signal output
rlabel metal2 s 28630 -400 28686 800 6 la_data_in_mprj[20]
port 172 nsew signal output
rlabel metal2 s 30010 -400 30066 800 6 la_data_in_mprj[21]
port 173 nsew signal output
rlabel metal2 s 31482 -400 31538 800 6 la_data_in_mprj[22]
port 174 nsew signal output
rlabel metal2 s 32862 -400 32918 800 6 la_data_in_mprj[23]
port 175 nsew signal output
rlabel metal2 s 34334 -400 34390 800 6 la_data_in_mprj[24]
port 176 nsew signal output
rlabel metal2 s 35714 -400 35770 800 6 la_data_in_mprj[25]
port 177 nsew signal output
rlabel metal2 s 37186 -400 37242 800 6 la_data_in_mprj[26]
port 178 nsew signal output
rlabel metal2 s 38566 -400 38622 800 6 la_data_in_mprj[27]
port 179 nsew signal output
rlabel metal2 s 40038 -400 40094 800 6 la_data_in_mprj[28]
port 180 nsew signal output
rlabel metal2 s 41418 -400 41474 800 6 la_data_in_mprj[29]
port 181 nsew signal output
rlabel metal2 s 2962 -400 3018 800 6 la_data_in_mprj[2]
port 182 nsew signal output
rlabel metal2 s 42890 -400 42946 800 6 la_data_in_mprj[30]
port 183 nsew signal output
rlabel metal2 s 44270 -400 44326 800 6 la_data_in_mprj[31]
port 184 nsew signal output
rlabel metal2 s 45742 -400 45798 800 6 la_data_in_mprj[32]
port 185 nsew signal output
rlabel metal2 s 47122 -400 47178 800 6 la_data_in_mprj[33]
port 186 nsew signal output
rlabel metal2 s 48594 -400 48650 800 6 la_data_in_mprj[34]
port 187 nsew signal output
rlabel metal2 s 49974 -400 50030 800 6 la_data_in_mprj[35]
port 188 nsew signal output
rlabel metal2 s 51446 -400 51502 800 6 la_data_in_mprj[36]
port 189 nsew signal output
rlabel metal2 s 52826 -400 52882 800 6 la_data_in_mprj[37]
port 190 nsew signal output
rlabel metal2 s 54298 -400 54354 800 6 la_data_in_mprj[38]
port 191 nsew signal output
rlabel metal2 s 55678 -400 55734 800 6 la_data_in_mprj[39]
port 192 nsew signal output
rlabel metal2 s 4342 -400 4398 800 6 la_data_in_mprj[3]
port 193 nsew signal output
rlabel metal2 s 57150 -400 57206 800 6 la_data_in_mprj[40]
port 194 nsew signal output
rlabel metal2 s 58530 -400 58586 800 6 la_data_in_mprj[41]
port 195 nsew signal output
rlabel metal2 s 60002 -400 60058 800 6 la_data_in_mprj[42]
port 196 nsew signal output
rlabel metal2 s 61382 -400 61438 800 6 la_data_in_mprj[43]
port 197 nsew signal output
rlabel metal2 s 62854 -400 62910 800 6 la_data_in_mprj[44]
port 198 nsew signal output
rlabel metal2 s 64234 -400 64290 800 6 la_data_in_mprj[45]
port 199 nsew signal output
rlabel metal2 s 65706 -400 65762 800 6 la_data_in_mprj[46]
port 200 nsew signal output
rlabel metal2 s 67086 -400 67142 800 6 la_data_in_mprj[47]
port 201 nsew signal output
rlabel metal2 s 68558 -400 68614 800 6 la_data_in_mprj[48]
port 202 nsew signal output
rlabel metal2 s 69938 -400 69994 800 6 la_data_in_mprj[49]
port 203 nsew signal output
rlabel metal2 s 5814 -400 5870 800 6 la_data_in_mprj[4]
port 204 nsew signal output
rlabel metal2 s 71410 -400 71466 800 6 la_data_in_mprj[50]
port 205 nsew signal output
rlabel metal2 s 72790 -400 72846 800 6 la_data_in_mprj[51]
port 206 nsew signal output
rlabel metal2 s 74262 -400 74318 800 6 la_data_in_mprj[52]
port 207 nsew signal output
rlabel metal2 s 75642 -400 75698 800 6 la_data_in_mprj[53]
port 208 nsew signal output
rlabel metal2 s 77114 -400 77170 800 6 la_data_in_mprj[54]
port 209 nsew signal output
rlabel metal2 s 78494 -400 78550 800 6 la_data_in_mprj[55]
port 210 nsew signal output
rlabel metal2 s 79966 -400 80022 800 6 la_data_in_mprj[56]
port 211 nsew signal output
rlabel metal2 s 81346 -400 81402 800 6 la_data_in_mprj[57]
port 212 nsew signal output
rlabel metal2 s 82818 -400 82874 800 6 la_data_in_mprj[58]
port 213 nsew signal output
rlabel metal2 s 84198 -400 84254 800 6 la_data_in_mprj[59]
port 214 nsew signal output
rlabel metal2 s 7194 -400 7250 800 6 la_data_in_mprj[5]
port 215 nsew signal output
rlabel metal2 s 85670 -400 85726 800 6 la_data_in_mprj[60]
port 216 nsew signal output
rlabel metal2 s 87050 -400 87106 800 6 la_data_in_mprj[61]
port 217 nsew signal output
rlabel metal2 s 88522 -400 88578 800 6 la_data_in_mprj[62]
port 218 nsew signal output
rlabel metal2 s 89902 -400 89958 800 6 la_data_in_mprj[63]
port 219 nsew signal output
rlabel metal2 s 91374 -400 91430 800 6 la_data_in_mprj[64]
port 220 nsew signal output
rlabel metal2 s 92754 -400 92810 800 6 la_data_in_mprj[65]
port 221 nsew signal output
rlabel metal2 s 94226 -400 94282 800 6 la_data_in_mprj[66]
port 222 nsew signal output
rlabel metal2 s 95606 -400 95662 800 6 la_data_in_mprj[67]
port 223 nsew signal output
rlabel metal2 s 97078 -400 97134 800 6 la_data_in_mprj[68]
port 224 nsew signal output
rlabel metal2 s 98458 -400 98514 800 6 la_data_in_mprj[69]
port 225 nsew signal output
rlabel metal2 s 8666 -400 8722 800 6 la_data_in_mprj[6]
port 226 nsew signal output
rlabel metal2 s 99930 -400 99986 800 6 la_data_in_mprj[70]
port 227 nsew signal output
rlabel metal2 s 101310 -400 101366 800 6 la_data_in_mprj[71]
port 228 nsew signal output
rlabel metal2 s 102782 -400 102838 800 6 la_data_in_mprj[72]
port 229 nsew signal output
rlabel metal2 s 104162 -400 104218 800 6 la_data_in_mprj[73]
port 230 nsew signal output
rlabel metal2 s 105634 -400 105690 800 6 la_data_in_mprj[74]
port 231 nsew signal output
rlabel metal2 s 107014 -400 107070 800 6 la_data_in_mprj[75]
port 232 nsew signal output
rlabel metal2 s 108486 -400 108542 800 6 la_data_in_mprj[76]
port 233 nsew signal output
rlabel metal2 s 109866 -400 109922 800 6 la_data_in_mprj[77]
port 234 nsew signal output
rlabel metal2 s 111338 -400 111394 800 6 la_data_in_mprj[78]
port 235 nsew signal output
rlabel metal2 s 112718 -400 112774 800 6 la_data_in_mprj[79]
port 236 nsew signal output
rlabel metal2 s 10046 -400 10102 800 6 la_data_in_mprj[7]
port 237 nsew signal output
rlabel metal2 s 114190 -400 114246 800 6 la_data_in_mprj[80]
port 238 nsew signal output
rlabel metal2 s 115570 -400 115626 800 6 la_data_in_mprj[81]
port 239 nsew signal output
rlabel metal2 s 117042 -400 117098 800 6 la_data_in_mprj[82]
port 240 nsew signal output
rlabel metal2 s 118422 -400 118478 800 6 la_data_in_mprj[83]
port 241 nsew signal output
rlabel metal2 s 119894 -400 119950 800 6 la_data_in_mprj[84]
port 242 nsew signal output
rlabel metal2 s 121274 -400 121330 800 6 la_data_in_mprj[85]
port 243 nsew signal output
rlabel metal2 s 122746 -400 122802 800 6 la_data_in_mprj[86]
port 244 nsew signal output
rlabel metal2 s 124126 -400 124182 800 6 la_data_in_mprj[87]
port 245 nsew signal output
rlabel metal2 s 125598 -400 125654 800 6 la_data_in_mprj[88]
port 246 nsew signal output
rlabel metal2 s 126978 -400 127034 800 6 la_data_in_mprj[89]
port 247 nsew signal output
rlabel metal2 s 11518 -400 11574 800 6 la_data_in_mprj[8]
port 248 nsew signal output
rlabel metal2 s 128450 -400 128506 800 6 la_data_in_mprj[90]
port 249 nsew signal output
rlabel metal2 s 129830 -400 129886 800 6 la_data_in_mprj[91]
port 250 nsew signal output
rlabel metal2 s 131302 -400 131358 800 6 la_data_in_mprj[92]
port 251 nsew signal output
rlabel metal2 s 132682 -400 132738 800 6 la_data_in_mprj[93]
port 252 nsew signal output
rlabel metal2 s 134154 -400 134210 800 6 la_data_in_mprj[94]
port 253 nsew signal output
rlabel metal2 s 135534 -400 135590 800 6 la_data_in_mprj[95]
port 254 nsew signal output
rlabel metal2 s 137006 -400 137062 800 6 la_data_in_mprj[96]
port 255 nsew signal output
rlabel metal2 s 138386 -400 138442 800 6 la_data_in_mprj[97]
port 256 nsew signal output
rlabel metal2 s 139858 -400 139914 800 6 la_data_in_mprj[98]
port 257 nsew signal output
rlabel metal2 s 141238 -400 141294 800 6 la_data_in_mprj[99]
port 258 nsew signal output
rlabel metal2 s 12898 -400 12954 800 6 la_data_in_mprj[9]
port 259 nsew signal output
rlabel metal2 s 47766 31200 47822 32400 6 la_data_out_core[0]
port 260 nsew signal input
rlabel metal2 s 181350 31200 181406 32400 6 la_data_out_core[100]
port 261 nsew signal input
rlabel metal2 s 182730 31200 182786 32400 6 la_data_out_core[101]
port 262 nsew signal input
rlabel metal2 s 184018 31200 184074 32400 6 la_data_out_core[102]
port 263 nsew signal input
rlabel metal2 s 185398 31200 185454 32400 6 la_data_out_core[103]
port 264 nsew signal input
rlabel metal2 s 186686 31200 186742 32400 6 la_data_out_core[104]
port 265 nsew signal input
rlabel metal2 s 188066 31200 188122 32400 6 la_data_out_core[105]
port 266 nsew signal input
rlabel metal2 s 189446 31200 189502 32400 6 la_data_out_core[106]
port 267 nsew signal input
rlabel metal2 s 190734 31200 190790 32400 6 la_data_out_core[107]
port 268 nsew signal input
rlabel metal2 s 192114 31200 192170 32400 6 la_data_out_core[108]
port 269 nsew signal input
rlabel metal2 s 193402 31200 193458 32400 6 la_data_out_core[109]
port 270 nsew signal input
rlabel metal2 s 61198 31200 61254 32400 6 la_data_out_core[10]
port 271 nsew signal input
rlabel metal2 s 194782 31200 194838 32400 6 la_data_out_core[110]
port 272 nsew signal input
rlabel metal2 s 196070 31200 196126 32400 6 la_data_out_core[111]
port 273 nsew signal input
rlabel metal2 s 197450 31200 197506 32400 6 la_data_out_core[112]
port 274 nsew signal input
rlabel metal2 s 198738 31200 198794 32400 6 la_data_out_core[113]
port 275 nsew signal input
rlabel metal2 s 200118 31200 200174 32400 6 la_data_out_core[114]
port 276 nsew signal input
rlabel metal2 s 201406 31200 201462 32400 6 la_data_out_core[115]
port 277 nsew signal input
rlabel metal2 s 202786 31200 202842 32400 6 la_data_out_core[116]
port 278 nsew signal input
rlabel metal2 s 204074 31200 204130 32400 6 la_data_out_core[117]
port 279 nsew signal input
rlabel metal2 s 205454 31200 205510 32400 6 la_data_out_core[118]
port 280 nsew signal input
rlabel metal2 s 206742 31200 206798 32400 6 la_data_out_core[119]
port 281 nsew signal input
rlabel metal2 s 62486 31200 62542 32400 6 la_data_out_core[11]
port 282 nsew signal input
rlabel metal2 s 208122 31200 208178 32400 6 la_data_out_core[120]
port 283 nsew signal input
rlabel metal2 s 209410 31200 209466 32400 6 la_data_out_core[121]
port 284 nsew signal input
rlabel metal2 s 210790 31200 210846 32400 6 la_data_out_core[122]
port 285 nsew signal input
rlabel metal2 s 212078 31200 212134 32400 6 la_data_out_core[123]
port 286 nsew signal input
rlabel metal2 s 213458 31200 213514 32400 6 la_data_out_core[124]
port 287 nsew signal input
rlabel metal2 s 214746 31200 214802 32400 6 la_data_out_core[125]
port 288 nsew signal input
rlabel metal2 s 216126 31200 216182 32400 6 la_data_out_core[126]
port 289 nsew signal input
rlabel metal2 s 217414 31200 217470 32400 6 la_data_out_core[127]
port 290 nsew signal input
rlabel metal2 s 63866 31200 63922 32400 6 la_data_out_core[12]
port 291 nsew signal input
rlabel metal2 s 65154 31200 65210 32400 6 la_data_out_core[13]
port 292 nsew signal input
rlabel metal2 s 66534 31200 66590 32400 6 la_data_out_core[14]
port 293 nsew signal input
rlabel metal2 s 67822 31200 67878 32400 6 la_data_out_core[15]
port 294 nsew signal input
rlabel metal2 s 69202 31200 69258 32400 6 la_data_out_core[16]
port 295 nsew signal input
rlabel metal2 s 70490 31200 70546 32400 6 la_data_out_core[17]
port 296 nsew signal input
rlabel metal2 s 71870 31200 71926 32400 6 la_data_out_core[18]
port 297 nsew signal input
rlabel metal2 s 73158 31200 73214 32400 6 la_data_out_core[19]
port 298 nsew signal input
rlabel metal2 s 49146 31200 49202 32400 6 la_data_out_core[1]
port 299 nsew signal input
rlabel metal2 s 74538 31200 74594 32400 6 la_data_out_core[20]
port 300 nsew signal input
rlabel metal2 s 75826 31200 75882 32400 6 la_data_out_core[21]
port 301 nsew signal input
rlabel metal2 s 77206 31200 77262 32400 6 la_data_out_core[22]
port 302 nsew signal input
rlabel metal2 s 78494 31200 78550 32400 6 la_data_out_core[23]
port 303 nsew signal input
rlabel metal2 s 79874 31200 79930 32400 6 la_data_out_core[24]
port 304 nsew signal input
rlabel metal2 s 81162 31200 81218 32400 6 la_data_out_core[25]
port 305 nsew signal input
rlabel metal2 s 82542 31200 82598 32400 6 la_data_out_core[26]
port 306 nsew signal input
rlabel metal2 s 83830 31200 83886 32400 6 la_data_out_core[27]
port 307 nsew signal input
rlabel metal2 s 85210 31200 85266 32400 6 la_data_out_core[28]
port 308 nsew signal input
rlabel metal2 s 86498 31200 86554 32400 6 la_data_out_core[29]
port 309 nsew signal input
rlabel metal2 s 50434 31200 50490 32400 6 la_data_out_core[2]
port 310 nsew signal input
rlabel metal2 s 87878 31200 87934 32400 6 la_data_out_core[30]
port 311 nsew signal input
rlabel metal2 s 89258 31200 89314 32400 6 la_data_out_core[31]
port 312 nsew signal input
rlabel metal2 s 90546 31200 90602 32400 6 la_data_out_core[32]
port 313 nsew signal input
rlabel metal2 s 91926 31200 91982 32400 6 la_data_out_core[33]
port 314 nsew signal input
rlabel metal2 s 93214 31200 93270 32400 6 la_data_out_core[34]
port 315 nsew signal input
rlabel metal2 s 94594 31200 94650 32400 6 la_data_out_core[35]
port 316 nsew signal input
rlabel metal2 s 95882 31200 95938 32400 6 la_data_out_core[36]
port 317 nsew signal input
rlabel metal2 s 97262 31200 97318 32400 6 la_data_out_core[37]
port 318 nsew signal input
rlabel metal2 s 98550 31200 98606 32400 6 la_data_out_core[38]
port 319 nsew signal input
rlabel metal2 s 99930 31200 99986 32400 6 la_data_out_core[39]
port 320 nsew signal input
rlabel metal2 s 51814 31200 51870 32400 6 la_data_out_core[3]
port 321 nsew signal input
rlabel metal2 s 101218 31200 101274 32400 6 la_data_out_core[40]
port 322 nsew signal input
rlabel metal2 s 102598 31200 102654 32400 6 la_data_out_core[41]
port 323 nsew signal input
rlabel metal2 s 103886 31200 103942 32400 6 la_data_out_core[42]
port 324 nsew signal input
rlabel metal2 s 105266 31200 105322 32400 6 la_data_out_core[43]
port 325 nsew signal input
rlabel metal2 s 106554 31200 106610 32400 6 la_data_out_core[44]
port 326 nsew signal input
rlabel metal2 s 107934 31200 107990 32400 6 la_data_out_core[45]
port 327 nsew signal input
rlabel metal2 s 109222 31200 109278 32400 6 la_data_out_core[46]
port 328 nsew signal input
rlabel metal2 s 110602 31200 110658 32400 6 la_data_out_core[47]
port 329 nsew signal input
rlabel metal2 s 111890 31200 111946 32400 6 la_data_out_core[48]
port 330 nsew signal input
rlabel metal2 s 113270 31200 113326 32400 6 la_data_out_core[49]
port 331 nsew signal input
rlabel metal2 s 53102 31200 53158 32400 6 la_data_out_core[4]
port 332 nsew signal input
rlabel metal2 s 114558 31200 114614 32400 6 la_data_out_core[50]
port 333 nsew signal input
rlabel metal2 s 115938 31200 115994 32400 6 la_data_out_core[51]
port 334 nsew signal input
rlabel metal2 s 117226 31200 117282 32400 6 la_data_out_core[52]
port 335 nsew signal input
rlabel metal2 s 118606 31200 118662 32400 6 la_data_out_core[53]
port 336 nsew signal input
rlabel metal2 s 119894 31200 119950 32400 6 la_data_out_core[54]
port 337 nsew signal input
rlabel metal2 s 121274 31200 121330 32400 6 la_data_out_core[55]
port 338 nsew signal input
rlabel metal2 s 122654 31200 122710 32400 6 la_data_out_core[56]
port 339 nsew signal input
rlabel metal2 s 123942 31200 123998 32400 6 la_data_out_core[57]
port 340 nsew signal input
rlabel metal2 s 125322 31200 125378 32400 6 la_data_out_core[58]
port 341 nsew signal input
rlabel metal2 s 126610 31200 126666 32400 6 la_data_out_core[59]
port 342 nsew signal input
rlabel metal2 s 54482 31200 54538 32400 6 la_data_out_core[5]
port 343 nsew signal input
rlabel metal2 s 127990 31200 128046 32400 6 la_data_out_core[60]
port 344 nsew signal input
rlabel metal2 s 129278 31200 129334 32400 6 la_data_out_core[61]
port 345 nsew signal input
rlabel metal2 s 130658 31200 130714 32400 6 la_data_out_core[62]
port 346 nsew signal input
rlabel metal2 s 131946 31200 132002 32400 6 la_data_out_core[63]
port 347 nsew signal input
rlabel metal2 s 133326 31200 133382 32400 6 la_data_out_core[64]
port 348 nsew signal input
rlabel metal2 s 134614 31200 134670 32400 6 la_data_out_core[65]
port 349 nsew signal input
rlabel metal2 s 135994 31200 136050 32400 6 la_data_out_core[66]
port 350 nsew signal input
rlabel metal2 s 137282 31200 137338 32400 6 la_data_out_core[67]
port 351 nsew signal input
rlabel metal2 s 138662 31200 138718 32400 6 la_data_out_core[68]
port 352 nsew signal input
rlabel metal2 s 139950 31200 140006 32400 6 la_data_out_core[69]
port 353 nsew signal input
rlabel metal2 s 55862 31200 55918 32400 6 la_data_out_core[6]
port 354 nsew signal input
rlabel metal2 s 141330 31200 141386 32400 6 la_data_out_core[70]
port 355 nsew signal input
rlabel metal2 s 142618 31200 142674 32400 6 la_data_out_core[71]
port 356 nsew signal input
rlabel metal2 s 143998 31200 144054 32400 6 la_data_out_core[72]
port 357 nsew signal input
rlabel metal2 s 145286 31200 145342 32400 6 la_data_out_core[73]
port 358 nsew signal input
rlabel metal2 s 146666 31200 146722 32400 6 la_data_out_core[74]
port 359 nsew signal input
rlabel metal2 s 147954 31200 148010 32400 6 la_data_out_core[75]
port 360 nsew signal input
rlabel metal2 s 149334 31200 149390 32400 6 la_data_out_core[76]
port 361 nsew signal input
rlabel metal2 s 150622 31200 150678 32400 6 la_data_out_core[77]
port 362 nsew signal input
rlabel metal2 s 152002 31200 152058 32400 6 la_data_out_core[78]
port 363 nsew signal input
rlabel metal2 s 153290 31200 153346 32400 6 la_data_out_core[79]
port 364 nsew signal input
rlabel metal2 s 57150 31200 57206 32400 6 la_data_out_core[7]
port 365 nsew signal input
rlabel metal2 s 154670 31200 154726 32400 6 la_data_out_core[80]
port 366 nsew signal input
rlabel metal2 s 156050 31200 156106 32400 6 la_data_out_core[81]
port 367 nsew signal input
rlabel metal2 s 157338 31200 157394 32400 6 la_data_out_core[82]
port 368 nsew signal input
rlabel metal2 s 158718 31200 158774 32400 6 la_data_out_core[83]
port 369 nsew signal input
rlabel metal2 s 160006 31200 160062 32400 6 la_data_out_core[84]
port 370 nsew signal input
rlabel metal2 s 161386 31200 161442 32400 6 la_data_out_core[85]
port 371 nsew signal input
rlabel metal2 s 162674 31200 162730 32400 6 la_data_out_core[86]
port 372 nsew signal input
rlabel metal2 s 164054 31200 164110 32400 6 la_data_out_core[87]
port 373 nsew signal input
rlabel metal2 s 165342 31200 165398 32400 6 la_data_out_core[88]
port 374 nsew signal input
rlabel metal2 s 166722 31200 166778 32400 6 la_data_out_core[89]
port 375 nsew signal input
rlabel metal2 s 58530 31200 58586 32400 6 la_data_out_core[8]
port 376 nsew signal input
rlabel metal2 s 168010 31200 168066 32400 6 la_data_out_core[90]
port 377 nsew signal input
rlabel metal2 s 169390 31200 169446 32400 6 la_data_out_core[91]
port 378 nsew signal input
rlabel metal2 s 170678 31200 170734 32400 6 la_data_out_core[92]
port 379 nsew signal input
rlabel metal2 s 172058 31200 172114 32400 6 la_data_out_core[93]
port 380 nsew signal input
rlabel metal2 s 173346 31200 173402 32400 6 la_data_out_core[94]
port 381 nsew signal input
rlabel metal2 s 174726 31200 174782 32400 6 la_data_out_core[95]
port 382 nsew signal input
rlabel metal2 s 176014 31200 176070 32400 6 la_data_out_core[96]
port 383 nsew signal input
rlabel metal2 s 177394 31200 177450 32400 6 la_data_out_core[97]
port 384 nsew signal input
rlabel metal2 s 178682 31200 178738 32400 6 la_data_out_core[98]
port 385 nsew signal input
rlabel metal2 s 180062 31200 180118 32400 6 la_data_out_core[99]
port 386 nsew signal input
rlabel metal2 s 59818 31200 59874 32400 6 la_data_out_core[9]
port 387 nsew signal input
rlabel metal2 s 386 -400 442 800 6 la_data_out_mprj[0]
port 388 nsew signal input
rlabel metal2 s 142986 -400 143042 800 6 la_data_out_mprj[100]
port 389 nsew signal input
rlabel metal2 s 144458 -400 144514 800 6 la_data_out_mprj[101]
port 390 nsew signal input
rlabel metal2 s 145838 -400 145894 800 6 la_data_out_mprj[102]
port 391 nsew signal input
rlabel metal2 s 147310 -400 147366 800 6 la_data_out_mprj[103]
port 392 nsew signal input
rlabel metal2 s 148690 -400 148746 800 6 la_data_out_mprj[104]
port 393 nsew signal input
rlabel metal2 s 150162 -400 150218 800 6 la_data_out_mprj[105]
port 394 nsew signal input
rlabel metal2 s 151542 -400 151598 800 6 la_data_out_mprj[106]
port 395 nsew signal input
rlabel metal2 s 153014 -400 153070 800 6 la_data_out_mprj[107]
port 396 nsew signal input
rlabel metal2 s 154394 -400 154450 800 6 la_data_out_mprj[108]
port 397 nsew signal input
rlabel metal2 s 155866 -400 155922 800 6 la_data_out_mprj[109]
port 398 nsew signal input
rlabel metal2 s 14646 -400 14702 800 6 la_data_out_mprj[10]
port 399 nsew signal input
rlabel metal2 s 157246 -400 157302 800 6 la_data_out_mprj[110]
port 400 nsew signal input
rlabel metal2 s 158718 -400 158774 800 6 la_data_out_mprj[111]
port 401 nsew signal input
rlabel metal2 s 160098 -400 160154 800 6 la_data_out_mprj[112]
port 402 nsew signal input
rlabel metal2 s 161570 -400 161626 800 6 la_data_out_mprj[113]
port 403 nsew signal input
rlabel metal2 s 162950 -400 163006 800 6 la_data_out_mprj[114]
port 404 nsew signal input
rlabel metal2 s 164422 -400 164478 800 6 la_data_out_mprj[115]
port 405 nsew signal input
rlabel metal2 s 165802 -400 165858 800 6 la_data_out_mprj[116]
port 406 nsew signal input
rlabel metal2 s 167274 -400 167330 800 6 la_data_out_mprj[117]
port 407 nsew signal input
rlabel metal2 s 168654 -400 168710 800 6 la_data_out_mprj[118]
port 408 nsew signal input
rlabel metal2 s 170126 -400 170182 800 6 la_data_out_mprj[119]
port 409 nsew signal input
rlabel metal2 s 16118 -400 16174 800 6 la_data_out_mprj[11]
port 410 nsew signal input
rlabel metal2 s 171506 -400 171562 800 6 la_data_out_mprj[120]
port 411 nsew signal input
rlabel metal2 s 172978 -400 173034 800 6 la_data_out_mprj[121]
port 412 nsew signal input
rlabel metal2 s 174358 -400 174414 800 6 la_data_out_mprj[122]
port 413 nsew signal input
rlabel metal2 s 175830 -400 175886 800 6 la_data_out_mprj[123]
port 414 nsew signal input
rlabel metal2 s 177210 -400 177266 800 6 la_data_out_mprj[124]
port 415 nsew signal input
rlabel metal2 s 178682 -400 178738 800 6 la_data_out_mprj[125]
port 416 nsew signal input
rlabel metal2 s 180062 -400 180118 800 6 la_data_out_mprj[126]
port 417 nsew signal input
rlabel metal2 s 181534 -400 181590 800 6 la_data_out_mprj[127]
port 418 nsew signal input
rlabel metal2 s 17498 -400 17554 800 6 la_data_out_mprj[12]
port 419 nsew signal input
rlabel metal2 s 18970 -400 19026 800 6 la_data_out_mprj[13]
port 420 nsew signal input
rlabel metal2 s 20350 -400 20406 800 6 la_data_out_mprj[14]
port 421 nsew signal input
rlabel metal2 s 21822 -400 21878 800 6 la_data_out_mprj[15]
port 422 nsew signal input
rlabel metal2 s 23202 -400 23258 800 6 la_data_out_mprj[16]
port 423 nsew signal input
rlabel metal2 s 24674 -400 24730 800 6 la_data_out_mprj[17]
port 424 nsew signal input
rlabel metal2 s 26054 -400 26110 800 6 la_data_out_mprj[18]
port 425 nsew signal input
rlabel metal2 s 27526 -400 27582 800 6 la_data_out_mprj[19]
port 426 nsew signal input
rlabel metal2 s 1858 -400 1914 800 6 la_data_out_mprj[1]
port 427 nsew signal input
rlabel metal2 s 28906 -400 28962 800 6 la_data_out_mprj[20]
port 428 nsew signal input
rlabel metal2 s 30378 -400 30434 800 6 la_data_out_mprj[21]
port 429 nsew signal input
rlabel metal2 s 31758 -400 31814 800 6 la_data_out_mprj[22]
port 430 nsew signal input
rlabel metal2 s 33230 -400 33286 800 6 la_data_out_mprj[23]
port 431 nsew signal input
rlabel metal2 s 34610 -400 34666 800 6 la_data_out_mprj[24]
port 432 nsew signal input
rlabel metal2 s 36082 -400 36138 800 6 la_data_out_mprj[25]
port 433 nsew signal input
rlabel metal2 s 37462 -400 37518 800 6 la_data_out_mprj[26]
port 434 nsew signal input
rlabel metal2 s 38934 -400 38990 800 6 la_data_out_mprj[27]
port 435 nsew signal input
rlabel metal2 s 40314 -400 40370 800 6 la_data_out_mprj[28]
port 436 nsew signal input
rlabel metal2 s 41786 -400 41842 800 6 la_data_out_mprj[29]
port 437 nsew signal input
rlabel metal2 s 3238 -400 3294 800 6 la_data_out_mprj[2]
port 438 nsew signal input
rlabel metal2 s 43166 -400 43222 800 6 la_data_out_mprj[30]
port 439 nsew signal input
rlabel metal2 s 44638 -400 44694 800 6 la_data_out_mprj[31]
port 440 nsew signal input
rlabel metal2 s 46018 -400 46074 800 6 la_data_out_mprj[32]
port 441 nsew signal input
rlabel metal2 s 47490 -400 47546 800 6 la_data_out_mprj[33]
port 442 nsew signal input
rlabel metal2 s 48870 -400 48926 800 6 la_data_out_mprj[34]
port 443 nsew signal input
rlabel metal2 s 50342 -400 50398 800 6 la_data_out_mprj[35]
port 444 nsew signal input
rlabel metal2 s 51722 -400 51778 800 6 la_data_out_mprj[36]
port 445 nsew signal input
rlabel metal2 s 53194 -400 53250 800 6 la_data_out_mprj[37]
port 446 nsew signal input
rlabel metal2 s 54574 -400 54630 800 6 la_data_out_mprj[38]
port 447 nsew signal input
rlabel metal2 s 56046 -400 56102 800 6 la_data_out_mprj[39]
port 448 nsew signal input
rlabel metal2 s 4710 -400 4766 800 6 la_data_out_mprj[3]
port 449 nsew signal input
rlabel metal2 s 57426 -400 57482 800 6 la_data_out_mprj[40]
port 450 nsew signal input
rlabel metal2 s 58898 -400 58954 800 6 la_data_out_mprj[41]
port 451 nsew signal input
rlabel metal2 s 60278 -400 60334 800 6 la_data_out_mprj[42]
port 452 nsew signal input
rlabel metal2 s 61750 -400 61806 800 6 la_data_out_mprj[43]
port 453 nsew signal input
rlabel metal2 s 63130 -400 63186 800 6 la_data_out_mprj[44]
port 454 nsew signal input
rlabel metal2 s 64602 -400 64658 800 6 la_data_out_mprj[45]
port 455 nsew signal input
rlabel metal2 s 65982 -400 66038 800 6 la_data_out_mprj[46]
port 456 nsew signal input
rlabel metal2 s 67454 -400 67510 800 6 la_data_out_mprj[47]
port 457 nsew signal input
rlabel metal2 s 68834 -400 68890 800 6 la_data_out_mprj[48]
port 458 nsew signal input
rlabel metal2 s 70306 -400 70362 800 6 la_data_out_mprj[49]
port 459 nsew signal input
rlabel metal2 s 6090 -400 6146 800 6 la_data_out_mprj[4]
port 460 nsew signal input
rlabel metal2 s 71686 -400 71742 800 6 la_data_out_mprj[50]
port 461 nsew signal input
rlabel metal2 s 73158 -400 73214 800 6 la_data_out_mprj[51]
port 462 nsew signal input
rlabel metal2 s 74538 -400 74594 800 6 la_data_out_mprj[52]
port 463 nsew signal input
rlabel metal2 s 76010 -400 76066 800 6 la_data_out_mprj[53]
port 464 nsew signal input
rlabel metal2 s 77390 -400 77446 800 6 la_data_out_mprj[54]
port 465 nsew signal input
rlabel metal2 s 78862 -400 78918 800 6 la_data_out_mprj[55]
port 466 nsew signal input
rlabel metal2 s 80242 -400 80298 800 6 la_data_out_mprj[56]
port 467 nsew signal input
rlabel metal2 s 81714 -400 81770 800 6 la_data_out_mprj[57]
port 468 nsew signal input
rlabel metal2 s 83094 -400 83150 800 6 la_data_out_mprj[58]
port 469 nsew signal input
rlabel metal2 s 84566 -400 84622 800 6 la_data_out_mprj[59]
port 470 nsew signal input
rlabel metal2 s 7562 -400 7618 800 6 la_data_out_mprj[5]
port 471 nsew signal input
rlabel metal2 s 85946 -400 86002 800 6 la_data_out_mprj[60]
port 472 nsew signal input
rlabel metal2 s 87418 -400 87474 800 6 la_data_out_mprj[61]
port 473 nsew signal input
rlabel metal2 s 88798 -400 88854 800 6 la_data_out_mprj[62]
port 474 nsew signal input
rlabel metal2 s 90270 -400 90326 800 6 la_data_out_mprj[63]
port 475 nsew signal input
rlabel metal2 s 91650 -400 91706 800 6 la_data_out_mprj[64]
port 476 nsew signal input
rlabel metal2 s 93122 -400 93178 800 6 la_data_out_mprj[65]
port 477 nsew signal input
rlabel metal2 s 94502 -400 94558 800 6 la_data_out_mprj[66]
port 478 nsew signal input
rlabel metal2 s 95974 -400 96030 800 6 la_data_out_mprj[67]
port 479 nsew signal input
rlabel metal2 s 97354 -400 97410 800 6 la_data_out_mprj[68]
port 480 nsew signal input
rlabel metal2 s 98826 -400 98882 800 6 la_data_out_mprj[69]
port 481 nsew signal input
rlabel metal2 s 8942 -400 8998 800 6 la_data_out_mprj[6]
port 482 nsew signal input
rlabel metal2 s 100206 -400 100262 800 6 la_data_out_mprj[70]
port 483 nsew signal input
rlabel metal2 s 101678 -400 101734 800 6 la_data_out_mprj[71]
port 484 nsew signal input
rlabel metal2 s 103058 -400 103114 800 6 la_data_out_mprj[72]
port 485 nsew signal input
rlabel metal2 s 104530 -400 104586 800 6 la_data_out_mprj[73]
port 486 nsew signal input
rlabel metal2 s 105910 -400 105966 800 6 la_data_out_mprj[74]
port 487 nsew signal input
rlabel metal2 s 107382 -400 107438 800 6 la_data_out_mprj[75]
port 488 nsew signal input
rlabel metal2 s 108762 -400 108818 800 6 la_data_out_mprj[76]
port 489 nsew signal input
rlabel metal2 s 110234 -400 110290 800 6 la_data_out_mprj[77]
port 490 nsew signal input
rlabel metal2 s 111614 -400 111670 800 6 la_data_out_mprj[78]
port 491 nsew signal input
rlabel metal2 s 113086 -400 113142 800 6 la_data_out_mprj[79]
port 492 nsew signal input
rlabel metal2 s 10414 -400 10470 800 6 la_data_out_mprj[7]
port 493 nsew signal input
rlabel metal2 s 114466 -400 114522 800 6 la_data_out_mprj[80]
port 494 nsew signal input
rlabel metal2 s 115938 -400 115994 800 6 la_data_out_mprj[81]
port 495 nsew signal input
rlabel metal2 s 117318 -400 117374 800 6 la_data_out_mprj[82]
port 496 nsew signal input
rlabel metal2 s 118790 -400 118846 800 6 la_data_out_mprj[83]
port 497 nsew signal input
rlabel metal2 s 120170 -400 120226 800 6 la_data_out_mprj[84]
port 498 nsew signal input
rlabel metal2 s 121642 -400 121698 800 6 la_data_out_mprj[85]
port 499 nsew signal input
rlabel metal2 s 123022 -400 123078 800 6 la_data_out_mprj[86]
port 500 nsew signal input
rlabel metal2 s 124494 -400 124550 800 6 la_data_out_mprj[87]
port 501 nsew signal input
rlabel metal2 s 125874 -400 125930 800 6 la_data_out_mprj[88]
port 502 nsew signal input
rlabel metal2 s 127346 -400 127402 800 6 la_data_out_mprj[89]
port 503 nsew signal input
rlabel metal2 s 11794 -400 11850 800 6 la_data_out_mprj[8]
port 504 nsew signal input
rlabel metal2 s 128726 -400 128782 800 6 la_data_out_mprj[90]
port 505 nsew signal input
rlabel metal2 s 130198 -400 130254 800 6 la_data_out_mprj[91]
port 506 nsew signal input
rlabel metal2 s 131578 -400 131634 800 6 la_data_out_mprj[92]
port 507 nsew signal input
rlabel metal2 s 133050 -400 133106 800 6 la_data_out_mprj[93]
port 508 nsew signal input
rlabel metal2 s 134430 -400 134486 800 6 la_data_out_mprj[94]
port 509 nsew signal input
rlabel metal2 s 135902 -400 135958 800 6 la_data_out_mprj[95]
port 510 nsew signal input
rlabel metal2 s 137282 -400 137338 800 6 la_data_out_mprj[96]
port 511 nsew signal input
rlabel metal2 s 138754 -400 138810 800 6 la_data_out_mprj[97]
port 512 nsew signal input
rlabel metal2 s 140134 -400 140190 800 6 la_data_out_mprj[98]
port 513 nsew signal input
rlabel metal2 s 141606 -400 141662 800 6 la_data_out_mprj[99]
port 514 nsew signal input
rlabel metal2 s 13266 -400 13322 800 6 la_data_out_mprj[9]
port 515 nsew signal input
rlabel metal2 s 754 -400 810 800 6 la_iena_mprj[0]
port 516 nsew signal input
rlabel metal2 s 143354 -400 143410 800 6 la_iena_mprj[100]
port 517 nsew signal input
rlabel metal2 s 144826 -400 144882 800 6 la_iena_mprj[101]
port 518 nsew signal input
rlabel metal2 s 146206 -400 146262 800 6 la_iena_mprj[102]
port 519 nsew signal input
rlabel metal2 s 147678 -400 147734 800 6 la_iena_mprj[103]
port 520 nsew signal input
rlabel metal2 s 149058 -400 149114 800 6 la_iena_mprj[104]
port 521 nsew signal input
rlabel metal2 s 150530 -400 150586 800 6 la_iena_mprj[105]
port 522 nsew signal input
rlabel metal2 s 151910 -400 151966 800 6 la_iena_mprj[106]
port 523 nsew signal input
rlabel metal2 s 153382 -400 153438 800 6 la_iena_mprj[107]
port 524 nsew signal input
rlabel metal2 s 154762 -400 154818 800 6 la_iena_mprj[108]
port 525 nsew signal input
rlabel metal2 s 156234 -400 156290 800 6 la_iena_mprj[109]
port 526 nsew signal input
rlabel metal2 s 15014 -400 15070 800 6 la_iena_mprj[10]
port 527 nsew signal input
rlabel metal2 s 157614 -400 157670 800 6 la_iena_mprj[110]
port 528 nsew signal input
rlabel metal2 s 159086 -400 159142 800 6 la_iena_mprj[111]
port 529 nsew signal input
rlabel metal2 s 160466 -400 160522 800 6 la_iena_mprj[112]
port 530 nsew signal input
rlabel metal2 s 161938 -400 161994 800 6 la_iena_mprj[113]
port 531 nsew signal input
rlabel metal2 s 163318 -400 163374 800 6 la_iena_mprj[114]
port 532 nsew signal input
rlabel metal2 s 164790 -400 164846 800 6 la_iena_mprj[115]
port 533 nsew signal input
rlabel metal2 s 166170 -400 166226 800 6 la_iena_mprj[116]
port 534 nsew signal input
rlabel metal2 s 167642 -400 167698 800 6 la_iena_mprj[117]
port 535 nsew signal input
rlabel metal2 s 169022 -400 169078 800 6 la_iena_mprj[118]
port 536 nsew signal input
rlabel metal2 s 170494 -400 170550 800 6 la_iena_mprj[119]
port 537 nsew signal input
rlabel metal2 s 16486 -400 16542 800 6 la_iena_mprj[11]
port 538 nsew signal input
rlabel metal2 s 171874 -400 171930 800 6 la_iena_mprj[120]
port 539 nsew signal input
rlabel metal2 s 173346 -400 173402 800 6 la_iena_mprj[121]
port 540 nsew signal input
rlabel metal2 s 174726 -400 174782 800 6 la_iena_mprj[122]
port 541 nsew signal input
rlabel metal2 s 176198 -400 176254 800 6 la_iena_mprj[123]
port 542 nsew signal input
rlabel metal2 s 177578 -400 177634 800 6 la_iena_mprj[124]
port 543 nsew signal input
rlabel metal2 s 179050 -400 179106 800 6 la_iena_mprj[125]
port 544 nsew signal input
rlabel metal2 s 180430 -400 180486 800 6 la_iena_mprj[126]
port 545 nsew signal input
rlabel metal2 s 181902 -400 181958 800 6 la_iena_mprj[127]
port 546 nsew signal input
rlabel metal2 s 17866 -400 17922 800 6 la_iena_mprj[12]
port 547 nsew signal input
rlabel metal2 s 19338 -400 19394 800 6 la_iena_mprj[13]
port 548 nsew signal input
rlabel metal2 s 20718 -400 20774 800 6 la_iena_mprj[14]
port 549 nsew signal input
rlabel metal2 s 22190 -400 22246 800 6 la_iena_mprj[15]
port 550 nsew signal input
rlabel metal2 s 23570 -400 23626 800 6 la_iena_mprj[16]
port 551 nsew signal input
rlabel metal2 s 25042 -400 25098 800 6 la_iena_mprj[17]
port 552 nsew signal input
rlabel metal2 s 26422 -400 26478 800 6 la_iena_mprj[18]
port 553 nsew signal input
rlabel metal2 s 27894 -400 27950 800 6 la_iena_mprj[19]
port 554 nsew signal input
rlabel metal2 s 2226 -400 2282 800 6 la_iena_mprj[1]
port 555 nsew signal input
rlabel metal2 s 29274 -400 29330 800 6 la_iena_mprj[20]
port 556 nsew signal input
rlabel metal2 s 30746 -400 30802 800 6 la_iena_mprj[21]
port 557 nsew signal input
rlabel metal2 s 32126 -400 32182 800 6 la_iena_mprj[22]
port 558 nsew signal input
rlabel metal2 s 33598 -400 33654 800 6 la_iena_mprj[23]
port 559 nsew signal input
rlabel metal2 s 34978 -400 35034 800 6 la_iena_mprj[24]
port 560 nsew signal input
rlabel metal2 s 36450 -400 36506 800 6 la_iena_mprj[25]
port 561 nsew signal input
rlabel metal2 s 37830 -400 37886 800 6 la_iena_mprj[26]
port 562 nsew signal input
rlabel metal2 s 39302 -400 39358 800 6 la_iena_mprj[27]
port 563 nsew signal input
rlabel metal2 s 40682 -400 40738 800 6 la_iena_mprj[28]
port 564 nsew signal input
rlabel metal2 s 42154 -400 42210 800 6 la_iena_mprj[29]
port 565 nsew signal input
rlabel metal2 s 3606 -400 3662 800 6 la_iena_mprj[2]
port 566 nsew signal input
rlabel metal2 s 43534 -400 43590 800 6 la_iena_mprj[30]
port 567 nsew signal input
rlabel metal2 s 45006 -400 45062 800 6 la_iena_mprj[31]
port 568 nsew signal input
rlabel metal2 s 46386 -400 46442 800 6 la_iena_mprj[32]
port 569 nsew signal input
rlabel metal2 s 47858 -400 47914 800 6 la_iena_mprj[33]
port 570 nsew signal input
rlabel metal2 s 49238 -400 49294 800 6 la_iena_mprj[34]
port 571 nsew signal input
rlabel metal2 s 50710 -400 50766 800 6 la_iena_mprj[35]
port 572 nsew signal input
rlabel metal2 s 52090 -400 52146 800 6 la_iena_mprj[36]
port 573 nsew signal input
rlabel metal2 s 53562 -400 53618 800 6 la_iena_mprj[37]
port 574 nsew signal input
rlabel metal2 s 54942 -400 54998 800 6 la_iena_mprj[38]
port 575 nsew signal input
rlabel metal2 s 56414 -400 56470 800 6 la_iena_mprj[39]
port 576 nsew signal input
rlabel metal2 s 5078 -400 5134 800 6 la_iena_mprj[3]
port 577 nsew signal input
rlabel metal2 s 57794 -400 57850 800 6 la_iena_mprj[40]
port 578 nsew signal input
rlabel metal2 s 59266 -400 59322 800 6 la_iena_mprj[41]
port 579 nsew signal input
rlabel metal2 s 60646 -400 60702 800 6 la_iena_mprj[42]
port 580 nsew signal input
rlabel metal2 s 62118 -400 62174 800 6 la_iena_mprj[43]
port 581 nsew signal input
rlabel metal2 s 63498 -400 63554 800 6 la_iena_mprj[44]
port 582 nsew signal input
rlabel metal2 s 64970 -400 65026 800 6 la_iena_mprj[45]
port 583 nsew signal input
rlabel metal2 s 66350 -400 66406 800 6 la_iena_mprj[46]
port 584 nsew signal input
rlabel metal2 s 67822 -400 67878 800 6 la_iena_mprj[47]
port 585 nsew signal input
rlabel metal2 s 69202 -400 69258 800 6 la_iena_mprj[48]
port 586 nsew signal input
rlabel metal2 s 70674 -400 70730 800 6 la_iena_mprj[49]
port 587 nsew signal input
rlabel metal2 s 6458 -400 6514 800 6 la_iena_mprj[4]
port 588 nsew signal input
rlabel metal2 s 72054 -400 72110 800 6 la_iena_mprj[50]
port 589 nsew signal input
rlabel metal2 s 73526 -400 73582 800 6 la_iena_mprj[51]
port 590 nsew signal input
rlabel metal2 s 74906 -400 74962 800 6 la_iena_mprj[52]
port 591 nsew signal input
rlabel metal2 s 76378 -400 76434 800 6 la_iena_mprj[53]
port 592 nsew signal input
rlabel metal2 s 77758 -400 77814 800 6 la_iena_mprj[54]
port 593 nsew signal input
rlabel metal2 s 79230 -400 79286 800 6 la_iena_mprj[55]
port 594 nsew signal input
rlabel metal2 s 80610 -400 80666 800 6 la_iena_mprj[56]
port 595 nsew signal input
rlabel metal2 s 82082 -400 82138 800 6 la_iena_mprj[57]
port 596 nsew signal input
rlabel metal2 s 83462 -400 83518 800 6 la_iena_mprj[58]
port 597 nsew signal input
rlabel metal2 s 84934 -400 84990 800 6 la_iena_mprj[59]
port 598 nsew signal input
rlabel metal2 s 7930 -400 7986 800 6 la_iena_mprj[5]
port 599 nsew signal input
rlabel metal2 s 86314 -400 86370 800 6 la_iena_mprj[60]
port 600 nsew signal input
rlabel metal2 s 87786 -400 87842 800 6 la_iena_mprj[61]
port 601 nsew signal input
rlabel metal2 s 89166 -400 89222 800 6 la_iena_mprj[62]
port 602 nsew signal input
rlabel metal2 s 90638 -400 90694 800 6 la_iena_mprj[63]
port 603 nsew signal input
rlabel metal2 s 92018 -400 92074 800 6 la_iena_mprj[64]
port 604 nsew signal input
rlabel metal2 s 93490 -400 93546 800 6 la_iena_mprj[65]
port 605 nsew signal input
rlabel metal2 s 94870 -400 94926 800 6 la_iena_mprj[66]
port 606 nsew signal input
rlabel metal2 s 96342 -400 96398 800 6 la_iena_mprj[67]
port 607 nsew signal input
rlabel metal2 s 97722 -400 97778 800 6 la_iena_mprj[68]
port 608 nsew signal input
rlabel metal2 s 99194 -400 99250 800 6 la_iena_mprj[69]
port 609 nsew signal input
rlabel metal2 s 9310 -400 9366 800 6 la_iena_mprj[6]
port 610 nsew signal input
rlabel metal2 s 100574 -400 100630 800 6 la_iena_mprj[70]
port 611 nsew signal input
rlabel metal2 s 102046 -400 102102 800 6 la_iena_mprj[71]
port 612 nsew signal input
rlabel metal2 s 103426 -400 103482 800 6 la_iena_mprj[72]
port 613 nsew signal input
rlabel metal2 s 104898 -400 104954 800 6 la_iena_mprj[73]
port 614 nsew signal input
rlabel metal2 s 106278 -400 106334 800 6 la_iena_mprj[74]
port 615 nsew signal input
rlabel metal2 s 107750 -400 107806 800 6 la_iena_mprj[75]
port 616 nsew signal input
rlabel metal2 s 109130 -400 109186 800 6 la_iena_mprj[76]
port 617 nsew signal input
rlabel metal2 s 110602 -400 110658 800 6 la_iena_mprj[77]
port 618 nsew signal input
rlabel metal2 s 111982 -400 112038 800 6 la_iena_mprj[78]
port 619 nsew signal input
rlabel metal2 s 113454 -400 113510 800 6 la_iena_mprj[79]
port 620 nsew signal input
rlabel metal2 s 10782 -400 10838 800 6 la_iena_mprj[7]
port 621 nsew signal input
rlabel metal2 s 114834 -400 114890 800 6 la_iena_mprj[80]
port 622 nsew signal input
rlabel metal2 s 116306 -400 116362 800 6 la_iena_mprj[81]
port 623 nsew signal input
rlabel metal2 s 117686 -400 117742 800 6 la_iena_mprj[82]
port 624 nsew signal input
rlabel metal2 s 119158 -400 119214 800 6 la_iena_mprj[83]
port 625 nsew signal input
rlabel metal2 s 120538 -400 120594 800 6 la_iena_mprj[84]
port 626 nsew signal input
rlabel metal2 s 122010 -400 122066 800 6 la_iena_mprj[85]
port 627 nsew signal input
rlabel metal2 s 123390 -400 123446 800 6 la_iena_mprj[86]
port 628 nsew signal input
rlabel metal2 s 124862 -400 124918 800 6 la_iena_mprj[87]
port 629 nsew signal input
rlabel metal2 s 126242 -400 126298 800 6 la_iena_mprj[88]
port 630 nsew signal input
rlabel metal2 s 127714 -400 127770 800 6 la_iena_mprj[89]
port 631 nsew signal input
rlabel metal2 s 12162 -400 12218 800 6 la_iena_mprj[8]
port 632 nsew signal input
rlabel metal2 s 129094 -400 129150 800 6 la_iena_mprj[90]
port 633 nsew signal input
rlabel metal2 s 130566 -400 130622 800 6 la_iena_mprj[91]
port 634 nsew signal input
rlabel metal2 s 131946 -400 132002 800 6 la_iena_mprj[92]
port 635 nsew signal input
rlabel metal2 s 133418 -400 133474 800 6 la_iena_mprj[93]
port 636 nsew signal input
rlabel metal2 s 134798 -400 134854 800 6 la_iena_mprj[94]
port 637 nsew signal input
rlabel metal2 s 136270 -400 136326 800 6 la_iena_mprj[95]
port 638 nsew signal input
rlabel metal2 s 137650 -400 137706 800 6 la_iena_mprj[96]
port 639 nsew signal input
rlabel metal2 s 139122 -400 139178 800 6 la_iena_mprj[97]
port 640 nsew signal input
rlabel metal2 s 140502 -400 140558 800 6 la_iena_mprj[98]
port 641 nsew signal input
rlabel metal2 s 141974 -400 142030 800 6 la_iena_mprj[99]
port 642 nsew signal input
rlabel metal2 s 13634 -400 13690 800 6 la_iena_mprj[9]
port 643 nsew signal input
rlabel metal2 s 48226 31200 48282 32400 6 la_oenb_core[0]
port 644 nsew signal output
rlabel metal2 s 181810 31200 181866 32400 6 la_oenb_core[100]
port 645 nsew signal output
rlabel metal2 s 183190 31200 183246 32400 6 la_oenb_core[101]
port 646 nsew signal output
rlabel metal2 s 184478 31200 184534 32400 6 la_oenb_core[102]
port 647 nsew signal output
rlabel metal2 s 185858 31200 185914 32400 6 la_oenb_core[103]
port 648 nsew signal output
rlabel metal2 s 187146 31200 187202 32400 6 la_oenb_core[104]
port 649 nsew signal output
rlabel metal2 s 188526 31200 188582 32400 6 la_oenb_core[105]
port 650 nsew signal output
rlabel metal2 s 189814 31200 189870 32400 6 la_oenb_core[106]
port 651 nsew signal output
rlabel metal2 s 191194 31200 191250 32400 6 la_oenb_core[107]
port 652 nsew signal output
rlabel metal2 s 192482 31200 192538 32400 6 la_oenb_core[108]
port 653 nsew signal output
rlabel metal2 s 193862 31200 193918 32400 6 la_oenb_core[109]
port 654 nsew signal output
rlabel metal2 s 61566 31200 61622 32400 6 la_oenb_core[10]
port 655 nsew signal output
rlabel metal2 s 195150 31200 195206 32400 6 la_oenb_core[110]
port 656 nsew signal output
rlabel metal2 s 196530 31200 196586 32400 6 la_oenb_core[111]
port 657 nsew signal output
rlabel metal2 s 197818 31200 197874 32400 6 la_oenb_core[112]
port 658 nsew signal output
rlabel metal2 s 199198 31200 199254 32400 6 la_oenb_core[113]
port 659 nsew signal output
rlabel metal2 s 200578 31200 200634 32400 6 la_oenb_core[114]
port 660 nsew signal output
rlabel metal2 s 201866 31200 201922 32400 6 la_oenb_core[115]
port 661 nsew signal output
rlabel metal2 s 203246 31200 203302 32400 6 la_oenb_core[116]
port 662 nsew signal output
rlabel metal2 s 204534 31200 204590 32400 6 la_oenb_core[117]
port 663 nsew signal output
rlabel metal2 s 205914 31200 205970 32400 6 la_oenb_core[118]
port 664 nsew signal output
rlabel metal2 s 207202 31200 207258 32400 6 la_oenb_core[119]
port 665 nsew signal output
rlabel metal2 s 62946 31200 63002 32400 6 la_oenb_core[11]
port 666 nsew signal output
rlabel metal2 s 208582 31200 208638 32400 6 la_oenb_core[120]
port 667 nsew signal output
rlabel metal2 s 209870 31200 209926 32400 6 la_oenb_core[121]
port 668 nsew signal output
rlabel metal2 s 211250 31200 211306 32400 6 la_oenb_core[122]
port 669 nsew signal output
rlabel metal2 s 212538 31200 212594 32400 6 la_oenb_core[123]
port 670 nsew signal output
rlabel metal2 s 213918 31200 213974 32400 6 la_oenb_core[124]
port 671 nsew signal output
rlabel metal2 s 215206 31200 215262 32400 6 la_oenb_core[125]
port 672 nsew signal output
rlabel metal2 s 216586 31200 216642 32400 6 la_oenb_core[126]
port 673 nsew signal output
rlabel metal2 s 217874 31200 217930 32400 6 la_oenb_core[127]
port 674 nsew signal output
rlabel metal2 s 64234 31200 64290 32400 6 la_oenb_core[12]
port 675 nsew signal output
rlabel metal2 s 65614 31200 65670 32400 6 la_oenb_core[13]
port 676 nsew signal output
rlabel metal2 s 66994 31200 67050 32400 6 la_oenb_core[14]
port 677 nsew signal output
rlabel metal2 s 68282 31200 68338 32400 6 la_oenb_core[15]
port 678 nsew signal output
rlabel metal2 s 69662 31200 69718 32400 6 la_oenb_core[16]
port 679 nsew signal output
rlabel metal2 s 70950 31200 71006 32400 6 la_oenb_core[17]
port 680 nsew signal output
rlabel metal2 s 72330 31200 72386 32400 6 la_oenb_core[18]
port 681 nsew signal output
rlabel metal2 s 73618 31200 73674 32400 6 la_oenb_core[19]
port 682 nsew signal output
rlabel metal2 s 49606 31200 49662 32400 6 la_oenb_core[1]
port 683 nsew signal output
rlabel metal2 s 74998 31200 75054 32400 6 la_oenb_core[20]
port 684 nsew signal output
rlabel metal2 s 76286 31200 76342 32400 6 la_oenb_core[21]
port 685 nsew signal output
rlabel metal2 s 77666 31200 77722 32400 6 la_oenb_core[22]
port 686 nsew signal output
rlabel metal2 s 78954 31200 79010 32400 6 la_oenb_core[23]
port 687 nsew signal output
rlabel metal2 s 80334 31200 80390 32400 6 la_oenb_core[24]
port 688 nsew signal output
rlabel metal2 s 81622 31200 81678 32400 6 la_oenb_core[25]
port 689 nsew signal output
rlabel metal2 s 83002 31200 83058 32400 6 la_oenb_core[26]
port 690 nsew signal output
rlabel metal2 s 84290 31200 84346 32400 6 la_oenb_core[27]
port 691 nsew signal output
rlabel metal2 s 85670 31200 85726 32400 6 la_oenb_core[28]
port 692 nsew signal output
rlabel metal2 s 86958 31200 87014 32400 6 la_oenb_core[29]
port 693 nsew signal output
rlabel metal2 s 50894 31200 50950 32400 6 la_oenb_core[2]
port 694 nsew signal output
rlabel metal2 s 88338 31200 88394 32400 6 la_oenb_core[30]
port 695 nsew signal output
rlabel metal2 s 89626 31200 89682 32400 6 la_oenb_core[31]
port 696 nsew signal output
rlabel metal2 s 91006 31200 91062 32400 6 la_oenb_core[32]
port 697 nsew signal output
rlabel metal2 s 92294 31200 92350 32400 6 la_oenb_core[33]
port 698 nsew signal output
rlabel metal2 s 93674 31200 93730 32400 6 la_oenb_core[34]
port 699 nsew signal output
rlabel metal2 s 94962 31200 95018 32400 6 la_oenb_core[35]
port 700 nsew signal output
rlabel metal2 s 96342 31200 96398 32400 6 la_oenb_core[36]
port 701 nsew signal output
rlabel metal2 s 97630 31200 97686 32400 6 la_oenb_core[37]
port 702 nsew signal output
rlabel metal2 s 99010 31200 99066 32400 6 la_oenb_core[38]
port 703 nsew signal output
rlabel metal2 s 100390 31200 100446 32400 6 la_oenb_core[39]
port 704 nsew signal output
rlabel metal2 s 52274 31200 52330 32400 6 la_oenb_core[3]
port 705 nsew signal output
rlabel metal2 s 101678 31200 101734 32400 6 la_oenb_core[40]
port 706 nsew signal output
rlabel metal2 s 103058 31200 103114 32400 6 la_oenb_core[41]
port 707 nsew signal output
rlabel metal2 s 104346 31200 104402 32400 6 la_oenb_core[42]
port 708 nsew signal output
rlabel metal2 s 105726 31200 105782 32400 6 la_oenb_core[43]
port 709 nsew signal output
rlabel metal2 s 107014 31200 107070 32400 6 la_oenb_core[44]
port 710 nsew signal output
rlabel metal2 s 108394 31200 108450 32400 6 la_oenb_core[45]
port 711 nsew signal output
rlabel metal2 s 109682 31200 109738 32400 6 la_oenb_core[46]
port 712 nsew signal output
rlabel metal2 s 111062 31200 111118 32400 6 la_oenb_core[47]
port 713 nsew signal output
rlabel metal2 s 112350 31200 112406 32400 6 la_oenb_core[48]
port 714 nsew signal output
rlabel metal2 s 113730 31200 113786 32400 6 la_oenb_core[49]
port 715 nsew signal output
rlabel metal2 s 53562 31200 53618 32400 6 la_oenb_core[4]
port 716 nsew signal output
rlabel metal2 s 115018 31200 115074 32400 6 la_oenb_core[50]
port 717 nsew signal output
rlabel metal2 s 116398 31200 116454 32400 6 la_oenb_core[51]
port 718 nsew signal output
rlabel metal2 s 117686 31200 117742 32400 6 la_oenb_core[52]
port 719 nsew signal output
rlabel metal2 s 119066 31200 119122 32400 6 la_oenb_core[53]
port 720 nsew signal output
rlabel metal2 s 120354 31200 120410 32400 6 la_oenb_core[54]
port 721 nsew signal output
rlabel metal2 s 121734 31200 121790 32400 6 la_oenb_core[55]
port 722 nsew signal output
rlabel metal2 s 123022 31200 123078 32400 6 la_oenb_core[56]
port 723 nsew signal output
rlabel metal2 s 124402 31200 124458 32400 6 la_oenb_core[57]
port 724 nsew signal output
rlabel metal2 s 125690 31200 125746 32400 6 la_oenb_core[58]
port 725 nsew signal output
rlabel metal2 s 127070 31200 127126 32400 6 la_oenb_core[59]
port 726 nsew signal output
rlabel metal2 s 54942 31200 54998 32400 6 la_oenb_core[5]
port 727 nsew signal output
rlabel metal2 s 128358 31200 128414 32400 6 la_oenb_core[60]
port 728 nsew signal output
rlabel metal2 s 129738 31200 129794 32400 6 la_oenb_core[61]
port 729 nsew signal output
rlabel metal2 s 131026 31200 131082 32400 6 la_oenb_core[62]
port 730 nsew signal output
rlabel metal2 s 132406 31200 132462 32400 6 la_oenb_core[63]
port 731 nsew signal output
rlabel metal2 s 133786 31200 133842 32400 6 la_oenb_core[64]
port 732 nsew signal output
rlabel metal2 s 135074 31200 135130 32400 6 la_oenb_core[65]
port 733 nsew signal output
rlabel metal2 s 136454 31200 136510 32400 6 la_oenb_core[66]
port 734 nsew signal output
rlabel metal2 s 137742 31200 137798 32400 6 la_oenb_core[67]
port 735 nsew signal output
rlabel metal2 s 139122 31200 139178 32400 6 la_oenb_core[68]
port 736 nsew signal output
rlabel metal2 s 140410 31200 140466 32400 6 la_oenb_core[69]
port 737 nsew signal output
rlabel metal2 s 56230 31200 56286 32400 6 la_oenb_core[6]
port 738 nsew signal output
rlabel metal2 s 141790 31200 141846 32400 6 la_oenb_core[70]
port 739 nsew signal output
rlabel metal2 s 143078 31200 143134 32400 6 la_oenb_core[71]
port 740 nsew signal output
rlabel metal2 s 144458 31200 144514 32400 6 la_oenb_core[72]
port 741 nsew signal output
rlabel metal2 s 145746 31200 145802 32400 6 la_oenb_core[73]
port 742 nsew signal output
rlabel metal2 s 147126 31200 147182 32400 6 la_oenb_core[74]
port 743 nsew signal output
rlabel metal2 s 148414 31200 148470 32400 6 la_oenb_core[75]
port 744 nsew signal output
rlabel metal2 s 149794 31200 149850 32400 6 la_oenb_core[76]
port 745 nsew signal output
rlabel metal2 s 151082 31200 151138 32400 6 la_oenb_core[77]
port 746 nsew signal output
rlabel metal2 s 152462 31200 152518 32400 6 la_oenb_core[78]
port 747 nsew signal output
rlabel metal2 s 153750 31200 153806 32400 6 la_oenb_core[79]
port 748 nsew signal output
rlabel metal2 s 57610 31200 57666 32400 6 la_oenb_core[7]
port 749 nsew signal output
rlabel metal2 s 155130 31200 155186 32400 6 la_oenb_core[80]
port 750 nsew signal output
rlabel metal2 s 156418 31200 156474 32400 6 la_oenb_core[81]
port 751 nsew signal output
rlabel metal2 s 157798 31200 157854 32400 6 la_oenb_core[82]
port 752 nsew signal output
rlabel metal2 s 159086 31200 159142 32400 6 la_oenb_core[83]
port 753 nsew signal output
rlabel metal2 s 160466 31200 160522 32400 6 la_oenb_core[84]
port 754 nsew signal output
rlabel metal2 s 161754 31200 161810 32400 6 la_oenb_core[85]
port 755 nsew signal output
rlabel metal2 s 163134 31200 163190 32400 6 la_oenb_core[86]
port 756 nsew signal output
rlabel metal2 s 164422 31200 164478 32400 6 la_oenb_core[87]
port 757 nsew signal output
rlabel metal2 s 165802 31200 165858 32400 6 la_oenb_core[88]
port 758 nsew signal output
rlabel metal2 s 167182 31200 167238 32400 6 la_oenb_core[89]
port 759 nsew signal output
rlabel metal2 s 58898 31200 58954 32400 6 la_oenb_core[8]
port 760 nsew signal output
rlabel metal2 s 168470 31200 168526 32400 6 la_oenb_core[90]
port 761 nsew signal output
rlabel metal2 s 169850 31200 169906 32400 6 la_oenb_core[91]
port 762 nsew signal output
rlabel metal2 s 171138 31200 171194 32400 6 la_oenb_core[92]
port 763 nsew signal output
rlabel metal2 s 172518 31200 172574 32400 6 la_oenb_core[93]
port 764 nsew signal output
rlabel metal2 s 173806 31200 173862 32400 6 la_oenb_core[94]
port 765 nsew signal output
rlabel metal2 s 175186 31200 175242 32400 6 la_oenb_core[95]
port 766 nsew signal output
rlabel metal2 s 176474 31200 176530 32400 6 la_oenb_core[96]
port 767 nsew signal output
rlabel metal2 s 177854 31200 177910 32400 6 la_oenb_core[97]
port 768 nsew signal output
rlabel metal2 s 179142 31200 179198 32400 6 la_oenb_core[98]
port 769 nsew signal output
rlabel metal2 s 180522 31200 180578 32400 6 la_oenb_core[99]
port 770 nsew signal output
rlabel metal2 s 60278 31200 60334 32400 6 la_oenb_core[9]
port 771 nsew signal output
rlabel metal2 s 1122 -400 1178 800 6 la_oenb_mprj[0]
port 772 nsew signal input
rlabel metal2 s 143722 -400 143778 800 6 la_oenb_mprj[100]
port 773 nsew signal input
rlabel metal2 s 145194 -400 145250 800 6 la_oenb_mprj[101]
port 774 nsew signal input
rlabel metal2 s 146574 -400 146630 800 6 la_oenb_mprj[102]
port 775 nsew signal input
rlabel metal2 s 148046 -400 148102 800 6 la_oenb_mprj[103]
port 776 nsew signal input
rlabel metal2 s 149426 -400 149482 800 6 la_oenb_mprj[104]
port 777 nsew signal input
rlabel metal2 s 150898 -400 150954 800 6 la_oenb_mprj[105]
port 778 nsew signal input
rlabel metal2 s 152278 -400 152334 800 6 la_oenb_mprj[106]
port 779 nsew signal input
rlabel metal2 s 153750 -400 153806 800 6 la_oenb_mprj[107]
port 780 nsew signal input
rlabel metal2 s 155130 -400 155186 800 6 la_oenb_mprj[108]
port 781 nsew signal input
rlabel metal2 s 156602 -400 156658 800 6 la_oenb_mprj[109]
port 782 nsew signal input
rlabel metal2 s 15382 -400 15438 800 6 la_oenb_mprj[10]
port 783 nsew signal input
rlabel metal2 s 157982 -400 158038 800 6 la_oenb_mprj[110]
port 784 nsew signal input
rlabel metal2 s 159454 -400 159510 800 6 la_oenb_mprj[111]
port 785 nsew signal input
rlabel metal2 s 160834 -400 160890 800 6 la_oenb_mprj[112]
port 786 nsew signal input
rlabel metal2 s 162306 -400 162362 800 6 la_oenb_mprj[113]
port 787 nsew signal input
rlabel metal2 s 163686 -400 163742 800 6 la_oenb_mprj[114]
port 788 nsew signal input
rlabel metal2 s 165158 -400 165214 800 6 la_oenb_mprj[115]
port 789 nsew signal input
rlabel metal2 s 166538 -400 166594 800 6 la_oenb_mprj[116]
port 790 nsew signal input
rlabel metal2 s 168010 -400 168066 800 6 la_oenb_mprj[117]
port 791 nsew signal input
rlabel metal2 s 169390 -400 169446 800 6 la_oenb_mprj[118]
port 792 nsew signal input
rlabel metal2 s 170862 -400 170918 800 6 la_oenb_mprj[119]
port 793 nsew signal input
rlabel metal2 s 16854 -400 16910 800 6 la_oenb_mprj[11]
port 794 nsew signal input
rlabel metal2 s 172242 -400 172298 800 6 la_oenb_mprj[120]
port 795 nsew signal input
rlabel metal2 s 173714 -400 173770 800 6 la_oenb_mprj[121]
port 796 nsew signal input
rlabel metal2 s 175094 -400 175150 800 6 la_oenb_mprj[122]
port 797 nsew signal input
rlabel metal2 s 176566 -400 176622 800 6 la_oenb_mprj[123]
port 798 nsew signal input
rlabel metal2 s 177946 -400 178002 800 6 la_oenb_mprj[124]
port 799 nsew signal input
rlabel metal2 s 179418 -400 179474 800 6 la_oenb_mprj[125]
port 800 nsew signal input
rlabel metal2 s 180798 -400 180854 800 6 la_oenb_mprj[126]
port 801 nsew signal input
rlabel metal2 s 182270 -400 182326 800 6 la_oenb_mprj[127]
port 802 nsew signal input
rlabel metal2 s 18234 -400 18290 800 6 la_oenb_mprj[12]
port 803 nsew signal input
rlabel metal2 s 19706 -400 19762 800 6 la_oenb_mprj[13]
port 804 nsew signal input
rlabel metal2 s 21086 -400 21142 800 6 la_oenb_mprj[14]
port 805 nsew signal input
rlabel metal2 s 22558 -400 22614 800 6 la_oenb_mprj[15]
port 806 nsew signal input
rlabel metal2 s 23938 -400 23994 800 6 la_oenb_mprj[16]
port 807 nsew signal input
rlabel metal2 s 25410 -400 25466 800 6 la_oenb_mprj[17]
port 808 nsew signal input
rlabel metal2 s 26790 -400 26846 800 6 la_oenb_mprj[18]
port 809 nsew signal input
rlabel metal2 s 28262 -400 28318 800 6 la_oenb_mprj[19]
port 810 nsew signal input
rlabel metal2 s 2594 -400 2650 800 6 la_oenb_mprj[1]
port 811 nsew signal input
rlabel metal2 s 29642 -400 29698 800 6 la_oenb_mprj[20]
port 812 nsew signal input
rlabel metal2 s 31114 -400 31170 800 6 la_oenb_mprj[21]
port 813 nsew signal input
rlabel metal2 s 32494 -400 32550 800 6 la_oenb_mprj[22]
port 814 nsew signal input
rlabel metal2 s 33966 -400 34022 800 6 la_oenb_mprj[23]
port 815 nsew signal input
rlabel metal2 s 35346 -400 35402 800 6 la_oenb_mprj[24]
port 816 nsew signal input
rlabel metal2 s 36818 -400 36874 800 6 la_oenb_mprj[25]
port 817 nsew signal input
rlabel metal2 s 38198 -400 38254 800 6 la_oenb_mprj[26]
port 818 nsew signal input
rlabel metal2 s 39670 -400 39726 800 6 la_oenb_mprj[27]
port 819 nsew signal input
rlabel metal2 s 41050 -400 41106 800 6 la_oenb_mprj[28]
port 820 nsew signal input
rlabel metal2 s 42522 -400 42578 800 6 la_oenb_mprj[29]
port 821 nsew signal input
rlabel metal2 s 3974 -400 4030 800 6 la_oenb_mprj[2]
port 822 nsew signal input
rlabel metal2 s 43902 -400 43958 800 6 la_oenb_mprj[30]
port 823 nsew signal input
rlabel metal2 s 45374 -400 45430 800 6 la_oenb_mprj[31]
port 824 nsew signal input
rlabel metal2 s 46754 -400 46810 800 6 la_oenb_mprj[32]
port 825 nsew signal input
rlabel metal2 s 48226 -400 48282 800 6 la_oenb_mprj[33]
port 826 nsew signal input
rlabel metal2 s 49606 -400 49662 800 6 la_oenb_mprj[34]
port 827 nsew signal input
rlabel metal2 s 51078 -400 51134 800 6 la_oenb_mprj[35]
port 828 nsew signal input
rlabel metal2 s 52458 -400 52514 800 6 la_oenb_mprj[36]
port 829 nsew signal input
rlabel metal2 s 53930 -400 53986 800 6 la_oenb_mprj[37]
port 830 nsew signal input
rlabel metal2 s 55310 -400 55366 800 6 la_oenb_mprj[38]
port 831 nsew signal input
rlabel metal2 s 56782 -400 56838 800 6 la_oenb_mprj[39]
port 832 nsew signal input
rlabel metal2 s 5446 -400 5502 800 6 la_oenb_mprj[3]
port 833 nsew signal input
rlabel metal2 s 58162 -400 58218 800 6 la_oenb_mprj[40]
port 834 nsew signal input
rlabel metal2 s 59634 -400 59690 800 6 la_oenb_mprj[41]
port 835 nsew signal input
rlabel metal2 s 61014 -400 61070 800 6 la_oenb_mprj[42]
port 836 nsew signal input
rlabel metal2 s 62486 -400 62542 800 6 la_oenb_mprj[43]
port 837 nsew signal input
rlabel metal2 s 63866 -400 63922 800 6 la_oenb_mprj[44]
port 838 nsew signal input
rlabel metal2 s 65338 -400 65394 800 6 la_oenb_mprj[45]
port 839 nsew signal input
rlabel metal2 s 66718 -400 66774 800 6 la_oenb_mprj[46]
port 840 nsew signal input
rlabel metal2 s 68190 -400 68246 800 6 la_oenb_mprj[47]
port 841 nsew signal input
rlabel metal2 s 69570 -400 69626 800 6 la_oenb_mprj[48]
port 842 nsew signal input
rlabel metal2 s 71042 -400 71098 800 6 la_oenb_mprj[49]
port 843 nsew signal input
rlabel metal2 s 6826 -400 6882 800 6 la_oenb_mprj[4]
port 844 nsew signal input
rlabel metal2 s 72422 -400 72478 800 6 la_oenb_mprj[50]
port 845 nsew signal input
rlabel metal2 s 73894 -400 73950 800 6 la_oenb_mprj[51]
port 846 nsew signal input
rlabel metal2 s 75274 -400 75330 800 6 la_oenb_mprj[52]
port 847 nsew signal input
rlabel metal2 s 76746 -400 76802 800 6 la_oenb_mprj[53]
port 848 nsew signal input
rlabel metal2 s 78126 -400 78182 800 6 la_oenb_mprj[54]
port 849 nsew signal input
rlabel metal2 s 79598 -400 79654 800 6 la_oenb_mprj[55]
port 850 nsew signal input
rlabel metal2 s 80978 -400 81034 800 6 la_oenb_mprj[56]
port 851 nsew signal input
rlabel metal2 s 82450 -400 82506 800 6 la_oenb_mprj[57]
port 852 nsew signal input
rlabel metal2 s 83830 -400 83886 800 6 la_oenb_mprj[58]
port 853 nsew signal input
rlabel metal2 s 85302 -400 85358 800 6 la_oenb_mprj[59]
port 854 nsew signal input
rlabel metal2 s 8298 -400 8354 800 6 la_oenb_mprj[5]
port 855 nsew signal input
rlabel metal2 s 86682 -400 86738 800 6 la_oenb_mprj[60]
port 856 nsew signal input
rlabel metal2 s 88154 -400 88210 800 6 la_oenb_mprj[61]
port 857 nsew signal input
rlabel metal2 s 89534 -400 89590 800 6 la_oenb_mprj[62]
port 858 nsew signal input
rlabel metal2 s 91006 -400 91062 800 6 la_oenb_mprj[63]
port 859 nsew signal input
rlabel metal2 s 92386 -400 92442 800 6 la_oenb_mprj[64]
port 860 nsew signal input
rlabel metal2 s 93858 -400 93914 800 6 la_oenb_mprj[65]
port 861 nsew signal input
rlabel metal2 s 95238 -400 95294 800 6 la_oenb_mprj[66]
port 862 nsew signal input
rlabel metal2 s 96710 -400 96766 800 6 la_oenb_mprj[67]
port 863 nsew signal input
rlabel metal2 s 98090 -400 98146 800 6 la_oenb_mprj[68]
port 864 nsew signal input
rlabel metal2 s 99562 -400 99618 800 6 la_oenb_mprj[69]
port 865 nsew signal input
rlabel metal2 s 9678 -400 9734 800 6 la_oenb_mprj[6]
port 866 nsew signal input
rlabel metal2 s 100942 -400 100998 800 6 la_oenb_mprj[70]
port 867 nsew signal input
rlabel metal2 s 102414 -400 102470 800 6 la_oenb_mprj[71]
port 868 nsew signal input
rlabel metal2 s 103794 -400 103850 800 6 la_oenb_mprj[72]
port 869 nsew signal input
rlabel metal2 s 105266 -400 105322 800 6 la_oenb_mprj[73]
port 870 nsew signal input
rlabel metal2 s 106646 -400 106702 800 6 la_oenb_mprj[74]
port 871 nsew signal input
rlabel metal2 s 108118 -400 108174 800 6 la_oenb_mprj[75]
port 872 nsew signal input
rlabel metal2 s 109498 -400 109554 800 6 la_oenb_mprj[76]
port 873 nsew signal input
rlabel metal2 s 110970 -400 111026 800 6 la_oenb_mprj[77]
port 874 nsew signal input
rlabel metal2 s 112350 -400 112406 800 6 la_oenb_mprj[78]
port 875 nsew signal input
rlabel metal2 s 113822 -400 113878 800 6 la_oenb_mprj[79]
port 876 nsew signal input
rlabel metal2 s 11150 -400 11206 800 6 la_oenb_mprj[7]
port 877 nsew signal input
rlabel metal2 s 115202 -400 115258 800 6 la_oenb_mprj[80]
port 878 nsew signal input
rlabel metal2 s 116674 -400 116730 800 6 la_oenb_mprj[81]
port 879 nsew signal input
rlabel metal2 s 118054 -400 118110 800 6 la_oenb_mprj[82]
port 880 nsew signal input
rlabel metal2 s 119526 -400 119582 800 6 la_oenb_mprj[83]
port 881 nsew signal input
rlabel metal2 s 120906 -400 120962 800 6 la_oenb_mprj[84]
port 882 nsew signal input
rlabel metal2 s 122378 -400 122434 800 6 la_oenb_mprj[85]
port 883 nsew signal input
rlabel metal2 s 123758 -400 123814 800 6 la_oenb_mprj[86]
port 884 nsew signal input
rlabel metal2 s 125230 -400 125286 800 6 la_oenb_mprj[87]
port 885 nsew signal input
rlabel metal2 s 126610 -400 126666 800 6 la_oenb_mprj[88]
port 886 nsew signal input
rlabel metal2 s 128082 -400 128138 800 6 la_oenb_mprj[89]
port 887 nsew signal input
rlabel metal2 s 12530 -400 12586 800 6 la_oenb_mprj[8]
port 888 nsew signal input
rlabel metal2 s 129462 -400 129518 800 6 la_oenb_mprj[90]
port 889 nsew signal input
rlabel metal2 s 130934 -400 130990 800 6 la_oenb_mprj[91]
port 890 nsew signal input
rlabel metal2 s 132314 -400 132370 800 6 la_oenb_mprj[92]
port 891 nsew signal input
rlabel metal2 s 133786 -400 133842 800 6 la_oenb_mprj[93]
port 892 nsew signal input
rlabel metal2 s 135166 -400 135222 800 6 la_oenb_mprj[94]
port 893 nsew signal input
rlabel metal2 s 136638 -400 136694 800 6 la_oenb_mprj[95]
port 894 nsew signal input
rlabel metal2 s 138018 -400 138074 800 6 la_oenb_mprj[96]
port 895 nsew signal input
rlabel metal2 s 139490 -400 139546 800 6 la_oenb_mprj[97]
port 896 nsew signal input
rlabel metal2 s 140870 -400 140926 800 6 la_oenb_mprj[98]
port 897 nsew signal input
rlabel metal2 s 142342 -400 142398 800 6 la_oenb_mprj[99]
port 898 nsew signal input
rlabel metal2 s 14002 -400 14058 800 6 la_oenb_mprj[9]
port 899 nsew signal input
rlabel metal2 s 182638 -400 182694 800 6 mprj_ack_i_core
port 900 nsew signal output
rlabel metal2 s 1030 31200 1086 32400 6 mprj_ack_i_user
port 901 nsew signal input
rlabel metal2 s 184018 -400 184074 800 6 mprj_adr_o_core[0]
port 902 nsew signal input
rlabel metal2 s 196162 -400 196218 800 6 mprj_adr_o_core[10]
port 903 nsew signal input
rlabel metal2 s 197174 -400 197230 800 6 mprj_adr_o_core[11]
port 904 nsew signal input
rlabel metal2 s 198278 -400 198334 800 6 mprj_adr_o_core[12]
port 905 nsew signal input
rlabel metal2 s 199382 -400 199438 800 6 mprj_adr_o_core[13]
port 906 nsew signal input
rlabel metal2 s 200394 -400 200450 800 6 mprj_adr_o_core[14]
port 907 nsew signal input
rlabel metal2 s 201498 -400 201554 800 6 mprj_adr_o_core[15]
port 908 nsew signal input
rlabel metal2 s 202602 -400 202658 800 6 mprj_adr_o_core[16]
port 909 nsew signal input
rlabel metal2 s 203614 -400 203670 800 6 mprj_adr_o_core[17]
port 910 nsew signal input
rlabel metal2 s 204718 -400 204774 800 6 mprj_adr_o_core[18]
port 911 nsew signal input
rlabel metal2 s 205730 -400 205786 800 6 mprj_adr_o_core[19]
port 912 nsew signal input
rlabel metal2 s 185490 -400 185546 800 6 mprj_adr_o_core[1]
port 913 nsew signal input
rlabel metal2 s 206834 -400 206890 800 6 mprj_adr_o_core[20]
port 914 nsew signal input
rlabel metal2 s 207938 -400 207994 800 6 mprj_adr_o_core[21]
port 915 nsew signal input
rlabel metal2 s 208950 -400 209006 800 6 mprj_adr_o_core[22]
port 916 nsew signal input
rlabel metal2 s 210054 -400 210110 800 6 mprj_adr_o_core[23]
port 917 nsew signal input
rlabel metal2 s 211158 -400 211214 800 6 mprj_adr_o_core[24]
port 918 nsew signal input
rlabel metal2 s 212170 -400 212226 800 6 mprj_adr_o_core[25]
port 919 nsew signal input
rlabel metal2 s 213274 -400 213330 800 6 mprj_adr_o_core[26]
port 920 nsew signal input
rlabel metal2 s 214286 -400 214342 800 6 mprj_adr_o_core[27]
port 921 nsew signal input
rlabel metal2 s 215390 -400 215446 800 6 mprj_adr_o_core[28]
port 922 nsew signal input
rlabel metal2 s 216494 -400 216550 800 6 mprj_adr_o_core[29]
port 923 nsew signal input
rlabel metal2 s 186870 -400 186926 800 6 mprj_adr_o_core[2]
port 924 nsew signal input
rlabel metal2 s 217506 -400 217562 800 6 mprj_adr_o_core[30]
port 925 nsew signal input
rlabel metal2 s 218610 -400 218666 800 6 mprj_adr_o_core[31]
port 926 nsew signal input
rlabel metal2 s 188342 -400 188398 800 6 mprj_adr_o_core[3]
port 927 nsew signal input
rlabel metal2 s 189722 -400 189778 800 6 mprj_adr_o_core[4]
port 928 nsew signal input
rlabel metal2 s 190826 -400 190882 800 6 mprj_adr_o_core[5]
port 929 nsew signal input
rlabel metal2 s 191838 -400 191894 800 6 mprj_adr_o_core[6]
port 930 nsew signal input
rlabel metal2 s 192942 -400 192998 800 6 mprj_adr_o_core[7]
port 931 nsew signal input
rlabel metal2 s 194046 -400 194102 800 6 mprj_adr_o_core[8]
port 932 nsew signal input
rlabel metal2 s 195058 -400 195114 800 6 mprj_adr_o_core[9]
port 933 nsew signal input
rlabel metal2 s 2870 31200 2926 32400 6 mprj_adr_o_user[0]
port 934 nsew signal output
rlabel metal2 s 17958 31200 18014 32400 6 mprj_adr_o_user[10]
port 935 nsew signal output
rlabel metal2 s 19338 31200 19394 32400 6 mprj_adr_o_user[11]
port 936 nsew signal output
rlabel metal2 s 20626 31200 20682 32400 6 mprj_adr_o_user[12]
port 937 nsew signal output
rlabel metal2 s 22006 31200 22062 32400 6 mprj_adr_o_user[13]
port 938 nsew signal output
rlabel metal2 s 23294 31200 23350 32400 6 mprj_adr_o_user[14]
port 939 nsew signal output
rlabel metal2 s 24674 31200 24730 32400 6 mprj_adr_o_user[15]
port 940 nsew signal output
rlabel metal2 s 25962 31200 26018 32400 6 mprj_adr_o_user[16]
port 941 nsew signal output
rlabel metal2 s 27342 31200 27398 32400 6 mprj_adr_o_user[17]
port 942 nsew signal output
rlabel metal2 s 28630 31200 28686 32400 6 mprj_adr_o_user[18]
port 943 nsew signal output
rlabel metal2 s 30010 31200 30066 32400 6 mprj_adr_o_user[19]
port 944 nsew signal output
rlabel metal2 s 4618 31200 4674 32400 6 mprj_adr_o_user[1]
port 945 nsew signal output
rlabel metal2 s 31298 31200 31354 32400 6 mprj_adr_o_user[20]
port 946 nsew signal output
rlabel metal2 s 32678 31200 32734 32400 6 mprj_adr_o_user[21]
port 947 nsew signal output
rlabel metal2 s 33966 31200 34022 32400 6 mprj_adr_o_user[22]
port 948 nsew signal output
rlabel metal2 s 35346 31200 35402 32400 6 mprj_adr_o_user[23]
port 949 nsew signal output
rlabel metal2 s 36634 31200 36690 32400 6 mprj_adr_o_user[24]
port 950 nsew signal output
rlabel metal2 s 38014 31200 38070 32400 6 mprj_adr_o_user[25]
port 951 nsew signal output
rlabel metal2 s 39302 31200 39358 32400 6 mprj_adr_o_user[26]
port 952 nsew signal output
rlabel metal2 s 40682 31200 40738 32400 6 mprj_adr_o_user[27]
port 953 nsew signal output
rlabel metal2 s 41970 31200 42026 32400 6 mprj_adr_o_user[28]
port 954 nsew signal output
rlabel metal2 s 43350 31200 43406 32400 6 mprj_adr_o_user[29]
port 955 nsew signal output
rlabel metal2 s 6366 31200 6422 32400 6 mprj_adr_o_user[2]
port 956 nsew signal output
rlabel metal2 s 44730 31200 44786 32400 6 mprj_adr_o_user[30]
port 957 nsew signal output
rlabel metal2 s 46018 31200 46074 32400 6 mprj_adr_o_user[31]
port 958 nsew signal output
rlabel metal2 s 8206 31200 8262 32400 6 mprj_adr_o_user[3]
port 959 nsew signal output
rlabel metal2 s 9954 31200 10010 32400 6 mprj_adr_o_user[4]
port 960 nsew signal output
rlabel metal2 s 11334 31200 11390 32400 6 mprj_adr_o_user[5]
port 961 nsew signal output
rlabel metal2 s 12622 31200 12678 32400 6 mprj_adr_o_user[6]
port 962 nsew signal output
rlabel metal2 s 14002 31200 14058 32400 6 mprj_adr_o_user[7]
port 963 nsew signal output
rlabel metal2 s 15290 31200 15346 32400 6 mprj_adr_o_user[8]
port 964 nsew signal output
rlabel metal2 s 16670 31200 16726 32400 6 mprj_adr_o_user[9]
port 965 nsew signal output
rlabel metal2 s 182914 -400 182970 800 6 mprj_cyc_o_core
port 966 nsew signal input
rlabel metal2 s 1490 31200 1546 32400 6 mprj_cyc_o_user
port 967 nsew signal output
rlabel metal2 s 184386 -400 184442 800 6 mprj_dat_i_core[0]
port 968 nsew signal output
rlabel metal2 s 196530 -400 196586 800 6 mprj_dat_i_core[10]
port 969 nsew signal output
rlabel metal2 s 197542 -400 197598 800 6 mprj_dat_i_core[11]
port 970 nsew signal output
rlabel metal2 s 198646 -400 198702 800 6 mprj_dat_i_core[12]
port 971 nsew signal output
rlabel metal2 s 199750 -400 199806 800 6 mprj_dat_i_core[13]
port 972 nsew signal output
rlabel metal2 s 200762 -400 200818 800 6 mprj_dat_i_core[14]
port 973 nsew signal output
rlabel metal2 s 201866 -400 201922 800 6 mprj_dat_i_core[15]
port 974 nsew signal output
rlabel metal2 s 202878 -400 202934 800 6 mprj_dat_i_core[16]
port 975 nsew signal output
rlabel metal2 s 203982 -400 204038 800 6 mprj_dat_i_core[17]
port 976 nsew signal output
rlabel metal2 s 205086 -400 205142 800 6 mprj_dat_i_core[18]
port 977 nsew signal output
rlabel metal2 s 206098 -400 206154 800 6 mprj_dat_i_core[19]
port 978 nsew signal output
rlabel metal2 s 185766 -400 185822 800 6 mprj_dat_i_core[1]
port 979 nsew signal output
rlabel metal2 s 207202 -400 207258 800 6 mprj_dat_i_core[20]
port 980 nsew signal output
rlabel metal2 s 208306 -400 208362 800 6 mprj_dat_i_core[21]
port 981 nsew signal output
rlabel metal2 s 209318 -400 209374 800 6 mprj_dat_i_core[22]
port 982 nsew signal output
rlabel metal2 s 210422 -400 210478 800 6 mprj_dat_i_core[23]
port 983 nsew signal output
rlabel metal2 s 211434 -400 211490 800 6 mprj_dat_i_core[24]
port 984 nsew signal output
rlabel metal2 s 212538 -400 212594 800 6 mprj_dat_i_core[25]
port 985 nsew signal output
rlabel metal2 s 213642 -400 213698 800 6 mprj_dat_i_core[26]
port 986 nsew signal output
rlabel metal2 s 214654 -400 214710 800 6 mprj_dat_i_core[27]
port 987 nsew signal output
rlabel metal2 s 215758 -400 215814 800 6 mprj_dat_i_core[28]
port 988 nsew signal output
rlabel metal2 s 216862 -400 216918 800 6 mprj_dat_i_core[29]
port 989 nsew signal output
rlabel metal2 s 187238 -400 187294 800 6 mprj_dat_i_core[2]
port 990 nsew signal output
rlabel metal2 s 217874 -400 217930 800 6 mprj_dat_i_core[30]
port 991 nsew signal output
rlabel metal2 s 218978 -400 219034 800 6 mprj_dat_i_core[31]
port 992 nsew signal output
rlabel metal2 s 188618 -400 188674 800 6 mprj_dat_i_core[3]
port 993 nsew signal output
rlabel metal2 s 190090 -400 190146 800 6 mprj_dat_i_core[4]
port 994 nsew signal output
rlabel metal2 s 191194 -400 191250 800 6 mprj_dat_i_core[5]
port 995 nsew signal output
rlabel metal2 s 192206 -400 192262 800 6 mprj_dat_i_core[6]
port 996 nsew signal output
rlabel metal2 s 193310 -400 193366 800 6 mprj_dat_i_core[7]
port 997 nsew signal output
rlabel metal2 s 194322 -400 194378 800 6 mprj_dat_i_core[8]
port 998 nsew signal output
rlabel metal2 s 195426 -400 195482 800 6 mprj_dat_i_core[9]
port 999 nsew signal output
rlabel metal2 s 3238 31200 3294 32400 6 mprj_dat_i_user[0]
port 1000 nsew signal input
rlabel metal2 s 18418 31200 18474 32400 6 mprj_dat_i_user[10]
port 1001 nsew signal input
rlabel metal2 s 19706 31200 19762 32400 6 mprj_dat_i_user[11]
port 1002 nsew signal input
rlabel metal2 s 21086 31200 21142 32400 6 mprj_dat_i_user[12]
port 1003 nsew signal input
rlabel metal2 s 22466 31200 22522 32400 6 mprj_dat_i_user[13]
port 1004 nsew signal input
rlabel metal2 s 23754 31200 23810 32400 6 mprj_dat_i_user[14]
port 1005 nsew signal input
rlabel metal2 s 25134 31200 25190 32400 6 mprj_dat_i_user[15]
port 1006 nsew signal input
rlabel metal2 s 26422 31200 26478 32400 6 mprj_dat_i_user[16]
port 1007 nsew signal input
rlabel metal2 s 27802 31200 27858 32400 6 mprj_dat_i_user[17]
port 1008 nsew signal input
rlabel metal2 s 29090 31200 29146 32400 6 mprj_dat_i_user[18]
port 1009 nsew signal input
rlabel metal2 s 30470 31200 30526 32400 6 mprj_dat_i_user[19]
port 1010 nsew signal input
rlabel metal2 s 5078 31200 5134 32400 6 mprj_dat_i_user[1]
port 1011 nsew signal input
rlabel metal2 s 31758 31200 31814 32400 6 mprj_dat_i_user[20]
port 1012 nsew signal input
rlabel metal2 s 33138 31200 33194 32400 6 mprj_dat_i_user[21]
port 1013 nsew signal input
rlabel metal2 s 34426 31200 34482 32400 6 mprj_dat_i_user[22]
port 1014 nsew signal input
rlabel metal2 s 35806 31200 35862 32400 6 mprj_dat_i_user[23]
port 1015 nsew signal input
rlabel metal2 s 37094 31200 37150 32400 6 mprj_dat_i_user[24]
port 1016 nsew signal input
rlabel metal2 s 38474 31200 38530 32400 6 mprj_dat_i_user[25]
port 1017 nsew signal input
rlabel metal2 s 39762 31200 39818 32400 6 mprj_dat_i_user[26]
port 1018 nsew signal input
rlabel metal2 s 41142 31200 41198 32400 6 mprj_dat_i_user[27]
port 1019 nsew signal input
rlabel metal2 s 42430 31200 42486 32400 6 mprj_dat_i_user[28]
port 1020 nsew signal input
rlabel metal2 s 43810 31200 43866 32400 6 mprj_dat_i_user[29]
port 1021 nsew signal input
rlabel metal2 s 6826 31200 6882 32400 6 mprj_dat_i_user[2]
port 1022 nsew signal input
rlabel metal2 s 45098 31200 45154 32400 6 mprj_dat_i_user[30]
port 1023 nsew signal input
rlabel metal2 s 46478 31200 46534 32400 6 mprj_dat_i_user[31]
port 1024 nsew signal input
rlabel metal2 s 8574 31200 8630 32400 6 mprj_dat_i_user[3]
port 1025 nsew signal input
rlabel metal2 s 10414 31200 10470 32400 6 mprj_dat_i_user[4]
port 1026 nsew signal input
rlabel metal2 s 11702 31200 11758 32400 6 mprj_dat_i_user[5]
port 1027 nsew signal input
rlabel metal2 s 13082 31200 13138 32400 6 mprj_dat_i_user[6]
port 1028 nsew signal input
rlabel metal2 s 14370 31200 14426 32400 6 mprj_dat_i_user[7]
port 1029 nsew signal input
rlabel metal2 s 15750 31200 15806 32400 6 mprj_dat_i_user[8]
port 1030 nsew signal input
rlabel metal2 s 17038 31200 17094 32400 6 mprj_dat_i_user[9]
port 1031 nsew signal input
rlabel metal2 s 184754 -400 184810 800 6 mprj_dat_o_core[0]
port 1032 nsew signal input
rlabel metal2 s 196898 -400 196954 800 6 mprj_dat_o_core[10]
port 1033 nsew signal input
rlabel metal2 s 197910 -400 197966 800 6 mprj_dat_o_core[11]
port 1034 nsew signal input
rlabel metal2 s 199014 -400 199070 800 6 mprj_dat_o_core[12]
port 1035 nsew signal input
rlabel metal2 s 200026 -400 200082 800 6 mprj_dat_o_core[13]
port 1036 nsew signal input
rlabel metal2 s 201130 -400 201186 800 6 mprj_dat_o_core[14]
port 1037 nsew signal input
rlabel metal2 s 202234 -400 202290 800 6 mprj_dat_o_core[15]
port 1038 nsew signal input
rlabel metal2 s 203246 -400 203302 800 6 mprj_dat_o_core[16]
port 1039 nsew signal input
rlabel metal2 s 204350 -400 204406 800 6 mprj_dat_o_core[17]
port 1040 nsew signal input
rlabel metal2 s 205454 -400 205510 800 6 mprj_dat_o_core[18]
port 1041 nsew signal input
rlabel metal2 s 206466 -400 206522 800 6 mprj_dat_o_core[19]
port 1042 nsew signal input
rlabel metal2 s 186134 -400 186190 800 6 mprj_dat_o_core[1]
port 1043 nsew signal input
rlabel metal2 s 207570 -400 207626 800 6 mprj_dat_o_core[20]
port 1044 nsew signal input
rlabel metal2 s 208582 -400 208638 800 6 mprj_dat_o_core[21]
port 1045 nsew signal input
rlabel metal2 s 209686 -400 209742 800 6 mprj_dat_o_core[22]
port 1046 nsew signal input
rlabel metal2 s 210790 -400 210846 800 6 mprj_dat_o_core[23]
port 1047 nsew signal input
rlabel metal2 s 211802 -400 211858 800 6 mprj_dat_o_core[24]
port 1048 nsew signal input
rlabel metal2 s 212906 -400 212962 800 6 mprj_dat_o_core[25]
port 1049 nsew signal input
rlabel metal2 s 214010 -400 214066 800 6 mprj_dat_o_core[26]
port 1050 nsew signal input
rlabel metal2 s 215022 -400 215078 800 6 mprj_dat_o_core[27]
port 1051 nsew signal input
rlabel metal2 s 216126 -400 216182 800 6 mprj_dat_o_core[28]
port 1052 nsew signal input
rlabel metal2 s 217138 -400 217194 800 6 mprj_dat_o_core[29]
port 1053 nsew signal input
rlabel metal2 s 187606 -400 187662 800 6 mprj_dat_o_core[2]
port 1054 nsew signal input
rlabel metal2 s 218242 -400 218298 800 6 mprj_dat_o_core[30]
port 1055 nsew signal input
rlabel metal2 s 219346 -400 219402 800 6 mprj_dat_o_core[31]
port 1056 nsew signal input
rlabel metal2 s 188986 -400 189042 800 6 mprj_dat_o_core[3]
port 1057 nsew signal input
rlabel metal2 s 190458 -400 190514 800 6 mprj_dat_o_core[4]
port 1058 nsew signal input
rlabel metal2 s 191470 -400 191526 800 6 mprj_dat_o_core[5]
port 1059 nsew signal input
rlabel metal2 s 192574 -400 192630 800 6 mprj_dat_o_core[6]
port 1060 nsew signal input
rlabel metal2 s 193678 -400 193734 800 6 mprj_dat_o_core[7]
port 1061 nsew signal input
rlabel metal2 s 194690 -400 194746 800 6 mprj_dat_o_core[8]
port 1062 nsew signal input
rlabel metal2 s 195794 -400 195850 800 6 mprj_dat_o_core[9]
port 1063 nsew signal input
rlabel metal2 s 3698 31200 3754 32400 6 mprj_dat_o_user[0]
port 1064 nsew signal output
rlabel metal2 s 18878 31200 18934 32400 6 mprj_dat_o_user[10]
port 1065 nsew signal output
rlabel metal2 s 20166 31200 20222 32400 6 mprj_dat_o_user[11]
port 1066 nsew signal output
rlabel metal2 s 21546 31200 21602 32400 6 mprj_dat_o_user[12]
port 1067 nsew signal output
rlabel metal2 s 22834 31200 22890 32400 6 mprj_dat_o_user[13]
port 1068 nsew signal output
rlabel metal2 s 24214 31200 24270 32400 6 mprj_dat_o_user[14]
port 1069 nsew signal output
rlabel metal2 s 25502 31200 25558 32400 6 mprj_dat_o_user[15]
port 1070 nsew signal output
rlabel metal2 s 26882 31200 26938 32400 6 mprj_dat_o_user[16]
port 1071 nsew signal output
rlabel metal2 s 28170 31200 28226 32400 6 mprj_dat_o_user[17]
port 1072 nsew signal output
rlabel metal2 s 29550 31200 29606 32400 6 mprj_dat_o_user[18]
port 1073 nsew signal output
rlabel metal2 s 30838 31200 30894 32400 6 mprj_dat_o_user[19]
port 1074 nsew signal output
rlabel metal2 s 5538 31200 5594 32400 6 mprj_dat_o_user[1]
port 1075 nsew signal output
rlabel metal2 s 32218 31200 32274 32400 6 mprj_dat_o_user[20]
port 1076 nsew signal output
rlabel metal2 s 33598 31200 33654 32400 6 mprj_dat_o_user[21]
port 1077 nsew signal output
rlabel metal2 s 34886 31200 34942 32400 6 mprj_dat_o_user[22]
port 1078 nsew signal output
rlabel metal2 s 36266 31200 36322 32400 6 mprj_dat_o_user[23]
port 1079 nsew signal output
rlabel metal2 s 37554 31200 37610 32400 6 mprj_dat_o_user[24]
port 1080 nsew signal output
rlabel metal2 s 38934 31200 38990 32400 6 mprj_dat_o_user[25]
port 1081 nsew signal output
rlabel metal2 s 40222 31200 40278 32400 6 mprj_dat_o_user[26]
port 1082 nsew signal output
rlabel metal2 s 41602 31200 41658 32400 6 mprj_dat_o_user[27]
port 1083 nsew signal output
rlabel metal2 s 42890 31200 42946 32400 6 mprj_dat_o_user[28]
port 1084 nsew signal output
rlabel metal2 s 44270 31200 44326 32400 6 mprj_dat_o_user[29]
port 1085 nsew signal output
rlabel metal2 s 7286 31200 7342 32400 6 mprj_dat_o_user[2]
port 1086 nsew signal output
rlabel metal2 s 45558 31200 45614 32400 6 mprj_dat_o_user[30]
port 1087 nsew signal output
rlabel metal2 s 46938 31200 46994 32400 6 mprj_dat_o_user[31]
port 1088 nsew signal output
rlabel metal2 s 9034 31200 9090 32400 6 mprj_dat_o_user[3]
port 1089 nsew signal output
rlabel metal2 s 10874 31200 10930 32400 6 mprj_dat_o_user[4]
port 1090 nsew signal output
rlabel metal2 s 12162 31200 12218 32400 6 mprj_dat_o_user[5]
port 1091 nsew signal output
rlabel metal2 s 13542 31200 13598 32400 6 mprj_dat_o_user[6]
port 1092 nsew signal output
rlabel metal2 s 14830 31200 14886 32400 6 mprj_dat_o_user[7]
port 1093 nsew signal output
rlabel metal2 s 16210 31200 16266 32400 6 mprj_dat_o_user[8]
port 1094 nsew signal output
rlabel metal2 s 17498 31200 17554 32400 6 mprj_dat_o_user[9]
port 1095 nsew signal output
rlabel metal2 s 219714 -400 219770 800 6 mprj_iena_wb
port 1096 nsew signal input
rlabel metal2 s 185122 -400 185178 800 6 mprj_sel_o_core[0]
port 1097 nsew signal input
rlabel metal2 s 186502 -400 186558 800 6 mprj_sel_o_core[1]
port 1098 nsew signal input
rlabel metal2 s 187974 -400 188030 800 6 mprj_sel_o_core[2]
port 1099 nsew signal input
rlabel metal2 s 189354 -400 189410 800 6 mprj_sel_o_core[3]
port 1100 nsew signal input
rlabel metal2 s 4158 31200 4214 32400 6 mprj_sel_o_user[0]
port 1101 nsew signal output
rlabel metal2 s 5906 31200 5962 32400 6 mprj_sel_o_user[1]
port 1102 nsew signal output
rlabel metal2 s 7746 31200 7802 32400 6 mprj_sel_o_user[2]
port 1103 nsew signal output
rlabel metal2 s 9494 31200 9550 32400 6 mprj_sel_o_user[3]
port 1104 nsew signal output
rlabel metal2 s 183282 -400 183338 800 6 mprj_stb_o_core
port 1105 nsew signal input
rlabel metal2 s 1950 31200 2006 32400 6 mprj_stb_o_user
port 1106 nsew signal output
rlabel metal2 s 183650 -400 183706 800 6 mprj_we_o_core
port 1107 nsew signal input
rlabel metal2 s 2410 31200 2466 32400 6 mprj_we_o_user
port 1108 nsew signal output
rlabel metal3 s 219200 1504 220400 1624 6 user1_vcc_powergood
port 1109 nsew signal output
rlabel metal3 s 219200 4632 220400 4752 6 user1_vdd_powergood
port 1110 nsew signal output
rlabel metal3 s 219200 7896 220400 8016 6 user2_vcc_powergood
port 1111 nsew signal output
rlabel metal3 s 219200 11024 220400 11144 6 user2_vdd_powergood
port 1112 nsew signal output
rlabel metal2 s 202 31200 258 32400 6 user_clock
port 1113 nsew signal output
rlabel metal2 s 218334 31200 218390 32400 6 user_clock2
port 1114 nsew signal output
rlabel metal3 s 219200 14288 220400 14408 6 user_irq[0]
port 1115 nsew signal output
rlabel metal3 s 219200 17416 220400 17536 6 user_irq[1]
port 1116 nsew signal output
rlabel metal3 s 219200 20680 220400 20800 6 user_irq[2]
port 1117 nsew signal output
rlabel metal2 s 218794 31200 218850 32400 6 user_irq_core[0]
port 1118 nsew signal input
rlabel metal2 s 219254 31200 219310 32400 6 user_irq_core[1]
port 1119 nsew signal input
rlabel metal2 s 219714 31200 219770 32400 6 user_irq_core[2]
port 1120 nsew signal input
rlabel metal3 s 219200 23808 220400 23928 6 user_irq_ena[0]
port 1121 nsew signal input
rlabel metal3 s 219200 27072 220400 27192 6 user_irq_ena[1]
port 1122 nsew signal input
rlabel metal3 s 219200 30200 220400 30320 6 user_irq_ena[2]
port 1123 nsew signal input
rlabel metal2 s 570 31200 626 32400 6 user_reset
port 1124 nsew signal output
rlabel metal4 s 4014 1040 4194 30512 6 vccd
port 1125 nsew power input
rlabel metal4 s 34114 1040 34294 30512 6 vccd
port 1125 nsew power input
rlabel metal4 s 64214 1040 64394 30512 6 vccd
port 1125 nsew power input
rlabel metal4 s 94314 1040 94494 30512 6 vccd
port 1125 nsew power input
rlabel metal4 s 124414 1040 124594 30512 6 vccd
port 1125 nsew power input
rlabel metal4 s 154514 1040 154694 30512 6 vccd
port 1125 nsew power input
rlabel metal4 s 184614 1040 184794 30512 6 vccd
port 1125 nsew power input
rlabel metal4 s 214714 1040 214894 30512 6 vccd
port 1125 nsew power input
rlabel metal4 s 4834 1088 5014 30464 6 vccd1
port 1126 nsew power input
rlabel metal4 s 34934 1088 35114 30464 6 vccd1
port 1126 nsew power input
rlabel metal4 s 65034 1088 65214 30464 6 vccd1
port 1126 nsew power input
rlabel metal4 s 95134 1088 95314 30464 6 vccd1
port 1126 nsew power input
rlabel metal4 s 125234 1088 125414 30464 6 vccd1
port 1126 nsew power input
rlabel metal4 s 155334 1088 155514 30464 6 vccd1
port 1126 nsew power input
rlabel metal4 s 185434 1088 185614 30464 6 vccd1
port 1126 nsew power input
rlabel metal4 s 215534 1088 215714 30464 6 vccd1
port 1126 nsew power input
rlabel metal4 s 5654 1088 5834 30464 6 vccd2
port 1127 nsew power input
rlabel metal4 s 35754 1088 35934 30464 6 vccd2
port 1127 nsew power input
rlabel metal4 s 65854 1088 66034 30464 6 vccd2
port 1127 nsew power input
rlabel metal4 s 95954 1088 96134 30464 6 vccd2
port 1127 nsew power input
rlabel metal4 s 126054 1088 126234 30464 6 vccd2
port 1127 nsew power input
rlabel metal4 s 156154 1088 156334 30464 6 vccd2
port 1127 nsew power input
rlabel metal4 s 186254 1088 186434 30464 6 vccd2
port 1127 nsew power input
rlabel metal4 s 216354 1088 216534 30464 6 vccd2
port 1127 nsew power input
rlabel metal4 s 186814 1088 186994 30464 6 vdda1
port 1128 nsew power input
rlabel metal4 s 216914 1088 217094 30464 6 vdda1
port 1128 nsew power input
rlabel metal4 s 187414 1088 187594 30464 6 vdda2
port 1129 nsew power input
rlabel metal4 s 217514 1088 217694 30464 6 vdda2
port 1129 nsew power input
rlabel metal4 s 201864 1088 202044 30464 6 vssa1
port 1130 nsew ground input
rlabel metal4 s 202464 1088 202644 30464 6 vssa2
port 1131 nsew ground input
rlabel metal4 s 19064 1040 19244 30512 6 vssd
port 1132 nsew ground input
rlabel metal4 s 49164 1040 49344 30512 6 vssd
port 1132 nsew ground input
rlabel metal4 s 79264 1040 79444 30512 6 vssd
port 1132 nsew ground input
rlabel metal4 s 109364 1040 109544 30512 6 vssd
port 1132 nsew ground input
rlabel metal4 s 139464 1040 139644 30512 6 vssd
port 1132 nsew ground input
rlabel metal4 s 169564 1040 169744 30512 6 vssd
port 1132 nsew ground input
rlabel metal4 s 199664 1040 199844 30512 6 vssd
port 1132 nsew ground input
rlabel metal4 s 19884 1088 20064 30464 6 vssd1
port 1133 nsew ground input
rlabel metal4 s 49984 1088 50164 30464 6 vssd1
port 1133 nsew ground input
rlabel metal4 s 80084 1088 80264 30464 6 vssd1
port 1133 nsew ground input
rlabel metal4 s 110184 1088 110364 30464 6 vssd1
port 1133 nsew ground input
rlabel metal4 s 140284 1088 140464 30464 6 vssd1
port 1133 nsew ground input
rlabel metal4 s 170384 1088 170564 30464 6 vssd1
port 1133 nsew ground input
rlabel metal4 s 200484 1088 200664 30464 6 vssd1
port 1133 nsew ground input
rlabel metal4 s 20704 1088 20884 30464 6 vssd2
port 1134 nsew ground input
rlabel metal4 s 50804 1088 50984 30464 6 vssd2
port 1134 nsew ground input
rlabel metal4 s 80904 1088 81084 30464 6 vssd2
port 1134 nsew ground input
rlabel metal4 s 111004 1088 111184 30464 6 vssd2
port 1134 nsew ground input
rlabel metal4 s 141104 1088 141284 30464 6 vssd2
port 1134 nsew ground input
rlabel metal4 s 171204 1088 171384 30464 6 vssd2
port 1134 nsew ground input
rlabel metal4 s 201304 1088 201484 30464 6 vssd2
port 1134 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 220000 32000
string LEFview TRUE
string GDS_FILE /home/marwan/caravel/openlane/mgmt_protect/runs/mgmt_protect/results/magic/mgmt_protect.gds
string GDS_END 8991246
string GDS_START 298528
<< end >>

