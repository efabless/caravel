VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mgmt_protect_hv
  CLASS BLOCK ;
  FOREIGN mgmt_protect_hv ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 20.000 ;
  PIN mprj2_vdd_logic1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.510 4.000 5.110 ;
    END
  END mprj2_vdd_logic1
  PIN mprj_vdd_logic1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.130 4.000 14.730 ;
    END
  END mprj_vdd_logic1
  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 94.650 3.815 94.950 16.535 ;
    END
  END vccd
  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 14.650 3.815 14.950 16.535 ;
    END
  END vccd
  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 4.800 15.465 149.760 15.765 ;
    END
  END vccd
  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 4.800 4.665 149.760 4.965 ;
    END
  END vccd
  PIN vssd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 134.650 3.815 134.950 16.535 ;
    END
  END vssd
  PIN vssd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 54.650 3.815 54.950 16.535 ;
    END
  END vssd
  PIN vssd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 4.800 10.065 149.760 10.365 ;
    END
  END vssd
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 96.650 4.070 96.950 16.280 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 16.650 4.070 16.950 16.280 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 4.800 6.920 149.760 7.220 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 136.650 4.070 136.950 16.280 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 56.650 4.070 56.950 16.280 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 4.800 12.320 149.760 12.620 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 98.650 4.070 98.950 16.280 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 18.650 4.070 18.950 16.280 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 4.800 8.920 149.760 9.220 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 138.650 4.070 138.950 16.280 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 58.650 4.070 58.950 16.280 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 4.800 14.320 149.760 14.620 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 4.800 3.985 149.760 16.365 ;
      LAYER met1 ;
        RECT 3.920 3.815 149.760 16.535 ;
      LAYER met2 ;
        RECT 3.940 4.625 14.370 14.855 ;
        RECT 15.230 4.625 16.370 14.855 ;
        RECT 17.230 4.625 18.370 14.855 ;
        RECT 19.230 4.625 54.370 14.855 ;
        RECT 55.230 4.625 56.370 14.855 ;
        RECT 57.230 4.625 58.370 14.855 ;
        RECT 59.230 4.625 94.370 14.855 ;
        RECT 95.230 4.625 96.370 14.855 ;
        RECT 97.230 4.625 98.370 14.855 ;
        RECT 99.230 4.625 134.370 14.855 ;
        RECT 135.230 4.625 136.370 14.855 ;
        RECT 137.230 4.625 138.370 14.855 ;
        RECT 139.230 4.625 146.560 14.855 ;
      LAYER met3 ;
        RECT 4.000 15.130 4.400 15.780 ;
        RECT 4.400 15.020 146.585 15.065 ;
        RECT 4.400 13.730 146.585 13.920 ;
        RECT 4.000 13.020 146.585 13.730 ;
        RECT 4.000 11.920 4.400 13.020 ;
        RECT 4.000 10.765 146.585 11.920 ;
        RECT 4.000 9.665 4.400 10.765 ;
        RECT 4.000 9.620 146.585 9.665 ;
        RECT 4.000 8.520 4.400 9.620 ;
        RECT 4.000 7.620 146.585 8.520 ;
        RECT 4.000 6.520 4.400 7.620 ;
        RECT 4.000 5.510 146.585 6.520 ;
        RECT 4.400 5.365 146.585 5.510 ;
  END
END mgmt_protect_hv
END LIBRARY

