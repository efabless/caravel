magic
tech sky130A
magscale 1 2
timestamp 1666117611
<< metal1 >>
rect 366174 1027828 366180 1027880
rect 366232 1027868 366238 1027880
rect 366542 1027868 366548 1027880
rect 366232 1027840 366548 1027868
rect 366232 1027828 366238 1027840
rect 366542 1027828 366548 1027840
rect 366600 1027828 366606 1027880
rect 366174 1024360 366180 1024412
rect 366232 1024400 366238 1024412
rect 366542 1024400 366548 1024412
rect 366232 1024372 366548 1024400
rect 366232 1024360 366238 1024372
rect 366542 1024360 366548 1024372
rect 366600 1024360 366606 1024412
rect 426342 1007088 426348 1007140
rect 426400 1007128 426406 1007140
rect 437474 1007128 437480 1007140
rect 426400 1007100 437480 1007128
rect 426400 1007088 426406 1007100
rect 437474 1007088 437480 1007100
rect 437532 1007088 437538 1007140
rect 358538 1006952 358544 1007004
rect 358596 1006992 358602 1007004
rect 373258 1006992 373264 1007004
rect 358596 1006964 373264 1006992
rect 358596 1006952 358602 1006964
rect 373258 1006952 373264 1006964
rect 373316 1006952 373322 1007004
rect 553946 1006952 553952 1007004
rect 554004 1006992 554010 1007004
rect 562318 1006992 562324 1007004
rect 554004 1006964 562324 1006992
rect 554004 1006952 554010 1006964
rect 562318 1006952 562324 1006964
rect 562376 1006952 562382 1007004
rect 505002 1006884 505008 1006936
rect 505060 1006924 505066 1006936
rect 513374 1006924 513380 1006936
rect 505060 1006896 513380 1006924
rect 505060 1006884 505066 1006896
rect 513374 1006884 513380 1006896
rect 513432 1006884 513438 1006936
rect 359366 1006816 359372 1006868
rect 359424 1006856 359430 1006868
rect 380158 1006856 380164 1006868
rect 359424 1006828 380164 1006856
rect 359424 1006816 359430 1006828
rect 380158 1006816 380164 1006828
rect 380216 1006816 380222 1006868
rect 555970 1006816 555976 1006868
rect 556028 1006856 556034 1006868
rect 569402 1006856 569408 1006868
rect 556028 1006828 569408 1006856
rect 556028 1006816 556034 1006828
rect 569402 1006816 569408 1006828
rect 569460 1006816 569466 1006868
rect 429194 1006748 429200 1006800
rect 429252 1006788 429258 1006800
rect 429252 1006760 441614 1006788
rect 429252 1006748 429258 1006760
rect 144178 1006680 144184 1006732
rect 144236 1006720 144242 1006732
rect 150250 1006720 150256 1006732
rect 144236 1006692 150256 1006720
rect 144236 1006680 144242 1006692
rect 150250 1006680 150256 1006692
rect 150308 1006680 150314 1006732
rect 161934 1006680 161940 1006732
rect 161992 1006720 161998 1006732
rect 164878 1006720 164884 1006732
rect 161992 1006692 164884 1006720
rect 161992 1006680 161998 1006692
rect 164878 1006680 164884 1006692
rect 164936 1006680 164942 1006732
rect 360194 1006680 360200 1006732
rect 360252 1006720 360258 1006732
rect 360252 1006692 372108 1006720
rect 360252 1006680 360258 1006692
rect 94498 1006544 94504 1006596
rect 94556 1006584 94562 1006596
rect 101950 1006584 101956 1006596
rect 94556 1006556 101956 1006584
rect 94556 1006544 94562 1006556
rect 101950 1006544 101956 1006556
rect 102008 1006544 102014 1006596
rect 145742 1006544 145748 1006596
rect 145800 1006584 145806 1006596
rect 153746 1006584 153752 1006596
rect 145800 1006556 153752 1006584
rect 145800 1006544 145806 1006556
rect 153746 1006544 153752 1006556
rect 153804 1006544 153810 1006596
rect 157426 1006544 157432 1006596
rect 157484 1006584 157490 1006596
rect 166258 1006584 166264 1006596
rect 157484 1006556 166264 1006584
rect 157484 1006544 157490 1006556
rect 166258 1006544 166264 1006556
rect 166316 1006544 166322 1006596
rect 173158 1006584 173164 1006596
rect 171106 1006556 173164 1006584
rect 93118 1006408 93124 1006460
rect 93176 1006448 93182 1006460
rect 98270 1006448 98276 1006460
rect 93176 1006420 98276 1006448
rect 93176 1006408 93182 1006420
rect 98270 1006408 98276 1006420
rect 98328 1006408 98334 1006460
rect 145558 1006408 145564 1006460
rect 145616 1006448 145622 1006460
rect 152918 1006448 152924 1006460
rect 145616 1006420 152924 1006448
rect 145616 1006408 145622 1006420
rect 152918 1006408 152924 1006420
rect 152976 1006408 152982 1006460
rect 160278 1006408 160284 1006460
rect 160336 1006448 160342 1006460
rect 161934 1006448 161940 1006460
rect 160336 1006420 161940 1006448
rect 160336 1006408 160342 1006420
rect 161934 1006408 161940 1006420
rect 161992 1006408 161998 1006460
rect 162762 1006408 162768 1006460
rect 162820 1006448 162826 1006460
rect 171106 1006448 171134 1006556
rect 173158 1006544 173164 1006556
rect 173216 1006544 173222 1006596
rect 364886 1006544 364892 1006596
rect 364944 1006584 364950 1006596
rect 371878 1006584 371884 1006596
rect 364944 1006556 371884 1006584
rect 364944 1006544 364950 1006556
rect 371878 1006544 371884 1006556
rect 371936 1006544 371942 1006596
rect 162820 1006420 171134 1006448
rect 162820 1006408 162826 1006420
rect 247678 1006408 247684 1006460
rect 247736 1006448 247742 1006460
rect 256142 1006448 256148 1006460
rect 247736 1006420 256148 1006448
rect 247736 1006408 247742 1006420
rect 256142 1006408 256148 1006420
rect 256200 1006408 256206 1006460
rect 354858 1006408 354864 1006460
rect 354916 1006448 354922 1006460
rect 363598 1006448 363604 1006460
rect 354916 1006420 363604 1006448
rect 354916 1006408 354922 1006420
rect 363598 1006408 363604 1006420
rect 363656 1006408 363662 1006460
rect 372080 1006448 372108 1006692
rect 431678 1006652 431684 1006664
rect 412606 1006624 431684 1006652
rect 374638 1006448 374644 1006460
rect 372080 1006420 374644 1006448
rect 374638 1006408 374644 1006420
rect 374696 1006408 374702 1006460
rect 101398 1006272 101404 1006324
rect 101456 1006312 101462 1006324
rect 103974 1006312 103980 1006324
rect 101456 1006284 103980 1006312
rect 101456 1006272 101462 1006284
rect 103974 1006272 103980 1006284
rect 104032 1006272 104038 1006324
rect 108482 1006272 108488 1006324
rect 108540 1006312 108546 1006324
rect 126238 1006312 126244 1006324
rect 108540 1006284 126244 1006312
rect 108540 1006272 108546 1006284
rect 126238 1006272 126244 1006284
rect 126296 1006272 126302 1006324
rect 152090 1006312 152096 1006324
rect 151786 1006284 152096 1006312
rect 144362 1006204 144368 1006256
rect 144420 1006244 144426 1006256
rect 151262 1006244 151268 1006256
rect 144420 1006216 151268 1006244
rect 144420 1006204 144426 1006216
rect 151262 1006204 151268 1006216
rect 151320 1006204 151326 1006256
rect 92474 1006136 92480 1006188
rect 92532 1006176 92538 1006188
rect 92532 1006148 99696 1006176
rect 92532 1006136 92538 1006148
rect 94682 1006000 94688 1006052
rect 94740 1006040 94746 1006052
rect 99466 1006040 99472 1006052
rect 94740 1006012 99472 1006040
rect 94740 1006000 94746 1006012
rect 99466 1006000 99472 1006012
rect 99524 1006000 99530 1006052
rect 99668 1006040 99696 1006148
rect 101582 1006136 101588 1006188
rect 101640 1006176 101646 1006188
rect 104802 1006176 104808 1006188
rect 101640 1006148 104808 1006176
rect 101640 1006136 101646 1006148
rect 104802 1006136 104808 1006148
rect 104860 1006136 104866 1006188
rect 106826 1006136 106832 1006188
rect 106884 1006176 106890 1006188
rect 113818 1006176 113824 1006188
rect 106884 1006148 113824 1006176
rect 106884 1006136 106890 1006148
rect 113818 1006136 113824 1006148
rect 113876 1006136 113882 1006188
rect 148870 1006068 148876 1006120
rect 148928 1006108 148934 1006120
rect 150066 1006108 150072 1006120
rect 148928 1006080 150072 1006108
rect 148928 1006068 148934 1006080
rect 150066 1006068 150072 1006080
rect 150124 1006068 150130 1006120
rect 150250 1006068 150256 1006120
rect 150308 1006108 150314 1006120
rect 151786 1006108 151814 1006284
rect 152090 1006272 152096 1006284
rect 152148 1006272 152154 1006324
rect 158254 1006272 158260 1006324
rect 158312 1006312 158318 1006324
rect 171778 1006312 171784 1006324
rect 158312 1006284 171784 1006312
rect 158312 1006272 158318 1006284
rect 171778 1006272 171784 1006284
rect 171836 1006272 171842 1006324
rect 255958 1006272 255964 1006324
rect 256016 1006312 256022 1006324
rect 258994 1006312 259000 1006324
rect 256016 1006284 259000 1006312
rect 256016 1006272 256022 1006284
rect 258994 1006272 259000 1006284
rect 259052 1006272 259058 1006324
rect 301498 1006272 301504 1006324
rect 301556 1006312 301562 1006324
rect 307754 1006312 307760 1006324
rect 301556 1006284 307760 1006312
rect 301556 1006272 301562 1006284
rect 307754 1006272 307760 1006284
rect 307812 1006272 307818 1006324
rect 314654 1006272 314660 1006324
rect 314712 1006312 314718 1006324
rect 320818 1006312 320824 1006324
rect 314712 1006284 320824 1006312
rect 314712 1006272 314718 1006284
rect 320818 1006272 320824 1006284
rect 320876 1006272 320882 1006324
rect 361390 1006272 361396 1006324
rect 361448 1006312 361454 1006324
rect 361448 1006284 369256 1006312
rect 361448 1006272 361454 1006284
rect 158622 1006136 158628 1006188
rect 158680 1006176 158686 1006188
rect 162762 1006176 162768 1006188
rect 158680 1006148 162768 1006176
rect 158680 1006136 158686 1006148
rect 162762 1006136 162768 1006148
rect 162820 1006136 162826 1006188
rect 166258 1006136 166264 1006188
rect 166316 1006176 166322 1006188
rect 175918 1006176 175924 1006188
rect 166316 1006148 175924 1006176
rect 166316 1006136 166322 1006148
rect 175918 1006136 175924 1006148
rect 175976 1006136 175982 1006188
rect 210418 1006136 210424 1006188
rect 210476 1006176 210482 1006188
rect 228358 1006176 228364 1006188
rect 210476 1006148 228364 1006176
rect 210476 1006136 210482 1006148
rect 228358 1006136 228364 1006148
rect 228416 1006136 228422 1006188
rect 249058 1006136 249064 1006188
rect 249116 1006176 249122 1006188
rect 257338 1006176 257344 1006188
rect 249116 1006148 257344 1006176
rect 249116 1006136 249122 1006148
rect 257338 1006136 257344 1006148
rect 257396 1006136 257402 1006188
rect 262674 1006136 262680 1006188
rect 262732 1006176 262738 1006188
rect 269758 1006176 269764 1006188
rect 262732 1006148 269764 1006176
rect 262732 1006136 262738 1006148
rect 269758 1006136 269764 1006148
rect 269816 1006136 269822 1006188
rect 298738 1006136 298744 1006188
rect 298796 1006176 298802 1006188
rect 304902 1006176 304908 1006188
rect 298796 1006148 304908 1006176
rect 298796 1006136 298802 1006148
rect 304902 1006136 304908 1006148
rect 304960 1006136 304966 1006188
rect 360562 1006136 360568 1006188
rect 360620 1006176 360626 1006188
rect 360620 1006148 363000 1006176
rect 360620 1006136 360626 1006148
rect 150308 1006080 151814 1006108
rect 150308 1006068 150314 1006080
rect 103146 1006040 103152 1006052
rect 99668 1006012 103152 1006040
rect 103146 1006000 103152 1006012
rect 103204 1006000 103210 1006052
rect 105998 1006000 106004 1006052
rect 106056 1006040 106062 1006052
rect 124858 1006040 124864 1006052
rect 106056 1006012 124864 1006040
rect 106056 1006000 106062 1006012
rect 124858 1006000 124864 1006012
rect 124916 1006000 124922 1006052
rect 153930 1006000 153936 1006052
rect 153988 1006040 153994 1006052
rect 158254 1006040 158260 1006052
rect 153988 1006012 158260 1006040
rect 153988 1006000 153994 1006012
rect 158254 1006000 158260 1006012
rect 158312 1006000 158318 1006052
rect 159450 1006000 159456 1006052
rect 159508 1006040 159514 1006052
rect 177298 1006040 177304 1006052
rect 159508 1006012 177304 1006040
rect 159508 1006000 159514 1006012
rect 177298 1006000 177304 1006012
rect 177356 1006000 177362 1006052
rect 195146 1006000 195152 1006052
rect 195204 1006040 195210 1006052
rect 201034 1006040 201040 1006052
rect 195204 1006012 201040 1006040
rect 195204 1006000 195210 1006012
rect 201034 1006000 201040 1006012
rect 201092 1006000 201098 1006052
rect 208394 1006000 208400 1006052
rect 208452 1006040 208458 1006052
rect 229738 1006040 229744 1006052
rect 208452 1006012 229744 1006040
rect 208452 1006000 208458 1006012
rect 229738 1006000 229744 1006012
rect 229796 1006000 229802 1006052
rect 257338 1006000 257344 1006052
rect 257396 1006040 257402 1006052
rect 258166 1006040 258172 1006052
rect 257396 1006012 258172 1006040
rect 257396 1006000 257402 1006012
rect 258166 1006000 258172 1006012
rect 258224 1006000 258230 1006052
rect 261846 1006000 261852 1006052
rect 261904 1006040 261910 1006052
rect 279418 1006040 279424 1006052
rect 261904 1006012 279424 1006040
rect 261904 1006000 261910 1006012
rect 279418 1006000 279424 1006012
rect 279476 1006000 279482 1006052
rect 298922 1006000 298928 1006052
rect 298980 1006040 298986 1006052
rect 298980 1006012 303108 1006040
rect 298980 1006000 298986 1006012
rect 303080 1005904 303108 1006012
rect 303246 1006000 303252 1006052
rect 303304 1006040 303310 1006052
rect 304074 1006040 304080 1006052
rect 303304 1006012 304080 1006040
rect 303304 1006000 303310 1006012
rect 304074 1006000 304080 1006012
rect 304132 1006000 304138 1006052
rect 311802 1006040 311808 1006052
rect 304276 1006012 311808 1006040
rect 304276 1005904 304304 1006012
rect 311802 1006000 311808 1006012
rect 311860 1006000 311866 1006052
rect 314654 1006000 314660 1006052
rect 314712 1006040 314718 1006052
rect 319438 1006040 319444 1006052
rect 314712 1006012 319444 1006040
rect 314712 1006000 314718 1006012
rect 319438 1006000 319444 1006012
rect 319496 1006000 319502 1006052
rect 358538 1006000 358544 1006052
rect 358596 1006040 358602 1006052
rect 362218 1006040 362224 1006052
rect 358596 1006012 362224 1006040
rect 358596 1006000 358602 1006012
rect 362218 1006000 362224 1006012
rect 362276 1006000 362282 1006052
rect 362972 1006040 363000 1006148
rect 363414 1006136 363420 1006188
rect 363472 1006176 363478 1006188
rect 369228 1006176 369256 1006284
rect 402238 1006272 402244 1006324
rect 402296 1006312 402302 1006324
rect 412606 1006312 412634 1006624
rect 431678 1006612 431684 1006624
rect 431736 1006612 431742 1006664
rect 441586 1006584 441614 1006760
rect 507854 1006680 507860 1006732
rect 507912 1006720 507918 1006732
rect 520918 1006720 520924 1006732
rect 507912 1006692 520924 1006720
rect 507912 1006680 507918 1006692
rect 520918 1006680 520924 1006692
rect 520976 1006680 520982 1006732
rect 556798 1006680 556804 1006732
rect 556856 1006720 556862 1006732
rect 564434 1006720 564440 1006732
rect 556856 1006692 564440 1006720
rect 556856 1006680 556862 1006692
rect 564434 1006680 564440 1006692
rect 564492 1006680 564498 1006732
rect 469858 1006584 469864 1006596
rect 441586 1006556 469864 1006584
rect 469858 1006544 469864 1006556
rect 469916 1006544 469922 1006596
rect 505370 1006544 505376 1006596
rect 505428 1006584 505434 1006596
rect 518158 1006584 518164 1006596
rect 505428 1006556 518164 1006584
rect 505428 1006544 505434 1006556
rect 518158 1006544 518164 1006556
rect 518216 1006544 518222 1006596
rect 428366 1006476 428372 1006528
rect 428424 1006516 428430 1006528
rect 440878 1006516 440884 1006528
rect 428424 1006488 440884 1006516
rect 428424 1006476 428430 1006488
rect 440878 1006476 440884 1006488
rect 440936 1006476 440942 1006528
rect 506198 1006408 506204 1006460
rect 506256 1006448 506262 1006460
rect 506256 1006420 518894 1006448
rect 506256 1006408 506262 1006420
rect 402296 1006284 412634 1006312
rect 402296 1006272 402302 1006284
rect 427538 1006272 427544 1006324
rect 427596 1006312 427602 1006324
rect 427596 1006284 437474 1006312
rect 427596 1006272 427602 1006284
rect 377398 1006176 377404 1006188
rect 363472 1006148 369164 1006176
rect 369228 1006148 377404 1006176
rect 363472 1006136 363478 1006148
rect 364886 1006040 364892 1006052
rect 362972 1006012 364892 1006040
rect 364886 1006000 364892 1006012
rect 364944 1006000 364950 1006052
rect 365070 1006000 365076 1006052
rect 365128 1006040 365134 1006052
rect 367738 1006040 367744 1006052
rect 365128 1006012 367744 1006040
rect 365128 1006000 365134 1006012
rect 367738 1006000 367744 1006012
rect 367796 1006000 367802 1006052
rect 369136 1006040 369164 1006148
rect 377398 1006136 377404 1006148
rect 377456 1006136 377462 1006188
rect 429194 1006176 429200 1006188
rect 412606 1006148 429200 1006176
rect 382826 1006040 382832 1006052
rect 369136 1006012 382832 1006040
rect 382826 1006000 382832 1006012
rect 382884 1006000 382890 1006052
rect 400858 1006000 400864 1006052
rect 400916 1006040 400922 1006052
rect 412606 1006040 412634 1006148
rect 429194 1006136 429200 1006148
rect 429252 1006136 429258 1006188
rect 437446 1006176 437474 1006284
rect 451918 1006176 451924 1006188
rect 437446 1006148 451924 1006176
rect 451918 1006136 451924 1006148
rect 451976 1006136 451982 1006188
rect 400916 1006012 412634 1006040
rect 400916 1006000 400922 1006012
rect 425146 1006000 425152 1006052
rect 425204 1006040 425210 1006052
rect 429746 1006040 429752 1006052
rect 425204 1006012 429752 1006040
rect 425204 1006000 425210 1006012
rect 429746 1006000 429752 1006012
rect 429804 1006000 429810 1006052
rect 431678 1006000 431684 1006052
rect 431736 1006040 431742 1006052
rect 471238 1006040 471244 1006052
rect 431736 1006012 471244 1006040
rect 431736 1006000 431742 1006012
rect 471238 1006000 471244 1006012
rect 471296 1006000 471302 1006052
rect 496722 1006000 496728 1006052
rect 496780 1006040 496786 1006052
rect 498838 1006040 498844 1006052
rect 496780 1006012 498844 1006040
rect 496780 1006000 496786 1006012
rect 498838 1006000 498844 1006012
rect 498896 1006000 498902 1006052
rect 518866 1006040 518894 1006420
rect 555142 1006408 555148 1006460
rect 555200 1006448 555206 1006460
rect 570322 1006448 570328 1006460
rect 555200 1006420 570328 1006448
rect 555200 1006408 555206 1006420
rect 570322 1006408 570328 1006420
rect 570380 1006408 570386 1006460
rect 551462 1006272 551468 1006324
rect 551520 1006312 551526 1006324
rect 556798 1006312 556804 1006324
rect 551520 1006284 556804 1006312
rect 551520 1006272 551526 1006284
rect 556798 1006272 556804 1006284
rect 556856 1006272 556862 1006324
rect 555418 1006136 555424 1006188
rect 555476 1006176 555482 1006188
rect 558822 1006176 558828 1006188
rect 555476 1006148 558828 1006176
rect 555476 1006136 555482 1006148
rect 558822 1006136 558828 1006148
rect 558880 1006136 558886 1006188
rect 562318 1006136 562324 1006188
rect 562376 1006176 562382 1006188
rect 567838 1006176 567844 1006188
rect 562376 1006148 567844 1006176
rect 562376 1006136 562382 1006148
rect 567838 1006136 567844 1006148
rect 567896 1006136 567902 1006188
rect 522298 1006040 522304 1006052
rect 518866 1006012 522304 1006040
rect 522298 1006000 522304 1006012
rect 522356 1006000 522362 1006052
rect 549162 1006000 549168 1006052
rect 549220 1006040 549226 1006052
rect 550266 1006040 550272 1006052
rect 549220 1006012 550272 1006040
rect 549220 1006000 549226 1006012
rect 550266 1006000 550272 1006012
rect 550324 1006000 550330 1006052
rect 554774 1006000 554780 1006052
rect 554832 1006040 554838 1006052
rect 573542 1006040 573548 1006052
rect 554832 1006012 573548 1006040
rect 554832 1006000 554838 1006012
rect 573542 1006000 573548 1006012
rect 573600 1006000 573606 1006052
rect 303080 1005876 304304 1005904
rect 428366 1005796 428372 1005848
rect 428424 1005836 428430 1005848
rect 454678 1005836 454684 1005848
rect 428424 1005808 454684 1005836
rect 428424 1005796 428430 1005808
rect 454678 1005796 454684 1005808
rect 454736 1005796 454742 1005848
rect 423490 1005660 423496 1005712
rect 423548 1005700 423554 1005712
rect 432414 1005700 432420 1005712
rect 423548 1005672 432420 1005700
rect 423548 1005660 423554 1005672
rect 432414 1005660 432420 1005672
rect 432472 1005660 432478 1005712
rect 445018 1005700 445024 1005712
rect 432616 1005672 445024 1005700
rect 421834 1005524 421840 1005576
rect 421892 1005564 421898 1005576
rect 425698 1005564 425704 1005576
rect 421892 1005536 425704 1005564
rect 421892 1005524 421898 1005536
rect 425698 1005524 425704 1005536
rect 425756 1005524 425762 1005576
rect 432616 1005564 432644 1005672
rect 445018 1005660 445024 1005672
rect 445076 1005660 445082 1005712
rect 427004 1005536 432644 1005564
rect 360562 1005388 360568 1005440
rect 360620 1005428 360626 1005440
rect 378778 1005428 378784 1005440
rect 360620 1005400 378784 1005428
rect 360620 1005388 360626 1005400
rect 378778 1005388 378784 1005400
rect 378836 1005388 378842 1005440
rect 423490 1005388 423496 1005440
rect 423548 1005428 423554 1005440
rect 427004 1005428 427032 1005536
rect 437474 1005524 437480 1005576
rect 437532 1005564 437538 1005576
rect 467098 1005564 467104 1005576
rect 437532 1005536 467104 1005564
rect 437532 1005524 437538 1005536
rect 467098 1005524 467104 1005536
rect 467156 1005524 467162 1005576
rect 423548 1005400 427032 1005428
rect 423548 1005388 423554 1005400
rect 432414 1005388 432420 1005440
rect 432472 1005428 432478 1005440
rect 457438 1005428 457444 1005440
rect 432472 1005400 457444 1005428
rect 432472 1005388 432478 1005400
rect 457438 1005388 457444 1005400
rect 457496 1005388 457502 1005440
rect 499482 1005388 499488 1005440
rect 499540 1005428 499546 1005440
rect 500494 1005428 500500 1005440
rect 499540 1005400 500500 1005428
rect 499540 1005388 499546 1005400
rect 500494 1005388 500500 1005400
rect 500552 1005388 500558 1005440
rect 564434 1005388 564440 1005440
rect 564492 1005428 564498 1005440
rect 570598 1005428 570604 1005440
rect 564492 1005400 570604 1005428
rect 564492 1005388 564498 1005400
rect 570598 1005388 570604 1005400
rect 570656 1005388 570662 1005440
rect 427170 1005320 427176 1005372
rect 427228 1005360 427234 1005372
rect 427228 1005332 427814 1005360
rect 427228 1005320 427234 1005332
rect 102778 1005252 102784 1005304
rect 102836 1005292 102842 1005304
rect 108850 1005292 108856 1005304
rect 102836 1005264 108856 1005292
rect 102836 1005252 102842 1005264
rect 108850 1005252 108856 1005264
rect 108908 1005252 108914 1005304
rect 204898 1005252 204904 1005304
rect 204956 1005292 204962 1005304
rect 212074 1005292 212080 1005304
rect 204956 1005264 212080 1005292
rect 204956 1005252 204962 1005264
rect 212074 1005252 212080 1005264
rect 212132 1005252 212138 1005304
rect 355686 1005252 355692 1005304
rect 355744 1005292 355750 1005304
rect 376018 1005292 376024 1005304
rect 355744 1005264 376024 1005292
rect 355744 1005252 355750 1005264
rect 376018 1005252 376024 1005264
rect 376076 1005252 376082 1005304
rect 427786 1005292 427814 1005332
rect 463694 1005292 463700 1005304
rect 427786 1005264 463700 1005292
rect 463694 1005252 463700 1005264
rect 463752 1005252 463758 1005304
rect 498838 1005252 498844 1005304
rect 498896 1005292 498902 1005304
rect 516778 1005292 516784 1005304
rect 498896 1005264 516784 1005292
rect 498896 1005252 498902 1005264
rect 516778 1005252 516784 1005264
rect 516836 1005252 516842 1005304
rect 551462 1005252 551468 1005304
rect 551520 1005292 551526 1005304
rect 569218 1005292 569224 1005304
rect 551520 1005264 569224 1005292
rect 551520 1005252 551526 1005264
rect 569218 1005252 569224 1005264
rect 569276 1005252 569282 1005304
rect 304258 1005184 304264 1005236
rect 304316 1005224 304322 1005236
rect 307294 1005224 307300 1005236
rect 304316 1005196 307300 1005224
rect 304316 1005184 304322 1005196
rect 307294 1005184 307300 1005196
rect 307352 1005184 307358 1005236
rect 151078 1005048 151084 1005100
rect 151136 1005088 151142 1005100
rect 153746 1005088 153752 1005100
rect 151136 1005060 153752 1005088
rect 151136 1005048 151142 1005060
rect 153746 1005048 153752 1005060
rect 153804 1005048 153810 1005100
rect 365070 1005048 365076 1005100
rect 365128 1005088 365134 1005100
rect 370498 1005088 370504 1005100
rect 365128 1005060 370504 1005088
rect 365128 1005048 365134 1005060
rect 370498 1005048 370504 1005060
rect 370556 1005048 370562 1005100
rect 425514 1005048 425520 1005100
rect 425572 1005088 425578 1005100
rect 431218 1005088 431224 1005100
rect 425572 1005060 431224 1005088
rect 425572 1005048 425578 1005060
rect 431218 1005048 431224 1005060
rect 431276 1005048 431282 1005100
rect 439498 1005088 439504 1005100
rect 437446 1005060 439504 1005088
rect 149698 1004912 149704 1004964
rect 149756 1004952 149762 1004964
rect 152918 1004952 152924 1004964
rect 149756 1004924 152924 1004952
rect 149756 1004912 149762 1004924
rect 152918 1004912 152924 1004924
rect 152976 1004912 152982 1004964
rect 209222 1004912 209228 1004964
rect 209280 1004952 209286 1004964
rect 211798 1004952 211804 1004964
rect 209280 1004924 211804 1004952
rect 209280 1004912 209286 1004924
rect 211798 1004912 211804 1004924
rect 211856 1004912 211862 1004964
rect 263042 1004912 263048 1004964
rect 263100 1004952 263106 1004964
rect 268378 1004952 268384 1004964
rect 263100 1004924 268384 1004952
rect 263100 1004912 263106 1004924
rect 268378 1004912 268384 1004924
rect 268436 1004912 268442 1004964
rect 303614 1004912 303620 1004964
rect 303672 1004952 303678 1004964
rect 306926 1004952 306932 1004964
rect 303672 1004924 306932 1004952
rect 303672 1004912 303678 1004924
rect 306926 1004912 306932 1004924
rect 306984 1004912 306990 1004964
rect 354582 1004912 354588 1004964
rect 354640 1004952 354646 1004964
rect 356514 1004952 356520 1004964
rect 354640 1004924 356520 1004952
rect 354640 1004912 354646 1004924
rect 356514 1004912 356520 1004924
rect 356572 1004912 356578 1004964
rect 361390 1004912 361396 1004964
rect 361448 1004952 361454 1004964
rect 364978 1004952 364984 1004964
rect 361448 1004924 364984 1004952
rect 361448 1004912 361454 1004924
rect 364978 1004912 364984 1004924
rect 365036 1004912 365042 1004964
rect 427998 1004912 428004 1004964
rect 428056 1004952 428062 1004964
rect 437446 1004952 437474 1005060
rect 439498 1005048 439504 1005060
rect 439556 1005048 439562 1005100
rect 428056 1004924 437474 1004952
rect 428056 1004912 428062 1004924
rect 498102 1004912 498108 1004964
rect 498160 1004952 498166 1004964
rect 500494 1004952 500500 1004964
rect 498160 1004924 500500 1004952
rect 498160 1004912 498166 1004924
rect 500494 1004912 500500 1004924
rect 500552 1004912 500558 1004964
rect 557166 1004912 557172 1004964
rect 557224 1004952 557230 1004964
rect 558914 1004952 558920 1004964
rect 557224 1004924 558920 1004952
rect 557224 1004912 557230 1004924
rect 558914 1004912 558920 1004924
rect 558972 1004912 558978 1004964
rect 151262 1004776 151268 1004828
rect 151320 1004816 151326 1004828
rect 154114 1004816 154120 1004828
rect 151320 1004788 154120 1004816
rect 151320 1004776 151326 1004788
rect 154114 1004776 154120 1004788
rect 154172 1004776 154178 1004828
rect 160646 1004776 160652 1004828
rect 160704 1004816 160710 1004828
rect 163130 1004816 163136 1004828
rect 160704 1004788 163136 1004816
rect 160704 1004776 160710 1004788
rect 163130 1004776 163136 1004788
rect 163188 1004776 163194 1004828
rect 211246 1004776 211252 1004828
rect 211304 1004816 211310 1004828
rect 215938 1004816 215944 1004828
rect 211304 1004788 215944 1004816
rect 211304 1004776 211310 1004788
rect 215938 1004776 215944 1004788
rect 215996 1004776 216002 1004828
rect 258166 1004776 258172 1004828
rect 258224 1004816 258230 1004828
rect 259454 1004816 259460 1004828
rect 258224 1004788 259460 1004816
rect 258224 1004776 258230 1004788
rect 259454 1004776 259460 1004788
rect 259512 1004776 259518 1004828
rect 305822 1004776 305828 1004828
rect 305880 1004816 305886 1004828
rect 308950 1004816 308956 1004828
rect 305880 1004788 308956 1004816
rect 305880 1004776 305886 1004788
rect 308950 1004776 308956 1004788
rect 309008 1004776 309014 1004828
rect 313826 1004776 313832 1004828
rect 313884 1004816 313890 1004828
rect 316034 1004816 316040 1004828
rect 313884 1004788 316040 1004816
rect 313884 1004776 313890 1004788
rect 316034 1004776 316040 1004788
rect 316092 1004776 316098 1004828
rect 353202 1004776 353208 1004828
rect 353260 1004816 353266 1004828
rect 355686 1004816 355692 1004828
rect 353260 1004788 355692 1004816
rect 353260 1004776 353266 1004788
rect 355686 1004776 355692 1004788
rect 355744 1004776 355750 1004828
rect 362586 1004776 362592 1004828
rect 362644 1004816 362650 1004828
rect 365162 1004816 365168 1004828
rect 362644 1004788 365168 1004816
rect 362644 1004776 362650 1004788
rect 365162 1004776 365168 1004788
rect 365220 1004776 365226 1004828
rect 420454 1004776 420460 1004828
rect 420512 1004816 420518 1004828
rect 422662 1004816 422668 1004828
rect 420512 1004788 422668 1004816
rect 420512 1004776 420518 1004788
rect 422662 1004776 422668 1004788
rect 422720 1004776 422726 1004828
rect 497918 1004776 497924 1004828
rect 497976 1004816 497982 1004828
rect 499666 1004816 499672 1004828
rect 497976 1004788 499672 1004816
rect 497976 1004776 497982 1004788
rect 499666 1004776 499672 1004788
rect 499724 1004776 499730 1004828
rect 555970 1004776 555976 1004828
rect 556028 1004816 556034 1004828
rect 558178 1004816 558184 1004828
rect 556028 1004788 558184 1004816
rect 556028 1004776 556034 1004788
rect 558178 1004776 558184 1004788
rect 558236 1004776 558242 1004828
rect 106182 1004640 106188 1004692
rect 106240 1004680 106246 1004692
rect 108482 1004680 108488 1004692
rect 106240 1004652 108488 1004680
rect 106240 1004640 106246 1004652
rect 108482 1004640 108488 1004652
rect 108540 1004640 108546 1004692
rect 149882 1004640 149888 1004692
rect 149940 1004680 149946 1004692
rect 151722 1004680 151728 1004692
rect 149940 1004652 151728 1004680
rect 149940 1004640 149946 1004652
rect 151722 1004640 151728 1004652
rect 151780 1004640 151786 1004692
rect 161106 1004640 161112 1004692
rect 161164 1004680 161170 1004692
rect 162946 1004680 162952 1004692
rect 161164 1004652 162952 1004680
rect 161164 1004640 161170 1004652
rect 162946 1004640 162952 1004652
rect 163004 1004640 163010 1004692
rect 209222 1004640 209228 1004692
rect 209280 1004680 209286 1004692
rect 211154 1004680 211160 1004692
rect 209280 1004652 211160 1004680
rect 209280 1004640 209286 1004652
rect 211154 1004640 211160 1004652
rect 211212 1004640 211218 1004692
rect 305638 1004640 305644 1004692
rect 305696 1004680 305702 1004692
rect 308122 1004680 308128 1004692
rect 305696 1004652 308128 1004680
rect 305696 1004640 305702 1004652
rect 308122 1004640 308128 1004652
rect 308180 1004640 308186 1004692
rect 315482 1004640 315488 1004692
rect 315540 1004680 315546 1004692
rect 318058 1004680 318064 1004692
rect 315540 1004652 318064 1004680
rect 315540 1004640 315546 1004652
rect 318058 1004640 318064 1004652
rect 318116 1004640 318122 1004692
rect 364242 1004640 364248 1004692
rect 364300 1004680 364306 1004692
rect 366358 1004680 366364 1004692
rect 364300 1004652 366364 1004680
rect 364300 1004640 364306 1004652
rect 366358 1004640 366364 1004652
rect 366416 1004640 366422 1004692
rect 432874 1004640 432880 1004692
rect 432932 1004680 432938 1004692
rect 438118 1004680 438124 1004692
rect 432932 1004652 438124 1004680
rect 432932 1004640 432938 1004652
rect 438118 1004640 438124 1004652
rect 438176 1004640 438182 1004692
rect 557626 1004640 557632 1004692
rect 557684 1004680 557690 1004692
rect 559558 1004680 559564 1004692
rect 557684 1004652 559564 1004680
rect 557684 1004640 557690 1004652
rect 559558 1004640 559564 1004652
rect 559616 1004640 559622 1004692
rect 560846 1004640 560852 1004692
rect 560904 1004680 560910 1004692
rect 566458 1004680 566464 1004692
rect 560904 1004652 566464 1004680
rect 560904 1004640 560910 1004652
rect 566458 1004640 566464 1004652
rect 566516 1004640 566522 1004692
rect 570322 1004096 570328 1004148
rect 570380 1004136 570386 1004148
rect 573358 1004136 573364 1004148
rect 570380 1004108 573364 1004136
rect 570380 1004096 570386 1004108
rect 573358 1004096 573364 1004108
rect 573416 1004096 573422 1004148
rect 513374 1004028 513380 1004080
rect 513432 1004068 513438 1004080
rect 518894 1004068 518900 1004080
rect 513432 1004040 518900 1004068
rect 513432 1004028 513438 1004040
rect 518894 1004028 518900 1004040
rect 518952 1004028 518958 1004080
rect 247126 1003892 247132 1003944
rect 247184 1003932 247190 1003944
rect 255314 1003932 255320 1003944
rect 247184 1003904 255320 1003932
rect 247184 1003892 247190 1003904
rect 255314 1003892 255320 1003904
rect 255372 1003892 255378 1003944
rect 424318 1003892 424324 1003944
rect 424376 1003932 424382 1003944
rect 443638 1003932 443644 1003944
rect 424376 1003904 443644 1003932
rect 424376 1003892 424382 1003904
rect 443638 1003892 443644 1003904
rect 443696 1003892 443702 1003944
rect 558914 1003892 558920 1003944
rect 558972 1003932 558978 1003944
rect 570782 1003932 570788 1003944
rect 558972 1003904 570788 1003932
rect 558972 1003892 558978 1003904
rect 570782 1003892 570788 1003904
rect 570840 1003892 570846 1003944
rect 300302 1003280 300308 1003332
rect 300360 1003320 300366 1003332
rect 305270 1003320 305276 1003332
rect 300360 1003292 305276 1003320
rect 300360 1003280 300366 1003292
rect 305270 1003280 305276 1003292
rect 305328 1003280 305334 1003332
rect 553394 1003280 553400 1003332
rect 553452 1003320 553458 1003332
rect 554590 1003320 554596 1003332
rect 553452 1003292 554596 1003320
rect 553452 1003280 553458 1003292
rect 554590 1003280 554596 1003292
rect 554648 1003280 554654 1003332
rect 299290 1003144 299296 1003196
rect 299348 1003184 299354 1003196
rect 308950 1003184 308956 1003196
rect 299348 1003156 308956 1003184
rect 299348 1003144 299354 1003156
rect 308950 1003144 308956 1003156
rect 309008 1003144 309014 1003196
rect 253106 1002668 253112 1002720
rect 253164 1002708 253170 1002720
rect 256142 1002708 256148 1002720
rect 253164 1002680 256148 1002708
rect 253164 1002668 253170 1002680
rect 256142 1002668 256148 1002680
rect 256200 1002668 256206 1002720
rect 424686 1002668 424692 1002720
rect 424744 1002708 424750 1002720
rect 448974 1002708 448980 1002720
rect 424744 1002680 448980 1002708
rect 424744 1002668 424750 1002680
rect 448974 1002668 448980 1002680
rect 449032 1002668 449038 1002720
rect 97258 1002600 97264 1002652
rect 97316 1002640 97322 1002652
rect 100294 1002640 100300 1002652
rect 97316 1002612 100300 1002640
rect 97316 1002600 97322 1002612
rect 100294 1002600 100300 1002612
rect 100352 1002600 100358 1002652
rect 553118 1002600 553124 1002652
rect 553176 1002640 553182 1002652
rect 553762 1002640 553768 1002652
rect 553176 1002612 553768 1002640
rect 553176 1002600 553182 1002612
rect 553762 1002600 553768 1002612
rect 553820 1002600 553826 1002652
rect 558822 1002600 558828 1002652
rect 558880 1002640 558886 1002652
rect 562502 1002640 562508 1002652
rect 558880 1002612 562508 1002640
rect 558880 1002600 558886 1002612
rect 562502 1002600 562508 1002612
rect 562560 1002600 562566 1002652
rect 246574 1002532 246580 1002584
rect 246632 1002572 246638 1002584
rect 254118 1002572 254124 1002584
rect 246632 1002544 254124 1002572
rect 246632 1002532 246638 1002544
rect 254118 1002532 254124 1002544
rect 254176 1002532 254182 1002584
rect 429746 1002532 429752 1002584
rect 429804 1002572 429810 1002584
rect 464982 1002572 464988 1002584
rect 429804 1002544 464988 1002572
rect 429804 1002532 429810 1002544
rect 464982 1002532 464988 1002544
rect 465040 1002532 465046 1002584
rect 98638 1002464 98644 1002516
rect 98696 1002504 98702 1002516
rect 101950 1002504 101956 1002516
rect 98696 1002476 101956 1002504
rect 98696 1002464 98702 1002476
rect 101950 1002464 101956 1002476
rect 102008 1002464 102014 1002516
rect 202874 1002464 202880 1002516
rect 202932 1002504 202938 1002516
rect 206370 1002504 206376 1002516
rect 202932 1002476 206376 1002504
rect 202932 1002464 202938 1002476
rect 206370 1002464 206376 1002476
rect 206428 1002464 206434 1002516
rect 509878 1002464 509884 1002516
rect 509936 1002504 509942 1002516
rect 515398 1002504 515404 1002516
rect 509936 1002476 515404 1002504
rect 509936 1002464 509942 1002476
rect 515398 1002464 515404 1002476
rect 515456 1002464 515462 1002516
rect 560846 1002464 560852 1002516
rect 560904 1002504 560910 1002516
rect 565078 1002504 565084 1002516
rect 560904 1002476 565084 1002504
rect 560904 1002464 560910 1002476
rect 565078 1002464 565084 1002476
rect 565136 1002464 565142 1002516
rect 97442 1002328 97448 1002380
rect 97500 1002368 97506 1002380
rect 100294 1002368 100300 1002380
rect 97500 1002340 100300 1002368
rect 97500 1002328 97506 1002340
rect 100294 1002328 100300 1002340
rect 100352 1002328 100358 1002380
rect 100478 1002328 100484 1002380
rect 100536 1002368 100542 1002380
rect 103146 1002368 103152 1002380
rect 100536 1002340 103152 1002368
rect 100536 1002328 100542 1002340
rect 103146 1002328 103152 1002340
rect 103204 1002328 103210 1002380
rect 107654 1002328 107660 1002380
rect 107712 1002368 107718 1002380
rect 109494 1002368 109500 1002380
rect 107712 1002340 109500 1002368
rect 107712 1002328 107718 1002340
rect 109494 1002328 109500 1002340
rect 109552 1002328 109558 1002380
rect 148502 1002328 148508 1002380
rect 148560 1002368 148566 1002380
rect 150894 1002368 150900 1002380
rect 148560 1002340 150900 1002368
rect 148560 1002328 148566 1002340
rect 150894 1002328 150900 1002340
rect 150952 1002328 150958 1002380
rect 251818 1002328 251824 1002380
rect 251876 1002368 251882 1002380
rect 254486 1002368 254492 1002380
rect 251876 1002340 254492 1002368
rect 251876 1002328 251882 1002340
rect 254486 1002328 254492 1002340
rect 254544 1002328 254550 1002380
rect 261018 1002328 261024 1002380
rect 261076 1002368 261082 1002380
rect 264238 1002368 264244 1002380
rect 261076 1002340 264244 1002368
rect 261076 1002328 261082 1002340
rect 264238 1002328 264244 1002340
rect 264296 1002328 264302 1002380
rect 357710 1002328 357716 1002380
rect 357768 1002368 357774 1002380
rect 360838 1002368 360844 1002380
rect 357768 1002340 360844 1002368
rect 357768 1002328 357774 1002340
rect 360838 1002328 360844 1002340
rect 360896 1002328 360902 1002380
rect 501690 1002328 501696 1002380
rect 501748 1002368 501754 1002380
rect 503714 1002368 503720 1002380
rect 501748 1002340 503720 1002368
rect 501748 1002328 501754 1002340
rect 503714 1002328 503720 1002340
rect 503772 1002328 503778 1002380
rect 560478 1002328 560484 1002380
rect 560536 1002368 560542 1002380
rect 563054 1002368 563060 1002380
rect 560536 1002340 563060 1002368
rect 560536 1002328 560542 1002340
rect 563054 1002328 563060 1002340
rect 563112 1002328 563118 1002380
rect 98822 1002192 98828 1002244
rect 98880 1002232 98886 1002244
rect 101122 1002232 101128 1002244
rect 98880 1002204 101128 1002232
rect 98880 1002192 98886 1002204
rect 101122 1002192 101128 1002204
rect 101180 1002192 101186 1002244
rect 105630 1002192 105636 1002244
rect 105688 1002232 105694 1002244
rect 107838 1002232 107844 1002244
rect 105688 1002204 107844 1002232
rect 105688 1002192 105694 1002204
rect 107838 1002192 107844 1002204
rect 107896 1002192 107902 1002244
rect 108022 1002192 108028 1002244
rect 108080 1002232 108086 1002244
rect 110414 1002232 110420 1002244
rect 108080 1002204 110420 1002232
rect 108080 1002192 108086 1002204
rect 110414 1002192 110420 1002204
rect 110472 1002192 110478 1002244
rect 155770 1002192 155776 1002244
rect 155828 1002232 155834 1002244
rect 157334 1002232 157340 1002244
rect 155828 1002204 157340 1002232
rect 155828 1002192 155834 1002204
rect 157334 1002192 157340 1002204
rect 157392 1002192 157398 1002244
rect 205082 1002192 205088 1002244
rect 205140 1002232 205146 1002244
rect 207198 1002232 207204 1002244
rect 205140 1002204 207204 1002232
rect 205140 1002192 205146 1002204
rect 207198 1002192 207204 1002204
rect 207256 1002192 207262 1002244
rect 254578 1002192 254584 1002244
rect 254636 1002232 254642 1002244
rect 256510 1002232 256516 1002244
rect 254636 1002204 256516 1002232
rect 254636 1002192 254642 1002204
rect 256510 1002192 256516 1002204
rect 256568 1002192 256574 1002244
rect 260190 1002192 260196 1002244
rect 260248 1002232 260254 1002244
rect 262858 1002232 262864 1002244
rect 260248 1002204 262864 1002232
rect 260248 1002192 260254 1002204
rect 262858 1002192 262864 1002204
rect 262916 1002192 262922 1002244
rect 303062 1002192 303068 1002244
rect 303120 1002232 303126 1002244
rect 306098 1002232 306104 1002244
rect 303120 1002204 306104 1002232
rect 303120 1002192 303126 1002204
rect 306098 1002192 306104 1002204
rect 306156 1002192 306162 1002244
rect 308398 1002192 308404 1002244
rect 308456 1002232 308462 1002244
rect 310606 1002232 310612 1002244
rect 308456 1002204 310612 1002232
rect 308456 1002192 308462 1002204
rect 310606 1002192 310612 1002204
rect 310664 1002192 310670 1002244
rect 500586 1002192 500592 1002244
rect 500644 1002232 500650 1002244
rect 503346 1002232 503352 1002244
rect 500644 1002204 503352 1002232
rect 500644 1002192 500650 1002204
rect 503346 1002192 503352 1002204
rect 503404 1002192 503410 1002244
rect 504174 1002192 504180 1002244
rect 504232 1002232 504238 1002244
rect 510062 1002232 510068 1002244
rect 504232 1002204 510068 1002232
rect 504232 1002192 504238 1002204
rect 510062 1002192 510068 1002204
rect 510120 1002192 510126 1002244
rect 557994 1002192 558000 1002244
rect 558052 1002232 558058 1002244
rect 560938 1002232 560944 1002244
rect 558052 1002204 560944 1002232
rect 558052 1002192 558058 1002204
rect 560938 1002192 560944 1002204
rect 560996 1002192 561002 1002244
rect 553210 1002124 553216 1002176
rect 553268 1002164 553274 1002176
rect 553946 1002164 553952 1002176
rect 553268 1002136 553952 1002164
rect 553268 1002124 553274 1002136
rect 553946 1002124 553952 1002136
rect 554004 1002124 554010 1002176
rect 96062 1002056 96068 1002108
rect 96120 1002096 96126 1002108
rect 99098 1002096 99104 1002108
rect 96120 1002068 99104 1002096
rect 96120 1002056 96126 1002068
rect 99098 1002056 99104 1002068
rect 99156 1002056 99162 1002108
rect 100018 1002056 100024 1002108
rect 100076 1002096 100082 1002108
rect 102318 1002096 102324 1002108
rect 100076 1002068 102324 1002096
rect 100076 1002056 100082 1002068
rect 102318 1002056 102324 1002068
rect 102376 1002056 102382 1002108
rect 103974 1002056 103980 1002108
rect 104032 1002096 104038 1002108
rect 106458 1002096 106464 1002108
rect 104032 1002068 106464 1002096
rect 104032 1002056 104038 1002068
rect 106458 1002056 106464 1002068
rect 106516 1002056 106522 1002108
rect 106826 1002056 106832 1002108
rect 106884 1002096 106890 1002108
rect 109034 1002096 109040 1002108
rect 106884 1002068 109040 1002096
rect 106884 1002056 106890 1002068
rect 109034 1002056 109040 1002068
rect 109092 1002056 109098 1002108
rect 109678 1002056 109684 1002108
rect 109736 1002096 109742 1002108
rect 111794 1002096 111800 1002108
rect 109736 1002068 111800 1002096
rect 109736 1002056 109742 1002068
rect 111794 1002056 111800 1002068
rect 111852 1002056 111858 1002108
rect 148318 1002056 148324 1002108
rect 148376 1002096 148382 1002108
rect 150894 1002096 150900 1002108
rect 148376 1002068 150900 1002096
rect 148376 1002056 148382 1002068
rect 150894 1002056 150900 1002068
rect 150952 1002056 150958 1002108
rect 152458 1002056 152464 1002108
rect 152516 1002096 152522 1002108
rect 154574 1002096 154580 1002108
rect 152516 1002068 154580 1002096
rect 152516 1002056 152522 1002068
rect 154574 1002056 154580 1002068
rect 154632 1002056 154638 1002108
rect 157794 1002056 157800 1002108
rect 157852 1002096 157858 1002108
rect 160094 1002096 160100 1002108
rect 157852 1002068 160100 1002096
rect 157852 1002056 157858 1002068
rect 160094 1002056 160100 1002068
rect 160152 1002056 160158 1002108
rect 206738 1002056 206744 1002108
rect 206796 1002096 206802 1002108
rect 208578 1002096 208584 1002108
rect 206796 1002068 208584 1002096
rect 206796 1002056 206802 1002068
rect 208578 1002056 208584 1002068
rect 208636 1002056 208642 1002108
rect 210878 1002056 210884 1002108
rect 210936 1002096 210942 1002108
rect 213178 1002096 213184 1002108
rect 210936 1002068 213184 1002096
rect 210936 1002056 210942 1002068
rect 213178 1002056 213184 1002068
rect 213236 1002056 213242 1002108
rect 253382 1002056 253388 1002108
rect 253440 1002096 253446 1002108
rect 255314 1002096 255320 1002108
rect 253440 1002068 255320 1002096
rect 253440 1002056 253446 1002068
rect 255314 1002056 255320 1002068
rect 255372 1002056 255378 1002108
rect 259822 1002056 259828 1002108
rect 259880 1002096 259886 1002108
rect 262214 1002096 262220 1002108
rect 259880 1002068 262220 1002096
rect 259880 1002056 259886 1002068
rect 262214 1002056 262220 1002068
rect 262272 1002056 262278 1002108
rect 263870 1002056 263876 1002108
rect 263928 1002096 263934 1002108
rect 266998 1002096 267004 1002108
rect 263928 1002068 267004 1002096
rect 263928 1002056 263934 1002068
rect 266998 1002056 267004 1002068
rect 267056 1002056 267062 1002108
rect 300118 1002056 300124 1002108
rect 300176 1002096 300182 1002108
rect 304074 1002096 304080 1002108
rect 300176 1002068 304080 1002096
rect 300176 1002056 300182 1002068
rect 304074 1002056 304080 1002068
rect 304132 1002056 304138 1002108
rect 355778 1002056 355784 1002108
rect 355836 1002096 355842 1002108
rect 357710 1002096 357716 1002108
rect 355836 1002068 357716 1002096
rect 355836 1002056 355842 1002068
rect 357710 1002056 357716 1002068
rect 357768 1002056 357774 1002108
rect 423582 1002056 423588 1002108
rect 423640 1002096 423646 1002108
rect 426342 1002096 426348 1002108
rect 423640 1002068 426348 1002096
rect 423640 1002056 423646 1002068
rect 426342 1002056 426348 1002068
rect 426400 1002056 426406 1002108
rect 502518 1002056 502524 1002108
rect 502576 1002096 502582 1002108
rect 505738 1002096 505744 1002108
rect 502576 1002068 505744 1002096
rect 502576 1002056 502582 1002068
rect 505738 1002056 505744 1002068
rect 505796 1002056 505802 1002108
rect 560018 1002056 560024 1002108
rect 560076 1002096 560082 1002108
rect 562318 1002096 562324 1002108
rect 560076 1002068 562324 1002096
rect 560076 1002056 560082 1002068
rect 562318 1002056 562324 1002068
rect 562376 1002056 562382 1002108
rect 95878 1001920 95884 1001972
rect 95936 1001960 95942 1001972
rect 98270 1001960 98276 1001972
rect 95936 1001932 98276 1001960
rect 95936 1001920 95942 1001932
rect 98270 1001920 98276 1001932
rect 98328 1001920 98334 1001972
rect 99006 1001920 99012 1001972
rect 99064 1001960 99070 1001972
rect 101122 1001960 101128 1001972
rect 99064 1001932 101128 1001960
rect 99064 1001920 99070 1001932
rect 101122 1001920 101128 1001932
rect 101180 1001920 101186 1001972
rect 105998 1001920 106004 1001972
rect 106056 1001960 106062 1001972
rect 107746 1001960 107752 1001972
rect 106056 1001932 107752 1001960
rect 106056 1001920 106062 1001932
rect 107746 1001920 107752 1001932
rect 107804 1001920 107810 1001972
rect 146938 1001920 146944 1001972
rect 146996 1001960 147002 1001972
rect 149238 1001960 149244 1001972
rect 146996 1001932 149244 1001960
rect 146996 1001920 147002 1001932
rect 149238 1001920 149244 1001932
rect 149296 1001920 149302 1001972
rect 156598 1001920 156604 1001972
rect 156656 1001960 156662 1001972
rect 158714 1001960 158720 1001972
rect 156656 1001932 158720 1001960
rect 156656 1001920 156662 1001932
rect 158714 1001920 158720 1001932
rect 158772 1001920 158778 1001972
rect 202874 1001960 202880 1001972
rect 195164 1001932 202880 1001960
rect 195164 1001768 195192 1001932
rect 202874 1001920 202880 1001932
rect 202932 1001920 202938 1001972
rect 204162 1001920 204168 1001972
rect 204220 1001960 204226 1001972
rect 205542 1001960 205548 1001972
rect 204220 1001932 205548 1001960
rect 204220 1001920 204226 1001932
rect 205542 1001920 205548 1001932
rect 205600 1001920 205606 1001972
rect 206278 1001920 206284 1001972
rect 206336 1001960 206342 1001972
rect 207566 1001960 207572 1001972
rect 206336 1001932 207572 1001960
rect 206336 1001920 206342 1001932
rect 207566 1001920 207572 1001932
rect 207624 1001920 207630 1001972
rect 212534 1001920 212540 1001972
rect 212592 1001960 212598 1001972
rect 214558 1001960 214564 1001972
rect 212592 1001932 214564 1001960
rect 212592 1001920 212598 1001932
rect 214558 1001920 214564 1001932
rect 214616 1001920 214622 1001972
rect 254762 1001920 254768 1001972
rect 254820 1001960 254826 1001972
rect 256970 1001960 256976 1001972
rect 254820 1001932 256976 1001960
rect 254820 1001920 254826 1001932
rect 256970 1001920 256976 1001932
rect 257028 1001920 257034 1001972
rect 260190 1001920 260196 1001972
rect 260248 1001960 260254 1001972
rect 260926 1001960 260932 1001972
rect 260248 1001932 260932 1001960
rect 260248 1001920 260254 1001932
rect 260926 1001920 260932 1001932
rect 260984 1001920 260990 1001972
rect 263502 1001920 263508 1001972
rect 263560 1001960 263566 1001972
rect 265618 1001960 265624 1001972
rect 263560 1001932 265624 1001960
rect 263560 1001920 263566 1001932
rect 265618 1001920 265624 1001932
rect 265676 1001920 265682 1001972
rect 302878 1001920 302884 1001972
rect 302936 1001960 302942 1001972
rect 306098 1001960 306104 1001972
rect 302936 1001932 306104 1001960
rect 302936 1001920 302942 1001932
rect 306098 1001920 306104 1001932
rect 306156 1001920 306162 1001972
rect 310146 1001920 310152 1001972
rect 310204 1001960 310210 1001972
rect 311894 1001960 311900 1001972
rect 310204 1001932 311900 1001960
rect 310204 1001920 310210 1001932
rect 311894 1001920 311900 1001932
rect 311952 1001920 311958 1001972
rect 351822 1001920 351828 1001972
rect 351880 1001960 351886 1001972
rect 354030 1001960 354036 1001972
rect 351880 1001932 354036 1001960
rect 351880 1001920 351886 1001932
rect 354030 1001920 354036 1001932
rect 354088 1001920 354094 1001972
rect 365898 1001920 365904 1001972
rect 365956 1001960 365962 1001972
rect 369118 1001960 369124 1001972
rect 365956 1001932 369124 1001960
rect 365956 1001920 365962 1001932
rect 369118 1001920 369124 1001932
rect 369176 1001920 369182 1001972
rect 419442 1001920 419448 1001972
rect 419500 1001960 419506 1001972
rect 421466 1001960 421472 1001972
rect 419500 1001932 421472 1001960
rect 419500 1001920 419506 1001932
rect 421466 1001920 421472 1001932
rect 421524 1001920 421530 1001972
rect 425514 1001920 425520 1001972
rect 425572 1001960 425578 1001972
rect 425572 1001932 427814 1001960
rect 425572 1001920 425578 1001932
rect 427786 1001892 427814 1001932
rect 500770 1001920 500776 1001972
rect 500828 1001960 500834 1001972
rect 501322 1001960 501328 1001972
rect 500828 1001932 501328 1001960
rect 500828 1001920 500834 1001932
rect 501322 1001920 501328 1001932
rect 501380 1001920 501386 1001972
rect 504542 1001920 504548 1001972
rect 504600 1001960 504606 1001972
rect 506842 1001960 506848 1001972
rect 504600 1001932 506848 1001960
rect 504600 1001920 504606 1001932
rect 506842 1001920 506848 1001932
rect 506900 1001920 506906 1001972
rect 557994 1001920 558000 1001972
rect 558052 1001960 558058 1001972
rect 560294 1001960 560300 1001972
rect 558052 1001932 560300 1001960
rect 558052 1001920 558058 1001932
rect 560294 1001920 560300 1001932
rect 560352 1001920 560358 1001972
rect 561674 1001920 561680 1001972
rect 561732 1001960 561738 1001972
rect 563698 1001960 563704 1001972
rect 561732 1001932 563704 1001960
rect 561732 1001920 561738 1001932
rect 563698 1001920 563704 1001932
rect 563756 1001920 563762 1001972
rect 428182 1001892 428188 1001904
rect 427786 1001864 428188 1001892
rect 428182 1001852 428188 1001864
rect 428240 1001852 428246 1001904
rect 195146 1001716 195152 1001768
rect 195204 1001716 195210 1001768
rect 439498 1001444 439504 1001496
rect 439556 1001484 439562 1001496
rect 458174 1001484 458180 1001496
rect 439556 1001456 458180 1001484
rect 439556 1001444 439562 1001456
rect 458174 1001444 458180 1001456
rect 458232 1001444 458238 1001496
rect 425698 1001308 425704 1001360
rect 425756 1001348 425762 1001360
rect 446398 1001348 446404 1001360
rect 425756 1001320 446404 1001348
rect 425756 1001308 425762 1001320
rect 446398 1001308 446404 1001320
rect 446456 1001308 446462 1001360
rect 353202 1001172 353208 1001224
rect 353260 1001212 353266 1001224
rect 380894 1001212 380900 1001224
rect 353260 1001184 380900 1001212
rect 353260 1001172 353266 1001184
rect 380894 1001172 380900 1001184
rect 380952 1001172 380958 1001224
rect 423582 1001172 423588 1001224
rect 423640 1001212 423646 1001224
rect 462222 1001212 462228 1001224
rect 423640 1001184 462228 1001212
rect 423640 1001172 423646 1001184
rect 462222 1001172 462228 1001184
rect 462280 1001172 462286 1001224
rect 497918 1001172 497924 1001224
rect 497976 1001212 497982 1001224
rect 521286 1001212 521292 1001224
rect 497976 1001184 521292 1001212
rect 497976 1001172 497982 1001184
rect 521286 1001172 521292 1001184
rect 521344 1001172 521350 1001224
rect 550266 1001172 550272 1001224
rect 550324 1001212 550330 1001224
rect 574094 1001212 574100 1001224
rect 550324 1001184 574100 1001212
rect 550324 1001172 550330 1001184
rect 574094 1001172 574100 1001184
rect 574152 1001172 574158 1001224
rect 298462 1000492 298468 1000544
rect 298520 1000532 298526 1000544
rect 305822 1000532 305828 1000544
rect 298520 1000504 305828 1000532
rect 298520 1000492 298526 1000504
rect 305822 1000492 305828 1000504
rect 305880 1000492 305886 1000544
rect 499482 1000492 499488 1000544
rect 499540 1000532 499546 1000544
rect 500310 1000532 500316 1000544
rect 499540 1000504 500316 1000532
rect 499540 1000492 499546 1000504
rect 500310 1000492 500316 1000504
rect 500368 1000492 500374 1000544
rect 503714 1000492 503720 1000544
rect 503772 1000532 503778 1000544
rect 516870 1000532 516876 1000544
rect 503772 1000504 516876 1000532
rect 503772 1000492 503778 1000504
rect 516870 1000492 516876 1000504
rect 516928 1000492 516934 1000544
rect 617334 1000492 617340 1000544
rect 617392 1000532 617398 1000544
rect 625430 1000532 625436 1000544
rect 617392 1000504 625436 1000532
rect 617392 1000492 617398 1000504
rect 625430 1000492 625436 1000504
rect 625488 1000492 625494 1000544
rect 567838 1000084 567844 1000136
rect 567896 1000124 567902 1000136
rect 571334 1000124 571340 1000136
rect 567896 1000096 571340 1000124
rect 567896 1000084 567902 1000096
rect 571334 1000084 571340 1000096
rect 571392 1000084 571398 1000136
rect 558178 999948 558184 1000000
rect 558236 999988 558242 1000000
rect 565814 999988 565820 1000000
rect 558236 999960 565820 999988
rect 558236 999948 558242 999960
rect 565814 999948 565820 999960
rect 565872 999948 565878 1000000
rect 93302 999744 93308 999796
rect 93360 999784 93366 999796
rect 99006 999784 99012 999796
rect 93360 999756 99012 999784
rect 93360 999744 93366 999756
rect 99006 999744 99012 999756
rect 99064 999744 99070 999796
rect 246942 999744 246948 999796
rect 247000 999784 247006 999796
rect 254762 999784 254768 999796
rect 247000 999756 254768 999784
rect 247000 999744 247006 999756
rect 254762 999744 254768 999756
rect 254820 999744 254826 999796
rect 590930 999268 590936 999320
rect 590988 999308 590994 999320
rect 625062 999308 625068 999320
rect 590988 999280 625068 999308
rect 590988 999268 590994 999280
rect 625062 999268 625068 999280
rect 625120 999268 625126 999320
rect 618162 999132 618168 999184
rect 618220 999172 618226 999184
rect 625614 999172 625620 999184
rect 618220 999144 625620 999172
rect 618220 999132 618226 999144
rect 625614 999132 625620 999144
rect 625672 999132 625678 999184
rect 507394 999064 507400 999116
rect 507452 999104 507458 999116
rect 509234 999104 509240 999116
rect 507452 999076 509240 999104
rect 507452 999064 507458 999076
rect 509234 999064 509240 999076
rect 509292 999064 509298 999116
rect 553394 999064 553400 999116
rect 553452 999104 553458 999116
rect 556338 999104 556344 999116
rect 553452 999076 556344 999104
rect 553452 999064 553458 999076
rect 556338 999064 556344 999076
rect 556396 999064 556402 999116
rect 505370 998928 505376 998980
rect 505428 998968 505434 998980
rect 511442 998968 511448 998980
rect 505428 998940 511448 998968
rect 505428 998928 505434 998940
rect 511442 998928 511448 998940
rect 511500 998928 511506 998980
rect 382642 998900 382648 998912
rect 373966 998872 382648 998900
rect 200206 998792 200212 998844
rect 200264 998832 200270 998844
rect 203886 998832 203892 998844
rect 200264 998804 203892 998832
rect 200264 998792 200270 998804
rect 203886 998792 203892 998804
rect 203944 998792 203950 998844
rect 356054 998792 356060 998844
rect 356112 998832 356118 998844
rect 372154 998832 372160 998844
rect 356112 998804 372160 998832
rect 356112 998792 356118 998804
rect 372154 998792 372160 998804
rect 372212 998792 372218 998844
rect 373258 998792 373264 998844
rect 373316 998832 373322 998844
rect 373966 998832 373994 998872
rect 382642 998860 382648 998872
rect 382700 998860 382706 998912
rect 523862 998900 523868 998912
rect 518866 998872 523868 998900
rect 373316 998804 373994 998832
rect 373316 998792 373322 998804
rect 440878 998792 440884 998844
rect 440936 998832 440942 998844
rect 448514 998832 448520 998844
rect 440936 998804 448520 998832
rect 440936 998792 440942 998804
rect 448514 998792 448520 998804
rect 448572 998792 448578 998844
rect 458358 998832 458364 998844
rect 451246 998804 458364 998832
rect 378778 998724 378784 998776
rect 378836 998764 378842 998776
rect 383562 998764 383568 998776
rect 378836 998736 383568 998764
rect 378836 998724 378842 998736
rect 383562 998724 383568 998736
rect 383620 998724 383626 998776
rect 196802 998656 196808 998708
rect 196860 998696 196866 998708
rect 204346 998696 204352 998708
rect 196860 998668 204352 998696
rect 196860 998656 196866 998668
rect 204346 998656 204352 998668
rect 204404 998656 204410 998708
rect 351822 998656 351828 998708
rect 351880 998696 351886 998708
rect 378594 998696 378600 998708
rect 351880 998668 378600 998696
rect 351880 998656 351886 998668
rect 378594 998656 378600 998668
rect 378652 998656 378658 998708
rect 446398 998656 446404 998708
rect 446456 998696 446462 998708
rect 451246 998696 451274 998804
rect 458358 998792 458364 998804
rect 458416 998792 458422 998844
rect 462222 998792 462228 998844
rect 462280 998832 462286 998844
rect 472250 998832 472256 998844
rect 462280 998804 472256 998832
rect 462280 998792 462286 998804
rect 472250 998792 472256 998804
rect 472308 998792 472314 998844
rect 500954 998792 500960 998844
rect 501012 998832 501018 998844
rect 517514 998832 517520 998844
rect 501012 998804 517520 998832
rect 501012 998792 501018 998804
rect 517514 998792 517520 998804
rect 517572 998792 517578 998844
rect 446456 998668 451274 998696
rect 446456 998656 446462 998668
rect 458174 998656 458180 998708
rect 458232 998696 458238 998708
rect 472434 998696 472440 998708
rect 458232 998668 472440 998696
rect 458232 998656 458238 998668
rect 472434 998656 472440 998668
rect 472492 998656 472498 998708
rect 507026 998656 507032 998708
rect 507084 998696 507090 998708
rect 509878 998696 509884 998708
rect 507084 998668 509884 998696
rect 507084 998656 507090 998668
rect 509878 998656 509884 998668
rect 509936 998656 509942 998708
rect 510062 998656 510068 998708
rect 510120 998696 510126 998708
rect 518866 998696 518894 998872
rect 523862 998860 523868 998872
rect 523920 998860 523926 998912
rect 510120 998668 518894 998696
rect 510120 998656 510126 998668
rect 556798 998656 556804 998708
rect 556856 998696 556862 998708
rect 567470 998696 567476 998708
rect 556856 998668 567476 998696
rect 556856 998656 556862 998668
rect 567470 998656 567476 998668
rect 567528 998656 567534 998708
rect 92290 998520 92296 998572
rect 92348 998560 92354 998572
rect 92842 998560 92848 998572
rect 92348 998532 92848 998560
rect 92348 998520 92354 998532
rect 92842 998520 92848 998532
rect 92900 998520 92906 998572
rect 196618 998520 196624 998572
rect 196676 998560 196682 998572
rect 203518 998560 203524 998572
rect 196676 998532 203524 998560
rect 196676 998520 196682 998532
rect 203518 998520 203524 998532
rect 203576 998520 203582 998572
rect 355778 998520 355784 998572
rect 355836 998560 355842 998572
rect 383286 998560 383292 998572
rect 355836 998532 383292 998560
rect 355836 998520 355842 998532
rect 383286 998520 383292 998532
rect 383344 998520 383350 998572
rect 445018 998520 445024 998572
rect 445076 998560 445082 998572
rect 461578 998560 461584 998572
rect 445076 998532 461584 998560
rect 445076 998520 445082 998532
rect 461578 998520 461584 998532
rect 461636 998520 461642 998572
rect 463694 998520 463700 998572
rect 463752 998560 463758 998572
rect 472618 998560 472624 998572
rect 463752 998532 472624 998560
rect 463752 998520 463758 998532
rect 472618 998520 472624 998532
rect 472676 998520 472682 998572
rect 502150 998520 502156 998572
rect 502208 998560 502214 998572
rect 516686 998560 516692 998572
rect 502208 998532 516692 998560
rect 502208 998520 502214 998532
rect 516686 998520 516692 998532
rect 516744 998520 516750 998572
rect 516870 998520 516876 998572
rect 516928 998560 516934 998572
rect 524046 998560 524052 998572
rect 516928 998532 524052 998560
rect 516928 998520 516934 998532
rect 524046 998520 524052 998532
rect 524104 998520 524110 998572
rect 553762 998520 553768 998572
rect 553820 998560 553826 998572
rect 569126 998560 569132 998572
rect 553820 998532 569132 998560
rect 553820 998520 553826 998532
rect 569126 998520 569132 998532
rect 569184 998520 569190 998572
rect 247310 998452 247316 998504
rect 247368 998492 247374 998504
rect 247368 998464 253934 998492
rect 247368 998452 247374 998464
rect 92290 998384 92296 998436
rect 92348 998424 92354 998436
rect 100478 998424 100484 998436
rect 92348 998396 100484 998424
rect 92348 998384 92354 998396
rect 100478 998384 100484 998396
rect 100536 998384 100542 998436
rect 143994 998384 144000 998436
rect 144052 998424 144058 998436
rect 155954 998424 155960 998436
rect 144052 998396 155960 998424
rect 144052 998384 144058 998396
rect 155954 998384 155960 998396
rect 156012 998384 156018 998436
rect 195698 998384 195704 998436
rect 195756 998424 195762 998436
rect 204162 998424 204168 998436
rect 195756 998396 204168 998424
rect 195756 998384 195762 998396
rect 204162 998384 204168 998396
rect 204220 998384 204226 998436
rect 246758 998316 246764 998368
rect 246816 998356 246822 998368
rect 252462 998356 252468 998368
rect 246816 998328 252468 998356
rect 246816 998316 246822 998328
rect 252462 998316 252468 998328
rect 252520 998316 252526 998368
rect 200390 998180 200396 998232
rect 200448 998220 200454 998232
rect 203518 998220 203524 998232
rect 200448 998192 203524 998220
rect 200448 998180 200454 998192
rect 203518 998180 203524 998192
rect 203576 998180 203582 998232
rect 250438 998112 250444 998164
rect 250496 998152 250502 998164
rect 253658 998152 253664 998164
rect 250496 998124 253664 998152
rect 250496 998112 250502 998124
rect 253658 998112 253664 998124
rect 253716 998112 253722 998164
rect 199378 998044 199384 998096
rect 199436 998084 199442 998096
rect 202690 998084 202696 998096
rect 199436 998056 202696 998084
rect 199436 998044 199442 998056
rect 202690 998044 202696 998056
rect 202748 998044 202754 998096
rect 197538 997908 197544 997960
rect 197596 997948 197602 997960
rect 201862 997948 201868 997960
rect 197596 997920 201868 997948
rect 197596 997908 197602 997920
rect 201862 997908 201868 997920
rect 201920 997908 201926 997960
rect 202138 997908 202144 997960
rect 202196 997948 202202 997960
rect 205542 997948 205548 997960
rect 202196 997920 205548 997948
rect 202196 997908 202202 997920
rect 205542 997908 205548 997920
rect 205600 997908 205606 997960
rect 251174 997908 251180 997960
rect 251232 997948 251238 997960
rect 253658 997948 253664 997960
rect 251232 997920 253664 997948
rect 251232 997908 251238 997920
rect 253658 997908 253664 997920
rect 253716 997908 253722 997960
rect 92658 997772 92664 997824
rect 92716 997812 92722 997824
rect 121730 997812 121736 997824
rect 92716 997784 121736 997812
rect 92716 997772 92722 997784
rect 121730 997772 121736 997784
rect 121788 997772 121794 997824
rect 202322 997772 202328 997824
rect 202380 997812 202386 997824
rect 204714 997812 204720 997824
rect 202380 997784 204720 997812
rect 202380 997772 202386 997784
rect 204714 997772 204720 997784
rect 204772 997772 204778 997824
rect 247862 997772 247868 997824
rect 247920 997812 247926 997824
rect 252462 997812 252468 997824
rect 247920 997784 252468 997812
rect 247920 997772 247926 997784
rect 252462 997772 252468 997784
rect 252520 997772 252526 997824
rect 253906 997812 253934 998464
rect 354582 998384 354588 998436
rect 354640 998424 354646 998436
rect 383470 998424 383476 998436
rect 354640 998396 383476 998424
rect 354640 998384 354646 998396
rect 383470 998384 383476 998396
rect 383528 998384 383534 998436
rect 428182 998384 428188 998436
rect 428240 998424 428246 998436
rect 472066 998424 472072 998436
rect 428240 998396 472072 998424
rect 428240 998384 428246 998396
rect 472066 998384 472072 998396
rect 472124 998384 472130 998436
rect 500770 998384 500776 998436
rect 500828 998424 500834 998436
rect 523678 998424 523684 998436
rect 500828 998396 523684 998424
rect 500828 998384 500834 998396
rect 523678 998384 523684 998396
rect 523736 998384 523742 998436
rect 549162 998384 549168 998436
rect 549220 998424 549226 998436
rect 564434 998424 564440 998436
rect 549220 998396 564440 998424
rect 549220 998384 549226 998396
rect 564434 998384 564440 998396
rect 564492 998384 564498 998436
rect 591114 998384 591120 998436
rect 591172 998424 591178 998436
rect 617334 998424 617340 998436
rect 591172 998396 617340 998424
rect 591172 998384 591178 998396
rect 617334 998384 617340 998396
rect 617392 998384 617398 998436
rect 371878 998248 371884 998300
rect 371936 998288 371942 998300
rect 372982 998288 372988 998300
rect 371936 998260 372988 998288
rect 371936 998248 371942 998260
rect 372982 998248 372988 998260
rect 373040 998248 373046 998300
rect 378594 998248 378600 998300
rect 378652 998288 378658 998300
rect 382458 998288 382464 998300
rect 378652 998260 382464 998288
rect 378652 998248 378658 998260
rect 382458 998248 382464 998260
rect 382516 998248 382522 998300
rect 430850 998248 430856 998300
rect 430908 998288 430914 998300
rect 433978 998288 433984 998300
rect 430908 998260 433984 998288
rect 430908 998248 430914 998260
rect 433978 998248 433984 998260
rect 434036 998248 434042 998300
rect 509050 998248 509056 998300
rect 509108 998288 509114 998300
rect 514018 998288 514024 998300
rect 509108 998260 514024 998288
rect 509108 998248 509114 998260
rect 514018 998248 514024 998260
rect 514076 998248 514082 998300
rect 550542 998248 550548 998300
rect 550600 998288 550606 998300
rect 552934 998288 552940 998300
rect 550600 998260 552940 998288
rect 550600 998248 550606 998260
rect 552934 998248 552940 998260
rect 552992 998248 552998 998300
rect 430022 998112 430028 998164
rect 430080 998152 430086 998164
rect 432598 998152 432604 998164
rect 430080 998124 432604 998152
rect 430080 998112 430086 998124
rect 432598 998112 432604 998124
rect 432656 998112 432662 998164
rect 508222 998112 508228 998164
rect 508280 998152 508286 998164
rect 511258 998152 511264 998164
rect 508280 998124 511264 998152
rect 508280 998112 508286 998124
rect 511258 998112 511264 998124
rect 511316 998112 511322 998164
rect 432046 997976 432052 998028
rect 432104 998016 432110 998028
rect 436738 998016 436744 998028
rect 432104 997988 436744 998016
rect 432104 997976 432110 997988
rect 436738 997976 436744 997988
rect 436796 997976 436802 998028
rect 508222 997908 508228 997960
rect 508280 997948 508286 997960
rect 510706 997948 510712 997960
rect 508280 997920 510712 997948
rect 508280 997908 508286 997920
rect 510706 997908 510712 997920
rect 510764 997908 510770 997960
rect 430022 997840 430028 997892
rect 430080 997880 430086 997892
rect 432046 997880 432052 997892
rect 430080 997852 432052 997880
rect 430080 997840 430086 997852
rect 432046 997840 432052 997852
rect 432104 997840 432110 997892
rect 278222 997812 278228 997824
rect 253906 997784 278228 997812
rect 278222 997772 278228 997784
rect 278280 997772 278286 997824
rect 377398 997772 377404 997824
rect 377456 997812 377462 997824
rect 383102 997812 383108 997824
rect 377456 997784 383108 997812
rect 377456 997772 377462 997784
rect 383102 997772 383108 997784
rect 383160 997772 383166 997824
rect 591298 997772 591304 997824
rect 591356 997812 591362 997824
rect 625798 997812 625804 997824
rect 591356 997784 625804 997812
rect 591356 997772 591362 997784
rect 625798 997772 625804 997784
rect 625856 997772 625862 997824
rect 143810 997704 143816 997756
rect 143868 997744 143874 997756
rect 153930 997744 153936 997756
rect 143868 997716 153936 997744
rect 143868 997704 143874 997716
rect 153930 997704 153936 997716
rect 153988 997704 153994 997756
rect 298830 997704 298836 997756
rect 298888 997744 298894 997756
rect 311894 997744 311900 997756
rect 298888 997716 311900 997744
rect 298888 997704 298894 997716
rect 311894 997704 311900 997716
rect 311952 997704 311958 997756
rect 358814 997704 358820 997756
rect 358872 997744 358878 997756
rect 372338 997744 372344 997756
rect 358872 997716 372344 997744
rect 358872 997704 358878 997716
rect 372338 997704 372344 997716
rect 372396 997704 372402 997756
rect 431218 997704 431224 997756
rect 431276 997744 431282 997756
rect 439682 997744 439688 997756
rect 431276 997716 439688 997744
rect 431276 997704 431282 997716
rect 439682 997704 439688 997716
rect 439740 997704 439746 997756
rect 488902 997704 488908 997756
rect 488960 997744 488966 997756
rect 509234 997744 509240 997756
rect 488960 997716 509240 997744
rect 488960 997704 488966 997716
rect 509234 997704 509240 997716
rect 509292 997704 509298 997756
rect 509878 997704 509884 997756
rect 509936 997744 509942 997756
rect 516870 997744 516876 997756
rect 509936 997716 516876 997744
rect 509936 997704 509942 997716
rect 516870 997704 516876 997716
rect 516928 997704 516934 997756
rect 92474 997636 92480 997688
rect 92532 997676 92538 997688
rect 101582 997676 101588 997688
rect 92532 997648 101588 997676
rect 92532 997636 92538 997648
rect 101582 997636 101588 997648
rect 101640 997636 101646 997688
rect 109494 997636 109500 997688
rect 109552 997676 109558 997688
rect 117222 997676 117228 997688
rect 109552 997648 117228 997676
rect 109552 997636 109558 997648
rect 117222 997636 117228 997648
rect 117280 997636 117286 997688
rect 246666 997636 246672 997688
rect 246724 997676 246730 997688
rect 258074 997676 258080 997688
rect 246724 997648 258080 997676
rect 246724 997636 246730 997648
rect 258074 997636 258080 997648
rect 258132 997636 258138 997688
rect 569494 997636 569500 997688
rect 569552 997676 569558 997688
rect 623682 997676 623688 997688
rect 569552 997648 623688 997676
rect 569552 997636 569558 997648
rect 623682 997636 623688 997648
rect 623740 997636 623746 997688
rect 144822 997568 144828 997620
rect 144880 997608 144886 997620
rect 160094 997608 160100 997620
rect 144880 997580 160100 997608
rect 144880 997568 144886 997580
rect 160094 997568 160100 997580
rect 160152 997568 160158 997620
rect 299474 997568 299480 997620
rect 299532 997608 299538 997620
rect 310514 997608 310520 997620
rect 299532 997580 310520 997608
rect 299532 997568 299538 997580
rect 310514 997568 310520 997580
rect 310572 997568 310578 997620
rect 365162 997568 365168 997620
rect 365220 997608 365226 997620
rect 372522 997608 372528 997620
rect 365220 997580 372528 997608
rect 365220 997568 365226 997580
rect 372522 997568 372528 997580
rect 372580 997568 372586 997620
rect 433978 997568 433984 997620
rect 434036 997608 434042 997620
rect 439866 997608 439872 997620
rect 434036 997580 439872 997608
rect 434036 997568 434042 997580
rect 439866 997568 439872 997580
rect 439924 997568 439930 997620
rect 489086 997568 489092 997620
rect 489144 997608 489150 997620
rect 510706 997608 510712 997620
rect 489144 997580 510712 997608
rect 489144 997568 489150 997580
rect 510706 997568 510712 997580
rect 510764 997568 510770 997620
rect 113818 997500 113824 997552
rect 113876 997540 113882 997552
rect 116946 997540 116952 997552
rect 113876 997512 116952 997540
rect 113876 997500 113882 997512
rect 116946 997500 116952 997512
rect 117004 997500 117010 997552
rect 550542 997500 550548 997552
rect 550600 997540 550606 997552
rect 618162 997540 618168 997552
rect 550600 997512 618168 997540
rect 550600 997500 550606 997512
rect 618162 997500 618168 997512
rect 618220 997500 618226 997552
rect 432598 997432 432604 997484
rect 432656 997472 432662 997484
rect 440050 997472 440056 997484
rect 432656 997444 440056 997472
rect 432656 997432 432662 997444
rect 440050 997432 440056 997444
rect 440108 997432 440114 997484
rect 500586 997432 500592 997484
rect 500644 997472 500650 997484
rect 516686 997472 516692 997484
rect 500644 997444 516692 997472
rect 500644 997432 500650 997444
rect 516686 997432 516692 997444
rect 516744 997432 516750 997484
rect 540330 997364 540336 997416
rect 540388 997404 540394 997416
rect 555418 997404 555424 997416
rect 540388 997376 555424 997404
rect 540388 997364 540394 997376
rect 555418 997364 555424 997376
rect 555476 997364 555482 997416
rect 590378 997404 590384 997416
rect 560266 997376 590384 997404
rect 200206 997228 200212 997280
rect 200264 997268 200270 997280
rect 205082 997268 205088 997280
rect 200264 997240 205088 997268
rect 200264 997228 200270 997240
rect 205082 997228 205088 997240
rect 205140 997228 205146 997280
rect 552290 997228 552296 997280
rect 552348 997268 552354 997280
rect 560266 997268 560294 997376
rect 590378 997364 590384 997376
rect 590436 997364 590442 997416
rect 552348 997240 560294 997268
rect 552348 997228 552354 997240
rect 573542 997228 573548 997280
rect 573600 997268 573606 997280
rect 591298 997268 591304 997280
rect 573600 997240 591304 997268
rect 573600 997228 573606 997240
rect 591298 997228 591304 997240
rect 591356 997228 591362 997280
rect 160738 997160 160744 997212
rect 160796 997200 160802 997212
rect 162946 997200 162952 997212
rect 160796 997172 162952 997200
rect 160796 997160 160802 997172
rect 162946 997160 162952 997172
rect 163004 997160 163010 997212
rect 399938 997092 399944 997144
rect 399996 997132 400002 997144
rect 432046 997132 432052 997144
rect 399996 997104 432052 997132
rect 399996 997092 400002 997104
rect 432046 997092 432052 997104
rect 432104 997092 432110 997144
rect 571334 997092 571340 997144
rect 571392 997132 571398 997144
rect 591114 997132 591120 997144
rect 571392 997104 591120 997132
rect 571392 997092 571398 997104
rect 591114 997092 591120 997104
rect 591172 997092 591178 997144
rect 144638 997024 144644 997076
rect 144696 997064 144702 997076
rect 158714 997064 158720 997076
rect 144696 997036 158720 997064
rect 144696 997024 144702 997036
rect 158714 997024 158720 997036
rect 158772 997024 158778 997076
rect 197354 997024 197360 997076
rect 197412 997064 197418 997076
rect 226334 997064 226340 997076
rect 197412 997036 226340 997064
rect 197412 997024 197418 997036
rect 226334 997024 226340 997036
rect 226392 997024 226398 997076
rect 320818 997024 320824 997076
rect 320876 997064 320882 997076
rect 332594 997064 332600 997076
rect 320876 997036 332600 997064
rect 320876 997024 320882 997036
rect 332594 997024 332600 997036
rect 332652 997024 332658 997076
rect 448974 997024 448980 997076
rect 449032 997064 449038 997076
rect 470502 997064 470508 997076
rect 449032 997036 470508 997064
rect 449032 997024 449038 997036
rect 470502 997024 470508 997036
rect 470560 997024 470566 997076
rect 498194 997024 498200 997076
rect 498252 997064 498258 997076
rect 517698 997064 517704 997076
rect 498252 997036 517704 997064
rect 498252 997024 498258 997036
rect 517698 997024 517704 997036
rect 517756 997024 517762 997076
rect 565814 996888 565820 996940
rect 565872 996928 565878 996940
rect 590562 996928 590568 996940
rect 565872 996900 590568 996928
rect 565872 996888 565878 996900
rect 590562 996888 590568 996900
rect 590620 996888 590626 996940
rect 553210 996752 553216 996804
rect 553268 996792 553274 996804
rect 553268 996764 586514 996792
rect 553268 996752 553274 996764
rect 586486 996724 586514 996764
rect 590562 996724 590568 996736
rect 586486 996696 590568 996724
rect 590562 996684 590568 996696
rect 590620 996684 590626 996736
rect 564434 996616 564440 996668
rect 564492 996656 564498 996668
rect 568850 996656 568856 996668
rect 564492 996628 568856 996656
rect 564492 996616 564498 996628
rect 568850 996616 568856 996628
rect 568908 996616 568914 996668
rect 143718 996344 143724 996396
rect 143776 996384 143782 996396
rect 151262 996384 151268 996396
rect 143776 996356 151268 996384
rect 143776 996344 143782 996356
rect 151262 996344 151268 996356
rect 151320 996344 151326 996396
rect 298646 996344 298652 996396
rect 298704 996384 298710 996396
rect 365162 996384 365168 996396
rect 298704 996356 365168 996384
rect 298704 996344 298710 996356
rect 365162 996344 365168 996356
rect 365220 996344 365226 996396
rect 262858 996276 262864 996328
rect 262916 996316 262922 996328
rect 270402 996316 270408 996328
rect 262916 996288 270408 996316
rect 262916 996276 262922 996288
rect 270402 996276 270408 996288
rect 270460 996276 270466 996328
rect 556338 996276 556344 996328
rect 556396 996316 556402 996328
rect 590378 996316 590384 996328
rect 556396 996288 590384 996316
rect 556396 996276 556402 996288
rect 590378 996276 590384 996288
rect 590436 996276 590442 996328
rect 195606 996208 195612 996260
rect 195664 996248 195670 996260
rect 200666 996248 200672 996260
rect 195664 996220 200672 996248
rect 195664 996208 195670 996220
rect 200666 996208 200672 996220
rect 200724 996208 200730 996260
rect 195256 996152 195468 996180
rect 171778 996072 171784 996124
rect 171836 996112 171842 996124
rect 195256 996112 195284 996152
rect 171836 996084 195284 996112
rect 195440 996112 195468 996152
rect 567470 996140 567476 996192
rect 567528 996180 567534 996192
rect 590562 996180 590568 996192
rect 567528 996152 590568 996180
rect 567528 996140 567534 996152
rect 590562 996140 590568 996152
rect 590620 996140 590626 996192
rect 211154 996112 211160 996124
rect 195440 996084 211160 996112
rect 171836 996072 171842 996084
rect 211154 996072 211160 996084
rect 211212 996072 211218 996124
rect 229738 996072 229744 996124
rect 229796 996112 229802 996124
rect 262214 996112 262220 996124
rect 229796 996084 262220 996112
rect 229796 996072 229802 996084
rect 262214 996072 262220 996084
rect 262272 996072 262278 996124
rect 269758 996072 269764 996124
rect 269816 996112 269822 996124
rect 316034 996112 316040 996124
rect 269816 996084 316040 996112
rect 269816 996072 269822 996084
rect 316034 996072 316040 996084
rect 316092 996072 316098 996124
rect 366358 996072 366364 996124
rect 366416 996112 366422 996124
rect 402238 996112 402244 996124
rect 366416 996084 402244 996112
rect 366416 996072 366422 996084
rect 402238 996072 402244 996084
rect 402296 996072 402302 996124
rect 511258 996072 511264 996124
rect 511316 996112 511322 996124
rect 563054 996112 563060 996124
rect 511316 996084 563060 996112
rect 511316 996072 511322 996084
rect 563054 996072 563060 996084
rect 563112 996072 563118 996124
rect 170674 995936 170680 995988
rect 170732 995976 170738 995988
rect 171226 995976 171232 995988
rect 170732 995948 171232 995976
rect 170732 995936 170738 995948
rect 171226 995936 171232 995948
rect 171284 995936 171290 995988
rect 195882 995936 195888 995988
rect 195940 995976 195946 995988
rect 202506 995976 202512 995988
rect 195940 995948 202512 995976
rect 195940 995936 195946 995948
rect 202506 995936 202512 995948
rect 202564 995936 202570 995988
rect 213178 995936 213184 995988
rect 213236 995976 213242 995988
rect 261110 995976 261116 995988
rect 213236 995948 261116 995976
rect 213236 995936 213242 995948
rect 261110 995936 261116 995948
rect 261168 995936 261174 995988
rect 264238 995936 264244 995988
rect 264296 995976 264302 995988
rect 299198 995976 299204 995988
rect 264296 995948 299204 995976
rect 264296 995936 264302 995948
rect 299198 995936 299204 995948
rect 299256 995936 299262 995988
rect 364978 995936 364984 995988
rect 365036 995976 365042 995988
rect 400858 995976 400864 995988
rect 365036 995948 400864 995976
rect 365036 995936 365042 995948
rect 400858 995936 400864 995948
rect 400916 995936 400922 995988
rect 522298 995936 522304 995988
rect 522356 995976 522362 995988
rect 560294 995976 560300 995988
rect 522356 995948 560300 995976
rect 522356 995936 522362 995948
rect 560294 995936 560300 995948
rect 560352 995936 560358 995988
rect 92658 995800 92664 995852
rect 92716 995840 92722 995852
rect 97442 995840 97448 995852
rect 92716 995812 97448 995840
rect 92716 995800 92722 995812
rect 97442 995800 97448 995812
rect 97500 995800 97506 995852
rect 140774 995800 140780 995852
rect 140832 995840 140838 995852
rect 143994 995840 144000 995852
rect 140832 995812 144000 995840
rect 140832 995800 140838 995812
rect 143994 995800 144000 995812
rect 144052 995800 144058 995852
rect 169386 995800 169392 995852
rect 169444 995840 169450 995852
rect 171502 995840 171508 995852
rect 169444 995812 171508 995840
rect 169444 995800 169450 995812
rect 171502 995800 171508 995812
rect 171560 995800 171566 995852
rect 211798 995800 211804 995852
rect 211856 995840 211862 995852
rect 260926 995840 260932 995852
rect 211856 995812 260932 995840
rect 211856 995800 211862 995812
rect 260926 995800 260932 995812
rect 260984 995800 260990 995852
rect 360838 995800 360844 995852
rect 360896 995840 360902 995852
rect 399846 995840 399852 995852
rect 360896 995812 399852 995840
rect 360896 995800 360902 995812
rect 399846 995800 399852 995812
rect 399904 995800 399910 995852
rect 517514 995800 517520 995852
rect 517572 995840 517578 995852
rect 523310 995840 523316 995852
rect 517572 995812 523316 995840
rect 517572 995800 517578 995812
rect 523310 995800 523316 995812
rect 523368 995800 523374 995852
rect 92474 995528 92480 995580
rect 92532 995568 92538 995580
rect 98822 995568 98828 995580
rect 92532 995540 98828 995568
rect 92532 995528 92538 995540
rect 98822 995528 98828 995540
rect 98880 995528 98886 995580
rect 143718 995528 143724 995580
rect 143776 995568 143782 995580
rect 145742 995568 145748 995580
rect 143776 995540 145748 995568
rect 143776 995528 143782 995540
rect 145742 995528 145748 995540
rect 145800 995528 145806 995580
rect 171042 995528 171048 995580
rect 171100 995568 171106 995580
rect 171100 995540 171916 995568
rect 171100 995528 171106 995540
rect 171888 995415 171916 995540
rect 297818 995528 297824 995580
rect 297876 995568 297882 995580
rect 298462 995568 298468 995580
rect 297876 995540 298468 995568
rect 297876 995528 297882 995540
rect 298462 995528 298468 995540
rect 298520 995528 298526 995580
rect 383102 995528 383108 995580
rect 383160 995568 383166 995580
rect 385678 995568 385684 995580
rect 383160 995540 385684 995568
rect 383160 995528 383166 995540
rect 385678 995528 385684 995540
rect 385736 995528 385742 995580
rect 472434 995528 472440 995580
rect 472492 995568 472498 995580
rect 473354 995568 473360 995580
rect 472492 995540 473360 995568
rect 472492 995528 472498 995540
rect 473354 995528 473360 995540
rect 473412 995528 473418 995580
rect 623682 995528 623688 995580
rect 623740 995568 623746 995580
rect 626534 995568 626540 995580
rect 623740 995540 626540 995568
rect 623740 995528 623746 995540
rect 626534 995528 626540 995540
rect 626592 995528 626598 995580
rect 194870 995460 194876 995512
rect 194928 995500 194934 995512
rect 195698 995500 195704 995512
rect 194928 995472 195704 995500
rect 194928 995460 194934 995472
rect 195698 995460 195704 995472
rect 195756 995460 195762 995512
rect 246206 995460 246212 995512
rect 246264 995500 246270 995512
rect 247126 995500 247132 995512
rect 246264 995472 247132 995500
rect 246264 995460 246270 995472
rect 247126 995460 247132 995472
rect 247184 995460 247190 995512
rect 507026 995460 507032 995512
rect 507084 995500 507090 995512
rect 527910 995500 527916 995512
rect 507084 995472 527916 995500
rect 507084 995460 507090 995472
rect 527910 995460 527916 995472
rect 527968 995460 527974 995512
rect 629202 995460 629208 995512
rect 629260 995500 629266 995512
rect 631502 995500 631508 995512
rect 629260 995472 631508 995500
rect 629260 995460 629266 995472
rect 631502 995460 631508 995472
rect 631560 995460 631566 995512
rect 380158 995392 380164 995444
rect 380216 995432 380222 995444
rect 383102 995432 383108 995444
rect 380216 995404 383108 995432
rect 380216 995392 380222 995404
rect 383102 995392 383108 995404
rect 383160 995392 383166 995444
rect 383286 995392 383292 995444
rect 383344 995432 383350 995444
rect 388622 995432 388628 995444
rect 383344 995404 388628 995432
rect 383344 995392 383350 995404
rect 388622 995392 388628 995404
rect 388680 995392 388686 995444
rect 389082 995392 389088 995444
rect 389140 995432 389146 995444
rect 389726 995432 389732 995444
rect 389140 995404 389732 995432
rect 389140 995392 389146 995404
rect 389726 995392 389732 995404
rect 389784 995392 389790 995444
rect 415394 995392 415400 995444
rect 415452 995432 415458 995444
rect 415452 995404 415716 995432
rect 415452 995392 415458 995404
rect 415688 995387 415716 995404
rect 171686 995277 171692 995329
rect 171744 995277 171750 995329
rect 180702 995324 180708 995376
rect 180760 995364 180766 995376
rect 202138 995364 202144 995376
rect 180760 995336 202144 995364
rect 180760 995324 180766 995336
rect 202138 995324 202144 995336
rect 202196 995324 202202 995376
rect 236546 995324 236552 995376
rect 236604 995364 236610 995376
rect 251818 995364 251824 995376
rect 236604 995336 251824 995364
rect 236604 995324 236610 995336
rect 251818 995324 251824 995336
rect 251876 995324 251882 995376
rect 293586 995324 293592 995376
rect 293644 995364 293650 995376
rect 295978 995364 295984 995376
rect 293644 995336 295984 995364
rect 293644 995324 293650 995336
rect 295978 995324 295984 995336
rect 296036 995324 296042 995376
rect 296162 995324 296168 995376
rect 296220 995364 296226 995376
rect 298094 995364 298100 995376
rect 296220 995336 298100 995364
rect 296220 995324 296226 995336
rect 298094 995324 298100 995336
rect 298152 995324 298158 995376
rect 395246 995324 395252 995376
rect 395304 995364 395310 995376
rect 399846 995364 399852 995376
rect 395304 995336 399852 995364
rect 395304 995324 395310 995336
rect 399846 995324 399852 995336
rect 399904 995324 399910 995376
rect 415688 995359 415978 995387
rect 382182 995256 382188 995308
rect 382240 995296 382246 995308
rect 386322 995296 386328 995308
rect 382240 995268 386328 995296
rect 382240 995256 382246 995268
rect 386322 995256 386328 995268
rect 386380 995256 386386 995308
rect 386506 995256 386512 995308
rect 386564 995296 386570 995308
rect 386564 995268 391934 995296
rect 386564 995256 386570 995268
rect 171502 995165 171508 995217
rect 171560 995165 171566 995217
rect 182956 995188 182962 995240
rect 183014 995228 183020 995240
rect 208578 995228 208584 995240
rect 183014 995200 208584 995228
rect 183014 995188 183020 995200
rect 208578 995188 208584 995200
rect 208636 995188 208642 995240
rect 234384 995188 234390 995240
rect 234442 995228 234448 995240
rect 259454 995228 259460 995240
rect 234442 995200 259460 995228
rect 234442 995188 234448 995200
rect 259454 995188 259460 995200
rect 259512 995188 259518 995240
rect 285950 995188 285956 995240
rect 286008 995228 286014 995240
rect 309134 995228 309140 995240
rect 286008 995200 309140 995228
rect 286008 995188 286014 995200
rect 309134 995188 309140 995200
rect 309192 995188 309198 995240
rect 391906 995228 391934 995268
rect 398834 995228 398840 995240
rect 391906 995200 398840 995228
rect 398834 995188 398840 995200
rect 398892 995188 398898 995240
rect 416130 995235 416136 995287
rect 416188 995235 416194 995287
rect 362218 995120 362224 995172
rect 362276 995160 362282 995172
rect 388346 995160 388352 995172
rect 362276 995132 388352 995160
rect 362276 995120 362282 995132
rect 388346 995120 388352 995132
rect 388404 995120 388410 995172
rect 528922 995120 528928 995172
rect 528980 995160 528986 995172
rect 532878 995160 532884 995172
rect 528980 995132 532884 995160
rect 528980 995120 528986 995132
rect 532878 995120 532884 995132
rect 532936 995120 532942 995172
rect 533338 995120 533344 995172
rect 533396 995160 533402 995172
rect 534074 995160 534080 995172
rect 533396 995132 534080 995160
rect 533396 995120 533402 995132
rect 534074 995120 534080 995132
rect 534132 995120 534138 995172
rect 625246 995120 625252 995172
rect 625304 995160 625310 995172
rect 633986 995160 633992 995172
rect 625304 995132 633992 995160
rect 625304 995120 625310 995132
rect 633986 995120 633992 995132
rect 634044 995120 634050 995172
rect 660304 995147 660356 995153
rect 171232 995105 171284 995111
rect 171232 995047 171284 995053
rect 180150 995052 180156 995104
rect 180208 995092 180214 995104
rect 207014 995092 207020 995104
rect 180208 995064 207020 995092
rect 180208 995052 180214 995064
rect 207014 995052 207020 995064
rect 207072 995052 207078 995104
rect 231578 995052 231584 995104
rect 231636 995092 231642 995104
rect 257338 995092 257344 995104
rect 231636 995064 257344 995092
rect 231636 995052 231642 995064
rect 257338 995052 257344 995064
rect 257396 995052 257402 995104
rect 284110 995052 284116 995104
rect 284168 995092 284174 995104
rect 308398 995092 308404 995104
rect 284168 995064 308404 995092
rect 284168 995052 284174 995064
rect 308398 995052 308404 995064
rect 308456 995052 308462 995104
rect 454678 995052 454684 995104
rect 454736 995092 454742 995104
rect 485958 995092 485964 995104
rect 454736 995064 485964 995092
rect 454736 995052 454742 995064
rect 485958 995052 485964 995064
rect 486016 995052 486022 995104
rect 505738 995052 505744 995104
rect 505796 995092 505802 995104
rect 528738 995092 528744 995104
rect 505796 995064 528744 995092
rect 505796 995052 505802 995064
rect 528738 995052 528744 995064
rect 528796 995052 528802 995104
rect 569126 995052 569132 995104
rect 569184 995092 569190 995104
rect 625108 995092 625114 995104
rect 569184 995064 625114 995092
rect 569184 995052 569190 995064
rect 625108 995052 625114 995064
rect 625166 995052 625172 995104
rect 638862 995052 638868 995104
rect 638920 995092 638926 995104
rect 640794 995092 640800 995104
rect 638920 995064 640800 995092
rect 638920 995052 638926 995064
rect 640794 995052 640800 995064
rect 640852 995052 640858 995104
rect 660304 995089 660356 995095
rect 358078 994984 358084 995036
rect 358136 995024 358142 995036
rect 393314 995024 393320 995036
rect 358136 994996 393320 995024
rect 358136 994984 358142 994996
rect 393314 994984 393320 994996
rect 393372 994984 393378 995036
rect 641732 995023 660252 995024
rect 641732 994996 660606 995023
rect 171244 994881 171272 994967
rect 181438 994916 181444 994968
rect 181496 994956 181502 994968
rect 206278 994956 206284 994968
rect 181496 994928 206284 994956
rect 181496 994916 181502 994928
rect 206278 994916 206284 994928
rect 206336 994916 206342 994968
rect 232866 994916 232872 994968
rect 232924 994956 232930 994968
rect 255958 994956 255964 994968
rect 232924 994928 255964 994956
rect 232924 994916 232930 994928
rect 255958 994916 255964 994928
rect 256016 994916 256022 994968
rect 287146 994916 287152 994968
rect 287204 994956 287210 994968
rect 304258 994956 304264 994968
rect 287204 994928 304264 994956
rect 287204 994916 287210 994928
rect 304258 994916 304264 994928
rect 304316 994916 304322 994968
rect 420454 994916 420460 994968
rect 420512 994956 420518 994968
rect 641732 994956 641760 994996
rect 660224 994995 660606 994996
rect 420512 994928 641760 994956
rect 420512 994916 420518 994928
rect 80146 994780 80152 994832
rect 80204 994820 80210 994832
rect 106458 994820 106464 994832
rect 80204 994792 106464 994820
rect 80204 994780 80210 994792
rect 106458 994780 106464 994792
rect 106516 994780 106522 994832
rect 129734 994780 129740 994832
rect 129792 994820 129798 994832
rect 137094 994820 137100 994832
rect 129792 994792 137100 994820
rect 129792 994780 129798 994792
rect 137094 994780 137100 994792
rect 137152 994780 137158 994832
rect 137278 994780 137284 994832
rect 137336 994820 137342 994832
rect 137336 994792 151814 994820
rect 137336 994780 137342 994792
rect 77662 994644 77668 994696
rect 77720 994684 77726 994696
rect 100018 994684 100024 994696
rect 77720 994656 100024 994684
rect 77720 994644 77726 994656
rect 100018 994644 100024 994656
rect 100076 994644 100082 994696
rect 129090 994644 129096 994696
rect 129148 994684 129154 994696
rect 151078 994684 151084 994696
rect 129148 994656 151084 994684
rect 129148 994644 129154 994656
rect 151078 994644 151084 994656
rect 151136 994644 151142 994696
rect 151786 994684 151814 994792
rect 170490 994712 170496 994764
rect 170548 994752 170554 994764
rect 170876 994752 170904 994855
rect 171226 994829 171232 994881
rect 171284 994829 171290 994881
rect 363598 994848 363604 994900
rect 363656 994888 363662 994900
rect 397638 994888 397644 994900
rect 363656 994860 397644 994888
rect 363656 994848 363662 994860
rect 397638 994848 397644 994860
rect 397696 994848 397702 994900
rect 461578 994780 461584 994832
rect 461636 994820 461642 994832
rect 490006 994820 490012 994832
rect 461636 994792 490012 994820
rect 461636 994780 461642 994792
rect 490006 994780 490012 994792
rect 490064 994780 490070 994832
rect 496722 994780 496728 994832
rect 496780 994820 496786 994832
rect 513650 994820 513656 994832
rect 496780 994792 513656 994820
rect 496780 994780 496786 994792
rect 513650 994780 513656 994792
rect 513708 994780 513714 994832
rect 513834 994780 513840 994832
rect 513892 994820 513898 994832
rect 539226 994820 539232 994832
rect 513892 994792 539232 994820
rect 513892 994780 513898 994792
rect 539226 994780 539232 994792
rect 539284 994780 539290 994832
rect 551922 994780 551928 994832
rect 551980 994820 551986 994832
rect 634814 994820 634820 994832
rect 551980 994792 634820 994820
rect 551980 994780 551986 994792
rect 634814 994780 634820 994792
rect 634872 994780 634878 994832
rect 170548 994724 170904 994752
rect 170548 994712 170554 994724
rect 171042 994712 171048 994764
rect 171100 994752 171106 994764
rect 295058 994752 295064 994764
rect 171100 994724 295064 994752
rect 171100 994712 171106 994724
rect 295058 994712 295064 994724
rect 295116 994712 295122 994764
rect 376018 994712 376024 994764
rect 376076 994752 376082 994764
rect 393958 994752 393964 994764
rect 376076 994724 393964 994752
rect 376076 994712 376082 994724
rect 393958 994712 393964 994724
rect 394016 994712 394022 994764
rect 157334 994684 157340 994696
rect 151786 994656 157340 994684
rect 157334 994644 157340 994656
rect 157392 994644 157398 994696
rect 419442 994644 419448 994696
rect 419500 994684 419506 994696
rect 660298 994684 660304 994696
rect 419500 994656 660304 994684
rect 419500 994644 419506 994656
rect 660298 994644 660304 994656
rect 660356 994644 660362 994696
rect 660776 994628 660804 994897
rect 170674 994576 170680 994628
rect 170732 994616 170738 994628
rect 250438 994616 250444 994628
rect 170732 994588 250444 994616
rect 170732 994576 170738 994588
rect 250438 994576 250444 994588
rect 250496 994576 250502 994628
rect 283466 994576 283472 994628
rect 283524 994616 283530 994628
rect 305638 994616 305644 994628
rect 283524 994588 305644 994616
rect 283524 994576 283530 994588
rect 305638 994576 305644 994588
rect 305696 994576 305702 994628
rect 372982 994576 372988 994628
rect 373040 994616 373046 994628
rect 396994 994616 397000 994628
rect 373040 994588 397000 994616
rect 373040 994576 373046 994588
rect 396994 994576 397000 994588
rect 397052 994576 397058 994628
rect 660758 994576 660764 994628
rect 660816 994576 660822 994628
rect 660960 994560 660988 994785
rect 81342 994508 81348 994560
rect 81400 994548 81406 994560
rect 98638 994548 98644 994560
rect 81400 994520 98644 994548
rect 81400 994508 81406 994520
rect 98638 994508 98644 994520
rect 98696 994508 98702 994560
rect 132402 994508 132408 994560
rect 132460 994548 132466 994560
rect 149882 994548 149888 994560
rect 132460 994520 149888 994548
rect 132460 994508 132466 994520
rect 149882 994508 149888 994520
rect 149940 994508 149946 994560
rect 470502 994508 470508 994560
rect 470560 994548 470566 994560
rect 482278 994548 482284 994560
rect 470560 994520 482284 994548
rect 470560 994508 470566 994520
rect 482278 994508 482284 994520
rect 482336 994508 482342 994560
rect 482922 994508 482928 994560
rect 482980 994548 482986 994560
rect 489822 994548 489828 994560
rect 482980 994520 489828 994548
rect 482980 994508 482986 994520
rect 489822 994508 489828 994520
rect 489880 994508 489886 994560
rect 502334 994508 502340 994560
rect 502392 994548 502398 994560
rect 513834 994548 513840 994560
rect 502392 994520 513840 994548
rect 502392 994508 502398 994520
rect 513834 994508 513840 994520
rect 513892 994508 513898 994560
rect 514202 994508 514208 994560
rect 514260 994548 514266 994560
rect 523494 994548 523500 994560
rect 514260 994520 523500 994548
rect 514260 994508 514266 994520
rect 523494 994508 523500 994520
rect 523552 994508 523558 994560
rect 523678 994508 523684 994560
rect 523736 994548 523742 994560
rect 534350 994548 534356 994560
rect 523736 994520 534356 994548
rect 523736 994508 523742 994520
rect 534350 994508 534356 994520
rect 534408 994508 534414 994560
rect 573358 994508 573364 994560
rect 573416 994548 573422 994560
rect 590930 994548 590936 994560
rect 573416 994520 590936 994548
rect 573416 994508 573422 994520
rect 590930 994508 590936 994520
rect 590988 994508 590994 994560
rect 591298 994508 591304 994560
rect 591356 994548 591362 994560
rect 639046 994548 639052 994560
rect 591356 994520 639052 994548
rect 591356 994508 591362 994520
rect 639046 994508 639052 994520
rect 639104 994508 639110 994560
rect 660942 994508 660948 994560
rect 661000 994508 661006 994560
rect 170858 994440 170864 994492
rect 170916 994480 170922 994492
rect 298830 994480 298836 994492
rect 170916 994452 298836 994480
rect 170916 994440 170922 994452
rect 298830 994440 298836 994452
rect 298888 994440 298894 994492
rect 80698 994372 80704 994424
rect 80756 994412 80762 994424
rect 94498 994412 94504 994424
rect 80756 994384 94504 994412
rect 80756 994372 80762 994384
rect 94498 994372 94504 994384
rect 94556 994372 94562 994424
rect 128446 994372 128452 994424
rect 128504 994412 128510 994424
rect 137278 994412 137284 994424
rect 128504 994384 137284 994412
rect 128504 994372 128510 994384
rect 137278 994372 137284 994384
rect 137336 994372 137342 994424
rect 471422 994372 471428 994424
rect 471480 994412 471486 994424
rect 484578 994412 484584 994424
rect 471480 994384 484584 994412
rect 471480 994372 471486 994384
rect 484578 994372 484584 994384
rect 484636 994372 484642 994424
rect 500310 994372 500316 994424
rect 500368 994412 500374 994424
rect 534074 994412 534080 994424
rect 500368 994384 534080 994412
rect 500368 994372 500374 994384
rect 534074 994372 534080 994384
rect 534132 994372 534138 994424
rect 568850 994372 568856 994424
rect 568908 994412 568914 994424
rect 639506 994412 639512 994424
rect 568908 994384 639512 994412
rect 568908 994372 568914 994384
rect 639506 994372 639512 994384
rect 639564 994372 639570 994424
rect 184474 994304 184480 994356
rect 184532 994344 184538 994356
rect 191098 994344 191104 994356
rect 184532 994316 191104 994344
rect 184532 994304 184538 994316
rect 191098 994304 191104 994316
rect 191156 994304 191162 994356
rect 191742 994304 191748 994356
rect 191800 994344 191806 994356
rect 197354 994344 197360 994356
rect 191800 994316 197360 994344
rect 191800 994304 191806 994316
rect 197354 994304 197360 994316
rect 197412 994304 197418 994356
rect 137094 994236 137100 994288
rect 137152 994276 137158 994288
rect 144638 994276 144644 994288
rect 137152 994248 144644 994276
rect 137152 994236 137158 994248
rect 144638 994236 144644 994248
rect 144696 994236 144702 994288
rect 226334 994236 226340 994288
rect 226392 994276 226398 994288
rect 251450 994276 251456 994288
rect 226392 994248 251456 994276
rect 226392 994236 226398 994248
rect 251450 994236 251456 994248
rect 251508 994236 251514 994288
rect 278222 994236 278228 994288
rect 278280 994276 278286 994288
rect 316402 994276 316408 994288
rect 278280 994248 316408 994276
rect 278280 994236 278286 994248
rect 316402 994236 316408 994248
rect 316460 994236 316466 994288
rect 365162 994236 365168 994288
rect 365220 994276 365226 994288
rect 381170 994276 381176 994288
rect 365220 994248 381176 994276
rect 365220 994236 365226 994248
rect 381170 994236 381176 994248
rect 381228 994236 381234 994288
rect 414474 994236 414480 994288
rect 414532 994276 414538 994288
rect 446122 994276 446128 994288
rect 414532 994248 446128 994276
rect 414532 994236 414538 994248
rect 446122 994236 446128 994248
rect 446180 994236 446186 994288
rect 472066 994236 472072 994288
rect 472124 994276 472130 994288
rect 477954 994276 477960 994288
rect 472124 994248 477960 994276
rect 472124 994236 472130 994248
rect 477954 994236 477960 994248
rect 478012 994236 478018 994288
rect 513650 994236 513656 994288
rect 513708 994276 513714 994288
rect 514202 994276 514208 994288
rect 513708 994248 514208 994276
rect 513708 994236 513714 994248
rect 514202 994236 514208 994248
rect 514260 994236 514266 994288
rect 517698 994236 517704 994288
rect 517756 994276 517762 994288
rect 523678 994276 523684 994288
rect 517756 994248 523684 994276
rect 517756 994236 517762 994248
rect 523678 994236 523684 994248
rect 523736 994236 523742 994288
rect 538030 994276 538036 994288
rect 524386 994248 538036 994276
rect 139210 994100 139216 994152
rect 139268 994140 139274 994152
rect 142062 994140 142068 994152
rect 139268 994112 142068 994140
rect 139268 994100 139274 994112
rect 142062 994100 142068 994112
rect 142120 994100 142126 994152
rect 169386 994100 169392 994152
rect 169444 994140 169450 994152
rect 247862 994140 247868 994152
rect 169444 994112 247868 994140
rect 169444 994100 169450 994112
rect 247862 994100 247868 994112
rect 247920 994100 247926 994152
rect 295058 994100 295064 994152
rect 295116 994140 295122 994152
rect 300118 994140 300124 994152
rect 295116 994112 300124 994140
rect 295116 994100 295122 994112
rect 300118 994100 300124 994112
rect 300176 994100 300182 994152
rect 523494 994100 523500 994152
rect 523552 994140 523558 994152
rect 524386 994140 524414 994248
rect 538030 994236 538036 994248
rect 538088 994236 538094 994288
rect 570598 994236 570604 994288
rect 570656 994276 570662 994288
rect 591298 994276 591304 994288
rect 570656 994248 591304 994276
rect 570656 994236 570662 994248
rect 591298 994236 591304 994248
rect 591356 994236 591362 994288
rect 625430 994236 625436 994288
rect 625488 994276 625494 994288
rect 630858 994276 630864 994288
rect 625488 994248 630864 994276
rect 625488 994236 625494 994248
rect 630858 994236 630864 994248
rect 630916 994236 630922 994288
rect 523552 994112 524414 994140
rect 523552 994100 523558 994112
rect 574094 994032 574100 994084
rect 574152 994072 574158 994084
rect 661144 994072 661172 994673
rect 574152 994044 661172 994072
rect 574152 994032 574158 994044
rect 141878 993964 141884 994016
rect 141936 994004 141942 994016
rect 142338 994004 142344 994016
rect 141936 993976 142344 994004
rect 141936 993964 141942 993976
rect 142338 993964 142344 993976
rect 142396 993964 142402 994016
rect 191098 993964 191104 994016
rect 191156 994004 191162 994016
rect 196802 994004 196808 994016
rect 191156 993976 196808 994004
rect 191156 993964 191162 993976
rect 196802 993964 196808 993976
rect 196860 993964 196866 994016
rect 232222 993964 232228 994016
rect 232280 994004 232286 994016
rect 254578 994004 254584 994016
rect 232280 993976 254584 994004
rect 232280 993964 232286 993976
rect 254578 993964 254584 993976
rect 254636 993964 254642 994016
rect 569310 993896 569316 993948
rect 569368 993936 569374 993948
rect 661328 993936 661356 994561
rect 569368 993908 661356 993936
rect 569368 993896 569374 993908
rect 171226 993760 171232 993812
rect 171284 993800 171290 993812
rect 195514 993800 195520 993812
rect 171284 993772 195520 993800
rect 171284 993760 171290 993772
rect 195514 993760 195520 993772
rect 195572 993760 195578 993812
rect 521286 993760 521292 993812
rect 521344 993800 521350 993812
rect 660942 993800 660948 993812
rect 521344 993772 660948 993800
rect 521344 993760 521350 993772
rect 660942 993760 660948 993772
rect 661000 993760 661006 993812
rect 142154 993692 142160 993744
rect 142212 993732 142218 993744
rect 143902 993732 143908 993744
rect 142212 993704 143908 993732
rect 142212 993692 142218 993704
rect 143902 993692 143908 993704
rect 143960 993692 143966 993744
rect 170490 993624 170496 993676
rect 170548 993664 170554 993676
rect 197538 993664 197544 993676
rect 170548 993636 197544 993664
rect 170548 993624 170554 993636
rect 197538 993624 197544 993636
rect 197596 993624 197602 993676
rect 517054 993624 517060 993676
rect 517112 993664 517118 993676
rect 660758 993664 660764 993676
rect 517112 993636 660764 993664
rect 517112 993624 517118 993636
rect 660758 993624 660764 993636
rect 660816 993624 660822 993676
rect 188154 993488 188160 993540
rect 188212 993528 188218 993540
rect 195882 993528 195888 993540
rect 188212 993500 195888 993528
rect 188212 993488 188218 993500
rect 195882 993488 195888 993500
rect 195940 993488 195946 993540
rect 50338 993148 50344 993200
rect 50396 993188 50402 993200
rect 107746 993188 107752 993200
rect 50396 993160 107752 993188
rect 50396 993148 50402 993160
rect 107746 993148 107752 993160
rect 107804 993148 107810 993200
rect 44818 993012 44824 993064
rect 44876 993052 44882 993064
rect 109034 993052 109040 993064
rect 44876 993024 109040 993052
rect 44876 993012 44882 993024
rect 109034 993012 109040 993024
rect 109092 993012 109098 993064
rect 318058 993012 318064 993064
rect 318116 993052 318122 993064
rect 349154 993052 349160 993064
rect 318116 993024 349160 993052
rect 318116 993012 318122 993024
rect 349154 993012 349160 993024
rect 349212 993012 349218 993064
rect 562502 993012 562508 993064
rect 562560 993052 562566 993064
rect 660298 993052 660304 993064
rect 562560 993024 660304 993052
rect 562560 993012 562566 993024
rect 660298 993012 660304 993024
rect 660356 993012 660362 993064
rect 54478 992876 54484 992928
rect 54536 992916 54542 992928
rect 148318 992916 148324 992928
rect 54536 992888 148324 992916
rect 54536 992876 54542 992888
rect 148318 992876 148324 992888
rect 148376 992876 148382 992928
rect 319438 992876 319444 992928
rect 319496 992916 319502 992928
rect 364978 992916 364984 992928
rect 319496 992888 364984 992916
rect 319496 992876 319502 992888
rect 364978 992876 364984 992888
rect 365036 992876 365042 992928
rect 560938 992876 560944 992928
rect 560996 992916 561002 992928
rect 667198 992916 667204 992928
rect 560996 992888 667204 992916
rect 560996 992876 561002 992888
rect 667198 992876 667204 992888
rect 667256 992876 667262 992928
rect 47578 991720 47584 991772
rect 47636 991760 47642 991772
rect 96062 991760 96068 991772
rect 47636 991732 96068 991760
rect 47636 991720 47642 991732
rect 96062 991720 96068 991732
rect 96120 991720 96126 991772
rect 51718 991584 51724 991636
rect 51776 991624 51782 991636
rect 110414 991624 110420 991636
rect 51776 991596 110420 991624
rect 51776 991584 51782 991596
rect 110414 991584 110420 991596
rect 110472 991584 110478 991636
rect 138290 991584 138296 991636
rect 138348 991624 138354 991636
rect 163130 991624 163136 991636
rect 138348 991596 163136 991624
rect 138348 991584 138354 991596
rect 163130 991584 163136 991596
rect 163188 991584 163194 991636
rect 369118 991584 369124 991636
rect 369176 991624 369182 991636
rect 414106 991624 414112 991636
rect 369176 991596 414112 991624
rect 369176 991584 369182 991596
rect 414106 991584 414112 991596
rect 414164 991584 414170 991636
rect 55858 991448 55864 991500
rect 55916 991488 55922 991500
rect 146938 991488 146944 991500
rect 55916 991460 146944 991488
rect 55916 991448 55922 991460
rect 146938 991448 146944 991460
rect 146996 991448 147002 991500
rect 266998 991448 267004 991500
rect 267056 991488 267062 991500
rect 284294 991488 284300 991500
rect 267056 991460 284300 991488
rect 267056 991448 267062 991460
rect 284294 991448 284300 991460
rect 284352 991448 284358 991500
rect 367738 991448 367744 991500
rect 367796 991488 367802 991500
rect 430298 991488 430304 991500
rect 367796 991460 430304 991488
rect 367796 991448 367802 991460
rect 430298 991448 430304 991460
rect 430356 991448 430362 991500
rect 435358 991448 435364 991500
rect 435416 991488 435422 991500
rect 478966 991488 478972 991500
rect 435416 991460 478972 991488
rect 435416 991448 435422 991460
rect 478966 991448 478972 991460
rect 479024 991448 479030 991500
rect 559558 991448 559564 991500
rect 559616 991488 559622 991500
rect 658918 991488 658924 991500
rect 559616 991460 658924 991488
rect 559616 991448 559622 991460
rect 658918 991448 658924 991460
rect 658976 991448 658982 991500
rect 214558 991176 214564 991228
rect 214616 991216 214622 991228
rect 219434 991216 219440 991228
rect 214616 991188 219440 991216
rect 214616 991176 214622 991188
rect 219434 991176 219440 991188
rect 219492 991176 219498 991228
rect 164878 990836 164884 990888
rect 164936 990876 164942 990888
rect 170766 990876 170772 990888
rect 164936 990848 170772 990876
rect 164936 990836 164942 990848
rect 170766 990836 170772 990848
rect 170824 990836 170830 990888
rect 265618 990836 265624 990888
rect 265676 990876 265682 990888
rect 267642 990876 267648 990888
rect 265676 990848 267648 990876
rect 265676 990836 265682 990848
rect 267642 990836 267648 990848
rect 267700 990836 267706 990888
rect 572806 990836 572812 990888
rect 572864 990876 572870 990888
rect 576302 990876 576308 990888
rect 572864 990848 576308 990876
rect 572864 990836 572870 990848
rect 576302 990836 576308 990848
rect 576360 990836 576366 990888
rect 53282 990224 53288 990276
rect 53340 990264 53346 990276
rect 95878 990264 95884 990276
rect 53340 990236 95884 990264
rect 53340 990224 53346 990236
rect 95878 990224 95884 990236
rect 95936 990224 95942 990276
rect 48958 990088 48964 990140
rect 49016 990128 49022 990140
rect 108114 990128 108120 990140
rect 49016 990100 108120 990128
rect 49016 990088 49022 990100
rect 108114 990088 108120 990100
rect 108172 990088 108178 990140
rect 512638 990088 512644 990140
rect 512696 990128 512702 990140
rect 543826 990128 543832 990140
rect 512696 990100 543832 990128
rect 512696 990088 512702 990100
rect 543826 990088 543832 990100
rect 543884 990088 543890 990140
rect 562318 990088 562324 990140
rect 562376 990128 562382 990140
rect 668578 990128 668584 990140
rect 562376 990100 668584 990128
rect 562376 990088 562382 990100
rect 668578 990088 668584 990100
rect 668636 990088 668642 990140
rect 563698 987368 563704 987420
rect 563756 987408 563762 987420
rect 608778 987408 608784 987420
rect 563756 987380 608784 987408
rect 563756 987368 563762 987380
rect 608778 987368 608784 987380
rect 608836 987368 608842 987420
rect 203150 986620 203156 986672
rect 203208 986660 203214 986672
rect 204898 986660 204904 986672
rect 203208 986632 204904 986660
rect 203208 986620 203214 986632
rect 204898 986620 204904 986632
rect 204956 986620 204962 986672
rect 89622 986076 89628 986128
rect 89680 986116 89686 986128
rect 111794 986116 111800 986128
rect 89680 986088 111800 986116
rect 89680 986076 89686 986088
rect 111794 986076 111800 986088
rect 111852 986076 111858 986128
rect 438118 986076 438124 986128
rect 438176 986116 438182 986128
rect 462774 986116 462780 986128
rect 438176 986088 462780 986116
rect 438176 986076 438182 986088
rect 462774 986076 462780 986088
rect 462832 986076 462838 986128
rect 515398 986076 515404 986128
rect 515456 986116 515462 986128
rect 527634 986116 527640 986128
rect 515456 986088 527640 986116
rect 515456 986076 515462 986088
rect 527634 986076 527640 986088
rect 527692 986076 527698 986128
rect 566458 986076 566464 986128
rect 566516 986116 566522 986128
rect 592494 986116 592500 986128
rect 566516 986088 592500 986116
rect 566516 986076 566522 986088
rect 592494 986076 592500 986088
rect 592552 986076 592558 986128
rect 73430 985940 73436 985992
rect 73488 985980 73494 985992
rect 102778 985980 102784 985992
rect 73488 985952 102784 985980
rect 73488 985940 73494 985952
rect 102778 985940 102784 985952
rect 102836 985940 102842 985992
rect 215938 985940 215944 985992
rect 215996 985980 216002 985992
rect 235626 985980 235632 985992
rect 215996 985952 235632 985980
rect 215996 985940 216002 985952
rect 235626 985940 235632 985952
rect 235684 985940 235690 985992
rect 268378 985940 268384 985992
rect 268436 985980 268442 985992
rect 300486 985980 300492 985992
rect 268436 985952 300492 985980
rect 268436 985940 268442 985952
rect 300486 985940 300492 985952
rect 300544 985940 300550 985992
rect 370498 985940 370504 985992
rect 370556 985980 370562 985992
rect 397822 985980 397828 985992
rect 370556 985952 397828 985980
rect 370556 985940 370562 985952
rect 397822 985940 397828 985952
rect 397880 985940 397886 985992
rect 436738 985940 436744 985992
rect 436796 985980 436802 985992
rect 495158 985980 495164 985992
rect 436796 985952 495164 985980
rect 436796 985940 436802 985952
rect 495158 985940 495164 985952
rect 495216 985940 495222 985992
rect 514018 985940 514024 985992
rect 514076 985980 514082 985992
rect 560110 985980 560116 985992
rect 514076 985952 560116 985980
rect 514076 985940 514082 985952
rect 560110 985940 560116 985952
rect 560168 985940 560174 985992
rect 565078 985940 565084 985992
rect 565136 985980 565142 985992
rect 624970 985980 624976 985992
rect 565136 985952 624976 985980
rect 565136 985940 565142 985952
rect 624970 985940 624976 985952
rect 625028 985940 625034 985992
rect 154482 985668 154488 985720
rect 154540 985708 154546 985720
rect 160738 985708 160744 985720
rect 154540 985680 160744 985708
rect 154540 985668 154546 985680
rect 160738 985668 160744 985680
rect 160796 985668 160802 985720
rect 43438 975672 43444 975724
rect 43496 975712 43502 975724
rect 62114 975712 62120 975724
rect 43496 975684 62120 975712
rect 43496 975672 43502 975684
rect 62114 975672 62120 975684
rect 62172 975672 62178 975724
rect 651650 975672 651656 975724
rect 651708 975712 651714 975724
rect 664438 975712 664444 975724
rect 651708 975684 664444 975712
rect 651708 975672 651714 975684
rect 664438 975672 664444 975684
rect 664496 975672 664502 975724
rect 46198 961868 46204 961920
rect 46256 961908 46262 961920
rect 62114 961908 62120 961920
rect 46256 961880 62120 961908
rect 46256 961868 46262 961880
rect 62114 961868 62120 961880
rect 62172 961868 62178 961920
rect 651466 961868 651472 961920
rect 651524 961908 651530 961920
rect 665818 961908 665824 961920
rect 651524 961880 665824 961908
rect 651524 961868 651530 961880
rect 665818 961868 665824 961880
rect 665876 961868 665882 961920
rect 36538 952348 36544 952400
rect 36596 952388 36602 952400
rect 41690 952388 41696 952400
rect 36596 952360 41696 952388
rect 36596 952348 36602 952360
rect 41690 952348 41696 952360
rect 41748 952348 41754 952400
rect 33778 951464 33784 951516
rect 33836 951504 33842 951516
rect 41506 951504 41512 951516
rect 33836 951476 41512 951504
rect 33836 951464 33842 951476
rect 41506 951464 41512 951476
rect 41564 951464 41570 951516
rect 675846 949424 675852 949476
rect 675904 949464 675910 949476
rect 682378 949464 682384 949476
rect 675904 949436 682384 949464
rect 675904 949424 675910 949436
rect 682378 949424 682384 949436
rect 682436 949424 682442 949476
rect 652202 948064 652208 948116
rect 652260 948104 652266 948116
rect 663058 948104 663064 948116
rect 652260 948076 663064 948104
rect 652260 948064 652266 948076
rect 663058 948064 663064 948076
rect 663116 948064 663122 948116
rect 676030 947996 676036 948048
rect 676088 948036 676094 948048
rect 680998 948036 681004 948048
rect 676088 948008 681004 948036
rect 676088 947996 676094 948008
rect 680998 947996 681004 948008
rect 681056 947996 681062 948048
rect 45554 945956 45560 946008
rect 45612 945996 45618 946008
rect 62114 945996 62120 946008
rect 45612 945968 62120 945996
rect 45612 945956 45618 945968
rect 62114 945956 62120 945968
rect 62172 945956 62178 946008
rect 28718 945276 28724 945328
rect 28776 945316 28782 945328
rect 31754 945316 31760 945328
rect 28776 945288 31760 945316
rect 28776 945276 28782 945288
rect 31754 945276 31760 945288
rect 31812 945276 31818 945328
rect 35802 942556 35808 942608
rect 35860 942596 35866 942608
rect 41690 942596 41696 942608
rect 35860 942568 41696 942596
rect 35860 942556 35866 942568
rect 41690 942556 41696 942568
rect 41748 942556 41754 942608
rect 35802 941196 35808 941248
rect 35860 941236 35866 941248
rect 41414 941236 41420 941248
rect 35860 941208 41420 941236
rect 35860 941196 35866 941208
rect 41414 941196 41420 941208
rect 41472 941196 41478 941248
rect 35802 939768 35808 939820
rect 35860 939808 35866 939820
rect 41598 939808 41604 939820
rect 35860 939780 41604 939808
rect 35860 939768 35866 939780
rect 41598 939768 41604 939780
rect 41656 939768 41662 939820
rect 651466 936980 651472 937032
rect 651524 937020 651530 937032
rect 661678 937020 661684 937032
rect 651524 936992 661684 937020
rect 651524 936980 651530 936992
rect 661678 936980 661684 936992
rect 661736 936980 661742 937032
rect 675846 928752 675852 928804
rect 675904 928792 675910 928804
rect 683114 928792 683120 928804
rect 675904 928764 683120 928792
rect 675904 928752 675910 928764
rect 683114 928752 683120 928764
rect 683172 928752 683178 928804
rect 53098 923244 53104 923296
rect 53156 923284 53162 923296
rect 62114 923284 62120 923296
rect 53156 923256 62120 923284
rect 53156 923244 53162 923256
rect 62114 923244 62120 923256
rect 62172 923244 62178 923296
rect 651466 921816 651472 921868
rect 651524 921856 651530 921868
rect 661678 921856 661684 921868
rect 651524 921828 661684 921856
rect 651524 921816 651530 921828
rect 661678 921816 661684 921828
rect 661736 921816 661742 921868
rect 50338 909440 50344 909492
rect 50396 909480 50402 909492
rect 62114 909480 62120 909492
rect 50396 909452 62120 909480
rect 50396 909440 50402 909452
rect 62114 909440 62120 909452
rect 62172 909440 62178 909492
rect 652386 909440 652392 909492
rect 652444 909480 652450 909492
rect 663058 909480 663064 909492
rect 652444 909452 663064 909480
rect 652444 909440 652450 909452
rect 663058 909440 663064 909452
rect 663116 909440 663122 909492
rect 47762 896996 47768 897048
rect 47820 897036 47826 897048
rect 62114 897036 62120 897048
rect 47820 897008 62120 897036
rect 47820 896996 47826 897008
rect 62114 896996 62120 897008
rect 62172 896996 62178 897048
rect 651466 895636 651472 895688
rect 651524 895676 651530 895688
rect 671338 895676 671344 895688
rect 651524 895648 671344 895676
rect 651524 895636 651530 895648
rect 671338 895636 671344 895648
rect 671396 895636 671402 895688
rect 42846 892492 42898 892498
rect 42846 892434 42898 892440
rect 43070 892304 43076 892356
rect 43128 892304 43134 892356
rect 42938 892254 42990 892260
rect 42938 892196 42990 892202
rect 43088 892058 43116 892304
rect 44082 891936 44088 891948
rect 43180 891908 44088 891936
rect 43180 891854 43208 891908
rect 44082 891896 44088 891908
rect 44140 891896 44146 891948
rect 651650 881832 651656 881884
rect 651708 881872 651714 881884
rect 664438 881872 664444 881884
rect 651708 881844 664444 881872
rect 651708 881832 651714 881844
rect 664438 881832 664444 881844
rect 664496 881832 664502 881884
rect 46198 870816 46204 870868
rect 46256 870856 46262 870868
rect 62114 870856 62120 870868
rect 46256 870828 62120 870856
rect 46256 870816 46262 870828
rect 62114 870816 62120 870828
rect 62172 870816 62178 870868
rect 651466 869388 651472 869440
rect 651524 869428 651530 869440
rect 658918 869428 658924 869440
rect 651524 869400 658924 869428
rect 651524 869388 651530 869400
rect 658918 869388 658924 869400
rect 658976 869388 658982 869440
rect 652386 855584 652392 855636
rect 652444 855624 652450 855636
rect 664438 855624 664444 855636
rect 652444 855596 664444 855624
rect 652444 855584 652450 855596
rect 664438 855584 664444 855596
rect 664496 855584 664502 855636
rect 54478 844568 54484 844620
rect 54536 844608 54542 844620
rect 62114 844608 62120 844620
rect 54536 844580 62120 844608
rect 54536 844568 54542 844580
rect 62114 844568 62120 844580
rect 62172 844568 62178 844620
rect 55858 832124 55864 832176
rect 55916 832164 55922 832176
rect 62114 832164 62120 832176
rect 55916 832136 62120 832164
rect 55916 832124 55922 832136
rect 62114 832124 62120 832136
rect 62172 832124 62178 832176
rect 651466 829404 651472 829456
rect 651524 829444 651530 829456
rect 660298 829444 660304 829456
rect 651524 829416 660304 829444
rect 651524 829404 651530 829416
rect 660298 829404 660304 829416
rect 660356 829404 660362 829456
rect 47578 818320 47584 818372
rect 47636 818360 47642 818372
rect 62114 818360 62120 818372
rect 47636 818332 62120 818360
rect 47636 818320 47642 818332
rect 62114 818320 62120 818332
rect 62172 818320 62178 818372
rect 35802 817028 35808 817080
rect 35860 817068 35866 817080
rect 41690 817068 41696 817080
rect 35860 817040 41696 817068
rect 35860 817028 35866 817040
rect 41690 817028 41696 817040
rect 41748 817028 41754 817080
rect 35802 815600 35808 815652
rect 35860 815640 35866 815652
rect 41414 815640 41420 815652
rect 35860 815612 41420 815640
rect 35860 815600 35866 815612
rect 41414 815600 41420 815612
rect 41472 815600 41478 815652
rect 651466 815600 651472 815652
rect 651524 815640 651530 815652
rect 669958 815640 669964 815652
rect 651524 815612 669964 815640
rect 651524 815600 651530 815612
rect 669958 815600 669964 815612
rect 670016 815600 670022 815652
rect 35802 814240 35808 814292
rect 35860 814280 35866 814292
rect 41598 814280 41604 814292
rect 35860 814252 41604 814280
rect 35860 814240 35866 814252
rect 41598 814240 41604 814252
rect 41656 814240 41662 814292
rect 41322 811452 41328 811504
rect 41380 811492 41386 811504
rect 41690 811492 41696 811504
rect 41380 811464 41696 811492
rect 41380 811452 41386 811464
rect 41690 811452 41696 811464
rect 41748 811452 41754 811504
rect 40586 808256 40592 808308
rect 40644 808296 40650 808308
rect 41598 808296 41604 808308
rect 40644 808268 41604 808296
rect 40644 808256 40650 808268
rect 41598 808256 41604 808268
rect 41656 808256 41662 808308
rect 50338 805944 50344 805996
rect 50396 805984 50402 805996
rect 62114 805984 62120 805996
rect 50396 805956 62120 805984
rect 50396 805944 50402 805956
rect 62114 805944 62120 805956
rect 62172 805944 62178 805996
rect 651466 803224 651472 803276
rect 651524 803264 651530 803276
rect 651524 803236 654134 803264
rect 651524 803224 651530 803236
rect 654106 803196 654134 803236
rect 667198 803196 667204 803208
rect 654106 803168 667204 803196
rect 667198 803156 667204 803168
rect 667256 803156 667262 803208
rect 35158 802408 35164 802460
rect 35216 802448 35222 802460
rect 41690 802448 41696 802460
rect 35216 802420 41696 802448
rect 35216 802408 35222 802420
rect 41690 802408 41696 802420
rect 41748 802408 41754 802460
rect 35894 802272 35900 802324
rect 35952 802312 35958 802324
rect 41690 802312 41696 802324
rect 35952 802284 41696 802312
rect 35952 802272 35958 802284
rect 41690 802272 41696 802284
rect 41748 802272 41754 802324
rect 651466 789352 651472 789404
rect 651524 789392 651530 789404
rect 668578 789392 668584 789404
rect 651524 789364 668584 789392
rect 651524 789352 651530 789364
rect 668578 789352 668584 789364
rect 668636 789352 668642 789404
rect 651466 775548 651472 775600
rect 651524 775588 651530 775600
rect 668762 775588 668768 775600
rect 651524 775560 668768 775588
rect 651524 775548 651530 775560
rect 668762 775548 668768 775560
rect 668820 775548 668826 775600
rect 35802 772828 35808 772880
rect 35860 772868 35866 772880
rect 41690 772868 41696 772880
rect 35860 772840 41696 772868
rect 35860 772828 35866 772840
rect 41690 772828 41696 772840
rect 41748 772828 41754 772880
rect 35802 768952 35808 769004
rect 35860 768992 35866 769004
rect 41322 768992 41328 769004
rect 35860 768964 41328 768992
rect 35860 768952 35866 768964
rect 41322 768952 41328 768964
rect 41380 768952 41386 769004
rect 35618 768816 35624 768868
rect 35676 768856 35682 768868
rect 41690 768856 41696 768868
rect 35676 768828 41696 768856
rect 35676 768816 35682 768828
rect 41690 768816 41696 768828
rect 41748 768816 41754 768868
rect 35434 768680 35440 768732
rect 35492 768720 35498 768732
rect 40034 768720 40040 768732
rect 35492 768692 40040 768720
rect 35492 768680 35498 768692
rect 40034 768680 40040 768692
rect 40092 768680 40098 768732
rect 35802 767524 35808 767576
rect 35860 767564 35866 767576
rect 35860 767524 35894 767564
rect 35866 767496 35894 767524
rect 37918 767496 37924 767508
rect 35866 767468 37924 767496
rect 37918 767456 37924 767468
rect 37976 767456 37982 767508
rect 35802 767320 35808 767372
rect 35860 767360 35866 767372
rect 36538 767360 36544 767372
rect 35860 767332 36544 767360
rect 35860 767320 35866 767332
rect 36538 767320 36544 767332
rect 36596 767320 36602 767372
rect 48958 767320 48964 767372
rect 49016 767360 49022 767372
rect 62114 767360 62120 767372
rect 49016 767332 62120 767360
rect 49016 767320 49022 767332
rect 62114 767320 62120 767332
rect 62172 767320 62178 767372
rect 37090 763240 37096 763292
rect 37148 763280 37154 763292
rect 39298 763280 39304 763292
rect 37148 763252 39304 763280
rect 37148 763240 37154 763252
rect 39298 763240 39304 763252
rect 39356 763240 39362 763292
rect 651466 763240 651472 763292
rect 651524 763280 651530 763292
rect 651524 763252 654134 763280
rect 651524 763240 651530 763252
rect 654106 763212 654134 763252
rect 660298 763212 660304 763224
rect 654106 763184 660304 763212
rect 660298 763172 660304 763184
rect 660356 763172 660362 763224
rect 37918 759092 37924 759144
rect 37976 759132 37982 759144
rect 40862 759132 40868 759144
rect 37976 759104 40868 759132
rect 37976 759092 37982 759104
rect 40862 759092 40868 759104
rect 40920 759092 40926 759144
rect 35158 758956 35164 759008
rect 35216 758996 35222 759008
rect 40310 758996 40316 759008
rect 35216 758968 40316 758996
rect 35216 758956 35222 758968
rect 40310 758956 40316 758968
rect 40368 758956 40374 759008
rect 31018 758276 31024 758328
rect 31076 758316 31082 758328
rect 40586 758316 40592 758328
rect 31076 758288 40592 758316
rect 31076 758276 31082 758288
rect 40586 758276 40592 758288
rect 40644 758276 40650 758328
rect 676030 757120 676036 757172
rect 676088 757160 676094 757172
rect 683114 757160 683120 757172
rect 676088 757132 683120 757160
rect 676088 757120 676094 757132
rect 683114 757120 683120 757132
rect 683172 757120 683178 757172
rect 51718 753516 51724 753568
rect 51776 753556 51782 753568
rect 62114 753556 62120 753568
rect 51776 753528 62120 753556
rect 51776 753516 51782 753528
rect 62114 753516 62120 753528
rect 62172 753516 62178 753568
rect 651466 749368 651472 749420
rect 651524 749408 651530 749420
rect 665818 749408 665824 749420
rect 651524 749380 665824 749408
rect 651524 749368 651530 749380
rect 665818 749368 665824 749380
rect 665876 749368 665882 749420
rect 54478 741072 54484 741124
rect 54536 741112 54542 741124
rect 62114 741112 62120 741124
rect 54536 741084 62120 741112
rect 54536 741072 54542 741084
rect 62114 741072 62120 741084
rect 62172 741072 62178 741124
rect 652570 735564 652576 735616
rect 652628 735604 652634 735616
rect 671338 735604 671344 735616
rect 652628 735576 671344 735604
rect 652628 735564 652634 735576
rect 671338 735564 671344 735576
rect 671396 735564 671402 735616
rect 673546 732096 673552 732148
rect 673604 732136 673610 732148
rect 674006 732136 674012 732148
rect 673604 732108 674012 732136
rect 673604 732096 673610 732108
rect 674006 732096 674012 732108
rect 674064 732096 674070 732148
rect 35618 730192 35624 730244
rect 35676 730232 35682 730244
rect 41690 730232 41696 730244
rect 35676 730204 41696 730232
rect 35676 730192 35682 730204
rect 41690 730192 41696 730204
rect 41748 730192 41754 730244
rect 35802 730056 35808 730108
rect 35860 730096 35866 730108
rect 41506 730096 41512 730108
rect 35860 730068 41512 730096
rect 35860 730056 35866 730068
rect 41506 730056 41512 730068
rect 41564 730056 41570 730108
rect 674208 728640 674406 728668
rect 673822 728560 673828 728612
rect 673880 728600 673886 728612
rect 674208 728600 674236 728640
rect 673880 728572 674236 728600
rect 673880 728560 673886 728572
rect 673362 728424 673368 728476
rect 673420 728464 673426 728476
rect 673420 728436 674268 728464
rect 673420 728424 673426 728436
rect 674150 728136 674202 728142
rect 672994 728084 673000 728136
rect 673052 728124 673058 728136
rect 673052 728096 674058 728124
rect 673052 728084 673058 728096
rect 674150 728078 674202 728084
rect 41322 726044 41328 726096
rect 41380 726084 41386 726096
rect 41690 726084 41696 726096
rect 41380 726056 41696 726084
rect 41380 726044 41386 726056
rect 41690 726044 41696 726056
rect 41748 726044 41754 726096
rect 41322 724480 41328 724532
rect 41380 724520 41386 724532
rect 41690 724520 41696 724532
rect 41380 724492 41696 724520
rect 41380 724480 41386 724492
rect 41690 724480 41696 724492
rect 41748 724480 41754 724532
rect 677318 724208 677324 724260
rect 677376 724248 677382 724260
rect 683298 724248 683304 724260
rect 677376 724220 683304 724248
rect 677376 724208 677382 724220
rect 683298 724208 683304 724220
rect 683356 724208 683362 724260
rect 651466 723120 651472 723172
rect 651524 723160 651530 723172
rect 663058 723160 663064 723172
rect 651524 723132 663064 723160
rect 651524 723120 651530 723132
rect 663058 723120 663064 723132
rect 663116 723120 663122 723172
rect 31018 716864 31024 716916
rect 31076 716904 31082 716916
rect 41506 716904 41512 716916
rect 31076 716876 41512 716904
rect 31076 716864 31082 716876
rect 41506 716864 41512 716876
rect 41564 716864 41570 716916
rect 33778 715640 33784 715692
rect 33836 715680 33842 715692
rect 39850 715680 39856 715692
rect 33836 715652 39856 715680
rect 33836 715640 33842 715652
rect 39850 715640 39856 715652
rect 39908 715640 39914 715692
rect 33042 715504 33048 715556
rect 33100 715544 33106 715556
rect 40218 715544 40224 715556
rect 33100 715516 40224 715544
rect 33100 715504 33106 715516
rect 40218 715504 40224 715516
rect 40276 715504 40282 715556
rect 36538 715300 36544 715352
rect 36596 715340 36602 715352
rect 41690 715340 41696 715352
rect 36596 715312 41696 715340
rect 36596 715300 36602 715312
rect 41690 715300 41696 715312
rect 41748 715300 41754 715352
rect 50338 714824 50344 714876
rect 50396 714864 50402 714876
rect 62114 714864 62120 714876
rect 50396 714836 62120 714864
rect 50396 714824 50402 714836
rect 62114 714824 62120 714836
rect 62172 714824 62178 714876
rect 652570 709316 652576 709368
rect 652628 709356 652634 709368
rect 664438 709356 664444 709368
rect 652628 709328 664444 709356
rect 652628 709316 652634 709328
rect 664438 709316 664444 709328
rect 664496 709316 664502 709368
rect 672442 707208 672448 707260
rect 672500 707248 672506 707260
rect 672994 707248 673000 707260
rect 672500 707220 673000 707248
rect 672500 707208 672506 707220
rect 672994 707208 673000 707220
rect 673052 707208 673058 707260
rect 55858 701020 55864 701072
rect 55916 701060 55922 701072
rect 62114 701060 62120 701072
rect 55916 701032 62120 701060
rect 55916 701020 55922 701032
rect 62114 701020 62120 701032
rect 62172 701020 62178 701072
rect 652386 696940 652392 696992
rect 652444 696980 652450 696992
rect 661678 696980 661684 696992
rect 652444 696952 661684 696980
rect 652444 696940 652450 696952
rect 661678 696940 661684 696952
rect 661736 696940 661742 696992
rect 53098 688644 53104 688696
rect 53156 688684 53162 688696
rect 62114 688684 62120 688696
rect 53156 688656 62120 688684
rect 53156 688644 53162 688656
rect 62114 688644 62120 688656
rect 62172 688644 62178 688696
rect 35802 687216 35808 687268
rect 35860 687256 35866 687268
rect 41690 687256 41696 687268
rect 35860 687228 41696 687256
rect 35860 687216 35866 687228
rect 41690 687216 41696 687228
rect 41748 687216 41754 687268
rect 44542 685040 44548 685092
rect 44600 685080 44606 685092
rect 45370 685080 45376 685092
rect 44600 685052 45376 685080
rect 44600 685040 44606 685052
rect 45370 685040 45376 685052
rect 45428 685040 45434 685092
rect 35802 683136 35808 683188
rect 35860 683176 35866 683188
rect 41690 683176 41696 683188
rect 35860 683148 41696 683176
rect 35860 683136 35866 683148
rect 41690 683136 41696 683148
rect 41748 683136 41754 683188
rect 35618 681844 35624 681896
rect 35676 681884 35682 681896
rect 41690 681884 41696 681896
rect 35676 681856 41696 681884
rect 35676 681844 35682 681856
rect 41690 681844 41696 681856
rect 41748 681844 41754 681896
rect 35802 681708 35808 681760
rect 35860 681748 35866 681760
rect 41322 681748 41328 681760
rect 35860 681720 41328 681748
rect 35860 681708 35866 681720
rect 41322 681708 41328 681720
rect 41380 681708 41386 681760
rect 35434 681028 35440 681080
rect 35492 681068 35498 681080
rect 41598 681068 41604 681080
rect 35492 681040 41604 681068
rect 35492 681028 35498 681040
rect 41598 681028 41604 681040
rect 41656 681028 41662 681080
rect 35618 680620 35624 680672
rect 35676 680660 35682 680672
rect 36538 680660 36544 680672
rect 35676 680632 36544 680660
rect 35676 680620 35682 680632
rect 36538 680620 36544 680632
rect 36596 680620 36602 680672
rect 35802 680348 35808 680400
rect 35860 680388 35866 680400
rect 37918 680388 37924 680400
rect 35860 680360 37924 680388
rect 35860 680348 35866 680360
rect 37918 680348 37924 680360
rect 37976 680348 37982 680400
rect 51718 674840 51724 674892
rect 51776 674880 51782 674892
rect 62114 674880 62120 674892
rect 51776 674852 62120 674880
rect 51776 674840 51782 674852
rect 62114 674840 62120 674852
rect 62172 674840 62178 674892
rect 35158 672732 35164 672784
rect 35216 672772 35222 672784
rect 38930 672772 38936 672784
rect 35216 672744 38936 672772
rect 35216 672732 35222 672744
rect 38930 672732 38936 672744
rect 38988 672732 38994 672784
rect 36538 672052 36544 672104
rect 36596 672092 36602 672104
rect 39574 672092 39580 672104
rect 36596 672064 39580 672092
rect 36596 672052 36602 672064
rect 39574 672052 39580 672064
rect 39632 672052 39638 672104
rect 651466 669332 651472 669384
rect 651524 669372 651530 669384
rect 661862 669372 661868 669384
rect 651524 669344 661868 669372
rect 651524 669332 651530 669344
rect 661862 669332 661868 669344
rect 661920 669332 661926 669384
rect 671062 666204 671068 666256
rect 671120 666244 671126 666256
rect 673362 666244 673368 666256
rect 671120 666216 673368 666244
rect 671120 666204 671126 666216
rect 673362 666204 673368 666216
rect 673420 666204 673426 666256
rect 47578 662396 47584 662448
rect 47636 662436 47642 662448
rect 62114 662436 62120 662448
rect 47636 662408 62120 662436
rect 47636 662396 47642 662408
rect 62114 662396 62120 662408
rect 62172 662396 62178 662448
rect 651466 656888 651472 656940
rect 651524 656928 651530 656940
rect 670142 656928 670148 656940
rect 651524 656900 670148 656928
rect 651524 656888 651530 656900
rect 670142 656888 670148 656900
rect 670200 656888 670206 656940
rect 54478 647844 54484 647896
rect 54536 647884 54542 647896
rect 62114 647884 62120 647896
rect 54536 647856 62120 647884
rect 54536 647844 54542 647856
rect 62114 647844 62120 647856
rect 62172 647844 62178 647896
rect 651466 643084 651472 643136
rect 651524 643124 651530 643136
rect 668578 643124 668584 643136
rect 651524 643096 668584 643124
rect 651524 643084 651530 643096
rect 668578 643084 668584 643096
rect 668636 643084 668642 643136
rect 35802 639140 35808 639192
rect 35860 639180 35866 639192
rect 35860 639140 35894 639180
rect 35866 639112 35894 639140
rect 41690 639112 41696 639124
rect 35866 639084 41696 639112
rect 41690 639072 41696 639084
rect 41748 639072 41754 639124
rect 35802 638936 35808 638988
rect 35860 638976 35866 638988
rect 40034 638976 40040 638988
rect 35860 638948 40040 638976
rect 35860 638936 35866 638948
rect 40034 638936 40040 638948
rect 40092 638936 40098 638988
rect 35802 637576 35808 637628
rect 35860 637616 35866 637628
rect 41322 637616 41328 637628
rect 35860 637588 41328 637616
rect 35860 637576 35866 637588
rect 41322 637576 41328 637588
rect 41380 637576 41386 637628
rect 51718 636216 51724 636268
rect 51776 636256 51782 636268
rect 62114 636256 62120 636268
rect 51776 636228 62120 636256
rect 51776 636216 51782 636228
rect 62114 636216 62120 636228
rect 62172 636216 62178 636268
rect 44910 635944 44916 635996
rect 44968 635944 44974 635996
rect 44928 635712 44956 635944
rect 45094 635712 45100 635724
rect 44928 635684 45100 635712
rect 45094 635672 45100 635684
rect 45152 635672 45158 635724
rect 32398 629892 32404 629944
rect 32456 629932 32462 629944
rect 41690 629932 41696 629944
rect 32456 629904 41696 629932
rect 32456 629892 32462 629904
rect 41690 629892 41696 629904
rect 41748 629892 41754 629944
rect 651466 629280 651472 629332
rect 651524 629320 651530 629332
rect 667198 629320 667204 629332
rect 651524 629292 667204 629320
rect 651524 629280 651530 629292
rect 667198 629280 667204 629292
rect 667256 629280 667262 629332
rect 670970 627104 670976 627156
rect 671028 627144 671034 627156
rect 672166 627144 672172 627156
rect 671028 627116 672172 627144
rect 671028 627104 671034 627116
rect 672166 627104 672172 627116
rect 672224 627104 672230 627156
rect 672902 626696 672908 626748
rect 672960 626736 672966 626748
rect 673546 626736 673552 626748
rect 672960 626708 673552 626736
rect 672960 626696 672966 626708
rect 673546 626696 673552 626708
rect 673604 626696 673610 626748
rect 673086 626600 673092 626612
rect 672920 626572 673092 626600
rect 672920 626408 672948 626572
rect 673086 626560 673092 626572
rect 673144 626560 673150 626612
rect 675846 626560 675852 626612
rect 675904 626600 675910 626612
rect 676490 626600 676496 626612
rect 675904 626572 676496 626600
rect 675904 626560 675910 626572
rect 676490 626560 676496 626572
rect 676548 626560 676554 626612
rect 672902 626356 672908 626408
rect 672960 626356 672966 626408
rect 44082 626084 44088 626136
rect 44140 626124 44146 626136
rect 44910 626124 44916 626136
rect 44140 626096 44916 626124
rect 44140 626084 44146 626096
rect 44910 626084 44916 626096
rect 44968 626084 44974 626136
rect 48958 623772 48964 623824
rect 49016 623812 49022 623824
rect 62114 623812 62120 623824
rect 49016 623784 62120 623812
rect 49016 623772 49022 623784
rect 62114 623772 62120 623784
rect 62172 623772 62178 623824
rect 651466 616836 651472 616888
rect 651524 616876 651530 616888
rect 660298 616876 660304 616888
rect 651524 616848 660304 616876
rect 651524 616836 651530 616848
rect 660298 616836 660304 616848
rect 660356 616836 660362 616888
rect 671430 616156 671436 616208
rect 671488 616196 671494 616208
rect 671890 616196 671896 616208
rect 671488 616168 671896 616196
rect 671488 616156 671494 616168
rect 671890 616156 671896 616168
rect 671948 616156 671954 616208
rect 43530 612932 43536 612944
rect 43286 612904 43536 612932
rect 43530 612892 43536 612904
rect 43588 612892 43594 612944
rect 43371 612740 43423 612746
rect 43371 612682 43423 612688
rect 43714 612524 43720 612536
rect 43516 612496 43720 612524
rect 43714 612484 43720 612496
rect 43772 612484 43778 612536
rect 46382 612388 46388 612400
rect 43732 612360 46388 612388
rect 43582 612332 43634 612338
rect 43582 612274 43634 612280
rect 43732 612102 43760 612360
rect 46382 612348 46388 612360
rect 46440 612348 46446 612400
rect 45554 612184 45560 612196
rect 43824 612156 45560 612184
rect 43824 611898 43852 612156
rect 45554 612144 45560 612156
rect 45612 612144 45618 612196
rect 46934 611708 46940 611720
rect 43957 611680 46940 611708
rect 46934 611668 46940 611680
rect 46992 611668 46998 611720
rect 44174 611572 44180 611584
rect 44054 611544 44180 611572
rect 44054 611490 44082 611544
rect 44174 611532 44180 611544
rect 44232 611532 44238 611584
rect 45738 611300 45744 611312
rect 44181 611272 45744 611300
rect 45738 611260 45744 611272
rect 45796 611260 45802 611312
rect 47210 611096 47216 611108
rect 44298 611068 47216 611096
rect 47210 611056 47216 611068
rect 47268 611056 47274 611108
rect 45370 610892 45376 610904
rect 44405 610864 45376 610892
rect 45370 610852 45376 610864
rect 45428 610852 45434 610904
rect 44502 610632 44554 610638
rect 44502 610574 44554 610580
rect 56042 608608 56048 608660
rect 56100 608648 56106 608660
rect 62114 608648 62120 608660
rect 56100 608620 62120 608648
rect 56100 608608 56106 608620
rect 62114 608608 62120 608620
rect 62172 608608 62178 608660
rect 651466 603100 651472 603152
rect 651524 603140 651530 603152
rect 664622 603140 664628 603152
rect 651524 603112 664628 603140
rect 651524 603100 651530 603112
rect 664622 603100 664628 603112
rect 664680 603100 664686 603152
rect 48958 597524 48964 597576
rect 49016 597564 49022 597576
rect 62114 597564 62120 597576
rect 49016 597536 62120 597564
rect 49016 597524 49022 597536
rect 62114 597524 62120 597536
rect 62172 597524 62178 597576
rect 40310 596164 40316 596216
rect 40368 596204 40374 596216
rect 41690 596204 41696 596216
rect 40368 596176 41696 596204
rect 40368 596164 40374 596176
rect 41690 596164 41696 596176
rect 41748 596164 41754 596216
rect 40862 596028 40868 596080
rect 40920 596068 40926 596080
rect 41322 596068 41328 596080
rect 40920 596040 41328 596068
rect 40920 596028 40926 596040
rect 41322 596028 41328 596040
rect 41380 596028 41386 596080
rect 40678 593240 40684 593292
rect 40736 593280 40742 593292
rect 41598 593280 41604 593292
rect 40736 593252 41604 593280
rect 40736 593240 40742 593252
rect 41598 593240 41604 593252
rect 41656 593240 41662 593292
rect 40954 593036 40960 593088
rect 41012 593076 41018 593088
rect 41598 593076 41604 593088
rect 41012 593048 41604 593076
rect 41012 593036 41018 593048
rect 41598 593036 41604 593048
rect 41656 593036 41662 593088
rect 675938 591336 675944 591388
rect 675996 591376 676002 591388
rect 679618 591376 679624 591388
rect 675996 591348 679624 591376
rect 675996 591336 676002 591348
rect 679618 591336 679624 591348
rect 679676 591336 679682 591388
rect 676122 591200 676128 591252
rect 676180 591240 676186 591252
rect 682378 591240 682384 591252
rect 676180 591212 682384 591240
rect 676180 591200 676186 591212
rect 682378 591200 682384 591212
rect 682436 591200 682442 591252
rect 651466 590656 651472 590708
rect 651524 590696 651530 590708
rect 662046 590696 662052 590708
rect 651524 590668 662052 590696
rect 651524 590656 651530 590668
rect 662046 590656 662052 590668
rect 662104 590656 662110 590708
rect 35158 585896 35164 585948
rect 35216 585936 35222 585948
rect 40494 585936 40500 585948
rect 35216 585908 40500 585936
rect 35216 585896 35222 585908
rect 40494 585896 40500 585908
rect 40552 585896 40558 585948
rect 32398 585760 32404 585812
rect 32456 585800 32462 585812
rect 39482 585800 39488 585812
rect 32456 585772 39488 585800
rect 32456 585760 32462 585772
rect 39482 585760 39488 585772
rect 39540 585760 39546 585812
rect 36538 585148 36544 585200
rect 36596 585188 36602 585200
rect 41414 585188 41420 585200
rect 36596 585160 41420 585188
rect 36596 585148 36602 585160
rect 41414 585148 41420 585160
rect 41472 585148 41478 585200
rect 51718 583720 51724 583772
rect 51776 583760 51782 583772
rect 62114 583760 62120 583772
rect 51776 583732 62120 583760
rect 51776 583720 51782 583732
rect 62114 583720 62120 583732
rect 62172 583720 62178 583772
rect 672350 579504 672356 579556
rect 672408 579544 672414 579556
rect 672994 579544 673000 579556
rect 672408 579516 673000 579544
rect 672408 579504 672414 579516
rect 672994 579504 673000 579516
rect 673052 579504 673058 579556
rect 651466 576852 651472 576904
rect 651524 576892 651530 576904
rect 665818 576892 665824 576904
rect 651524 576864 665824 576892
rect 651524 576852 651530 576864
rect 665818 576852 665824 576864
rect 665876 576852 665882 576904
rect 672442 572704 672448 572756
rect 672500 572744 672506 572756
rect 672902 572744 672908 572756
rect 672500 572716 672908 572744
rect 672500 572704 672506 572716
rect 672902 572704 672908 572716
rect 672960 572704 672966 572756
rect 679618 571276 679624 571328
rect 679676 571316 679682 571328
rect 683114 571316 683120 571328
rect 679676 571288 683120 571316
rect 679676 571276 679682 571288
rect 683114 571276 683120 571288
rect 683172 571276 683178 571328
rect 672258 567264 672264 567316
rect 672316 567304 672322 567316
rect 672902 567304 672908 567316
rect 672316 567276 672908 567304
rect 672316 567264 672322 567276
rect 672902 567264 672908 567276
rect 672960 567264 672966 567316
rect 651650 563048 651656 563100
rect 651708 563088 651714 563100
rect 658918 563088 658924 563100
rect 651708 563060 658924 563088
rect 651708 563048 651714 563060
rect 658918 563048 658924 563060
rect 658976 563048 658982 563100
rect 55858 558084 55864 558136
rect 55916 558124 55922 558136
rect 62114 558124 62120 558136
rect 55916 558096 62120 558124
rect 55916 558084 55922 558096
rect 62114 558084 62120 558096
rect 62172 558084 62178 558136
rect 35802 557540 35808 557592
rect 35860 557580 35866 557592
rect 41506 557580 41512 557592
rect 35860 557552 41512 557580
rect 35860 557540 35866 557552
rect 41506 557540 41512 557552
rect 41564 557540 41570 557592
rect 35802 554752 35808 554804
rect 35860 554792 35866 554804
rect 41690 554792 41696 554804
rect 35860 554764 41696 554792
rect 35860 554752 35866 554764
rect 41690 554752 41696 554764
rect 41748 554752 41754 554804
rect 35802 553528 35808 553580
rect 35860 553568 35866 553580
rect 41414 553568 41420 553580
rect 35860 553540 41420 553568
rect 35860 553528 35866 553540
rect 41414 553528 41420 553540
rect 41472 553528 41478 553580
rect 35618 553392 35624 553444
rect 35676 553432 35682 553444
rect 41690 553432 41696 553444
rect 35676 553404 41696 553432
rect 35676 553392 35682 553404
rect 41690 553392 41696 553404
rect 41748 553392 41754 553444
rect 41046 552100 41052 552152
rect 41104 552140 41110 552152
rect 41104 552112 41414 552140
rect 41104 552100 41110 552112
rect 41386 552072 41414 552112
rect 41690 552072 41696 552084
rect 41386 552044 41696 552072
rect 41690 552032 41696 552044
rect 41748 552032 41754 552084
rect 41230 550604 41236 550656
rect 41288 550644 41294 550656
rect 41690 550644 41696 550656
rect 41288 550616 41696 550644
rect 41288 550604 41294 550616
rect 41690 550604 41696 550616
rect 41748 550604 41754 550656
rect 651466 550604 651472 550656
rect 651524 550644 651530 550656
rect 660298 550644 660304 550656
rect 651524 550616 660304 550644
rect 651524 550604 651530 550616
rect 660298 550604 660304 550616
rect 660356 550604 660362 550656
rect 41322 547884 41328 547936
rect 41380 547924 41386 547936
rect 41690 547924 41696 547936
rect 41380 547896 41696 547924
rect 41380 547884 41386 547896
rect 41690 547884 41696 547896
rect 41748 547884 41754 547936
rect 675846 547612 675852 547664
rect 675904 547652 675910 547664
rect 678238 547652 678244 547664
rect 675904 547624 678244 547652
rect 675904 547612 675910 547624
rect 678238 547612 678244 547624
rect 678296 547612 678302 547664
rect 31754 547408 31760 547460
rect 31812 547448 31818 547460
rect 37090 547448 37096 547460
rect 31812 547420 37096 547448
rect 31812 547408 31818 547420
rect 37090 547408 37096 547420
rect 37148 547408 37154 547460
rect 47578 545096 47584 545148
rect 47636 545136 47642 545148
rect 62114 545136 62120 545148
rect 47636 545108 62120 545136
rect 47636 545096 47642 545108
rect 62114 545096 62120 545108
rect 62172 545096 62178 545148
rect 33778 542988 33784 543040
rect 33836 543028 33842 543040
rect 41506 543028 41512 543040
rect 33836 543000 41512 543028
rect 33836 542988 33842 543000
rect 41506 542988 41512 543000
rect 41564 542988 41570 543040
rect 37090 542308 37096 542360
rect 37148 542348 37154 542360
rect 41690 542348 41696 542360
rect 37148 542320 41696 542348
rect 37148 542308 37154 542320
rect 41690 542308 41696 542320
rect 41748 542308 41754 542360
rect 651466 536800 651472 536852
rect 651524 536840 651530 536852
rect 669958 536840 669964 536852
rect 651524 536812 669964 536840
rect 651524 536800 651530 536812
rect 669958 536800 669964 536812
rect 670016 536800 670022 536852
rect 671246 533168 671252 533180
rect 670896 533140 671252 533168
rect 670896 532908 670924 533140
rect 671246 533128 671252 533140
rect 671304 533128 671310 533180
rect 670878 532856 670884 532908
rect 670936 532856 670942 532908
rect 50338 532720 50344 532772
rect 50396 532760 50402 532772
rect 62114 532760 62120 532772
rect 50396 532732 62120 532760
rect 50396 532720 50402 532732
rect 62114 532720 62120 532732
rect 62172 532720 62178 532772
rect 675846 532244 675852 532296
rect 675904 532284 675910 532296
rect 676582 532284 676588 532296
rect 675904 532256 676588 532284
rect 675904 532244 675910 532256
rect 676582 532244 676588 532256
rect 676640 532244 676646 532296
rect 651834 522996 651840 523048
rect 651892 523036 651898 523048
rect 661862 523036 661868 523048
rect 651892 523008 661868 523036
rect 651892 522996 651898 523008
rect 661862 522996 661868 523008
rect 661920 522996 661926 523048
rect 54478 518916 54484 518968
rect 54536 518956 54542 518968
rect 62114 518956 62120 518968
rect 54536 518928 62120 518956
rect 54536 518916 54542 518928
rect 62114 518916 62120 518928
rect 62172 518916 62178 518968
rect 675846 518780 675852 518832
rect 675904 518820 675910 518832
rect 677870 518820 677876 518832
rect 675904 518792 677876 518820
rect 675904 518780 675910 518792
rect 677870 518780 677876 518792
rect 677928 518780 677934 518832
rect 651466 510620 651472 510672
rect 651524 510660 651530 510672
rect 659102 510660 659108 510672
rect 651524 510632 659108 510660
rect 651524 510620 651530 510632
rect 659102 510620 659108 510632
rect 659160 510620 659166 510672
rect 46198 506472 46204 506524
rect 46256 506512 46262 506524
rect 62114 506512 62120 506524
rect 46256 506484 62120 506512
rect 46256 506472 46262 506484
rect 62114 506472 62120 506484
rect 62172 506472 62178 506524
rect 675846 503616 675852 503668
rect 675904 503656 675910 503668
rect 679618 503656 679624 503668
rect 675904 503628 679624 503656
rect 675904 503616 675910 503628
rect 679618 503616 679624 503628
rect 679676 503616 679682 503668
rect 676030 503480 676036 503532
rect 676088 503520 676094 503532
rect 682378 503520 682384 503532
rect 676088 503492 682384 503520
rect 676088 503480 676094 503492
rect 682378 503480 682384 503492
rect 682436 503480 682442 503532
rect 675846 502324 675852 502376
rect 675904 502364 675910 502376
rect 676858 502364 676864 502376
rect 675904 502336 676864 502364
rect 675904 502324 675910 502336
rect 676858 502324 676864 502336
rect 676916 502324 676922 502376
rect 676030 500896 676036 500948
rect 676088 500936 676094 500948
rect 680998 500936 681004 500948
rect 676088 500908 681004 500936
rect 676088 500896 676094 500908
rect 680998 500896 681004 500908
rect 681056 500896 681062 500948
rect 651466 496816 651472 496868
rect 651524 496856 651530 496868
rect 663242 496856 663248 496868
rect 651524 496828 663248 496856
rect 651524 496816 651530 496828
rect 663242 496816 663248 496828
rect 663300 496816 663306 496868
rect 676030 492668 676036 492720
rect 676088 492708 676094 492720
rect 683390 492708 683396 492720
rect 676088 492680 683396 492708
rect 676088 492668 676094 492680
rect 683390 492668 683396 492680
rect 683448 492668 683454 492720
rect 48958 491920 48964 491972
rect 49016 491960 49022 491972
rect 62114 491960 62120 491972
rect 49016 491932 62120 491960
rect 49016 491920 49022 491932
rect 62114 491920 62120 491932
rect 62172 491920 62178 491972
rect 651466 484440 651472 484492
rect 651524 484480 651530 484492
rect 651524 484452 654134 484480
rect 651524 484440 651530 484452
rect 654106 484412 654134 484452
rect 667198 484412 667204 484424
rect 654106 484384 667204 484412
rect 667198 484372 667204 484384
rect 667256 484372 667262 484424
rect 51718 480224 51724 480276
rect 51776 480264 51782 480276
rect 62114 480264 62120 480276
rect 51776 480236 62120 480264
rect 51776 480224 51782 480236
rect 62114 480224 62120 480236
rect 62172 480224 62178 480276
rect 651466 470568 651472 470620
rect 651524 470608 651530 470620
rect 665818 470608 665824 470620
rect 651524 470580 665824 470608
rect 651524 470568 651530 470580
rect 665818 470568 665824 470580
rect 665876 470568 665882 470620
rect 51902 466420 51908 466472
rect 51960 466460 51966 466472
rect 62114 466460 62120 466472
rect 51960 466432 62120 466460
rect 51960 466420 51966 466432
rect 62114 466420 62120 466432
rect 62172 466420 62178 466472
rect 652386 456764 652392 456816
rect 652444 456804 652450 456816
rect 661678 456804 661684 456816
rect 652444 456776 661684 456804
rect 652444 456764 652450 456776
rect 661678 456764 661684 456776
rect 661736 456764 661742 456816
rect 673942 456424 673948 456476
rect 674000 456424 674006 456476
rect 673960 456246 673988 456424
rect 673828 456068 673880 456074
rect 673828 456010 673880 456016
rect 673454 455812 673460 455864
rect 673512 455852 673518 455864
rect 673512 455824 673762 455852
rect 673512 455812 673518 455824
rect 673598 455660 673650 455666
rect 673598 455602 673650 455608
rect 673506 455388 673558 455394
rect 673506 455330 673558 455336
rect 673388 455184 673440 455190
rect 673388 455126 673440 455132
rect 671062 454996 671068 455048
rect 671120 455036 671126 455048
rect 671120 455008 673302 455036
rect 671120 454996 671126 455008
rect 673164 454844 673216 454850
rect 673164 454786 673216 454792
rect 673046 454640 673098 454646
rect 673046 454582 673098 454588
rect 672954 454368 673006 454374
rect 672954 454310 673006 454316
rect 672816 454096 672868 454102
rect 53098 454044 53104 454096
rect 53156 454084 53162 454096
rect 62114 454084 62120 454096
rect 53156 454056 62120 454084
rect 53156 454044 53162 454056
rect 62114 454044 62120 454056
rect 62172 454044 62178 454096
rect 672816 454038 672868 454044
rect 672258 453908 672264 453960
rect 672316 453948 672322 453960
rect 672316 453920 672750 453948
rect 672316 453908 672322 453920
rect 651466 444456 651472 444508
rect 651524 444496 651530 444508
rect 651524 444468 654134 444496
rect 651524 444456 651530 444468
rect 654106 444428 654134 444468
rect 668578 444428 668584 444440
rect 654106 444400 668584 444428
rect 668578 444388 668584 444400
rect 668636 444388 668642 444440
rect 50522 440240 50528 440292
rect 50580 440280 50586 440292
rect 62114 440280 62120 440292
rect 50580 440252 62120 440280
rect 50580 440240 50586 440252
rect 62114 440240 62120 440252
rect 62172 440240 62178 440292
rect 651466 430584 651472 430636
rect 651524 430624 651530 430636
rect 671338 430624 671344 430636
rect 651524 430596 671344 430624
rect 651524 430584 651530 430596
rect 671338 430584 671344 430596
rect 671396 430584 671402 430636
rect 54478 427796 54484 427848
rect 54536 427836 54542 427848
rect 62114 427836 62120 427848
rect 54536 427808 62120 427836
rect 54536 427796 54542 427808
rect 62114 427796 62120 427808
rect 62172 427796 62178 427848
rect 41322 423648 41328 423700
rect 41380 423688 41386 423700
rect 41690 423688 41696 423700
rect 41380 423660 41696 423688
rect 41380 423648 41386 423660
rect 41690 423648 41696 423660
rect 41748 423648 41754 423700
rect 651834 416780 651840 416832
rect 651892 416820 651898 416832
rect 663058 416820 663064 416832
rect 651892 416792 663064 416820
rect 651892 416780 651898 416792
rect 663058 416780 663064 416792
rect 663116 416780 663122 416832
rect 47578 415420 47584 415472
rect 47636 415460 47642 415472
rect 62114 415460 62120 415472
rect 47636 415432 62120 415460
rect 47636 415420 47642 415432
rect 62114 415420 62120 415432
rect 62172 415420 62178 415472
rect 36538 415352 36544 415404
rect 36596 415392 36602 415404
rect 41690 415392 41696 415404
rect 36596 415364 41696 415392
rect 36596 415352 36602 415364
rect 41690 415352 41696 415364
rect 41748 415352 41754 415404
rect 651466 404336 651472 404388
rect 651524 404376 651530 404388
rect 664438 404376 664444 404388
rect 651524 404348 664444 404376
rect 651524 404336 651530 404348
rect 664438 404336 664444 404348
rect 664496 404336 664502 404388
rect 55858 401616 55864 401668
rect 55916 401656 55922 401668
rect 62114 401656 62120 401668
rect 55916 401628 62120 401656
rect 55916 401616 55922 401628
rect 62114 401616 62120 401628
rect 62172 401616 62178 401668
rect 675846 395700 675852 395752
rect 675904 395740 675910 395752
rect 676398 395740 676404 395752
rect 675904 395712 676404 395740
rect 675904 395700 675910 395712
rect 676398 395700 676404 395712
rect 676456 395700 676462 395752
rect 652570 390532 652576 390584
rect 652628 390572 652634 390584
rect 658918 390572 658924 390584
rect 652628 390544 658924 390572
rect 652628 390532 652634 390544
rect 658918 390532 658924 390544
rect 658976 390532 658982 390584
rect 47762 389240 47768 389292
rect 47820 389280 47826 389292
rect 62114 389280 62120 389292
rect 47820 389252 62120 389280
rect 47820 389240 47826 389252
rect 62114 389240 62120 389252
rect 62172 389240 62178 389292
rect 41138 387064 41144 387116
rect 41196 387104 41202 387116
rect 41690 387104 41696 387116
rect 41196 387076 41696 387104
rect 41196 387064 41202 387076
rect 41690 387064 41696 387076
rect 41748 387064 41754 387116
rect 41322 382372 41328 382424
rect 41380 382412 41386 382424
rect 41506 382412 41512 382424
rect 41380 382384 41512 382412
rect 41380 382372 41386 382384
rect 41506 382372 41512 382384
rect 41564 382372 41570 382424
rect 35802 379516 35808 379568
rect 35860 379556 35866 379568
rect 41690 379556 41696 379568
rect 35860 379528 41696 379556
rect 35860 379516 35866 379528
rect 41690 379516 41696 379528
rect 41748 379516 41754 379568
rect 40218 378496 40224 378548
rect 40276 378536 40282 378548
rect 41690 378536 41696 378548
rect 40276 378508 41696 378536
rect 40276 378496 40282 378508
rect 41690 378496 41696 378508
rect 41748 378496 41754 378548
rect 35802 375368 35808 375420
rect 35860 375408 35866 375420
rect 41690 375408 41696 375420
rect 35860 375380 41696 375408
rect 35860 375368 35866 375380
rect 41690 375368 41696 375380
rect 41748 375368 41754 375420
rect 51718 375368 51724 375420
rect 51776 375408 51782 375420
rect 62114 375408 62120 375420
rect 51776 375380 62120 375408
rect 51776 375368 51782 375380
rect 62114 375368 62120 375380
rect 62172 375368 62178 375420
rect 37918 372580 37924 372632
rect 37976 372620 37982 372632
rect 41690 372620 41696 372632
rect 37976 372592 41696 372620
rect 37976 372580 37982 372592
rect 41690 372580 41696 372592
rect 41748 372580 41754 372632
rect 651650 364352 651656 364404
rect 651708 364392 651714 364404
rect 661862 364392 661868 364404
rect 651708 364364 661868 364392
rect 651708 364352 651714 364364
rect 661862 364352 661868 364364
rect 661920 364352 661926 364404
rect 46382 362924 46388 362976
rect 46440 362964 46446 362976
rect 62114 362964 62120 362976
rect 46440 362936 62120 362964
rect 46440 362924 46446 362936
rect 62114 362924 62120 362936
rect 62172 362924 62178 362976
rect 45002 355784 45008 355836
rect 45060 355824 45066 355836
rect 45646 355824 45652 355836
rect 45060 355796 45652 355824
rect 45060 355784 45066 355796
rect 45646 355784 45652 355796
rect 45704 355784 45710 355836
rect 44634 355648 44640 355700
rect 44692 355688 44698 355700
rect 44692 355660 45048 355688
rect 44692 355648 44698 355660
rect 44569 354832 44575 354884
rect 44627 354872 44633 354884
rect 44627 354844 44839 354872
rect 44627 354832 44633 354844
rect 44575 354680 44627 354686
rect 44575 354622 44627 354628
rect 44811 354600 44839 354844
rect 45020 354600 45048 355660
rect 44811 354572 44956 354600
rect 45020 354572 45063 354600
rect 44793 354424 44799 354476
rect 44851 354424 44857 354476
rect 44686 354340 44738 354346
rect 44811 354314 44839 354424
rect 44686 354282 44738 354288
rect 44928 354110 44956 354572
rect 45035 353906 45063 354572
rect 45646 354056 45652 354068
rect 45158 354028 45652 354056
rect 45158 353702 45186 354028
rect 45646 354016 45652 354028
rect 45704 354016 45710 354068
rect 45922 353784 45928 353796
rect 45250 353756 45928 353784
rect 45250 353498 45278 353756
rect 45922 353744 45928 353756
rect 45980 353744 45986 353796
rect 45554 353240 45560 353252
rect 45385 353212 45560 353240
rect 45554 353200 45560 353212
rect 45612 353200 45618 353252
rect 651466 350548 651472 350600
rect 651524 350588 651530 350600
rect 667382 350588 667388 350600
rect 651524 350560 667388 350588
rect 651524 350548 651530 350560
rect 667382 350548 667388 350560
rect 667440 350548 667446 350600
rect 28902 345040 28908 345092
rect 28960 345080 28966 345092
rect 40218 345080 40224 345092
rect 28960 345052 40224 345080
rect 28960 345040 28966 345052
rect 40218 345040 40224 345052
rect 40276 345040 40282 345092
rect 35802 339464 35808 339516
rect 35860 339504 35866 339516
rect 37918 339504 37924 339516
rect 35860 339476 37924 339504
rect 35860 339464 35866 339476
rect 37918 339464 37924 339476
rect 37976 339464 37982 339516
rect 35802 338104 35808 338156
rect 35860 338144 35866 338156
rect 36538 338144 36544 338156
rect 35860 338116 36544 338144
rect 35860 338104 35866 338116
rect 36538 338104 36544 338116
rect 36596 338104 36602 338156
rect 651466 338104 651472 338156
rect 651524 338144 651530 338156
rect 667566 338144 667572 338156
rect 651524 338116 667572 338144
rect 651524 338104 651530 338116
rect 667566 338104 667572 338116
rect 667624 338104 667630 338156
rect 46198 336744 46204 336796
rect 46256 336784 46262 336796
rect 62114 336784 62120 336796
rect 46256 336756 62120 336784
rect 46256 336744 46262 336756
rect 62114 336744 62120 336756
rect 62172 336744 62178 336796
rect 651466 324300 651472 324352
rect 651524 324340 651530 324352
rect 667014 324340 667020 324352
rect 651524 324312 667020 324340
rect 651524 324300 651530 324312
rect 667014 324300 667020 324312
rect 667072 324300 667078 324352
rect 53282 322940 53288 322992
rect 53340 322980 53346 322992
rect 62114 322980 62120 322992
rect 53340 322952 62120 322980
rect 53340 322940 53346 322952
rect 62114 322940 62120 322952
rect 62172 322940 62178 322992
rect 54478 310496 54484 310548
rect 54536 310536 54542 310548
rect 62114 310536 62120 310548
rect 54536 310508 62120 310536
rect 54536 310496 54542 310508
rect 62114 310496 62120 310508
rect 62172 310496 62178 310548
rect 651466 310496 651472 310548
rect 651524 310536 651530 310548
rect 667198 310536 667204 310548
rect 651524 310508 667204 310536
rect 651524 310496 651530 310508
rect 667198 310496 667204 310508
rect 667256 310496 667262 310548
rect 45462 298120 45468 298172
rect 45520 298160 45526 298172
rect 62114 298160 62120 298172
rect 45520 298132 62120 298160
rect 45520 298120 45526 298132
rect 62114 298120 62120 298132
rect 62172 298120 62178 298172
rect 675846 298052 675852 298104
rect 675904 298092 675910 298104
rect 678974 298092 678980 298104
rect 675904 298064 678980 298092
rect 675904 298052 675910 298064
rect 678974 298052 678980 298064
rect 679032 298052 679038 298104
rect 676122 297848 676128 297900
rect 676180 297888 676186 297900
rect 680998 297888 681004 297900
rect 676180 297860 681004 297888
rect 676180 297848 676186 297860
rect 680998 297848 681004 297860
rect 681056 297848 681062 297900
rect 41322 285064 41328 285116
rect 41380 285104 41386 285116
rect 41690 285104 41696 285116
rect 41380 285076 41696 285104
rect 41380 285064 41386 285076
rect 41690 285064 41696 285076
rect 41748 285064 41754 285116
rect 32398 284928 32404 284980
rect 32456 284968 32462 284980
rect 41690 284968 41696 284980
rect 32456 284940 41696 284968
rect 32456 284928 32462 284940
rect 41690 284928 41696 284940
rect 41748 284928 41754 284980
rect 651466 284316 651472 284368
rect 651524 284356 651530 284368
rect 667750 284356 667756 284368
rect 651524 284328 667756 284356
rect 651524 284316 651530 284328
rect 667750 284316 667756 284328
rect 667808 284316 667814 284368
rect 522390 276360 522396 276412
rect 522448 276400 522454 276412
rect 526898 276400 526904 276412
rect 522448 276372 526904 276400
rect 522448 276360 522454 276372
rect 526898 276360 526904 276372
rect 526956 276360 526962 276412
rect 522206 276224 522212 276276
rect 522264 276264 522270 276276
rect 530486 276264 530492 276276
rect 522264 276236 530492 276264
rect 522264 276224 522270 276236
rect 530486 276224 530492 276236
rect 530544 276224 530550 276276
rect 524874 276128 524880 276140
rect 524156 276100 524880 276128
rect 524156 276060 524184 276100
rect 524874 276088 524880 276100
rect 524932 276088 524938 276140
rect 524064 276032 524184 276060
rect 88334 275952 88340 276004
rect 88392 275992 88398 276004
rect 143350 275992 143356 276004
rect 88392 275964 143356 275992
rect 88392 275952 88398 275964
rect 143350 275952 143356 275964
rect 143408 275952 143414 276004
rect 156874 275952 156880 276004
rect 156932 275992 156938 276004
rect 193858 275992 193864 276004
rect 156932 275964 193864 275992
rect 156932 275952 156938 275964
rect 193858 275952 193864 275964
rect 193916 275952 193922 276004
rect 201770 275952 201776 276004
rect 201828 275992 201834 276004
rect 222102 275992 222108 276004
rect 201828 275964 222108 275992
rect 201828 275952 201834 275964
rect 222102 275952 222108 275964
rect 222160 275952 222166 276004
rect 389174 275952 389180 276004
rect 389232 275992 389238 276004
rect 393314 275992 393320 276004
rect 389232 275964 393320 275992
rect 389232 275952 389238 275964
rect 393314 275952 393320 275964
rect 393372 275952 393378 276004
rect 400582 275952 400588 276004
rect 400640 275992 400646 276004
rect 415762 275992 415768 276004
rect 400640 275964 415768 275992
rect 400640 275952 400646 275964
rect 415762 275952 415768 275964
rect 415820 275952 415826 276004
rect 427814 275952 427820 276004
rect 427872 275992 427878 276004
rect 442994 275992 443000 276004
rect 427872 275964 443000 275992
rect 427872 275952 427878 275964
rect 442994 275952 443000 275964
rect 443052 275952 443058 276004
rect 443730 275952 443736 276004
rect 443788 275992 443794 276004
rect 453574 275992 453580 276004
rect 443788 275964 453580 275992
rect 443788 275952 443794 275964
rect 453574 275952 453580 275964
rect 453632 275952 453638 276004
rect 456978 275952 456984 276004
rect 457036 275992 457042 276004
rect 486694 275992 486700 276004
rect 457036 275964 486700 275992
rect 457036 275952 457042 275964
rect 486694 275952 486700 275964
rect 486752 275952 486758 276004
rect 486878 275952 486884 276004
rect 486936 275992 486942 276004
rect 495158 275992 495164 276004
rect 486936 275964 495164 275992
rect 486936 275952 486942 275964
rect 495158 275952 495164 275964
rect 495216 275952 495222 276004
rect 495434 275952 495440 276004
rect 495492 275992 495498 276004
rect 504542 275992 504548 276004
rect 495492 275964 504548 275992
rect 495492 275952 495498 275964
rect 504542 275952 504548 275964
rect 504600 275952 504606 276004
rect 504910 275952 504916 276004
rect 504968 275992 504974 276004
rect 507026 275992 507032 276004
rect 504968 275964 507032 275992
rect 504968 275952 504974 275964
rect 507026 275952 507032 275964
rect 507084 275952 507090 276004
rect 508038 275952 508044 276004
rect 508096 275992 508102 276004
rect 514018 275992 514024 276004
rect 508096 275964 514024 275992
rect 508096 275952 508102 275964
rect 514018 275952 514024 275964
rect 514076 275952 514082 276004
rect 519814 275992 519820 276004
rect 514220 275964 519820 275992
rect 95418 275816 95424 275868
rect 95476 275856 95482 275868
rect 104802 275856 104808 275868
rect 95476 275828 104808 275856
rect 95476 275816 95482 275828
rect 104802 275816 104808 275828
rect 104860 275816 104866 275868
rect 113174 275816 113180 275868
rect 113232 275856 113238 275868
rect 169938 275856 169944 275868
rect 113232 275828 169944 275856
rect 113232 275816 113238 275828
rect 169938 275816 169944 275828
rect 169996 275816 170002 275868
rect 181714 275816 181720 275868
rect 181772 275856 181778 275868
rect 218882 275856 218888 275868
rect 181772 275828 218888 275856
rect 181772 275816 181778 275828
rect 218882 275816 218888 275828
rect 218940 275816 218946 275868
rect 393590 275816 393596 275868
rect 393648 275856 393654 275868
rect 412266 275856 412272 275868
rect 393648 275828 412272 275856
rect 393648 275816 393654 275828
rect 412266 275816 412272 275828
rect 412324 275816 412330 275868
rect 415302 275816 415308 275868
rect 415360 275856 415366 275868
rect 425238 275856 425244 275868
rect 415360 275828 425244 275856
rect 415360 275816 415366 275828
rect 425238 275816 425244 275828
rect 425296 275816 425302 275868
rect 432966 275816 432972 275868
rect 433024 275856 433030 275868
rect 487890 275856 487896 275868
rect 433024 275828 487896 275856
rect 433024 275816 433030 275828
rect 487890 275816 487896 275828
rect 487948 275816 487954 275868
rect 488902 275816 488908 275868
rect 488960 275856 488966 275868
rect 492582 275856 492588 275868
rect 488960 275828 492588 275856
rect 488960 275816 488966 275828
rect 492582 275816 492588 275828
rect 492640 275816 492646 275868
rect 498194 275816 498200 275868
rect 498252 275856 498258 275868
rect 505646 275856 505652 275868
rect 498252 275828 505652 275856
rect 498252 275816 498258 275828
rect 505646 275816 505652 275828
rect 505704 275816 505710 275868
rect 507210 275816 507216 275868
rect 507268 275856 507274 275868
rect 512730 275856 512736 275868
rect 507268 275828 512736 275856
rect 507268 275816 507274 275828
rect 512730 275816 512736 275828
rect 512788 275816 512794 275868
rect 512914 275816 512920 275868
rect 512972 275856 512978 275868
rect 514220 275856 514248 275964
rect 519814 275952 519820 275964
rect 519872 275952 519878 276004
rect 519998 275952 520004 276004
rect 520056 275992 520062 276004
rect 524064 275992 524092 276032
rect 604914 275992 604920 276004
rect 520056 275964 524092 275992
rect 524248 275964 604920 275992
rect 520056 275952 520062 275964
rect 512972 275828 514248 275856
rect 512972 275816 512978 275828
rect 515490 275816 515496 275868
rect 515548 275856 515554 275868
rect 515548 275828 516456 275856
rect 515548 275816 515554 275828
rect 81250 275680 81256 275732
rect 81308 275720 81314 275732
rect 88978 275720 88984 275732
rect 81308 275692 88984 275720
rect 81308 275680 81314 275692
rect 88978 275680 88984 275692
rect 89036 275680 89042 275732
rect 103698 275680 103704 275732
rect 103756 275720 103762 275732
rect 160094 275720 160100 275732
rect 103756 275692 160100 275720
rect 103756 275680 103762 275692
rect 160094 275680 160100 275692
rect 160152 275680 160158 275732
rect 178126 275680 178132 275732
rect 178184 275720 178190 275732
rect 216858 275720 216864 275732
rect 178184 275692 216864 275720
rect 178184 275680 178190 275692
rect 216858 275680 216864 275692
rect 216916 275680 216922 275732
rect 299934 275680 299940 275732
rect 299992 275720 299998 275732
rect 300762 275720 300768 275732
rect 299992 275692 300768 275720
rect 299992 275680 299998 275692
rect 300762 275680 300768 275692
rect 300820 275680 300826 275732
rect 370498 275680 370504 275732
rect 370556 275720 370562 275732
rect 388622 275720 388628 275732
rect 370556 275692 388628 275720
rect 370556 275680 370562 275692
rect 388622 275680 388628 275692
rect 388680 275680 388686 275732
rect 410058 275680 410064 275732
rect 410116 275720 410122 275732
rect 428826 275720 428832 275732
rect 410116 275692 428832 275720
rect 410116 275680 410122 275692
rect 428826 275680 428832 275692
rect 428884 275680 428890 275732
rect 429194 275680 429200 275732
rect 429252 275720 429258 275732
rect 446490 275720 446496 275732
rect 429252 275692 446496 275720
rect 429252 275680 429258 275692
rect 446490 275680 446496 275692
rect 446548 275680 446554 275732
rect 446766 275680 446772 275732
rect 446824 275720 446830 275732
rect 502058 275720 502064 275732
rect 446824 275692 502064 275720
rect 446824 275680 446830 275692
rect 502058 275680 502064 275692
rect 502116 275680 502122 275732
rect 509142 275720 509148 275732
rect 504284 275692 509148 275720
rect 76466 275544 76472 275596
rect 76524 275584 76530 275596
rect 86862 275584 86868 275596
rect 76524 275556 86868 275584
rect 76524 275544 76530 275556
rect 86862 275544 86868 275556
rect 86920 275544 86926 275596
rect 96614 275544 96620 275596
rect 96672 275584 96678 275596
rect 156598 275584 156604 275596
rect 96672 275556 156604 275584
rect 96672 275544 96678 275556
rect 156598 275544 156604 275556
rect 156656 275544 156662 275596
rect 163958 275544 163964 275596
rect 164016 275584 164022 275596
rect 202138 275584 202144 275596
rect 164016 275556 202144 275584
rect 164016 275544 164022 275556
rect 202138 275544 202144 275556
rect 202196 275544 202202 275596
rect 221918 275544 221924 275596
rect 221976 275584 221982 275596
rect 233878 275584 233884 275596
rect 221976 275556 233884 275584
rect 221976 275544 221982 275556
rect 233878 275544 233884 275556
rect 233936 275544 233942 275596
rect 236086 275544 236092 275596
rect 236144 275584 236150 275596
rect 251082 275584 251088 275596
rect 236144 275556 251088 275584
rect 236144 275544 236150 275556
rect 251082 275544 251088 275556
rect 251140 275544 251146 275596
rect 350718 275544 350724 275596
rect 350776 275584 350782 275596
rect 361390 275584 361396 275596
rect 350776 275556 361396 275584
rect 350776 275544 350782 275556
rect 361390 275544 361396 275556
rect 361448 275544 361454 275596
rect 362218 275544 362224 275596
rect 362276 275584 362282 275596
rect 385034 275584 385040 275596
rect 362276 275556 385040 275584
rect 362276 275544 362282 275556
rect 385034 275544 385040 275556
rect 385092 275544 385098 275596
rect 388162 275544 388168 275596
rect 388220 275584 388226 275596
rect 418154 275584 418160 275596
rect 388220 275556 418160 275584
rect 388220 275544 388226 275556
rect 418154 275544 418160 275556
rect 418212 275544 418218 275596
rect 418338 275544 418344 275596
rect 418396 275584 418402 275596
rect 435910 275584 435916 275596
rect 418396 275556 435916 275584
rect 418396 275544 418402 275556
rect 435910 275544 435916 275556
rect 435968 275544 435974 275596
rect 449158 275544 449164 275596
rect 449216 275584 449222 275596
rect 504284 275584 504312 275692
rect 509142 275680 509148 275692
rect 509200 275680 509206 275732
rect 512178 275680 512184 275732
rect 512236 275720 512242 275732
rect 516226 275720 516232 275732
rect 512236 275692 516232 275720
rect 512236 275680 512242 275692
rect 516226 275680 516232 275692
rect 516284 275680 516290 275732
rect 516428 275720 516456 275828
rect 516778 275816 516784 275868
rect 516836 275856 516842 275868
rect 524248 275856 524276 275964
rect 604914 275952 604920 275964
rect 604972 275952 604978 276004
rect 516836 275828 524276 275856
rect 516836 275816 516842 275828
rect 524874 275816 524880 275868
rect 524932 275856 524938 275868
rect 611998 275856 612004 275868
rect 524932 275828 612004 275856
rect 524932 275816 524938 275828
rect 611998 275816 612004 275828
rect 612056 275816 612062 275868
rect 519170 275720 519176 275732
rect 516428 275692 519176 275720
rect 519170 275680 519176 275692
rect 519228 275680 519234 275732
rect 519354 275680 519360 275732
rect 519412 275720 519418 275732
rect 522206 275720 522212 275732
rect 519412 275692 522212 275720
rect 519412 275680 519418 275692
rect 522206 275680 522212 275692
rect 522264 275680 522270 275732
rect 530302 275680 530308 275732
rect 530360 275720 530366 275732
rect 530360 275692 530716 275720
rect 530360 275680 530366 275692
rect 519538 275584 519544 275596
rect 449216 275556 504312 275584
rect 504376 275556 519544 275584
rect 449216 275544 449222 275556
rect 85942 275408 85948 275460
rect 86000 275448 86006 275460
rect 146754 275448 146760 275460
rect 86000 275420 146760 275448
rect 86000 275408 86006 275420
rect 146754 275408 146760 275420
rect 146812 275408 146818 275460
rect 160462 275408 160468 275460
rect 160520 275448 160526 275460
rect 167730 275448 167736 275460
rect 160520 275420 167736 275448
rect 160520 275408 160526 275420
rect 167730 275408 167736 275420
rect 167788 275408 167794 275460
rect 171042 275408 171048 275460
rect 171100 275448 171106 275460
rect 210786 275448 210792 275460
rect 171100 275420 210792 275448
rect 171100 275408 171106 275420
rect 210786 275408 210792 275420
rect 210844 275408 210850 275460
rect 218330 275408 218336 275460
rect 218388 275448 218394 275460
rect 237466 275448 237472 275460
rect 218388 275420 237472 275448
rect 218388 275408 218394 275420
rect 237466 275408 237472 275420
rect 237524 275408 237530 275460
rect 244366 275408 244372 275460
rect 244424 275448 244430 275460
rect 254578 275448 254584 275460
rect 244424 275420 254584 275448
rect 244424 275408 244430 275420
rect 254578 275408 254584 275420
rect 254636 275408 254642 275460
rect 260926 275408 260932 275460
rect 260984 275448 260990 275460
rect 273530 275448 273536 275460
rect 260984 275420 273536 275448
rect 260984 275408 260990 275420
rect 273530 275408 273536 275420
rect 273588 275408 273594 275460
rect 273898 275408 273904 275460
rect 273956 275448 273962 275460
rect 282914 275448 282920 275460
rect 273956 275420 282920 275448
rect 273956 275408 273962 275420
rect 282914 275408 282920 275420
rect 282972 275408 282978 275460
rect 326430 275408 326436 275460
rect 326488 275448 326494 275460
rect 335354 275448 335360 275460
rect 326488 275420 335360 275448
rect 326488 275408 326494 275420
rect 335354 275408 335360 275420
rect 335412 275408 335418 275460
rect 341518 275408 341524 275460
rect 341576 275448 341582 275460
rect 354306 275448 354312 275460
rect 341576 275420 354312 275448
rect 341576 275408 341582 275420
rect 354306 275408 354312 275420
rect 354364 275408 354370 275460
rect 360194 275448 360200 275460
rect 354646 275420 360200 275448
rect 298738 275340 298744 275392
rect 298796 275380 298802 275392
rect 300026 275380 300032 275392
rect 298796 275352 300032 275380
rect 298796 275340 298802 275352
rect 300026 275340 300032 275352
rect 300084 275340 300090 275392
rect 70578 275272 70584 275324
rect 70636 275312 70642 275324
rect 140130 275312 140136 275324
rect 70636 275284 140136 275312
rect 70636 275272 70642 275284
rect 140130 275272 140136 275284
rect 140188 275272 140194 275324
rect 142706 275272 142712 275324
rect 142764 275312 142770 275324
rect 183462 275312 183468 275324
rect 142764 275284 183468 275312
rect 142764 275272 142770 275284
rect 183462 275272 183468 275284
rect 183520 275272 183526 275324
rect 186406 275272 186412 275324
rect 186464 275312 186470 275324
rect 187786 275312 187792 275324
rect 186464 275284 187792 275312
rect 186464 275272 186470 275284
rect 187786 275272 187792 275284
rect 187844 275272 187850 275324
rect 188798 275272 188804 275324
rect 188856 275312 188862 275324
rect 222838 275312 222844 275324
rect 188856 275284 222844 275312
rect 188856 275272 188862 275284
rect 222838 275272 222844 275284
rect 222896 275272 222902 275324
rect 225414 275272 225420 275324
rect 225472 275312 225478 275324
rect 245102 275312 245108 275324
rect 225472 275284 245108 275312
rect 225472 275272 225478 275284
rect 245102 275272 245108 275284
rect 245160 275272 245166 275324
rect 250254 275272 250260 275324
rect 250312 275312 250318 275324
rect 266354 275312 266360 275324
rect 250312 275284 266360 275312
rect 250312 275272 250318 275284
rect 266354 275272 266360 275284
rect 266412 275272 266418 275324
rect 266814 275272 266820 275324
rect 266872 275312 266878 275324
rect 276658 275312 276664 275324
rect 266872 275284 276664 275312
rect 266872 275272 266878 275284
rect 276658 275272 276664 275284
rect 276716 275272 276722 275324
rect 284570 275272 284576 275324
rect 284628 275312 284634 275324
rect 290090 275312 290096 275324
rect 284628 275284 290096 275312
rect 284628 275272 284634 275284
rect 290090 275272 290096 275284
rect 290148 275272 290154 275324
rect 329466 275272 329472 275324
rect 329524 275312 329530 275324
rect 338942 275312 338948 275324
rect 329524 275284 338948 275312
rect 329524 275272 329530 275284
rect 338942 275272 338948 275284
rect 339000 275272 339006 275324
rect 353110 275312 353116 275324
rect 344986 275284 353116 275312
rect 74074 275136 74080 275188
rect 74132 275176 74138 275188
rect 77202 275176 77208 275188
rect 74132 275148 77208 275176
rect 74132 275136 74138 275148
rect 77202 275136 77208 275148
rect 77260 275136 77266 275188
rect 110782 275136 110788 275188
rect 110840 275176 110846 275188
rect 162118 275176 162124 275188
rect 110840 275148 162124 275176
rect 110840 275136 110846 275148
rect 162118 275136 162124 275148
rect 162176 275136 162182 275188
rect 338942 275136 338948 275188
rect 339000 275176 339006 275188
rect 344986 275176 345014 275284
rect 353110 275272 353116 275284
rect 353168 275272 353174 275324
rect 353938 275272 353944 275324
rect 353996 275312 354002 275324
rect 354646 275312 354674 275420
rect 360194 275408 360200 275420
rect 360252 275408 360258 275460
rect 363046 275408 363052 275460
rect 363104 275448 363110 275460
rect 367278 275448 367284 275460
rect 363104 275420 367284 275448
rect 363104 275408 363110 275420
rect 367278 275408 367284 275420
rect 367336 275408 367342 275460
rect 369118 275408 369124 275460
rect 369176 275448 369182 275460
rect 377950 275448 377956 275460
rect 369176 275420 377956 275448
rect 369176 275408 369182 275420
rect 377950 275408 377956 275420
rect 378008 275408 378014 275460
rect 381998 275408 382004 275460
rect 382056 275448 382062 275460
rect 414566 275448 414572 275460
rect 382056 275420 414572 275448
rect 382056 275408 382062 275420
rect 414566 275408 414572 275420
rect 414624 275408 414630 275460
rect 416406 275408 416412 275460
rect 416464 275448 416470 275460
rect 463050 275448 463056 275460
rect 416464 275420 463056 275448
rect 416464 275408 416470 275420
rect 463050 275408 463056 275420
rect 463108 275408 463114 275460
rect 467650 275408 467656 275460
rect 467708 275448 467714 275460
rect 504376 275448 504404 275556
rect 519538 275544 519544 275556
rect 519596 275544 519602 275596
rect 519722 275544 519728 275596
rect 519780 275584 519786 275596
rect 522390 275584 522396 275596
rect 519780 275556 522396 275584
rect 519780 275544 519786 275556
rect 522390 275544 522396 275556
rect 522448 275544 522454 275596
rect 530688 275584 530716 275692
rect 530854 275680 530860 275732
rect 530912 275720 530918 275732
rect 619082 275720 619088 275732
rect 530912 275692 619088 275720
rect 530912 275680 530918 275692
rect 619082 275680 619088 275692
rect 619140 275680 619146 275732
rect 536834 275584 536840 275596
rect 530688 275556 536840 275584
rect 536834 275544 536840 275556
rect 536892 275544 536898 275596
rect 537018 275544 537024 275596
rect 537076 275584 537082 275596
rect 537754 275584 537760 275596
rect 537076 275556 537760 275584
rect 537076 275544 537082 275556
rect 537754 275544 537760 275556
rect 537812 275544 537818 275596
rect 537938 275544 537944 275596
rect 537996 275584 538002 275596
rect 626166 275584 626172 275596
rect 537996 275556 626172 275584
rect 537996 275544 538002 275556
rect 626166 275544 626172 275556
rect 626224 275544 626230 275596
rect 467708 275420 504404 275448
rect 467708 275408 467714 275420
rect 504542 275408 504548 275460
rect 504600 275448 504606 275460
rect 538214 275448 538220 275460
rect 504600 275420 538220 275448
rect 504600 275408 504606 275420
rect 538214 275408 538220 275420
rect 538272 275408 538278 275460
rect 540974 275448 540980 275460
rect 538416 275420 540980 275448
rect 353996 275284 354674 275312
rect 353996 275272 354002 275284
rect 356330 275272 356336 275324
rect 356388 275312 356394 275324
rect 368474 275312 368480 275324
rect 356388 275284 368480 275312
rect 356388 275272 356394 275284
rect 368474 275272 368480 275284
rect 368532 275272 368538 275324
rect 375098 275272 375104 275324
rect 375156 275312 375162 275324
rect 403986 275312 403992 275324
rect 375156 275284 403992 275312
rect 375156 275272 375162 275284
rect 403986 275272 403992 275284
rect 404044 275272 404050 275324
rect 411254 275272 411260 275324
rect 411312 275312 411318 275324
rect 455966 275312 455972 275324
rect 411312 275284 455972 275312
rect 411312 275272 411318 275284
rect 455966 275272 455972 275284
rect 456024 275272 456030 275324
rect 512178 275312 512184 275324
rect 456168 275284 512184 275312
rect 339000 275148 345014 275176
rect 339000 275136 339006 275148
rect 420914 275136 420920 275188
rect 420972 275176 420978 275188
rect 434714 275176 434720 275188
rect 420972 275148 434720 275176
rect 420972 275136 420978 275148
rect 434714 275136 434720 275148
rect 434772 275136 434778 275188
rect 437474 275136 437480 275188
rect 437532 275176 437538 275188
rect 450078 275176 450084 275188
rect 437532 275148 450084 275176
rect 437532 275136 437538 275148
rect 450078 275136 450084 275148
rect 450136 275136 450142 275188
rect 455874 275136 455880 275188
rect 455932 275176 455938 275188
rect 456168 275176 456196 275284
rect 512178 275272 512184 275284
rect 512236 275272 512242 275324
rect 519354 275312 519360 275324
rect 512380 275284 519360 275312
rect 455932 275148 456196 275176
rect 455932 275136 455938 275148
rect 456794 275136 456800 275188
rect 456852 275176 456858 275188
rect 467834 275176 467840 275188
rect 456852 275148 467840 275176
rect 456852 275136 456858 275148
rect 467834 275136 467840 275148
rect 467892 275136 467898 275188
rect 468202 275136 468208 275188
rect 468260 275176 468266 275188
rect 494974 275176 494980 275188
rect 468260 275148 494980 275176
rect 468260 275136 468266 275148
rect 494974 275136 494980 275148
rect 495032 275136 495038 275188
rect 495158 275136 495164 275188
rect 495216 275176 495222 275188
rect 512380 275176 512408 275284
rect 519354 275272 519360 275284
rect 519412 275272 519418 275324
rect 519538 275272 519544 275324
rect 519596 275312 519602 275324
rect 537570 275312 537576 275324
rect 519596 275284 537576 275312
rect 519596 275272 519602 275284
rect 537570 275272 537576 275284
rect 537628 275272 537634 275324
rect 537754 275272 537760 275324
rect 537812 275312 537818 275324
rect 538416 275312 538444 275420
rect 540974 275408 540980 275420
rect 541032 275408 541038 275460
rect 541158 275408 541164 275460
rect 541216 275448 541222 275460
rect 544654 275448 544660 275460
rect 541216 275420 544660 275448
rect 541216 275408 541222 275420
rect 544654 275408 544660 275420
rect 544712 275408 544718 275460
rect 544838 275408 544844 275460
rect 544896 275448 544902 275460
rect 546034 275448 546040 275460
rect 544896 275420 546040 275448
rect 544896 275408 544902 275420
rect 546034 275408 546040 275420
rect 546092 275408 546098 275460
rect 546218 275408 546224 275460
rect 546276 275448 546282 275460
rect 641622 275448 641628 275460
rect 546276 275420 641628 275448
rect 546276 275408 546282 275420
rect 641622 275408 641628 275420
rect 641680 275408 641686 275460
rect 537812 275284 538444 275312
rect 537812 275272 537818 275284
rect 538674 275272 538680 275324
rect 538732 275312 538738 275324
rect 633342 275312 633348 275324
rect 538732 275284 633348 275312
rect 538732 275272 538738 275284
rect 633342 275272 633348 275284
rect 633400 275272 633406 275324
rect 590746 275176 590752 275188
rect 495216 275148 512408 275176
rect 512472 275148 590752 275176
rect 495216 275136 495222 275148
rect 224218 275068 224224 275120
rect 224276 275108 224282 275120
rect 226150 275108 226156 275120
rect 224276 275080 226156 275108
rect 224276 275068 224282 275080
rect 226150 275068 226156 275080
rect 226208 275068 226214 275120
rect 294046 275068 294052 275120
rect 294104 275108 294110 275120
rect 295150 275108 295156 275120
rect 294104 275080 295156 275108
rect 294104 275068 294110 275080
rect 295150 275068 295156 275080
rect 295208 275068 295214 275120
rect 135622 275000 135628 275052
rect 135680 275040 135686 275052
rect 182082 275040 182088 275052
rect 135680 275012 182088 275040
rect 135680 275000 135686 275012
rect 182082 275000 182088 275012
rect 182140 275000 182146 275052
rect 449894 275000 449900 275052
rect 449952 275040 449958 275052
rect 460658 275040 460664 275052
rect 449952 275012 460664 275040
rect 449952 275000 449958 275012
rect 460658 275000 460664 275012
rect 460716 275000 460722 275052
rect 494698 275000 494704 275052
rect 494756 275040 494762 275052
rect 498562 275040 498568 275052
rect 494756 275012 498568 275040
rect 494756 275000 494762 275012
rect 498562 275000 498568 275012
rect 498620 275000 498626 275052
rect 505094 275000 505100 275052
rect 505152 275040 505158 275052
rect 506842 275040 506848 275052
rect 505152 275012 506848 275040
rect 505152 275000 505158 275012
rect 506842 275000 506848 275012
rect 506900 275000 506906 275052
rect 507026 275000 507032 275052
rect 507084 275040 507090 275052
rect 512472 275040 512500 275148
rect 590746 275136 590752 275148
rect 590804 275136 590810 275188
rect 611354 275136 611360 275188
rect 611412 275176 611418 275188
rect 616782 275176 616788 275188
rect 611412 275148 616788 275176
rect 611412 275136 611418 275148
rect 616782 275136 616788 275148
rect 616840 275136 616846 275188
rect 619174 275136 619180 275188
rect 619232 275176 619238 275188
rect 623866 275176 623872 275188
rect 619232 275148 623872 275176
rect 619232 275136 619238 275148
rect 623866 275136 623872 275148
rect 623924 275136 623930 275188
rect 507084 275012 512500 275040
rect 507084 275000 507090 275012
rect 514018 275000 514024 275052
rect 514076 275040 514082 275052
rect 583662 275040 583668 275052
rect 514076 275012 583668 275040
rect 514076 275000 514082 275012
rect 583662 275000 583668 275012
rect 583720 275000 583726 275052
rect 71774 274932 71780 274984
rect 71832 274972 71838 274984
rect 73798 274972 73804 274984
rect 71832 274944 73804 274972
rect 71832 274932 71838 274944
rect 73798 274932 73804 274944
rect 73856 274932 73862 274984
rect 277486 274932 277492 274984
rect 277544 274972 277550 274984
rect 284294 274972 284300 274984
rect 277544 274944 284300 274972
rect 277544 274932 277550 274944
rect 284294 274932 284300 274944
rect 284352 274932 284358 274984
rect 129642 274864 129648 274916
rect 129700 274904 129706 274916
rect 136542 274904 136548 274916
rect 129700 274876 136548 274904
rect 129700 274864 129706 274876
rect 136542 274864 136548 274876
rect 136600 274864 136606 274916
rect 149790 274864 149796 274916
rect 149848 274904 149854 274916
rect 185578 274904 185584 274916
rect 149848 274876 185584 274904
rect 149848 274864 149854 274876
rect 185578 274864 185584 274876
rect 185636 274864 185642 274916
rect 289262 274864 289268 274916
rect 289320 274904 289326 274916
rect 293402 274904 293408 274916
rect 289320 274876 293408 274904
rect 289320 274864 289326 274876
rect 293402 274864 293408 274876
rect 293460 274864 293466 274916
rect 470962 274864 470968 274916
rect 471020 274904 471026 274916
rect 523126 274904 523132 274916
rect 471020 274876 523132 274904
rect 471020 274864 471026 274876
rect 523126 274864 523132 274876
rect 523184 274864 523190 274916
rect 523310 274864 523316 274916
rect 523368 274904 523374 274916
rect 597830 274904 597836 274916
rect 523368 274876 597836 274904
rect 523368 274864 523374 274876
rect 597830 274864 597836 274876
rect 597888 274864 597894 274916
rect 283374 274796 283380 274848
rect 283432 274836 283438 274848
rect 289078 274836 289084 274848
rect 283432 274808 289084 274836
rect 283432 274796 283438 274808
rect 289078 274796 289084 274808
rect 289136 274796 289142 274848
rect 403986 274796 403992 274848
rect 404044 274836 404050 274848
rect 407482 274836 407488 274848
rect 404044 274808 407488 274836
rect 404044 274796 404050 274808
rect 407482 274796 407488 274808
rect 407540 274796 407546 274848
rect 426250 274796 426256 274848
rect 426308 274836 426314 274848
rect 432322 274836 432328 274848
rect 426308 274808 432328 274836
rect 426308 274796 426314 274808
rect 432322 274796 432328 274808
rect 432380 274796 432386 274848
rect 105998 274728 106004 274780
rect 106056 274768 106062 274780
rect 110414 274768 110420 274780
rect 106056 274740 110420 274768
rect 106056 274728 106062 274740
rect 110414 274728 110420 274740
rect 110472 274728 110478 274780
rect 140314 274728 140320 274780
rect 140372 274768 140378 274780
rect 144638 274768 144644 274780
rect 140372 274740 144644 274768
rect 140372 274728 140378 274740
rect 144638 274728 144644 274740
rect 144696 274728 144702 274780
rect 146202 274728 146208 274780
rect 146260 274768 146266 274780
rect 149882 274768 149888 274780
rect 146260 274740 149888 274768
rect 146260 274728 146266 274740
rect 149882 274728 149888 274740
rect 149940 274728 149946 274780
rect 435634 274728 435640 274780
rect 435692 274768 435698 274780
rect 439406 274768 439412 274780
rect 435692 274740 439412 274768
rect 435692 274728 435698 274740
rect 439406 274728 439412 274740
rect 439464 274728 439470 274780
rect 453942 274728 453948 274780
rect 454000 274768 454006 274780
rect 457162 274768 457168 274780
rect 454000 274740 457168 274768
rect 454000 274728 454006 274740
rect 457162 274728 457168 274740
rect 457220 274728 457226 274780
rect 464154 274728 464160 274780
rect 464212 274768 464218 274780
rect 471330 274768 471336 274780
rect 464212 274740 471336 274768
rect 464212 274728 464218 274740
rect 471330 274728 471336 274740
rect 471388 274728 471394 274780
rect 482922 274728 482928 274780
rect 482980 274768 482986 274780
rect 538306 274768 538312 274780
rect 482980 274740 538312 274768
rect 482980 274728 482986 274740
rect 538306 274728 538312 274740
rect 538364 274728 538370 274780
rect 538490 274728 538496 274780
rect 538548 274768 538554 274780
rect 545850 274768 545856 274780
rect 538548 274740 545856 274768
rect 538548 274728 538554 274740
rect 545850 274728 545856 274740
rect 545908 274728 545914 274780
rect 546034 274728 546040 274780
rect 546092 274768 546098 274780
rect 558822 274768 558828 274780
rect 546092 274740 558828 274768
rect 546092 274728 546098 274740
rect 558822 274728 558828 274740
rect 558880 274728 558886 274780
rect 66990 274660 66996 274712
rect 67048 274700 67054 274712
rect 71038 274700 71044 274712
rect 67048 274672 71044 274700
rect 67048 274660 67054 274672
rect 71038 274660 71044 274672
rect 71096 274660 71102 274712
rect 90634 274660 90640 274712
rect 90692 274700 90698 274712
rect 95878 274700 95884 274712
rect 90692 274672 95884 274700
rect 90692 274660 90698 274672
rect 95878 274660 95884 274672
rect 95936 274660 95942 274712
rect 161566 274660 161572 274712
rect 161624 274700 161630 274712
rect 163130 274700 163136 274712
rect 161624 274672 163136 274700
rect 161624 274660 161630 274672
rect 163130 274660 163136 274672
rect 163188 274660 163194 274712
rect 170122 274660 170128 274712
rect 170180 274700 170186 274712
rect 173066 274700 173072 274712
rect 170180 274672 173072 274700
rect 170180 274660 170186 274672
rect 173066 274660 173072 274672
rect 173124 274660 173130 274712
rect 185210 274660 185216 274712
rect 185268 274700 185274 274712
rect 187142 274700 187148 274712
rect 185268 274672 187148 274700
rect 185268 274660 185274 274672
rect 187142 274660 187148 274672
rect 187200 274660 187206 274712
rect 238478 274660 238484 274712
rect 238536 274700 238542 274712
rect 239766 274700 239772 274712
rect 238536 274672 239772 274700
rect 238536 274660 238542 274672
rect 239766 274660 239772 274672
rect 239824 274660 239830 274712
rect 285766 274660 285772 274712
rect 285824 274700 285830 274712
rect 286962 274700 286968 274712
rect 285824 274672 286968 274700
rect 285824 274660 285830 274672
rect 286962 274660 286968 274672
rect 287020 274660 287026 274712
rect 290458 274660 290464 274712
rect 290516 274700 290522 274712
rect 294138 274700 294144 274712
rect 290516 274672 294144 274700
rect 290516 274660 290522 274672
rect 294138 274660 294144 274672
rect 294196 274660 294202 274712
rect 296346 274660 296352 274712
rect 296404 274700 296410 274712
rect 298370 274700 298376 274712
rect 296404 274672 298376 274700
rect 296404 274660 296410 274672
rect 298370 274660 298376 274672
rect 298428 274660 298434 274712
rect 360286 274660 360292 274712
rect 360344 274700 360350 274712
rect 363782 274700 363788 274712
rect 360344 274672 363788 274700
rect 360344 274660 360350 274672
rect 363782 274660 363788 274672
rect 363840 274660 363846 274712
rect 367094 274660 367100 274712
rect 367152 274700 367158 274712
rect 369670 274700 369676 274712
rect 367152 274672 369676 274700
rect 367152 274660 367158 274672
rect 369670 274660 369676 274672
rect 369728 274660 369734 274712
rect 386046 274660 386052 274712
rect 386104 274700 386110 274712
rect 389726 274700 389732 274712
rect 386104 274672 389732 274700
rect 386104 274660 386110 274672
rect 389726 274660 389732 274672
rect 389784 274660 389790 274712
rect 407114 274660 407120 274712
rect 407172 274700 407178 274712
rect 411070 274700 411076 274712
rect 407172 274672 411076 274700
rect 407172 274660 407178 274672
rect 411070 274660 411076 274672
rect 411128 274660 411134 274712
rect 104802 274592 104808 274644
rect 104860 274632 104866 274644
rect 157610 274632 157616 274644
rect 104860 274604 157616 274632
rect 104860 274592 104866 274604
rect 157610 274592 157616 274604
rect 157668 274592 157674 274644
rect 195882 274592 195888 274644
rect 195940 274632 195946 274644
rect 206278 274632 206284 274644
rect 195940 274604 206284 274632
rect 195940 274592 195946 274604
rect 206278 274592 206284 274604
rect 206336 274592 206342 274644
rect 424962 274592 424968 274644
rect 425020 274632 425026 274644
rect 474918 274632 474924 274644
rect 425020 274604 474924 274632
rect 425020 274592 425026 274604
rect 474918 274592 474924 274604
rect 474976 274592 474982 274644
rect 475378 274592 475384 274644
rect 475436 274632 475442 274644
rect 490558 274632 490564 274644
rect 475436 274604 490564 274632
rect 475436 274592 475442 274604
rect 490558 274592 490564 274604
rect 490616 274592 490622 274644
rect 490742 274592 490748 274644
rect 490800 274632 490806 274644
rect 496170 274632 496176 274644
rect 490800 274604 496176 274632
rect 490800 274592 490806 274604
rect 496170 274592 496176 274604
rect 496228 274592 496234 274644
rect 570690 274632 570696 274644
rect 499546 274604 570696 274632
rect 121362 274456 121368 274508
rect 121420 274496 121426 274508
rect 176746 274496 176752 274508
rect 121420 274468 176752 274496
rect 121420 274456 121426 274468
rect 176746 274456 176752 274468
rect 176804 274456 176810 274508
rect 182910 274456 182916 274508
rect 182968 274496 182974 274508
rect 199654 274496 199660 274508
rect 182968 274468 199660 274496
rect 182968 274456 182974 274468
rect 199654 274456 199660 274468
rect 199712 274456 199718 274508
rect 210050 274456 210056 274508
rect 210108 274496 210114 274508
rect 237834 274496 237840 274508
rect 210108 274468 237840 274496
rect 210108 274456 210114 274468
rect 237834 274456 237840 274468
rect 237892 274456 237898 274508
rect 392578 274456 392584 274508
rect 392636 274496 392642 274508
rect 402790 274496 402796 274508
rect 392636 274468 402796 274496
rect 392636 274456 392642 274468
rect 402790 274456 402796 274468
rect 402848 274456 402854 274508
rect 406838 274456 406844 274508
rect 406896 274496 406902 274508
rect 437474 274496 437480 274508
rect 406896 274468 437480 274496
rect 406896 274456 406902 274468
rect 437474 274456 437480 274468
rect 437532 274456 437538 274508
rect 440878 274456 440884 274508
rect 440936 274496 440942 274508
rect 488442 274496 488448 274508
rect 440936 274468 488448 274496
rect 440936 274456 440942 274468
rect 488442 274456 488448 274468
rect 488500 274456 488506 274508
rect 491018 274496 491024 274508
rect 488644 274468 491024 274496
rect 101306 274320 101312 274372
rect 101364 274360 101370 274372
rect 160922 274360 160928 274372
rect 101364 274332 160928 274360
rect 101364 274320 101370 274332
rect 160922 274320 160928 274332
rect 160980 274320 160986 274372
rect 187786 274320 187792 274372
rect 187844 274360 187850 274372
rect 220906 274360 220912 274372
rect 187844 274332 220912 274360
rect 187844 274320 187850 274332
rect 220906 274320 220912 274332
rect 220964 274320 220970 274372
rect 362862 274320 362868 274372
rect 362920 274360 362926 274372
rect 386230 274360 386236 274372
rect 362920 274332 386236 274360
rect 362920 274320 362926 274332
rect 386230 274320 386236 274332
rect 386288 274320 386294 274372
rect 395890 274320 395896 274372
rect 395948 274360 395954 274372
rect 420914 274360 420920 274372
rect 395948 274332 420920 274360
rect 395948 274320 395954 274332
rect 420914 274320 420920 274332
rect 420972 274320 420978 274372
rect 471238 274320 471244 274372
rect 471296 274360 471302 274372
rect 488644 274360 488672 274468
rect 491018 274456 491024 274468
rect 491076 274456 491082 274508
rect 491202 274456 491208 274508
rect 491260 274496 491266 274508
rect 499546 274496 499574 274604
rect 570690 274592 570696 274604
rect 570748 274592 570754 274644
rect 570874 274592 570880 274644
rect 570932 274632 570938 274644
rect 587158 274632 587164 274644
rect 570932 274604 587164 274632
rect 570932 274592 570938 274604
rect 587158 274592 587164 274604
rect 587216 274592 587222 274644
rect 491260 274468 499574 274496
rect 491260 274456 491266 274468
rect 501966 274456 501972 274508
rect 502024 274496 502030 274508
rect 502024 274468 504588 274496
rect 502024 274456 502030 274468
rect 471296 274332 488672 274360
rect 471296 274320 471302 274332
rect 490558 274320 490564 274372
rect 490616 274360 490622 274372
rect 504560 274360 504588 274468
rect 504726 274456 504732 274508
rect 504784 274496 504790 274508
rect 577774 274496 577780 274508
rect 504784 274468 577780 274496
rect 504784 274456 504790 274468
rect 577774 274456 577780 274468
rect 577832 274456 577838 274508
rect 585778 274456 585784 274508
rect 585836 274496 585842 274508
rect 585836 274468 586514 274496
rect 585836 274456 585842 274468
rect 586054 274360 586060 274372
rect 490616 274332 504496 274360
rect 504560 274332 586060 274360
rect 490616 274320 490622 274332
rect 82354 274184 82360 274236
rect 82412 274224 82418 274236
rect 145558 274224 145564 274236
rect 82412 274196 145564 274224
rect 82412 274184 82418 274196
rect 145558 274184 145564 274196
rect 145616 274184 145622 274236
rect 160094 274184 160100 274236
rect 160152 274224 160158 274236
rect 164234 274224 164240 274236
rect 160152 274196 164240 274224
rect 160152 274184 160158 274196
rect 164234 274184 164240 274196
rect 164292 274184 164298 274236
rect 176930 274184 176936 274236
rect 176988 274224 176994 274236
rect 214650 274224 214656 274236
rect 176988 274196 214656 274224
rect 176988 274184 176994 274196
rect 214650 274184 214656 274196
rect 214708 274184 214714 274236
rect 220538 274184 220544 274236
rect 220596 274224 220602 274236
rect 240594 274224 240600 274236
rect 220596 274196 240600 274224
rect 220596 274184 220602 274196
rect 240594 274184 240600 274196
rect 240652 274184 240658 274236
rect 342898 274184 342904 274236
rect 342956 274224 342962 274236
rect 347222 274224 347228 274236
rect 342956 274196 347228 274224
rect 342956 274184 342962 274196
rect 347222 274184 347228 274196
rect 347280 274184 347286 274236
rect 366910 274184 366916 274236
rect 366968 274224 366974 274236
rect 389174 274224 389180 274236
rect 366968 274196 389180 274224
rect 366968 274184 366974 274196
rect 389174 274184 389180 274196
rect 389232 274184 389238 274236
rect 390278 274184 390284 274236
rect 390336 274224 390342 274236
rect 426434 274224 426440 274236
rect 390336 274196 426440 274224
rect 390336 274184 390342 274196
rect 426434 274184 426440 274196
rect 426492 274184 426498 274236
rect 438762 274184 438768 274236
rect 438820 274224 438826 274236
rect 490742 274224 490748 274236
rect 438820 274196 490748 274224
rect 438820 274184 438826 274196
rect 490742 274184 490748 274196
rect 490800 274184 490806 274236
rect 490926 274184 490932 274236
rect 490984 274224 490990 274236
rect 493778 274224 493784 274236
rect 490984 274196 493784 274224
rect 490984 274184 490990 274196
rect 493778 274184 493784 274196
rect 493836 274184 493842 274236
rect 496262 274184 496268 274236
rect 496320 274224 496326 274236
rect 504174 274224 504180 274236
rect 496320 274196 504180 274224
rect 496320 274184 496326 274196
rect 504174 274184 504180 274196
rect 504232 274184 504238 274236
rect 504468 274224 504496 274332
rect 586054 274320 586060 274332
rect 586112 274320 586118 274372
rect 586486 274360 586514 274468
rect 601418 274360 601424 274372
rect 586486 274332 601424 274360
rect 601418 274320 601424 274332
rect 601476 274320 601482 274372
rect 504468 274196 518296 274224
rect 84746 274048 84752 274100
rect 84804 274088 84810 274100
rect 148318 274088 148324 274100
rect 84804 274060 148324 274088
rect 84804 274048 84810 274060
rect 148318 274048 148324 274060
rect 148376 274048 148382 274100
rect 158070 274048 158076 274100
rect 158128 274088 158134 274100
rect 200666 274088 200672 274100
rect 158128 274060 200672 274088
rect 158128 274048 158134 274060
rect 200666 274048 200672 274060
rect 200724 274048 200730 274100
rect 206554 274048 206560 274100
rect 206612 274088 206618 274100
rect 235442 274088 235448 274100
rect 206612 274060 235448 274088
rect 206612 274048 206618 274060
rect 235442 274048 235448 274060
rect 235500 274048 235506 274100
rect 239582 274048 239588 274100
rect 239640 274088 239646 274100
rect 258626 274088 258632 274100
rect 239640 274060 258632 274088
rect 239640 274048 239646 274060
rect 258626 274048 258632 274060
rect 258684 274048 258690 274100
rect 360102 274048 360108 274100
rect 360160 274088 360166 274100
rect 383838 274088 383844 274100
rect 360160 274060 383844 274088
rect 360160 274048 360166 274060
rect 383838 274048 383844 274060
rect 383896 274048 383902 274100
rect 384942 274048 384948 274100
rect 385000 274088 385006 274100
rect 419350 274088 419356 274100
rect 385000 274060 419356 274088
rect 385000 274048 385006 274060
rect 419350 274048 419356 274060
rect 419408 274048 419414 274100
rect 421558 274048 421564 274100
rect 421616 274088 421622 274100
rect 458358 274088 458364 274100
rect 421616 274060 458364 274088
rect 421616 274048 421622 274060
rect 458358 274048 458364 274060
rect 458416 274048 458422 274100
rect 459370 274048 459376 274100
rect 459428 274088 459434 274100
rect 516594 274088 516600 274100
rect 459428 274060 516600 274088
rect 459428 274048 459434 274060
rect 516594 274048 516600 274060
rect 516652 274048 516658 274100
rect 518268 274088 518296 274196
rect 518434 274184 518440 274236
rect 518492 274224 518498 274236
rect 602522 274224 602528 274236
rect 518492 274196 602528 274224
rect 518492 274184 518498 274196
rect 602522 274184 602528 274196
rect 602580 274184 602586 274236
rect 613378 274184 613384 274236
rect 613436 274224 613442 274236
rect 615586 274224 615592 274236
rect 613436 274196 615592 274224
rect 613436 274184 613442 274196
rect 615586 274184 615592 274196
rect 615644 274184 615650 274236
rect 527818 274088 527824 274100
rect 518268 274060 527824 274088
rect 527818 274048 527824 274060
rect 527876 274048 527882 274100
rect 528002 274048 528008 274100
rect 528060 274088 528066 274100
rect 619174 274088 619180 274100
rect 528060 274060 619180 274088
rect 528060 274048 528066 274060
rect 619174 274048 619180 274060
rect 619232 274048 619238 274100
rect 77202 273912 77208 273964
rect 77260 273952 77266 273964
rect 143534 273952 143540 273964
rect 77260 273924 143540 273952
rect 77260 273912 77266 273924
rect 143534 273912 143540 273924
rect 143592 273912 143598 273964
rect 145006 273912 145012 273964
rect 145064 273952 145070 273964
rect 192478 273952 192484 273964
rect 145064 273924 192484 273952
rect 145064 273912 145070 273924
rect 192478 273912 192484 273924
rect 192536 273912 192542 273964
rect 193490 273912 193496 273964
rect 193548 273952 193554 273964
rect 226334 273952 226340 273964
rect 193548 273924 226340 273952
rect 193548 273912 193554 273924
rect 226334 273912 226340 273924
rect 226392 273912 226398 273964
rect 234890 273912 234896 273964
rect 234948 273952 234954 273964
rect 255498 273952 255504 273964
rect 234948 273924 255504 273952
rect 234948 273912 234954 273924
rect 255498 273912 255504 273924
rect 255556 273912 255562 273964
rect 256142 273912 256148 273964
rect 256200 273952 256206 273964
rect 270586 273952 270592 273964
rect 256200 273924 270592 273952
rect 256200 273912 256206 273924
rect 270586 273912 270592 273924
rect 270644 273912 270650 273964
rect 271506 273912 271512 273964
rect 271564 273952 271570 273964
rect 280798 273952 280804 273964
rect 271564 273924 280804 273952
rect 271564 273912 271570 273924
rect 280798 273912 280804 273924
rect 280856 273912 280862 273964
rect 346302 273912 346308 273964
rect 346360 273952 346366 273964
rect 362586 273952 362592 273964
rect 346360 273924 362592 273952
rect 346360 273912 346366 273924
rect 362586 273912 362592 273924
rect 362644 273912 362650 273964
rect 377766 273912 377772 273964
rect 377824 273952 377830 273964
rect 408678 273952 408684 273964
rect 377824 273924 408684 273952
rect 377824 273912 377830 273924
rect 408678 273912 408684 273924
rect 408736 273912 408742 273964
rect 413922 273912 413928 273964
rect 413980 273952 413986 273964
rect 449894 273952 449900 273964
rect 413980 273924 449900 273952
rect 413980 273912 413986 273924
rect 449894 273912 449900 273924
rect 449952 273912 449958 273964
rect 451090 273912 451096 273964
rect 451148 273952 451154 273964
rect 513834 273952 513840 273964
rect 451148 273924 513840 273952
rect 451148 273912 451154 273924
rect 513834 273912 513840 273924
rect 513892 273912 513898 273964
rect 519722 273912 519728 273964
rect 519780 273952 519786 273964
rect 524230 273952 524236 273964
rect 519780 273924 524236 273952
rect 519780 273912 519786 273924
rect 524230 273912 524236 273924
rect 524288 273912 524294 273964
rect 524414 273912 524420 273964
rect 524472 273952 524478 273964
rect 613194 273952 613200 273964
rect 524472 273924 613200 273952
rect 524472 273912 524478 273924
rect 613194 273912 613200 273924
rect 613252 273912 613258 273964
rect 123754 273776 123760 273828
rect 123812 273816 123818 273828
rect 177482 273816 177488 273828
rect 123812 273788 177488 273816
rect 123812 273776 123818 273788
rect 177482 273776 177488 273788
rect 177540 273776 177546 273828
rect 426894 273776 426900 273828
rect 426952 273816 426958 273828
rect 477218 273816 477224 273828
rect 426952 273788 477224 273816
rect 426952 273776 426958 273788
rect 477218 273776 477224 273788
rect 477276 273776 477282 273828
rect 488442 273776 488448 273828
rect 488500 273816 488506 273828
rect 490926 273816 490932 273828
rect 488500 273788 490932 273816
rect 488500 273776 488506 273788
rect 490926 273776 490932 273788
rect 490984 273776 490990 273828
rect 492030 273776 492036 273828
rect 492088 273816 492094 273828
rect 571794 273816 571800 273828
rect 492088 273788 571800 273816
rect 492088 273776 492094 273788
rect 571794 273776 571800 273788
rect 571852 273776 571858 273828
rect 280982 273708 280988 273760
rect 281040 273748 281046 273760
rect 287514 273748 287520 273760
rect 281040 273720 287520 273748
rect 281040 273708 281046 273720
rect 287514 273708 287520 273720
rect 287572 273708 287578 273760
rect 134426 273640 134432 273692
rect 134484 273680 134490 273692
rect 185026 273680 185032 273692
rect 134484 273652 185032 273680
rect 134484 273640 134490 273652
rect 185026 273640 185032 273652
rect 185084 273640 185090 273692
rect 460014 273640 460020 273692
rect 460072 273680 460078 273692
rect 484302 273680 484308 273692
rect 460072 273652 484308 273680
rect 460072 273640 460078 273652
rect 484302 273640 484308 273652
rect 484360 273640 484366 273692
rect 487982 273640 487988 273692
rect 488040 273680 488046 273692
rect 565906 273680 565912 273692
rect 488040 273652 565912 273680
rect 488040 273640 488046 273652
rect 565906 273640 565912 273652
rect 565964 273640 565970 273692
rect 144638 273504 144644 273556
rect 144696 273544 144702 273556
rect 187786 273544 187792 273556
rect 144696 273516 187792 273544
rect 144696 273504 144702 273516
rect 187786 273504 187792 273516
rect 187844 273504 187850 273556
rect 429010 273504 429016 273556
rect 429068 273544 429074 273556
rect 482002 273544 482008 273556
rect 429068 273516 482008 273544
rect 429068 273504 429074 273516
rect 482002 273504 482008 273516
rect 482060 273504 482066 273556
rect 487062 273504 487068 273556
rect 487120 273544 487126 273556
rect 563514 273544 563520 273556
rect 487120 273516 563520 273544
rect 487120 273504 487126 273516
rect 563514 273504 563520 273516
rect 563572 273504 563578 273556
rect 481358 273368 481364 273420
rect 481416 273408 481422 273420
rect 556430 273408 556436 273420
rect 481416 273380 556436 273408
rect 481416 273368 481422 273380
rect 556430 273368 556436 273380
rect 556488 273368 556494 273420
rect 347038 273232 347044 273284
rect 347096 273272 347102 273284
rect 349614 273272 349620 273284
rect 347096 273244 349620 273272
rect 347096 273232 347102 273244
rect 349614 273232 349620 273244
rect 349672 273232 349678 273284
rect 350258 273232 350264 273284
rect 350316 273272 350322 273284
rect 356330 273272 356336 273284
rect 350316 273244 356336 273272
rect 350316 273232 350322 273244
rect 356330 273232 356336 273244
rect 356388 273232 356394 273284
rect 409138 273232 409144 273284
rect 409196 273272 409202 273284
rect 409874 273272 409880 273284
rect 409196 273244 409880 273272
rect 409196 273232 409202 273244
rect 409874 273232 409880 273244
rect 409932 273232 409938 273284
rect 114278 273164 114284 273216
rect 114336 273204 114342 273216
rect 169018 273204 169024 273216
rect 114336 273176 169024 273204
rect 114336 273164 114342 273176
rect 169018 273164 169024 273176
rect 169076 273164 169082 273216
rect 211982 273204 211988 273216
rect 200086 273176 211988 273204
rect 104986 273028 104992 273080
rect 105044 273068 105050 273080
rect 163314 273068 163320 273080
rect 105044 273040 163320 273068
rect 105044 273028 105050 273040
rect 163314 273028 163320 273040
rect 163372 273028 163378 273080
rect 167546 273028 167552 273080
rect 167604 273068 167610 273080
rect 184198 273068 184204 273080
rect 167604 273040 184204 273068
rect 167604 273028 167610 273040
rect 184198 273028 184204 273040
rect 184256 273028 184262 273080
rect 187602 273028 187608 273080
rect 187660 273068 187666 273080
rect 200086 273068 200114 273176
rect 211982 273164 211988 273176
rect 212040 273164 212046 273216
rect 419166 273164 419172 273216
rect 419224 273204 419230 273216
rect 456794 273204 456800 273216
rect 419224 273176 456800 273204
rect 419224 273164 419230 273176
rect 456794 273164 456800 273176
rect 456852 273164 456858 273216
rect 463142 273164 463148 273216
rect 463200 273204 463206 273216
rect 486878 273204 486884 273216
rect 463200 273176 486884 273204
rect 463200 273164 463206 273176
rect 486878 273164 486884 273176
rect 486936 273164 486942 273216
rect 493686 273164 493692 273216
rect 493744 273204 493750 273216
rect 574186 273204 574192 273216
rect 493744 273176 574192 273204
rect 493744 273164 493750 273176
rect 574186 273164 574192 273176
rect 574244 273164 574250 273216
rect 578878 273164 578884 273216
rect 578936 273204 578942 273216
rect 594334 273204 594340 273216
rect 578936 273176 594340 273204
rect 578936 273164 578942 273176
rect 594334 273164 594340 273176
rect 594392 273164 594398 273216
rect 187660 273040 200114 273068
rect 187660 273028 187666 273040
rect 211246 273028 211252 273080
rect 211304 273068 211310 273080
rect 220078 273068 220084 273080
rect 211304 273040 220084 273068
rect 211304 273028 211310 273040
rect 220078 273028 220084 273040
rect 220136 273028 220142 273080
rect 382918 273028 382924 273080
rect 382976 273068 382982 273080
rect 392118 273068 392124 273080
rect 382976 273040 392124 273068
rect 382976 273028 382982 273040
rect 392118 273028 392124 273040
rect 392176 273028 392182 273080
rect 404170 273028 404176 273080
rect 404228 273068 404234 273080
rect 429194 273068 429200 273080
rect 404228 273040 429200 273068
rect 404228 273028 404234 273040
rect 429194 273028 429200 273040
rect 429252 273028 429258 273080
rect 434622 273028 434628 273080
rect 434680 273068 434686 273080
rect 488718 273068 488724 273080
rect 434680 273040 488724 273068
rect 434680 273028 434686 273040
rect 488718 273028 488724 273040
rect 488776 273028 488782 273080
rect 496630 273028 496636 273080
rect 496688 273068 496694 273080
rect 578510 273068 578516 273080
rect 496688 273040 578516 273068
rect 496688 273028 496694 273040
rect 578510 273028 578516 273040
rect 578568 273028 578574 273080
rect 580258 273028 580264 273080
rect 580316 273068 580322 273080
rect 640426 273068 640432 273080
rect 580316 273040 640432 273068
rect 580316 273028 580322 273040
rect 640426 273028 640432 273040
rect 640484 273028 640490 273080
rect 78858 272892 78864 272944
rect 78916 272932 78922 272944
rect 138658 272932 138664 272944
rect 78916 272904 138664 272932
rect 78916 272892 78922 272904
rect 138658 272892 138664 272904
rect 138716 272892 138722 272944
rect 141786 272892 141792 272944
rect 141844 272932 141850 272944
rect 189810 272932 189816 272944
rect 141844 272904 189816 272932
rect 141844 272892 141850 272904
rect 189810 272892 189816 272904
rect 189868 272892 189874 272944
rect 191190 272892 191196 272944
rect 191248 272932 191254 272944
rect 224862 272932 224868 272944
rect 191248 272904 224868 272932
rect 191248 272892 191254 272904
rect 224862 272892 224868 272904
rect 224920 272892 224926 272944
rect 288066 272892 288072 272944
rect 288124 272932 288130 272944
rect 290458 272932 290464 272944
rect 288124 272904 290464 272932
rect 288124 272892 288130 272904
rect 290458 272892 290464 272904
rect 290516 272892 290522 272944
rect 373258 272892 373264 272944
rect 373316 272932 373322 272944
rect 382642 272932 382648 272944
rect 373316 272904 382648 272932
rect 373316 272892 373322 272904
rect 382642 272892 382648 272904
rect 382700 272892 382706 272944
rect 388622 272932 388628 272944
rect 383626 272904 388628 272932
rect 94222 272756 94228 272808
rect 94280 272796 94286 272808
rect 156046 272796 156052 272808
rect 94280 272768 156052 272796
rect 94280 272756 94286 272768
rect 156046 272756 156052 272768
rect 156104 272756 156110 272808
rect 180518 272756 180524 272808
rect 180576 272796 180582 272808
rect 217226 272796 217232 272808
rect 180576 272768 217232 272796
rect 180576 272756 180582 272768
rect 217226 272756 217232 272768
rect 217284 272756 217290 272808
rect 228818 272756 228824 272808
rect 228876 272796 228882 272808
rect 249058 272796 249064 272808
rect 228876 272768 249064 272796
rect 228876 272756 228882 272768
rect 249058 272756 249064 272768
rect 249116 272756 249122 272808
rect 352926 272756 352932 272808
rect 352984 272796 352990 272808
rect 372982 272796 372988 272808
rect 352984 272768 372988 272796
rect 352984 272756 352990 272768
rect 372982 272756 372988 272768
rect 373040 272756 373046 272808
rect 380710 272756 380716 272808
rect 380768 272796 380774 272808
rect 383626 272796 383654 272904
rect 388622 272892 388628 272904
rect 388680 272892 388686 272944
rect 391842 272892 391848 272944
rect 391900 272932 391906 272944
rect 410058 272932 410064 272944
rect 391900 272904 410064 272932
rect 391900 272892 391906 272904
rect 410058 272892 410064 272904
rect 410116 272892 410122 272944
rect 412450 272892 412456 272944
rect 412508 272932 412514 272944
rect 453942 272932 453948 272944
rect 412508 272904 453948 272932
rect 412508 272892 412514 272904
rect 453942 272892 453948 272904
rect 454000 272892 454006 272944
rect 458082 272892 458088 272944
rect 458140 272932 458146 272944
rect 521838 272932 521844 272944
rect 458140 272904 521844 272932
rect 458140 272892 458146 272904
rect 521838 272892 521844 272904
rect 521896 272892 521902 272944
rect 524368 272932 524374 272944
rect 523604 272904 524374 272932
rect 394510 272796 394516 272808
rect 380768 272768 383654 272796
rect 388456 272768 394516 272796
rect 380768 272756 380774 272768
rect 87138 272620 87144 272672
rect 87196 272660 87202 272672
rect 151998 272660 152004 272672
rect 87196 272632 152004 272660
rect 87196 272620 87202 272632
rect 151998 272620 152004 272632
rect 152056 272620 152062 272672
rect 168650 272620 168656 272672
rect 168708 272660 168714 272672
rect 208486 272660 208492 272672
rect 168708 272632 208492 272660
rect 168708 272620 168714 272632
rect 208486 272620 208492 272632
rect 208544 272620 208550 272672
rect 217410 272620 217416 272672
rect 217468 272660 217474 272672
rect 242158 272660 242164 272672
rect 217468 272632 242164 272660
rect 217468 272620 217474 272632
rect 242158 272620 242164 272632
rect 242216 272620 242222 272672
rect 242342 272620 242348 272672
rect 242400 272660 242406 272672
rect 259546 272660 259552 272672
rect 242400 272632 259552 272660
rect 242400 272620 242406 272632
rect 259546 272620 259552 272632
rect 259604 272620 259610 272672
rect 331030 272620 331036 272672
rect 331088 272660 331094 272672
rect 342438 272660 342444 272672
rect 331088 272632 342444 272660
rect 331088 272620 331094 272632
rect 342438 272620 342444 272632
rect 342496 272620 342502 272672
rect 368382 272620 368388 272672
rect 368440 272660 368446 272672
rect 388456 272660 388484 272768
rect 394510 272756 394516 272768
rect 394568 272756 394574 272808
rect 397270 272756 397276 272808
rect 397328 272796 397334 272808
rect 418338 272796 418344 272808
rect 397328 272768 418344 272796
rect 397328 272756 397334 272768
rect 418338 272756 418344 272768
rect 418396 272756 418402 272808
rect 426066 272756 426072 272808
rect 426124 272796 426130 272808
rect 478414 272796 478420 272808
rect 426124 272768 478420 272796
rect 426124 272756 426130 272768
rect 478414 272756 478420 272768
rect 478472 272756 478478 272808
rect 482738 272756 482744 272808
rect 482796 272796 482802 272808
rect 523604 272796 523632 272904
rect 524368 272892 524374 272904
rect 524426 272892 524432 272944
rect 524506 272892 524512 272944
rect 524564 272932 524570 272944
rect 611354 272932 611360 272944
rect 524564 272904 611360 272932
rect 524564 272892 524570 272904
rect 611354 272892 611360 272904
rect 611412 272892 611418 272944
rect 606110 272796 606116 272808
rect 482796 272768 523632 272796
rect 523696 272768 606116 272796
rect 482796 272756 482802 272768
rect 368440 272632 388484 272660
rect 368440 272620 368446 272632
rect 388622 272620 388628 272672
rect 388680 272660 388686 272672
rect 393590 272660 393596 272672
rect 388680 272632 393596 272660
rect 388680 272620 388686 272632
rect 393590 272620 393596 272632
rect 393648 272620 393654 272672
rect 393958 272620 393964 272672
rect 394016 272660 394022 272672
rect 406286 272660 406292 272672
rect 394016 272632 406292 272660
rect 394016 272620 394022 272632
rect 406286 272620 406292 272632
rect 406344 272620 406350 272672
rect 408402 272620 408408 272672
rect 408460 272660 408466 272672
rect 452470 272660 452476 272672
rect 408460 272632 452476 272660
rect 408460 272620 408466 272632
rect 452470 272620 452476 272632
rect 452528 272620 452534 272672
rect 453850 272620 453856 272672
rect 453908 272660 453914 272672
rect 516410 272660 516416 272672
rect 453908 272632 516416 272660
rect 453908 272620 453914 272632
rect 516410 272620 516416 272632
rect 516468 272620 516474 272672
rect 516594 272620 516600 272672
rect 516652 272660 516658 272672
rect 523696 272660 523724 272768
rect 606110 272756 606116 272768
rect 606168 272756 606174 272808
rect 516652 272632 523724 272660
rect 516652 272620 516658 272632
rect 524322 272620 524328 272672
rect 524380 272660 524386 272672
rect 524506 272660 524512 272672
rect 524380 272632 524512 272660
rect 524380 272620 524386 272632
rect 524506 272620 524512 272632
rect 524564 272620 524570 272672
rect 524874 272620 524880 272672
rect 524932 272660 524938 272672
rect 614390 272660 614396 272672
rect 524932 272632 614396 272660
rect 524932 272620 524938 272632
rect 614390 272620 614396 272632
rect 614448 272620 614454 272672
rect 77662 272484 77668 272536
rect 77720 272524 77726 272536
rect 145098 272524 145104 272536
rect 77720 272496 145104 272524
rect 77720 272484 77726 272496
rect 145098 272484 145104 272496
rect 145156 272484 145162 272536
rect 152182 272484 152188 272536
rect 152240 272524 152246 272536
rect 197538 272524 197544 272536
rect 152240 272496 197544 272524
rect 152240 272484 152246 272496
rect 197538 272484 197544 272496
rect 197596 272484 197602 272536
rect 199470 272484 199476 272536
rect 199528 272524 199534 272536
rect 230566 272524 230572 272536
rect 199528 272496 230572 272524
rect 199528 272484 199534 272496
rect 230566 272484 230572 272496
rect 230624 272484 230630 272536
rect 231394 272484 231400 272536
rect 231452 272524 231458 272536
rect 252738 272524 252744 272536
rect 231452 272496 252744 272524
rect 231452 272484 231458 272496
rect 252738 272484 252744 272496
rect 252796 272484 252802 272536
rect 252922 272484 252928 272536
rect 252980 272524 252986 272536
rect 267734 272524 267740 272536
rect 252980 272496 267740 272524
rect 252980 272484 252986 272496
rect 267734 272484 267740 272496
rect 267792 272484 267798 272536
rect 268010 272484 268016 272536
rect 268068 272524 268074 272536
rect 278774 272524 278780 272536
rect 268068 272496 278780 272524
rect 268068 272484 268074 272496
rect 278774 272484 278780 272496
rect 278832 272484 278838 272536
rect 279786 272484 279792 272536
rect 279844 272524 279850 272536
rect 287146 272524 287152 272536
rect 279844 272496 287152 272524
rect 279844 272484 279850 272496
rect 287146 272484 287152 272496
rect 287204 272484 287210 272536
rect 338022 272484 338028 272536
rect 338080 272524 338086 272536
rect 351914 272524 351920 272536
rect 338080 272496 351920 272524
rect 338080 272484 338086 272496
rect 351914 272484 351920 272496
rect 351972 272484 351978 272536
rect 358630 272484 358636 272536
rect 358688 272524 358694 272536
rect 380342 272524 380348 272536
rect 358688 272496 380348 272524
rect 358688 272484 358694 272496
rect 380342 272484 380348 272496
rect 380400 272484 380406 272536
rect 380526 272484 380532 272536
rect 380584 272524 380590 272536
rect 413370 272524 413376 272536
rect 380584 272496 413376 272524
rect 380584 272484 380590 272496
rect 413370 272484 413376 272496
rect 413428 272484 413434 272536
rect 415118 272484 415124 272536
rect 415176 272524 415182 272536
rect 461854 272524 461860 272536
rect 415176 272496 461860 272524
rect 415176 272484 415182 272496
rect 461854 272484 461860 272496
rect 461912 272484 461918 272536
rect 463510 272484 463516 272536
rect 463568 272524 463574 272536
rect 524598 272524 524604 272536
rect 463568 272496 524604 272524
rect 463568 272484 463574 272496
rect 524598 272484 524604 272496
rect 524656 272484 524662 272536
rect 525058 272484 525064 272536
rect 525116 272524 525122 272536
rect 533982 272524 533988 272536
rect 525116 272496 533988 272524
rect 525116 272484 525122 272496
rect 533982 272484 533988 272496
rect 534040 272484 534046 272536
rect 534166 272484 534172 272536
rect 534224 272524 534230 272536
rect 632146 272524 632152 272536
rect 534224 272496 632152 272524
rect 534224 272484 534230 272496
rect 632146 272484 632152 272496
rect 632204 272484 632210 272536
rect 127342 272348 127348 272400
rect 127400 272388 127406 272400
rect 179874 272388 179880 272400
rect 127400 272360 179880 272388
rect 127400 272348 127406 272360
rect 179874 272348 179880 272360
rect 179932 272348 179938 272400
rect 439314 272348 439320 272400
rect 439372 272388 439378 272400
rect 473722 272388 473728 272400
rect 439372 272360 473728 272388
rect 439372 272348 439378 272360
rect 473722 272348 473728 272360
rect 473780 272348 473786 272400
rect 474642 272348 474648 272400
rect 474700 272388 474706 272400
rect 495434 272388 495440 272400
rect 474700 272360 495440 272388
rect 474700 272348 474706 272360
rect 495434 272348 495440 272360
rect 495492 272348 495498 272400
rect 501598 272348 501604 272400
rect 501656 272388 501662 272400
rect 581270 272388 581276 272400
rect 501656 272360 581276 272388
rect 501656 272348 501662 272360
rect 581270 272348 581276 272360
rect 581328 272348 581334 272400
rect 139118 272212 139124 272264
rect 139176 272252 139182 272264
rect 141602 272252 141608 272264
rect 139176 272224 141608 272252
rect 139176 272212 139182 272224
rect 141602 272212 141608 272224
rect 141660 272212 141666 272264
rect 143902 272212 143908 272264
rect 143960 272252 143966 272264
rect 190730 272252 190736 272264
rect 143960 272224 190736 272252
rect 143960 272212 143966 272224
rect 190730 272212 190736 272224
rect 190788 272212 190794 272264
rect 451734 272212 451740 272264
rect 451792 272252 451798 272264
rect 480806 272252 480812 272264
rect 451792 272224 480812 272252
rect 451792 272212 451798 272224
rect 480806 272212 480812 272224
rect 480864 272212 480870 272264
rect 488350 272212 488356 272264
rect 488408 272252 488414 272264
rect 567102 272252 567108 272264
rect 488408 272224 567108 272252
rect 488408 272212 488414 272224
rect 567102 272212 567108 272224
rect 567160 272212 567166 272264
rect 153286 272076 153292 272128
rect 153344 272116 153350 272128
rect 171778 272116 171784 272128
rect 153344 272088 171784 272116
rect 153344 272076 153350 272088
rect 171778 272076 171784 272088
rect 171836 272076 171842 272128
rect 473078 272076 473084 272128
rect 473136 272116 473142 272128
rect 482922 272116 482928 272128
rect 473136 272088 482928 272116
rect 473136 272076 473142 272088
rect 482922 272076 482928 272088
rect 482980 272076 482986 272128
rect 483750 272076 483756 272128
rect 483808 272116 483814 272128
rect 560018 272116 560024 272128
rect 483808 272088 560024 272116
rect 483808 272076 483814 272088
rect 560018 272076 560024 272088
rect 560076 272076 560082 272128
rect 478690 271940 478696 271992
rect 478748 271980 478754 271992
rect 552474 271980 552480 271992
rect 478748 271952 552480 271980
rect 478748 271940 478754 271952
rect 552474 271940 552480 271952
rect 552532 271940 552538 271992
rect 552842 271940 552848 271992
rect 552900 271980 552906 271992
rect 580074 271980 580080 271992
rect 552900 271952 580080 271980
rect 552900 271940 552906 271952
rect 580074 271940 580080 271952
rect 580132 271940 580138 271992
rect 110414 271804 110420 271856
rect 110472 271844 110478 271856
rect 164970 271844 164976 271856
rect 110472 271816 164976 271844
rect 110472 271804 110478 271816
rect 164970 271804 164976 271816
rect 165028 271804 165034 271856
rect 175826 271804 175832 271856
rect 175884 271844 175890 271856
rect 207658 271844 207664 271856
rect 175884 271816 207664 271844
rect 175884 271804 175890 271816
rect 207658 271804 207664 271816
rect 207716 271804 207722 271856
rect 214834 271804 214840 271856
rect 214892 271844 214898 271856
rect 221458 271844 221464 271856
rect 214892 271816 221464 271844
rect 214892 271804 214898 271816
rect 221458 271804 221464 271816
rect 221516 271804 221522 271856
rect 222102 271804 222108 271856
rect 222160 271844 222166 271856
rect 232130 271844 232136 271856
rect 222160 271816 232136 271844
rect 222160 271804 222166 271816
rect 232130 271804 232136 271816
rect 232188 271804 232194 271856
rect 356514 271804 356520 271856
rect 356572 271844 356578 271856
rect 358998 271844 359004 271856
rect 356572 271816 359004 271844
rect 356572 271804 356578 271816
rect 358998 271804 359004 271816
rect 359056 271804 359062 271856
rect 394326 271804 394332 271856
rect 394384 271844 394390 271856
rect 426250 271844 426256 271856
rect 394384 271816 426256 271844
rect 394384 271804 394390 271816
rect 426250 271804 426256 271816
rect 426308 271804 426314 271856
rect 427078 271804 427084 271856
rect 427136 271844 427142 271856
rect 433518 271844 433524 271856
rect 427136 271816 433524 271844
rect 427136 271804 427142 271816
rect 433518 271804 433524 271816
rect 433576 271804 433582 271856
rect 447778 271804 447784 271856
rect 447836 271844 447842 271856
rect 503990 271844 503996 271856
rect 447836 271816 503996 271844
rect 447836 271804 447842 271816
rect 503990 271804 503996 271816
rect 504048 271804 504054 271856
rect 504726 271804 504732 271856
rect 504784 271844 504790 271856
rect 589550 271844 589556 271856
rect 504784 271816 589556 271844
rect 504784 271804 504790 271816
rect 589550 271804 589556 271816
rect 589608 271804 589614 271856
rect 596634 271844 596640 271856
rect 591316 271816 596640 271844
rect 318610 271736 318616 271788
rect 318668 271776 318674 271788
rect 324774 271776 324780 271788
rect 318668 271748 324780 271776
rect 318668 271736 318674 271748
rect 324774 271736 324780 271748
rect 324832 271736 324838 271788
rect 93026 271668 93032 271720
rect 93084 271708 93090 271720
rect 120718 271708 120724 271720
rect 93084 271680 120724 271708
rect 93084 271668 93090 271680
rect 120718 271668 120724 271680
rect 120776 271668 120782 271720
rect 120902 271668 120908 271720
rect 120960 271708 120966 271720
rect 175274 271708 175280 271720
rect 120960 271680 175280 271708
rect 120960 271668 120966 271680
rect 175274 271668 175280 271680
rect 175332 271668 175338 271720
rect 192294 271668 192300 271720
rect 192352 271708 192358 271720
rect 225506 271708 225512 271720
rect 192352 271680 225512 271708
rect 192352 271668 192358 271680
rect 225506 271668 225512 271680
rect 225564 271668 225570 271720
rect 237466 271668 237472 271720
rect 237524 271708 237530 271720
rect 243722 271708 243728 271720
rect 237524 271680 243728 271708
rect 237524 271668 237530 271680
rect 243722 271668 243728 271680
rect 243780 271668 243786 271720
rect 355318 271668 355324 271720
rect 355376 271708 355382 271720
rect 374362 271708 374368 271720
rect 355376 271680 374368 271708
rect 355376 271668 355382 271680
rect 374362 271668 374368 271680
rect 374420 271668 374426 271720
rect 387702 271668 387708 271720
rect 387760 271708 387766 271720
rect 421374 271708 421380 271720
rect 387760 271680 421380 271708
rect 387760 271668 387766 271680
rect 421374 271668 421380 271680
rect 421432 271668 421438 271720
rect 421742 271668 421748 271720
rect 421800 271708 421806 271720
rect 438210 271708 438216 271720
rect 421800 271680 438216 271708
rect 421800 271668 421806 271680
rect 438210 271668 438216 271680
rect 438268 271668 438274 271720
rect 442902 271668 442908 271720
rect 442960 271708 442966 271720
rect 500494 271708 500500 271720
rect 442960 271680 500500 271708
rect 442960 271668 442966 271680
rect 500494 271668 500500 271680
rect 500552 271668 500558 271720
rect 500862 271668 500868 271720
rect 500920 271708 500926 271720
rect 508038 271708 508044 271720
rect 500920 271680 508044 271708
rect 500920 271668 500926 271680
rect 508038 271668 508044 271680
rect 508096 271668 508102 271720
rect 508958 271668 508964 271720
rect 509016 271708 509022 271720
rect 591316 271708 591344 271816
rect 596634 271804 596640 271816
rect 596692 271804 596698 271856
rect 509016 271680 591344 271708
rect 509016 271668 509022 271680
rect 591482 271668 591488 271720
rect 591540 271708 591546 271720
rect 603718 271708 603724 271720
rect 591540 271680 603724 271708
rect 591540 271668 591546 271680
rect 603718 271668 603724 271680
rect 603776 271668 603782 271720
rect 111978 271532 111984 271584
rect 112036 271572 112042 271584
rect 168374 271572 168380 271584
rect 112036 271544 168380 271572
rect 112036 271532 112042 271544
rect 168374 271532 168380 271544
rect 168432 271532 168438 271584
rect 173434 271532 173440 271584
rect 173492 271572 173498 271584
rect 212626 271572 212632 271584
rect 173492 271544 212632 271572
rect 173492 271532 173498 271544
rect 212626 271532 212632 271544
rect 212684 271532 212690 271584
rect 226150 271532 226156 271584
rect 226208 271572 226214 271584
rect 247126 271572 247132 271584
rect 226208 271544 247132 271572
rect 226208 271532 226214 271544
rect 247126 271532 247132 271544
rect 247184 271532 247190 271584
rect 259730 271532 259736 271584
rect 259788 271572 259794 271584
rect 272610 271572 272616 271584
rect 259788 271544 272616 271572
rect 259788 271532 259794 271544
rect 272610 271532 272616 271544
rect 272668 271532 272674 271584
rect 372522 271532 372528 271584
rect 372580 271572 372586 271584
rect 400398 271572 400404 271584
rect 372580 271544 400404 271572
rect 372580 271532 372586 271544
rect 400398 271532 400404 271544
rect 400456 271532 400462 271584
rect 409782 271532 409788 271584
rect 409840 271572 409846 271584
rect 443730 271572 443736 271584
rect 409840 271544 443736 271572
rect 409840 271532 409846 271544
rect 443730 271532 443736 271544
rect 443788 271532 443794 271584
rect 453298 271532 453304 271584
rect 453356 271572 453362 271584
rect 511534 271572 511540 271584
rect 453356 271544 511540 271572
rect 453356 271532 453362 271544
rect 511534 271532 511540 271544
rect 511592 271532 511598 271584
rect 511902 271532 511908 271584
rect 511960 271572 511966 271584
rect 600222 271572 600228 271584
rect 511960 271544 600228 271572
rect 511960 271532 511966 271544
rect 600222 271532 600228 271544
rect 600280 271532 600286 271584
rect 607858 271532 607864 271584
rect 607916 271572 607922 271584
rect 643922 271572 643928 271584
rect 607916 271544 643928 271572
rect 607916 271532 607922 271544
rect 643922 271532 643928 271544
rect 643980 271532 643986 271584
rect 89714 271396 89720 271448
rect 89772 271436 89778 271448
rect 152642 271436 152648 271448
rect 89772 271408 152648 271436
rect 89772 271396 89778 271408
rect 152642 271396 152648 271408
rect 152700 271396 152706 271448
rect 165154 271396 165160 271448
rect 165212 271436 165218 271448
rect 205726 271436 205732 271448
rect 165212 271408 205732 271436
rect 165212 271396 165218 271408
rect 205726 271396 205732 271408
rect 205784 271396 205790 271448
rect 223574 271396 223580 271448
rect 223632 271436 223638 271448
rect 247310 271436 247316 271448
rect 223632 271408 247316 271436
rect 223632 271396 223638 271408
rect 247310 271396 247316 271408
rect 247368 271396 247374 271448
rect 247862 271396 247868 271448
rect 247920 271436 247926 271448
rect 264330 271436 264336 271448
rect 247920 271408 264336 271436
rect 247920 271396 247926 271408
rect 264330 271396 264336 271408
rect 264388 271396 264394 271448
rect 334618 271396 334624 271448
rect 334676 271436 334682 271448
rect 341334 271436 341340 271448
rect 334676 271408 341340 271436
rect 334676 271396 334682 271408
rect 341334 271396 341340 271408
rect 341392 271396 341398 271448
rect 342162 271396 342168 271448
rect 342220 271436 342226 271448
rect 356698 271436 356704 271448
rect 342220 271408 356704 271436
rect 342220 271396 342226 271408
rect 356698 271396 356704 271408
rect 356756 271396 356762 271448
rect 360838 271396 360844 271448
rect 360896 271436 360902 271448
rect 381538 271436 381544 271448
rect 360896 271408 381544 271436
rect 360896 271396 360902 271408
rect 381538 271396 381544 271408
rect 381596 271396 381602 271448
rect 398098 271396 398104 271448
rect 398156 271436 398162 271448
rect 427078 271436 427084 271448
rect 398156 271408 427084 271436
rect 398156 271396 398162 271408
rect 427078 271396 427084 271408
rect 427136 271396 427142 271448
rect 427262 271396 427268 271448
rect 427320 271436 427326 271448
rect 427320 271408 436784 271436
rect 427320 271396 427326 271408
rect 68186 271260 68192 271312
rect 68244 271300 68250 271312
rect 138474 271300 138480 271312
rect 68244 271272 138480 271300
rect 68244 271260 68250 271272
rect 138474 271260 138480 271272
rect 138532 271260 138538 271312
rect 150986 271260 150992 271312
rect 151044 271300 151050 271312
rect 195974 271300 195980 271312
rect 151044 271272 195980 271300
rect 151044 271260 151050 271272
rect 195974 271260 195980 271272
rect 196032 271260 196038 271312
rect 215938 271260 215944 271312
rect 215996 271300 216002 271312
rect 242066 271300 242072 271312
rect 215996 271272 242072 271300
rect 215996 271260 216002 271272
rect 242066 271260 242072 271272
rect 242124 271260 242130 271312
rect 243170 271260 243176 271312
rect 243228 271300 243234 271312
rect 261018 271300 261024 271312
rect 243228 271272 261024 271300
rect 243228 271260 243234 271272
rect 261018 271260 261024 271272
rect 261076 271260 261082 271312
rect 275094 271260 275100 271312
rect 275152 271300 275158 271312
rect 283466 271300 283472 271312
rect 275152 271272 283472 271300
rect 275152 271260 275158 271272
rect 283466 271260 283472 271272
rect 283524 271260 283530 271312
rect 315758 271260 315764 271312
rect 315816 271300 315822 271312
rect 319990 271300 319996 271312
rect 315816 271272 319996 271300
rect 315816 271260 315822 271272
rect 319990 271260 319996 271272
rect 320048 271260 320054 271312
rect 325510 271260 325516 271312
rect 325568 271300 325574 271312
rect 334158 271300 334164 271312
rect 325568 271272 334164 271300
rect 325568 271260 325574 271272
rect 334158 271260 334164 271272
rect 334216 271260 334222 271312
rect 340598 271260 340604 271312
rect 340656 271300 340662 271312
rect 355502 271300 355508 271312
rect 340656 271272 355508 271300
rect 340656 271260 340662 271272
rect 355502 271260 355508 271272
rect 355560 271260 355566 271312
rect 364150 271260 364156 271312
rect 364208 271300 364214 271312
rect 386046 271300 386052 271312
rect 364208 271272 386052 271300
rect 364208 271260 364214 271272
rect 386046 271260 386052 271272
rect 386104 271260 386110 271312
rect 400122 271260 400128 271312
rect 400180 271300 400186 271312
rect 435634 271300 435640 271312
rect 400180 271272 435640 271300
rect 400180 271260 400186 271272
rect 435634 271260 435640 271272
rect 435692 271260 435698 271312
rect 436756 271300 436784 271408
rect 436922 271396 436928 271448
rect 436980 271436 436986 271448
rect 454770 271436 454776 271448
rect 436980 271408 454776 271436
rect 436980 271396 436986 271408
rect 454770 271396 454776 271408
rect 454828 271396 454834 271448
rect 457438 271396 457444 271448
rect 457496 271436 457502 271448
rect 511718 271436 511724 271448
rect 457496 271408 511724 271436
rect 457496 271396 457502 271408
rect 511718 271396 511724 271408
rect 511776 271396 511782 271448
rect 515122 271436 515128 271448
rect 512196 271408 515128 271436
rect 448882 271300 448888 271312
rect 436756 271272 448888 271300
rect 448882 271260 448888 271272
rect 448940 271260 448946 271312
rect 454678 271260 454684 271312
rect 454736 271300 454742 271312
rect 512196 271300 512224 271408
rect 515122 271396 515128 271408
rect 515180 271396 515186 271448
rect 515306 271396 515312 271448
rect 515364 271436 515370 271448
rect 518618 271436 518624 271448
rect 515364 271408 518624 271436
rect 515364 271396 515370 271408
rect 518618 271396 518624 271408
rect 518676 271396 518682 271448
rect 520090 271396 520096 271448
rect 520148 271436 520154 271448
rect 523954 271436 523960 271448
rect 520148 271408 523960 271436
rect 520148 271396 520154 271408
rect 523954 271396 523960 271408
rect 524012 271396 524018 271448
rect 524138 271396 524144 271448
rect 524196 271436 524202 271448
rect 524196 271408 529244 271436
rect 524196 271396 524202 271408
rect 454736 271272 512224 271300
rect 454736 271260 454742 271272
rect 514478 271260 514484 271312
rect 514536 271300 514542 271312
rect 529014 271300 529020 271312
rect 514536 271272 529020 271300
rect 514536 271260 514542 271272
rect 529014 271260 529020 271272
rect 529072 271260 529078 271312
rect 529216 271300 529244 271408
rect 529382 271396 529388 271448
rect 529440 271436 529446 271448
rect 610802 271436 610808 271448
rect 529440 271408 610808 271436
rect 529440 271396 529446 271408
rect 610802 271396 610808 271408
rect 610860 271396 610866 271448
rect 617978 271300 617984 271312
rect 529216 271272 617984 271300
rect 617978 271260 617984 271272
rect 618036 271260 618042 271312
rect 72970 271124 72976 271176
rect 73028 271164 73034 271176
rect 142154 271164 142160 271176
rect 73028 271136 142160 271164
rect 73028 271124 73034 271136
rect 142154 271124 142160 271136
rect 142212 271124 142218 271176
rect 148594 271124 148600 271176
rect 148652 271164 148658 271176
rect 194778 271164 194784 271176
rect 148652 271136 194784 271164
rect 148652 271124 148658 271136
rect 194778 271124 194784 271136
rect 194836 271124 194842 271176
rect 208854 271124 208860 271176
rect 208912 271164 208918 271176
rect 237466 271164 237472 271176
rect 208912 271136 237472 271164
rect 208912 271124 208918 271136
rect 237466 271124 237472 271136
rect 237524 271124 237530 271176
rect 240778 271124 240784 271176
rect 240836 271164 240842 271176
rect 259822 271164 259828 271176
rect 240836 271136 259828 271164
rect 240836 271124 240842 271136
rect 259822 271124 259828 271136
rect 259880 271124 259886 271176
rect 262122 271124 262128 271176
rect 262180 271164 262186 271176
rect 274634 271164 274640 271176
rect 262180 271136 274640 271164
rect 262180 271124 262186 271136
rect 274634 271124 274640 271136
rect 274692 271124 274698 271176
rect 276290 271124 276296 271176
rect 276348 271164 276354 271176
rect 284478 271164 284484 271176
rect 276348 271136 284484 271164
rect 276348 271124 276354 271136
rect 284478 271124 284484 271136
rect 284536 271124 284542 271176
rect 333882 271124 333888 271176
rect 333940 271164 333946 271176
rect 344462 271164 344468 271176
rect 333940 271136 344468 271164
rect 333940 271124 333946 271136
rect 344462 271124 344468 271136
rect 344520 271124 344526 271176
rect 344646 271124 344652 271176
rect 344704 271164 344710 271176
rect 350718 271164 350724 271176
rect 344704 271136 350724 271164
rect 344704 271124 344710 271136
rect 350718 271124 350724 271136
rect 350776 271124 350782 271176
rect 351822 271124 351828 271176
rect 351880 271164 351886 271176
rect 372062 271164 372068 271176
rect 351880 271136 372068 271164
rect 351880 271124 351886 271136
rect 372062 271124 372068 271136
rect 372120 271124 372126 271176
rect 379422 271124 379428 271176
rect 379480 271164 379486 271176
rect 407114 271164 407120 271176
rect 379480 271136 407120 271164
rect 379480 271124 379486 271136
rect 407114 271124 407120 271136
rect 407172 271124 407178 271176
rect 416590 271124 416596 271176
rect 416648 271164 416654 271176
rect 463970 271164 463976 271176
rect 416648 271136 463976 271164
rect 416648 271124 416654 271136
rect 463970 271124 463976 271136
rect 464028 271124 464034 271176
rect 464522 271124 464528 271176
rect 464580 271164 464586 271176
rect 524598 271164 524604 271176
rect 464580 271136 524604 271164
rect 464580 271124 464586 271136
rect 524598 271124 524604 271136
rect 524656 271124 524662 271176
rect 524782 271124 524788 271176
rect 524840 271164 524846 271176
rect 529382 271164 529388 271176
rect 524840 271136 529388 271164
rect 524840 271124 524846 271136
rect 529382 271124 529388 271136
rect 529440 271124 529446 271176
rect 529566 271124 529572 271176
rect 529624 271164 529630 271176
rect 532786 271164 532792 271176
rect 529624 271136 532792 271164
rect 529624 271124 529630 271136
rect 532786 271124 532792 271136
rect 532844 271124 532850 271176
rect 533154 271124 533160 271176
rect 533212 271164 533218 271176
rect 621474 271164 621480 271176
rect 533212 271136 621480 271164
rect 533212 271124 533218 271136
rect 621474 271124 621480 271136
rect 621532 271124 621538 271176
rect 621658 271124 621664 271176
rect 621716 271164 621722 271176
rect 636838 271164 636844 271176
rect 621716 271136 636844 271164
rect 621716 271124 621722 271136
rect 636838 271124 636844 271136
rect 636896 271124 636902 271176
rect 128538 270988 128544 271040
rect 128596 271028 128602 271040
rect 181346 271028 181352 271040
rect 128596 271000 181352 271028
rect 128596 270988 128602 271000
rect 181346 270988 181352 271000
rect 181404 270988 181410 271040
rect 189994 270988 190000 271040
rect 190052 271028 190058 271040
rect 216122 271028 216128 271040
rect 190052 271000 216128 271028
rect 190052 270988 190058 271000
rect 216122 270988 216128 271000
rect 216180 270988 216186 271040
rect 381538 270988 381544 271040
rect 381596 271028 381602 271040
rect 399202 271028 399208 271040
rect 381596 271000 399208 271028
rect 381596 270988 381602 271000
rect 399202 270988 399208 271000
rect 399260 270988 399266 271040
rect 401318 270988 401324 271040
rect 401376 271028 401382 271040
rect 401376 271000 422294 271028
rect 401376 270988 401382 271000
rect 130838 270852 130844 270904
rect 130896 270892 130902 270904
rect 182450 270892 182456 270904
rect 130896 270864 182456 270892
rect 130896 270852 130902 270864
rect 182450 270852 182456 270864
rect 182508 270852 182514 270904
rect 200482 270852 200488 270904
rect 200540 270892 200546 270904
rect 224218 270892 224224 270904
rect 200540 270864 224224 270892
rect 200540 270852 200546 270864
rect 224218 270852 224224 270864
rect 224276 270852 224282 270904
rect 389082 270852 389088 270904
rect 389140 270892 389146 270904
rect 415302 270892 415308 270904
rect 389140 270864 415308 270892
rect 389140 270852 389146 270864
rect 415302 270852 415308 270864
rect 415360 270852 415366 270904
rect 422266 270892 422294 271000
rect 425698 270988 425704 271040
rect 425756 271028 425762 271040
rect 427262 271028 427268 271040
rect 425756 271000 427268 271028
rect 425756 270988 425762 271000
rect 427262 270988 427268 271000
rect 427320 270988 427326 271040
rect 431678 270988 431684 271040
rect 431736 271028 431742 271040
rect 485498 271028 485504 271040
rect 431736 271000 485504 271028
rect 431736 270988 431742 271000
rect 485498 270988 485504 271000
rect 485556 270988 485562 271040
rect 488534 270988 488540 271040
rect 488592 271028 488598 271040
rect 551738 271028 551744 271040
rect 488592 271000 551744 271028
rect 488592 270988 488598 271000
rect 551738 270988 551744 271000
rect 551796 270988 551802 271040
rect 552658 270988 552664 271040
rect 552716 271028 552722 271040
rect 591482 271028 591488 271040
rect 552716 271000 591488 271028
rect 552716 270988 552722 271000
rect 591482 270988 591488 271000
rect 591540 270988 591546 271040
rect 427814 270892 427820 270904
rect 422266 270864 427820 270892
rect 427814 270852 427820 270864
rect 427872 270852 427878 270904
rect 435358 270852 435364 270904
rect 435416 270892 435422 270904
rect 436922 270892 436928 270904
rect 435416 270864 436928 270892
rect 435416 270852 435422 270864
rect 436922 270852 436928 270864
rect 436980 270852 436986 270904
rect 445018 270852 445024 270904
rect 445076 270892 445082 270904
rect 497366 270892 497372 270904
rect 445076 270864 497372 270892
rect 445076 270852 445082 270864
rect 497366 270852 497372 270864
rect 497424 270852 497430 270904
rect 507670 270852 507676 270904
rect 507728 270892 507734 270904
rect 523954 270892 523960 270904
rect 507728 270864 523960 270892
rect 507728 270852 507734 270864
rect 523954 270852 523960 270864
rect 524012 270852 524018 270904
rect 524874 270852 524880 270904
rect 524932 270892 524938 270904
rect 593138 270892 593144 270904
rect 524932 270864 593144 270892
rect 524932 270852 524938 270864
rect 593138 270852 593144 270864
rect 593196 270852 593202 270904
rect 137922 270716 137928 270768
rect 137980 270756 137986 270768
rect 187878 270756 187884 270768
rect 137980 270728 187884 270756
rect 137980 270716 137986 270728
rect 187878 270716 187884 270728
rect 187936 270716 187942 270768
rect 433150 270716 433156 270768
rect 433208 270756 433214 270768
rect 456978 270756 456984 270768
rect 433208 270728 456984 270756
rect 433208 270716 433214 270728
rect 456978 270716 456984 270728
rect 457036 270716 457042 270768
rect 465718 270716 465724 270768
rect 465776 270756 465782 270768
rect 526254 270756 526260 270768
rect 465776 270728 526260 270756
rect 465776 270716 465782 270728
rect 526254 270716 526260 270728
rect 526312 270716 526318 270768
rect 526438 270716 526444 270768
rect 526496 270756 526502 270768
rect 528646 270756 528652 270768
rect 526496 270728 528652 270756
rect 526496 270716 526502 270728
rect 528646 270716 528652 270728
rect 528704 270716 528710 270768
rect 529014 270716 529020 270768
rect 529072 270756 529078 270768
rect 529072 270728 539088 270756
rect 529072 270716 529078 270728
rect 116670 270580 116676 270632
rect 116728 270620 116734 270632
rect 151078 270620 151084 270632
rect 116728 270592 151084 270620
rect 116728 270580 116734 270592
rect 151078 270580 151084 270592
rect 151136 270580 151142 270632
rect 237282 270580 237288 270632
rect 237340 270620 237346 270632
rect 237340 270592 237512 270620
rect 237340 270580 237346 270592
rect 115842 270444 115848 270496
rect 115900 270484 115906 270496
rect 171226 270484 171232 270496
rect 115900 270456 171232 270484
rect 115900 270444 115906 270456
rect 171226 270444 171232 270456
rect 171284 270444 171290 270496
rect 172422 270444 172428 270496
rect 172480 270484 172486 270496
rect 208670 270484 208676 270496
rect 172480 270456 208676 270484
rect 172480 270444 172486 270456
rect 208670 270444 208676 270456
rect 208728 270444 208734 270496
rect 210786 270444 210792 270496
rect 210844 270484 210850 270496
rect 211798 270484 211804 270496
rect 210844 270456 211804 270484
rect 210844 270444 210850 270456
rect 211798 270444 211804 270456
rect 211856 270444 211862 270496
rect 233142 270444 233148 270496
rect 233200 270484 233206 270496
rect 237282 270484 237288 270496
rect 233200 270456 237288 270484
rect 233200 270444 233206 270456
rect 237282 270444 237288 270456
rect 237340 270444 237346 270496
rect 237484 270484 237512 270592
rect 428458 270580 428464 270632
rect 428516 270620 428522 270632
rect 466638 270620 466644 270632
rect 428516 270592 466644 270620
rect 428516 270580 428522 270592
rect 466638 270580 466644 270592
rect 466696 270580 466702 270632
rect 478138 270580 478144 270632
rect 478196 270620 478202 270632
rect 538858 270620 538864 270632
rect 478196 270592 538864 270620
rect 478196 270580 478202 270592
rect 538858 270580 538864 270592
rect 538916 270580 538922 270632
rect 539060 270620 539088 270728
rect 540514 270716 540520 270768
rect 540572 270756 540578 270768
rect 543550 270756 543556 270768
rect 540572 270728 543556 270756
rect 540572 270716 540578 270728
rect 543550 270716 543556 270728
rect 543608 270716 543614 270768
rect 543688 270716 543694 270768
rect 543746 270756 543752 270768
rect 607306 270756 607312 270768
rect 543746 270728 607312 270756
rect 543746 270716 543752 270728
rect 607306 270716 607312 270728
rect 607364 270716 607370 270768
rect 552658 270620 552664 270632
rect 539060 270592 552664 270620
rect 552658 270580 552664 270592
rect 552716 270580 552722 270632
rect 252002 270484 252008 270496
rect 237484 270456 252008 270484
rect 252002 270444 252008 270456
rect 252060 270444 252066 270496
rect 292850 270444 292856 270496
rect 292908 270484 292914 270496
rect 296254 270484 296260 270496
rect 292908 270456 296260 270484
rect 292908 270444 292914 270456
rect 296254 270444 296260 270456
rect 296312 270444 296318 270496
rect 358998 270444 359004 270496
rect 359056 270484 359062 270496
rect 376754 270484 376760 270496
rect 359056 270456 376760 270484
rect 359056 270444 359062 270456
rect 376754 270444 376760 270456
rect 376812 270444 376818 270496
rect 377582 270444 377588 270496
rect 377640 270484 377646 270496
rect 394694 270484 394700 270496
rect 377640 270456 394700 270484
rect 377640 270444 377646 270456
rect 394694 270444 394700 270456
rect 394752 270444 394758 270496
rect 396258 270444 396264 270496
rect 396316 270484 396322 270496
rect 423674 270484 423680 270496
rect 396316 270456 423680 270484
rect 396316 270444 396322 270456
rect 423674 270444 423680 270456
rect 423732 270444 423738 270496
rect 424594 270444 424600 270496
rect 424652 270484 424658 270496
rect 476298 270484 476304 270496
rect 424652 270456 476304 270484
rect 424652 270444 424658 270456
rect 476298 270444 476304 270456
rect 476356 270444 476362 270496
rect 479242 270444 479248 270496
rect 479300 270484 479306 270496
rect 552198 270484 552204 270496
rect 479300 270456 552204 270484
rect 479300 270444 479306 270456
rect 552198 270444 552204 270456
rect 552256 270444 552262 270496
rect 552382 270444 552388 270496
rect 552440 270484 552446 270496
rect 564434 270484 564440 270496
rect 552440 270456 564440 270484
rect 552440 270444 552446 270456
rect 564434 270444 564440 270456
rect 564492 270444 564498 270496
rect 110230 270308 110236 270360
rect 110288 270348 110294 270360
rect 167914 270348 167920 270360
rect 110288 270320 167920 270348
rect 110288 270308 110294 270320
rect 167914 270308 167920 270320
rect 167972 270308 167978 270360
rect 173066 270308 173072 270360
rect 173124 270348 173130 270360
rect 210142 270348 210148 270360
rect 173124 270320 210148 270348
rect 173124 270308 173130 270320
rect 210142 270308 210148 270320
rect 210200 270308 210206 270360
rect 212442 270308 212448 270360
rect 212500 270348 212506 270360
rect 239950 270348 239956 270360
rect 212500 270320 239956 270348
rect 212500 270308 212506 270320
rect 239950 270308 239956 270320
rect 240008 270308 240014 270360
rect 253842 270308 253848 270360
rect 253900 270348 253906 270360
rect 265066 270348 265072 270360
rect 253900 270320 265072 270348
rect 253900 270308 253906 270320
rect 265066 270308 265072 270320
rect 265124 270308 265130 270360
rect 291654 270308 291660 270360
rect 291712 270348 291718 270360
rect 295518 270348 295524 270360
rect 291712 270320 295524 270348
rect 291712 270308 291718 270320
rect 295518 270308 295524 270320
rect 295576 270308 295582 270360
rect 356698 270308 356704 270360
rect 356756 270348 356762 270360
rect 378134 270348 378140 270360
rect 356756 270320 378140 270348
rect 356756 270308 356762 270320
rect 378134 270308 378140 270320
rect 378192 270308 378198 270360
rect 385678 270308 385684 270360
rect 385736 270348 385742 270360
rect 419534 270348 419540 270360
rect 385736 270320 419540 270348
rect 385736 270308 385742 270320
rect 419534 270308 419540 270320
rect 419592 270308 419598 270360
rect 429562 270308 429568 270360
rect 429620 270348 429626 270360
rect 483106 270348 483112 270360
rect 429620 270320 483112 270348
rect 429620 270308 429626 270320
rect 483106 270308 483112 270320
rect 483164 270308 483170 270360
rect 486694 270308 486700 270360
rect 486752 270348 486758 270360
rect 494330 270348 494336 270360
rect 486752 270320 494336 270348
rect 486752 270308 486758 270320
rect 494330 270308 494336 270320
rect 494388 270308 494394 270360
rect 494514 270308 494520 270360
rect 494572 270348 494578 270360
rect 560294 270348 560300 270360
rect 494572 270320 560300 270348
rect 494572 270308 494578 270320
rect 560294 270308 560300 270320
rect 560352 270308 560358 270360
rect 316954 270240 316960 270292
rect 317012 270280 317018 270292
rect 321554 270280 321560 270292
rect 317012 270252 321560 270280
rect 317012 270240 317018 270252
rect 321554 270240 321560 270252
rect 321612 270240 321618 270292
rect 97902 270172 97908 270224
rect 97960 270212 97966 270224
rect 158806 270212 158812 270224
rect 97960 270184 158812 270212
rect 97960 270172 97966 270184
rect 158806 270172 158812 270184
rect 158864 270172 158870 270224
rect 166902 270172 166908 270224
rect 166960 270212 166966 270224
rect 207382 270212 207388 270224
rect 166960 270184 207388 270212
rect 166960 270172 166966 270184
rect 207382 270172 207388 270184
rect 207440 270172 207446 270224
rect 213822 270172 213828 270224
rect 213880 270212 213886 270224
rect 240502 270212 240508 270224
rect 213880 270184 240508 270212
rect 213880 270172 213886 270184
rect 240502 270172 240508 270184
rect 240560 270172 240566 270224
rect 249610 270172 249616 270224
rect 249668 270212 249674 270224
rect 263318 270212 263324 270224
rect 249668 270184 263324 270212
rect 249668 270172 249674 270184
rect 263318 270172 263324 270184
rect 263376 270172 263382 270224
rect 269206 270172 269212 270224
rect 269264 270212 269270 270224
rect 279694 270212 279700 270224
rect 269264 270184 279700 270212
rect 269264 270172 269270 270184
rect 279694 270172 279700 270184
rect 279752 270172 279758 270224
rect 321922 270172 321928 270224
rect 321980 270212 321986 270224
rect 328454 270212 328460 270224
rect 321980 270184 328460 270212
rect 321980 270172 321986 270184
rect 328454 270172 328460 270184
rect 328512 270172 328518 270224
rect 348418 270172 348424 270224
rect 348476 270212 348482 270224
rect 363046 270212 363052 270224
rect 348476 270184 363052 270212
rect 348476 270172 348482 270184
rect 363046 270172 363052 270184
rect 363104 270172 363110 270224
rect 364978 270172 364984 270224
rect 365036 270212 365042 270224
rect 390554 270212 390560 270224
rect 365036 270184 390560 270212
rect 365036 270172 365042 270184
rect 390554 270172 390560 270184
rect 390612 270172 390618 270224
rect 392302 270172 392308 270224
rect 392360 270212 392366 270224
rect 429378 270212 429384 270224
rect 392360 270184 429384 270212
rect 392360 270172 392366 270184
rect 429378 270172 429384 270184
rect 429436 270172 429442 270224
rect 446950 270172 446956 270224
rect 447008 270212 447014 270224
rect 504174 270212 504180 270224
rect 447008 270184 504180 270212
rect 447008 270172 447014 270184
rect 504174 270172 504180 270184
rect 504232 270172 504238 270224
rect 504358 270172 504364 270224
rect 504416 270212 504422 270224
rect 528462 270212 528468 270224
rect 504416 270184 528468 270212
rect 504416 270172 504422 270184
rect 528462 270172 528468 270184
rect 528520 270172 528526 270224
rect 533890 270212 533896 270224
rect 528848 270184 533896 270212
rect 309778 270104 309784 270156
rect 309836 270144 309842 270156
rect 311342 270144 311348 270156
rect 309836 270116 311348 270144
rect 309836 270104 309842 270116
rect 311342 270104 311348 270116
rect 311400 270104 311406 270156
rect 339310 270104 339316 270156
rect 339368 270144 339374 270156
rect 341518 270144 341524 270156
rect 339368 270116 341524 270144
rect 339368 270104 339374 270116
rect 341518 270104 341524 270116
rect 341576 270104 341582 270156
rect 80054 270036 80060 270088
rect 80112 270076 80118 270088
rect 146386 270076 146392 270088
rect 80112 270048 146392 270076
rect 80112 270036 80118 270048
rect 146386 270036 146392 270048
rect 146444 270036 146450 270088
rect 146754 270036 146760 270088
rect 146812 270076 146818 270088
rect 151354 270076 151360 270088
rect 146812 270048 151360 270076
rect 146812 270036 146818 270048
rect 151354 270036 151360 270048
rect 151412 270036 151418 270088
rect 153838 270076 153844 270088
rect 151786 270048 153844 270076
rect 75822 269900 75828 269952
rect 75880 269940 75886 269952
rect 142614 269940 142620 269952
rect 75880 269912 142620 269940
rect 75880 269900 75886 269912
rect 142614 269900 142620 269912
rect 142672 269900 142678 269952
rect 143350 269900 143356 269952
rect 143408 269940 143414 269952
rect 151786 269940 151814 270048
rect 153838 270036 153844 270048
rect 153896 270036 153902 270088
rect 159910 270036 159916 270088
rect 159968 270076 159974 270088
rect 202690 270076 202696 270088
rect 159968 270048 202696 270076
rect 159968 270036 159974 270048
rect 202690 270036 202696 270048
rect 202748 270036 202754 270088
rect 205542 270036 205548 270088
rect 205600 270076 205606 270088
rect 234982 270076 234988 270088
rect 205600 270048 234988 270076
rect 205600 270036 205606 270048
rect 234982 270036 234988 270048
rect 235040 270036 235046 270088
rect 239766 270036 239772 270088
rect 239824 270076 239830 270088
rect 253198 270076 253204 270088
rect 239824 270048 253204 270076
rect 239824 270036 239830 270048
rect 253198 270036 253204 270048
rect 253256 270036 253262 270088
rect 266170 270036 266176 270088
rect 266228 270076 266234 270088
rect 277210 270076 277216 270088
rect 266228 270048 277216 270076
rect 266228 270036 266234 270048
rect 277210 270036 277216 270048
rect 277268 270036 277274 270088
rect 323578 270036 323584 270088
rect 323636 270076 323642 270088
rect 331214 270076 331220 270088
rect 323636 270048 331220 270076
rect 323636 270036 323642 270048
rect 331214 270036 331220 270048
rect 331272 270036 331278 270088
rect 332318 270036 332324 270088
rect 332376 270076 332382 270088
rect 336734 270076 336740 270088
rect 332376 270048 336740 270076
rect 332376 270036 332382 270048
rect 336734 270036 336740 270048
rect 336792 270036 336798 270088
rect 341794 270036 341800 270088
rect 341852 270076 341858 270088
rect 357434 270076 357440 270088
rect 341852 270048 357440 270076
rect 341852 270036 341858 270048
rect 357434 270036 357440 270048
rect 357492 270036 357498 270088
rect 369394 270036 369400 270088
rect 369452 270076 369458 270088
rect 396074 270076 396080 270088
rect 369452 270048 396080 270076
rect 369452 270036 369458 270048
rect 396074 270036 396080 270048
rect 396132 270036 396138 270088
rect 403066 270036 403072 270088
rect 403124 270076 403130 270088
rect 444374 270076 444380 270088
rect 403124 270048 444380 270076
rect 403124 270036 403130 270048
rect 444374 270036 444380 270048
rect 444432 270036 444438 270088
rect 465994 270036 466000 270088
rect 466052 270076 466058 270088
rect 528848 270076 528876 270184
rect 533890 270172 533896 270184
rect 533948 270172 533954 270224
rect 534028 270172 534034 270224
rect 534086 270212 534092 270224
rect 626534 270212 626540 270224
rect 534086 270184 626540 270212
rect 534086 270172 534092 270184
rect 626534 270172 626540 270184
rect 626592 270172 626598 270224
rect 466052 270048 528876 270076
rect 466052 270036 466058 270048
rect 529014 270036 529020 270088
rect 529072 270076 529078 270088
rect 538858 270076 538864 270088
rect 529072 270048 538864 270076
rect 529072 270036 529078 270048
rect 538858 270036 538864 270048
rect 538916 270036 538922 270088
rect 540974 270036 540980 270088
rect 541032 270076 541038 270088
rect 541802 270076 541808 270088
rect 541032 270048 541808 270076
rect 541032 270036 541038 270048
rect 541802 270036 541808 270048
rect 541860 270036 541866 270088
rect 541986 270036 541992 270088
rect 542044 270076 542050 270088
rect 633618 270076 633624 270088
rect 542044 270048 633624 270076
rect 542044 270036 542050 270048
rect 633618 270036 633624 270048
rect 633676 270036 633682 270088
rect 143408 269912 151814 269940
rect 143408 269900 143414 269912
rect 154482 269900 154488 269952
rect 154540 269940 154546 269952
rect 198182 269940 198188 269952
rect 154540 269912 198188 269940
rect 154540 269900 154546 269912
rect 198182 269900 198188 269912
rect 198240 269900 198246 269952
rect 198642 269900 198648 269952
rect 198700 269940 198706 269952
rect 230014 269940 230020 269952
rect 198700 269912 230020 269940
rect 198700 269900 198706 269912
rect 230014 269900 230020 269912
rect 230072 269900 230078 269952
rect 230382 269900 230388 269952
rect 230440 269940 230446 269952
rect 252370 269940 252376 269952
rect 230440 269912 252376 269940
rect 230440 269900 230446 269912
rect 252370 269900 252376 269912
rect 252428 269900 252434 269952
rect 258442 269900 258448 269952
rect 258500 269940 258506 269952
rect 272242 269940 272248 269952
rect 258500 269912 272248 269940
rect 258500 269900 258506 269912
rect 272242 269900 272248 269912
rect 272300 269900 272306 269952
rect 273070 269900 273076 269952
rect 273128 269940 273134 269952
rect 282178 269940 282184 269952
rect 273128 269912 282184 269940
rect 273128 269900 273134 269912
rect 282178 269900 282184 269912
rect 282236 269900 282242 269952
rect 286778 269900 286784 269952
rect 286836 269940 286842 269952
rect 292114 269940 292120 269952
rect 286836 269912 292120 269940
rect 286836 269900 286842 269912
rect 292114 269900 292120 269912
rect 292172 269900 292178 269952
rect 326890 269900 326896 269952
rect 326948 269940 326954 269952
rect 335906 269940 335912 269952
rect 326948 269912 335912 269940
rect 326948 269900 326954 269912
rect 335906 269900 335912 269912
rect 335964 269900 335970 269952
rect 336826 269900 336832 269952
rect 336884 269940 336890 269952
rect 350534 269940 350540 269952
rect 336884 269912 350540 269940
rect 336884 269900 336890 269912
rect 350534 269900 350540 269912
rect 350592 269900 350598 269952
rect 354214 269900 354220 269952
rect 354272 269940 354278 269952
rect 375374 269940 375380 269952
rect 354272 269912 375380 269940
rect 354272 269900 354278 269912
rect 375374 269900 375380 269912
rect 375432 269900 375438 269952
rect 376570 269900 376576 269952
rect 376628 269940 376634 269952
rect 403986 269940 403992 269952
rect 376628 269912 403992 269940
rect 376628 269900 376634 269912
rect 403986 269900 403992 269912
rect 404044 269900 404050 269952
rect 413002 269900 413008 269952
rect 413060 269940 413066 269952
rect 459554 269940 459560 269952
rect 413060 269912 459560 269940
rect 413060 269900 413066 269912
rect 459554 269900 459560 269912
rect 459612 269900 459618 269952
rect 461854 269900 461860 269952
rect 461912 269940 461918 269952
rect 529198 269940 529204 269952
rect 461912 269912 529204 269940
rect 461912 269900 461918 269912
rect 529198 269900 529204 269912
rect 529256 269900 529262 269952
rect 529750 269900 529756 269952
rect 529808 269940 529814 269952
rect 530302 269940 530308 269952
rect 529808 269912 530308 269940
rect 529808 269900 529814 269912
rect 530302 269900 530308 269912
rect 530360 269900 530366 269952
rect 530578 269900 530584 269952
rect 530636 269940 530642 269952
rect 532878 269940 532884 269952
rect 530636 269912 532884 269940
rect 530636 269900 530642 269912
rect 532878 269900 532884 269912
rect 532936 269900 532942 269952
rect 533062 269900 533068 269952
rect 533120 269940 533126 269952
rect 630674 269940 630680 269952
rect 533120 269912 630680 269940
rect 533120 269900 533126 269912
rect 630674 269900 630680 269912
rect 630732 269900 630738 269952
rect 69382 269764 69388 269816
rect 69440 269804 69446 269816
rect 139762 269804 139768 269816
rect 69440 269776 139768 269804
rect 69440 269764 69446 269776
rect 139762 269764 139768 269776
rect 139820 269764 139826 269816
rect 139946 269764 139952 269816
rect 140004 269804 140010 269816
rect 181162 269804 181168 269816
rect 140004 269776 181168 269804
rect 140004 269764 140010 269776
rect 181162 269764 181168 269776
rect 181220 269764 181226 269816
rect 182082 269764 182088 269816
rect 182140 269804 182146 269816
rect 186958 269804 186964 269816
rect 182140 269776 186964 269804
rect 182140 269764 182146 269776
rect 186958 269764 186964 269776
rect 187016 269764 187022 269816
rect 187326 269764 187332 269816
rect 187384 269804 187390 269816
rect 191926 269804 191932 269816
rect 187384 269776 191932 269804
rect 187384 269764 187390 269776
rect 191926 269764 191932 269776
rect 191984 269764 191990 269816
rect 194594 269764 194600 269816
rect 194652 269804 194658 269816
rect 227254 269804 227260 269816
rect 194652 269776 227260 269804
rect 194652 269764 194658 269776
rect 227254 269764 227260 269776
rect 227312 269764 227318 269816
rect 249886 269804 249892 269816
rect 229066 269776 249892 269804
rect 84102 269628 84108 269680
rect 84160 269668 84166 269680
rect 119798 269668 119804 269680
rect 84160 269640 119804 269668
rect 84160 269628 84166 269640
rect 119798 269628 119804 269640
rect 119856 269628 119862 269680
rect 173710 269668 173716 269680
rect 122806 269640 173716 269668
rect 119062 269492 119068 269544
rect 119120 269532 119126 269544
rect 122806 269532 122834 269640
rect 173710 269628 173716 269640
rect 173768 269628 173774 269680
rect 184750 269628 184756 269680
rect 184808 269668 184814 269680
rect 213822 269668 213828 269680
rect 184808 269640 213828 269668
rect 184808 269628 184814 269640
rect 213822 269628 213828 269640
rect 213880 269628 213886 269680
rect 226610 269628 226616 269680
rect 226668 269668 226674 269680
rect 229066 269668 229094 269776
rect 249886 269764 249892 269776
rect 249944 269764 249950 269816
rect 251450 269764 251456 269816
rect 251508 269804 251514 269816
rect 267274 269804 267280 269816
rect 251508 269776 267280 269804
rect 251508 269764 251514 269776
rect 267274 269764 267280 269776
rect 267332 269764 267338 269816
rect 270310 269764 270316 269816
rect 270368 269804 270374 269816
rect 280522 269804 280528 269816
rect 270368 269776 280528 269804
rect 270368 269764 270374 269776
rect 280522 269764 280528 269776
rect 280580 269764 280586 269816
rect 314470 269764 314476 269816
rect 314528 269804 314534 269816
rect 318978 269804 318984 269816
rect 314528 269776 318984 269804
rect 314528 269764 314534 269776
rect 318978 269764 318984 269776
rect 319036 269764 319042 269816
rect 329650 269764 329656 269816
rect 329708 269804 329714 269816
rect 339494 269804 339500 269816
rect 329708 269776 339500 269804
rect 329708 269764 329714 269776
rect 339494 269764 339500 269776
rect 339552 269764 339558 269816
rect 347590 269764 347596 269816
rect 347648 269804 347654 269816
rect 365714 269804 365720 269816
rect 347648 269776 365720 269804
rect 347648 269764 347654 269776
rect 365714 269764 365720 269776
rect 365772 269764 365778 269816
rect 372338 269764 372344 269816
rect 372396 269804 372402 269816
rect 401778 269804 401784 269816
rect 372396 269776 401784 269804
rect 372396 269764 372402 269776
rect 401778 269764 401784 269776
rect 401836 269764 401842 269816
rect 457714 269764 457720 269816
rect 457772 269804 457778 269816
rect 470962 269804 470968 269816
rect 457772 269776 470968 269804
rect 457772 269764 457778 269776
rect 470962 269764 470968 269776
rect 471020 269764 471026 269816
rect 471606 269764 471612 269816
rect 471664 269804 471670 269816
rect 537938 269804 537944 269816
rect 471664 269776 537944 269804
rect 471664 269764 471670 269776
rect 537938 269764 537944 269776
rect 537996 269764 538002 269816
rect 538858 269764 538864 269816
rect 538916 269804 538922 269816
rect 552290 269804 552296 269816
rect 538916 269776 552296 269804
rect 538916 269764 538922 269776
rect 552290 269764 552296 269776
rect 552348 269764 552354 269816
rect 552474 269764 552480 269816
rect 552532 269804 552538 269816
rect 641898 269804 641904 269816
rect 552532 269776 641904 269804
rect 552532 269764 552538 269776
rect 641898 269764 641904 269776
rect 641956 269764 641962 269816
rect 226668 269640 229094 269668
rect 226668 269628 226674 269640
rect 253198 269628 253204 269680
rect 253256 269668 253262 269680
rect 258166 269668 258172 269680
rect 253256 269640 258172 269668
rect 253256 269628 253262 269640
rect 258166 269628 258172 269640
rect 258224 269628 258230 269680
rect 351638 269628 351644 269680
rect 351696 269668 351702 269680
rect 364334 269668 364340 269680
rect 351696 269640 364340 269668
rect 351696 269628 351702 269640
rect 364334 269628 364340 269640
rect 364392 269628 364398 269680
rect 384022 269628 384028 269680
rect 384080 269668 384086 269680
rect 388162 269668 388168 269680
rect 384080 269640 388168 269668
rect 384080 269628 384086 269640
rect 388162 269628 388168 269640
rect 388220 269628 388226 269680
rect 404354 269628 404360 269680
rect 404412 269668 404418 269680
rect 426618 269668 426624 269680
rect 404412 269640 426624 269668
rect 404412 269628 404418 269640
rect 426618 269628 426624 269640
rect 426676 269628 426682 269680
rect 427354 269628 427360 269680
rect 427412 269668 427418 269680
rect 478874 269668 478880 269680
rect 427412 269640 478880 269668
rect 427412 269628 427418 269640
rect 478874 269628 478880 269640
rect 478932 269628 478938 269680
rect 484210 269628 484216 269680
rect 484268 269668 484274 269680
rect 494514 269668 494520 269680
rect 484268 269640 494520 269668
rect 484268 269628 484274 269640
rect 494514 269628 494520 269640
rect 494572 269628 494578 269680
rect 494882 269628 494888 269680
rect 494940 269668 494946 269680
rect 504358 269668 504364 269680
rect 494940 269640 504364 269668
rect 494940 269628 494946 269640
rect 504358 269628 504364 269640
rect 504416 269628 504422 269680
rect 504542 269628 504548 269680
rect 504600 269668 504606 269680
rect 553026 269668 553032 269680
rect 504600 269640 553032 269668
rect 504600 269628 504606 269640
rect 553026 269628 553032 269640
rect 553084 269628 553090 269680
rect 558914 269628 558920 269680
rect 558972 269668 558978 269680
rect 572714 269668 572720 269680
rect 558972 269640 572720 269668
rect 558972 269628 558978 269640
rect 572714 269628 572720 269640
rect 572772 269628 572778 269680
rect 119120 269504 122834 269532
rect 119120 269492 119126 269504
rect 126882 269492 126888 269544
rect 126940 269532 126946 269544
rect 178678 269532 178684 269544
rect 126940 269504 178684 269532
rect 126940 269492 126946 269504
rect 178678 269492 178684 269504
rect 178736 269492 178742 269544
rect 183462 269492 183468 269544
rect 183520 269532 183526 269544
rect 187326 269532 187332 269544
rect 183520 269504 187332 269532
rect 183520 269492 183526 269504
rect 187326 269492 187332 269504
rect 187384 269492 187390 269544
rect 208302 269492 208308 269544
rect 208360 269532 208366 269544
rect 230750 269532 230756 269544
rect 208360 269504 230756 269532
rect 208360 269492 208366 269504
rect 230750 269492 230756 269504
rect 230808 269492 230814 269544
rect 394694 269492 394700 269544
rect 394752 269532 394758 269544
rect 416774 269532 416780 269544
rect 394752 269504 416780 269532
rect 394752 269492 394758 269504
rect 416774 269492 416780 269504
rect 416832 269492 416838 269544
rect 419626 269492 419632 269544
rect 419684 269532 419690 269544
rect 468018 269532 468024 269544
rect 419684 269504 468024 269532
rect 419684 269492 419690 269504
rect 468018 269492 468024 269504
rect 468076 269492 468082 269544
rect 474274 269492 474280 269544
rect 474332 269532 474338 269544
rect 474332 269504 537340 269532
rect 474332 269492 474338 269504
rect 335630 269424 335636 269476
rect 335688 269464 335694 269476
rect 343818 269464 343824 269476
rect 335688 269436 343824 269464
rect 335688 269424 335694 269436
rect 343818 269424 343824 269436
rect 343876 269424 343882 269476
rect 118602 269356 118608 269408
rect 118660 269396 118666 269408
rect 166902 269396 166908 269408
rect 118660 269368 166908 269396
rect 118660 269356 118666 269368
rect 166902 269356 166908 269368
rect 166960 269356 166966 269408
rect 401594 269356 401600 269408
rect 401652 269396 401658 269408
rect 430574 269396 430580 269408
rect 401652 269368 430580 269396
rect 401652 269356 401658 269368
rect 430574 269356 430580 269368
rect 430632 269356 430638 269408
rect 449894 269356 449900 269408
rect 449952 269396 449958 269408
rect 471974 269396 471980 269408
rect 449952 269368 471980 269396
rect 449952 269356 449958 269368
rect 471974 269356 471980 269368
rect 472032 269356 472038 269408
rect 476758 269356 476764 269408
rect 476816 269396 476822 269408
rect 537312 269396 537340 269504
rect 537938 269492 537944 269544
rect 537996 269532 538002 269544
rect 540974 269532 540980 269544
rect 537996 269504 540980 269532
rect 537996 269492 538002 269504
rect 540974 269492 540980 269504
rect 541032 269492 541038 269544
rect 541342 269492 541348 269544
rect 541400 269532 541406 269544
rect 552382 269532 552388 269544
rect 541400 269504 552388 269532
rect 541400 269492 541406 269504
rect 552382 269492 552388 269504
rect 552440 269492 552446 269544
rect 568574 269532 568580 269544
rect 552768 269504 568580 269532
rect 552768 269464 552796 269504
rect 568574 269492 568580 269504
rect 568632 269492 568638 269544
rect 552584 269436 552796 269464
rect 546218 269396 546224 269408
rect 476816 269368 537248 269396
rect 537312 269368 546224 269396
rect 476816 269356 476822 269368
rect 136818 269220 136824 269272
rect 136876 269260 136882 269272
rect 182174 269260 182180 269272
rect 136876 269232 182180 269260
rect 136876 269220 136882 269232
rect 182174 269220 182180 269232
rect 182232 269220 182238 269272
rect 264882 269220 264888 269272
rect 264940 269260 264946 269272
rect 269114 269260 269120 269272
rect 264940 269232 269120 269260
rect 264940 269220 264946 269232
rect 269114 269220 269120 269232
rect 269172 269220 269178 269272
rect 321094 269220 321100 269272
rect 321152 269260 321158 269272
rect 327902 269260 327908 269272
rect 321152 269232 327908 269260
rect 321152 269220 321158 269232
rect 327902 269220 327908 269232
rect 327960 269220 327966 269272
rect 417142 269220 417148 269272
rect 417200 269260 417206 269272
rect 465074 269260 465080 269272
rect 417200 269232 465080 269260
rect 417200 269220 417206 269232
rect 465074 269220 465080 269232
rect 465132 269220 465138 269272
rect 468754 269220 468760 269272
rect 468812 269260 468818 269272
rect 537018 269260 537024 269272
rect 468812 269232 537024 269260
rect 468812 269220 468818 269232
rect 537018 269220 537024 269232
rect 537076 269220 537082 269272
rect 537220 269260 537248 269368
rect 546218 269356 546224 269368
rect 546276 269356 546282 269408
rect 546402 269356 546408 269408
rect 546460 269396 546466 269408
rect 551922 269396 551928 269408
rect 546460 269368 551928 269396
rect 546460 269356 546466 269368
rect 551922 269356 551928 269368
rect 551980 269356 551986 269408
rect 552584 269396 552612 269436
rect 552124 269368 552612 269396
rect 549438 269260 549444 269272
rect 537220 269232 549444 269260
rect 549438 269220 549444 269232
rect 549496 269220 549502 269272
rect 549622 269220 549628 269272
rect 549680 269260 549686 269272
rect 552124 269260 552152 269368
rect 553026 269356 553032 269408
rect 553084 269396 553090 269408
rect 557534 269396 557540 269408
rect 553084 269368 557540 269396
rect 553084 269356 553090 269368
rect 557534 269356 557540 269368
rect 557592 269356 557598 269408
rect 549680 269232 552152 269260
rect 549680 269220 549686 269232
rect 552290 269220 552296 269272
rect 552348 269260 552354 269272
rect 607582 269260 607588 269272
rect 552348 269232 607588 269260
rect 552348 269220 552354 269232
rect 607582 269220 607588 269232
rect 607640 269220 607646 269272
rect 282730 269084 282736 269136
rect 282788 269124 282794 269136
rect 288802 269124 288808 269136
rect 282788 269096 288808 269124
rect 282788 269084 282794 269096
rect 288802 269084 288808 269096
rect 288860 269084 288866 269136
rect 295334 269084 295340 269136
rect 295392 269124 295398 269136
rect 297542 269124 297548 269136
rect 295392 269096 297548 269124
rect 295392 269084 295398 269096
rect 297542 269084 297548 269096
rect 297600 269084 297606 269136
rect 319438 269084 319444 269136
rect 319496 269124 319502 269136
rect 325694 269124 325700 269136
rect 319496 269096 325700 269124
rect 319496 269084 319502 269096
rect 325694 269084 325700 269096
rect 325752 269084 325758 269136
rect 434438 269084 434444 269136
rect 434496 269124 434502 269136
rect 490190 269124 490196 269136
rect 434496 269096 490196 269124
rect 434496 269084 434502 269096
rect 490190 269084 490196 269096
rect 490248 269084 490254 269136
rect 108942 269016 108948 269068
rect 109000 269056 109006 269068
rect 166258 269056 166264 269068
rect 109000 269028 166264 269056
rect 109000 269016 109006 269028
rect 166258 269016 166264 269028
rect 166316 269016 166322 269068
rect 185578 269016 185584 269068
rect 185636 269056 185642 269068
rect 196894 269056 196900 269068
rect 185636 269028 196900 269056
rect 185636 269016 185642 269028
rect 196894 269016 196900 269028
rect 196952 269016 196958 269068
rect 251082 269016 251088 269068
rect 251140 269056 251146 269068
rect 256510 269056 256516 269068
rect 251140 269028 256516 269056
rect 251140 269016 251146 269028
rect 256510 269016 256516 269028
rect 256568 269016 256574 269068
rect 422294 269056 422300 269068
rect 412606 269028 422300 269056
rect 86862 268880 86868 268932
rect 86920 268920 86926 268932
rect 144730 268920 144736 268932
rect 86920 268892 144736 268920
rect 86920 268880 86926 268892
rect 144730 268880 144736 268892
rect 144788 268880 144794 268932
rect 179322 268880 179328 268932
rect 179380 268920 179386 268932
rect 215938 268920 215944 268932
rect 179380 268892 215944 268920
rect 179380 268880 179386 268892
rect 215938 268880 215944 268892
rect 215996 268880 216002 268932
rect 382366 268880 382372 268932
rect 382424 268920 382430 268932
rect 400582 268920 400588 268932
rect 382424 268892 400588 268920
rect 382424 268880 382430 268892
rect 400582 268880 400588 268892
rect 400640 268880 400646 268932
rect 102502 268744 102508 268796
rect 102560 268784 102566 268796
rect 162946 268784 162952 268796
rect 102560 268756 162952 268784
rect 102560 268744 102566 268756
rect 162946 268744 162952 268756
rect 163004 268744 163010 268796
rect 163130 268744 163136 268796
rect 163188 268784 163194 268796
rect 203518 268784 203524 268796
rect 163188 268756 203524 268784
rect 163188 268744 163194 268756
rect 203518 268744 203524 268756
rect 203576 268744 203582 268796
rect 203886 268744 203892 268796
rect 203944 268784 203950 268796
rect 227714 268784 227720 268796
rect 203944 268756 227720 268784
rect 203944 268744 203950 268756
rect 227714 268744 227720 268756
rect 227772 268744 227778 268796
rect 227898 268744 227904 268796
rect 227956 268784 227962 268796
rect 250714 268784 250720 268796
rect 227956 268756 250720 268784
rect 227956 268744 227962 268756
rect 250714 268744 250720 268756
rect 250772 268744 250778 268796
rect 387334 268744 387340 268796
rect 387392 268784 387398 268796
rect 412606 268784 412634 269028
rect 422294 269016 422300 269028
rect 422352 269016 422358 269068
rect 499114 269016 499120 269068
rect 499172 269056 499178 269068
rect 582374 269056 582380 269068
rect 499172 269028 582380 269056
rect 499172 269016 499178 269028
rect 582374 269016 582380 269028
rect 582432 269016 582438 269068
rect 590654 269016 590660 269068
rect 590712 269056 590718 269068
rect 590712 269028 596174 269056
rect 590712 269016 590718 269028
rect 418982 268880 418988 268932
rect 419040 268920 419046 268932
rect 440234 268920 440240 268932
rect 419040 268892 440240 268920
rect 419040 268880 419046 268892
rect 440234 268880 440240 268892
rect 440292 268880 440298 268932
rect 443638 268880 443644 268932
rect 443696 268920 443702 268932
rect 502518 268920 502524 268932
rect 443696 268892 502524 268920
rect 443696 268880 443702 268892
rect 502518 268880 502524 268892
rect 502576 268880 502582 268932
rect 503070 268880 503076 268932
rect 503128 268920 503134 268932
rect 505094 268920 505100 268932
rect 503128 268892 505100 268920
rect 503128 268880 503134 268892
rect 505094 268880 505100 268892
rect 505152 268880 505158 268932
rect 508222 268880 508228 268932
rect 508280 268920 508286 268932
rect 594794 268920 594800 268932
rect 508280 268892 594800 268920
rect 508280 268880 508286 268892
rect 594794 268880 594800 268892
rect 594852 268880 594858 268932
rect 387392 268756 412634 268784
rect 387392 268744 387398 268756
rect 422294 268744 422300 268796
rect 422352 268784 422358 268796
rect 436094 268784 436100 268796
rect 422352 268756 436100 268784
rect 422352 268744 422358 268756
rect 436094 268744 436100 268756
rect 436152 268744 436158 268796
rect 441154 268744 441160 268796
rect 441212 268784 441218 268796
rect 499574 268784 499580 268796
rect 441212 268756 499580 268784
rect 441212 268744 441218 268756
rect 499574 268744 499580 268756
rect 499632 268744 499638 268796
rect 504082 268744 504088 268796
rect 504140 268784 504146 268796
rect 509326 268784 509332 268796
rect 504140 268756 509332 268784
rect 504140 268744 504146 268756
rect 509326 268744 509332 268756
rect 509384 268744 509390 268796
rect 510706 268744 510712 268796
rect 510764 268784 510770 268796
rect 510764 268756 513972 268784
rect 510764 268744 510770 268756
rect 513944 268716 513972 268756
rect 514294 268744 514300 268796
rect 514352 268784 514358 268796
rect 581638 268784 581644 268796
rect 514352 268756 581644 268784
rect 514352 268744 514358 268756
rect 581638 268744 581644 268756
rect 581696 268744 581702 268796
rect 581822 268744 581828 268796
rect 581880 268784 581886 268796
rect 596146 268784 596174 269028
rect 598842 268784 598848 268796
rect 581880 268756 590884 268784
rect 596146 268756 598848 268784
rect 581880 268744 581886 268756
rect 590856 268716 590884 268756
rect 598842 268744 598848 268756
rect 598900 268744 598906 268796
rect 513944 268688 514156 268716
rect 590856 268688 590976 268716
rect 99282 268608 99288 268660
rect 99340 268648 99346 268660
rect 160462 268648 160468 268660
rect 99340 268620 160468 268648
rect 99340 268608 99346 268620
rect 160462 268608 160468 268620
rect 160520 268608 160526 268660
rect 162762 268608 162768 268660
rect 162820 268648 162826 268660
rect 205174 268648 205180 268660
rect 162820 268620 205180 268648
rect 162820 268608 162826 268620
rect 205174 268608 205180 268620
rect 205232 268608 205238 268660
rect 219526 268608 219532 268660
rect 219584 268648 219590 268660
rect 244918 268648 244924 268660
rect 219584 268620 244924 268648
rect 219584 268608 219590 268620
rect 244918 268608 244924 268620
rect 244976 268608 244982 268660
rect 363046 268608 363052 268660
rect 363104 268648 363110 268660
rect 386414 268648 386420 268660
rect 363104 268620 386420 268648
rect 363104 268608 363110 268620
rect 386414 268608 386420 268620
rect 386472 268608 386478 268660
rect 402238 268608 402244 268660
rect 402296 268648 402302 268660
rect 443270 268648 443276 268660
rect 402296 268620 443276 268648
rect 402296 268608 402302 268620
rect 443270 268608 443276 268620
rect 443328 268608 443334 268660
rect 446122 268608 446128 268660
rect 446180 268648 446186 268660
rect 503070 268648 503076 268660
rect 446180 268620 503076 268648
rect 446180 268608 446186 268620
rect 503070 268608 503076 268620
rect 503128 268608 503134 268660
rect 503254 268608 503260 268660
rect 503312 268648 503318 268660
rect 513742 268648 513748 268660
rect 503312 268620 513748 268648
rect 503312 268608 503318 268620
rect 513742 268608 513748 268620
rect 513800 268608 513806 268660
rect 514128 268648 514156 268688
rect 590654 268648 590660 268660
rect 514128 268620 590660 268648
rect 590654 268608 590660 268620
rect 590712 268608 590718 268660
rect 590948 268648 590976 268688
rect 608686 268648 608692 268660
rect 590948 268620 608692 268648
rect 608686 268608 608692 268620
rect 608744 268608 608750 268660
rect 92382 268472 92388 268524
rect 92440 268512 92446 268524
rect 155494 268512 155500 268524
rect 92440 268484 155500 268512
rect 92440 268472 92446 268484
rect 155494 268472 155500 268484
rect 155552 268472 155558 268524
rect 155862 268472 155868 268524
rect 155920 268512 155926 268524
rect 200206 268512 200212 268524
rect 155920 268484 200212 268512
rect 155920 268472 155926 268484
rect 200206 268472 200212 268484
rect 200264 268472 200270 268524
rect 202966 268472 202972 268524
rect 203024 268512 203030 268524
rect 233326 268512 233332 268524
rect 203024 268484 233332 268512
rect 203024 268472 203030 268484
rect 233326 268472 233332 268484
rect 233384 268472 233390 268524
rect 245562 268472 245568 268524
rect 245620 268512 245626 268524
rect 263134 268512 263140 268524
rect 245620 268484 263140 268512
rect 245620 268472 245626 268484
rect 263134 268472 263140 268484
rect 263192 268472 263198 268524
rect 263502 268472 263508 268524
rect 263560 268512 263566 268524
rect 275554 268512 275560 268524
rect 263560 268484 275560 268512
rect 263560 268472 263566 268484
rect 275554 268472 275560 268484
rect 275612 268472 275618 268524
rect 333514 268472 333520 268524
rect 333572 268512 333578 268524
rect 345106 268512 345112 268524
rect 333572 268484 345112 268512
rect 333572 268472 333578 268484
rect 345106 268472 345112 268484
rect 345164 268472 345170 268524
rect 345934 268472 345940 268524
rect 345992 268512 345998 268524
rect 360286 268512 360292 268524
rect 345992 268484 360292 268512
rect 345992 268472 345998 268484
rect 360286 268472 360292 268484
rect 360344 268472 360350 268524
rect 361022 268472 361028 268524
rect 361080 268512 361086 268524
rect 369854 268512 369860 268524
rect 361080 268484 369860 268512
rect 361080 268472 361086 268484
rect 369854 268472 369860 268484
rect 369912 268472 369918 268524
rect 370314 268472 370320 268524
rect 370372 268512 370378 268524
rect 397454 268512 397460 268524
rect 370372 268484 397460 268512
rect 370372 268472 370378 268484
rect 397454 268472 397460 268484
rect 397512 268472 397518 268524
rect 400582 268472 400588 268524
rect 400640 268512 400646 268524
rect 441614 268512 441620 268524
rect 400640 268484 441620 268512
rect 400640 268472 400646 268484
rect 441614 268472 441620 268484
rect 441672 268472 441678 268524
rect 442718 268472 442724 268524
rect 442776 268512 442782 268524
rect 446766 268512 446772 268524
rect 442776 268484 446772 268512
rect 442776 268472 442782 268484
rect 446766 268472 446772 268484
rect 446824 268472 446830 268524
rect 448606 268472 448612 268524
rect 448664 268512 448670 268524
rect 504082 268512 504088 268524
rect 448664 268484 504088 268512
rect 448664 268472 448670 268484
rect 504082 268472 504088 268484
rect 504140 268472 504146 268524
rect 504266 268472 504272 268524
rect 504324 268512 504330 268524
rect 504324 268484 519124 268512
rect 504324 268472 504330 268484
rect 66254 268336 66260 268388
rect 66312 268376 66318 268388
rect 137278 268376 137284 268388
rect 66312 268348 137284 268376
rect 66312 268336 66318 268348
rect 137278 268336 137284 268348
rect 137336 268336 137342 268388
rect 147582 268336 147588 268388
rect 147640 268376 147646 268388
rect 193582 268376 193588 268388
rect 147640 268348 193588 268376
rect 147640 268336 147646 268348
rect 193582 268336 193588 268348
rect 193640 268336 193646 268388
rect 197262 268336 197268 268388
rect 197320 268376 197326 268388
rect 229186 268376 229192 268388
rect 197320 268348 229192 268376
rect 197320 268336 197326 268348
rect 229186 268336 229192 268348
rect 229244 268336 229250 268388
rect 233694 268336 233700 268388
rect 233752 268376 233758 268388
rect 254854 268376 254860 268388
rect 233752 268348 254860 268376
rect 233752 268336 233758 268348
rect 254854 268336 254860 268348
rect 254912 268336 254918 268388
rect 255314 268336 255320 268388
rect 255372 268376 255378 268388
rect 269758 268376 269764 268388
rect 255372 268348 269764 268376
rect 255372 268336 255378 268348
rect 269758 268336 269764 268348
rect 269816 268336 269822 268388
rect 322750 268336 322756 268388
rect 322808 268376 322814 268388
rect 329834 268376 329840 268388
rect 322808 268348 329840 268376
rect 322808 268336 322814 268348
rect 329834 268336 329840 268348
rect 329892 268336 329898 268388
rect 335170 268336 335176 268388
rect 335228 268376 335234 268388
rect 347774 268376 347780 268388
rect 335228 268348 347780 268376
rect 335228 268336 335234 268348
rect 347774 268336 347780 268348
rect 347832 268336 347838 268388
rect 350074 268336 350080 268388
rect 350132 268376 350138 268388
rect 367094 268376 367100 268388
rect 350132 268348 367100 268376
rect 350132 268336 350138 268348
rect 367094 268336 367100 268348
rect 367152 268336 367158 268388
rect 374914 268336 374920 268388
rect 374972 268376 374978 268388
rect 404538 268376 404544 268388
rect 374972 268348 404544 268376
rect 374972 268336 374978 268348
rect 404538 268336 404544 268348
rect 404596 268336 404602 268388
rect 407206 268336 407212 268388
rect 407264 268376 407270 268388
rect 451458 268376 451464 268388
rect 407264 268348 451464 268376
rect 407264 268336 407270 268348
rect 451458 268336 451464 268348
rect 451516 268336 451522 268388
rect 461026 268336 461032 268388
rect 461084 268376 461090 268388
rect 518802 268376 518808 268388
rect 461084 268348 518808 268376
rect 461084 268336 461090 268348
rect 518802 268336 518808 268348
rect 518860 268336 518866 268388
rect 519096 268376 519124 268484
rect 519354 268472 519360 268524
rect 519412 268512 519418 268524
rect 533890 268512 533896 268524
rect 519412 268484 533896 268512
rect 519412 268472 519418 268484
rect 533890 268472 533896 268484
rect 533948 268472 533954 268524
rect 534028 268472 534034 268524
rect 534086 268512 534092 268524
rect 619634 268512 619640 268524
rect 534086 268484 619640 268512
rect 534086 268472 534092 268484
rect 619634 268472 619640 268484
rect 619692 268472 619698 268524
rect 520274 268376 520280 268388
rect 519096 268348 520280 268376
rect 520274 268336 520280 268348
rect 520332 268336 520338 268388
rect 520458 268336 520464 268388
rect 520516 268376 520522 268388
rect 526990 268376 526996 268388
rect 520516 268348 526996 268376
rect 520516 268336 520522 268348
rect 526990 268336 526996 268348
rect 527048 268336 527054 268388
rect 527174 268336 527180 268388
rect 527232 268376 527238 268388
rect 547506 268376 547512 268388
rect 527232 268348 547512 268376
rect 527232 268336 527238 268348
rect 547506 268336 547512 268348
rect 547564 268336 547570 268388
rect 547690 268336 547696 268388
rect 547748 268376 547754 268388
rect 638954 268376 638960 268388
rect 547748 268348 638960 268376
rect 547748 268336 547754 268348
rect 638954 268336 638960 268348
rect 639012 268336 639018 268388
rect 122742 268200 122748 268252
rect 122800 268240 122806 268252
rect 176194 268240 176200 268252
rect 122800 268212 176200 268240
rect 122800 268200 122806 268212
rect 176194 268200 176200 268212
rect 176252 268200 176258 268252
rect 436186 268200 436192 268252
rect 436244 268240 436250 268252
rect 488902 268240 488908 268252
rect 436244 268212 488908 268240
rect 436244 268200 436250 268212
rect 488902 268200 488908 268212
rect 488960 268200 488966 268252
rect 504266 268240 504272 268252
rect 489886 268212 504272 268240
rect 133782 268064 133788 268116
rect 133840 268104 133846 268116
rect 183646 268104 183652 268116
rect 133840 268076 183652 268104
rect 133840 268064 133846 268076
rect 183646 268064 183652 268076
rect 183704 268064 183710 268116
rect 420454 268064 420460 268116
rect 420512 268104 420518 268116
rect 469030 268104 469036 268116
rect 420512 268076 469036 268104
rect 420512 268064 420518 268076
rect 469030 268064 469036 268076
rect 469088 268064 469094 268116
rect 469214 268064 469220 268116
rect 469272 268104 469278 268116
rect 489886 268104 489914 268212
rect 504266 268200 504272 268212
rect 504324 268200 504330 268252
rect 505738 268200 505744 268252
rect 505796 268240 505802 268252
rect 591022 268240 591028 268252
rect 505796 268212 591028 268240
rect 505796 268200 505802 268212
rect 591022 268200 591028 268212
rect 591080 268200 591086 268252
rect 469272 268076 489914 268104
rect 469272 268064 469278 268076
rect 492766 268064 492772 268116
rect 492824 268104 492830 268116
rect 498194 268104 498200 268116
rect 492824 268076 498200 268104
rect 492824 268064 492830 268076
rect 498194 268064 498200 268076
rect 498252 268064 498258 268116
rect 500678 268064 500684 268116
rect 500736 268104 500742 268116
rect 580442 268104 580448 268116
rect 500736 268076 580448 268104
rect 500736 268064 500742 268076
rect 580442 268064 580448 268076
rect 580500 268064 580506 268116
rect 581638 268064 581644 268116
rect 581696 268104 581702 268116
rect 587894 268104 587900 268116
rect 581696 268076 587900 268104
rect 581696 268064 581702 268076
rect 587894 268064 587900 268076
rect 587952 268064 587958 268116
rect 125502 267928 125508 267980
rect 125560 267968 125566 267980
rect 147582 267968 147588 267980
rect 125560 267940 147588 267968
rect 125560 267928 125566 267940
rect 147582 267928 147588 267940
rect 147640 267928 147646 267980
rect 437842 267928 437848 267980
rect 437900 267968 437906 267980
rect 468202 267968 468208 267980
rect 437900 267940 468208 267968
rect 437900 267928 437906 267940
rect 468202 267928 468208 267940
rect 468260 267928 468266 267980
rect 533890 267968 533896 267980
rect 470566 267940 533896 267968
rect 431954 267792 431960 267844
rect 432012 267832 432018 267844
rect 447134 267832 447140 267844
rect 432012 267804 447140 267832
rect 432012 267792 432018 267804
rect 447134 267792 447140 267804
rect 447192 267792 447198 267844
rect 470566 267764 470594 267940
rect 533890 267928 533896 267940
rect 533948 267928 533954 267980
rect 534028 267928 534034 267980
rect 534086 267968 534092 267980
rect 581822 267968 581828 267980
rect 534086 267940 581828 267968
rect 534086 267928 534092 267940
rect 581822 267928 581828 267940
rect 581880 267928 581886 267980
rect 488534 267832 488540 267844
rect 467852 267736 470594 267764
rect 481560 267804 488540 267832
rect 88978 267656 88984 267708
rect 89036 267696 89042 267708
rect 144546 267696 144552 267708
rect 89036 267668 144552 267696
rect 89036 267656 89042 267668
rect 144546 267656 144552 267668
rect 144604 267656 144610 267708
rect 144914 267656 144920 267708
rect 144972 267696 144978 267708
rect 150526 267696 150532 267708
rect 144972 267668 150532 267696
rect 144972 267656 144978 267668
rect 150526 267656 150532 267668
rect 150584 267656 150590 267708
rect 171778 267656 171784 267708
rect 171836 267696 171842 267708
rect 199378 267696 199384 267708
rect 171836 267668 199384 267696
rect 171836 267656 171842 267668
rect 199378 267656 199384 267668
rect 199436 267656 199442 267708
rect 207658 267656 207664 267708
rect 207716 267696 207722 267708
rect 213454 267696 213460 267708
rect 207716 267668 213460 267696
rect 207716 267656 207722 267668
rect 213454 267656 213460 267668
rect 213512 267656 213518 267708
rect 368198 267656 368204 267708
rect 368256 267696 368262 267708
rect 377582 267696 377588 267708
rect 368256 267668 377588 267696
rect 368256 267656 368262 267668
rect 377582 267656 377588 267668
rect 377640 267656 377646 267708
rect 383194 267656 383200 267708
rect 383252 267696 383258 267708
rect 394694 267696 394700 267708
rect 383252 267668 394700 267696
rect 383252 267656 383258 267668
rect 394694 267656 394700 267668
rect 394752 267656 394758 267708
rect 398466 267656 398472 267708
rect 398524 267696 398530 267708
rect 421742 267696 421748 267708
rect 398524 267668 421748 267696
rect 398524 267656 398530 267668
rect 421742 267656 421748 267668
rect 421800 267656 421806 267708
rect 435634 267656 435640 267708
rect 435692 267696 435698 267708
rect 465534 267696 465540 267708
rect 435692 267668 465540 267696
rect 435692 267656 435698 267668
rect 465534 267656 465540 267668
rect 465592 267656 465598 267708
rect 466822 267656 466828 267708
rect 466880 267696 466886 267708
rect 467852 267696 467880 267736
rect 466880 267668 467880 267696
rect 466880 267656 466886 267668
rect 477586 267656 477592 267708
rect 477644 267696 477650 267708
rect 481560 267696 481588 267804
rect 488534 267792 488540 267804
rect 488592 267792 488598 267844
rect 489178 267792 489184 267844
rect 489236 267832 489242 267844
rect 567286 267832 567292 267844
rect 489236 267804 567292 267832
rect 489236 267792 489242 267804
rect 567286 267792 567292 267804
rect 567344 267792 567350 267844
rect 580442 267792 580448 267844
rect 580500 267832 580506 267844
rect 584030 267832 584036 267844
rect 580500 267804 584036 267832
rect 580500 267792 580506 267804
rect 584030 267792 584036 267804
rect 584088 267792 584094 267844
rect 492766 267696 492772 267708
rect 477644 267668 481588 267696
rect 485056 267668 492772 267696
rect 477644 267656 477650 267668
rect 95878 267520 95884 267572
rect 95936 267560 95942 267572
rect 154666 267560 154672 267572
rect 95936 267532 154672 267560
rect 95936 267520 95942 267532
rect 154666 267520 154672 267532
rect 154724 267520 154730 267572
rect 162118 267520 162124 267572
rect 162176 267560 162182 267572
rect 169570 267560 169576 267572
rect 162176 267532 169576 267560
rect 162176 267520 162182 267532
rect 169570 267520 169576 267532
rect 169628 267520 169634 267572
rect 187142 267520 187148 267572
rect 187200 267560 187206 267572
rect 221734 267560 221740 267572
rect 187200 267532 221740 267560
rect 187200 267520 187206 267532
rect 221734 267520 221740 267532
rect 221792 267520 221798 267572
rect 227714 267520 227720 267572
rect 227772 267560 227778 267572
rect 234154 267560 234160 267572
rect 227772 267532 234160 267560
rect 227772 267520 227778 267532
rect 234154 267520 234160 267532
rect 234212 267520 234218 267572
rect 370774 267520 370780 267572
rect 370832 267560 370838 267572
rect 381538 267560 381544 267572
rect 370832 267532 381544 267560
rect 370832 267520 370838 267532
rect 381538 267520 381544 267532
rect 381596 267520 381602 267572
rect 390646 267520 390652 267572
rect 390704 267560 390710 267572
rect 404354 267560 404360 267572
rect 390704 267532 404360 267560
rect 390704 267520 390710 267532
rect 404354 267520 404360 267532
rect 404412 267520 404418 267572
rect 409598 267520 409604 267572
rect 409656 267560 409662 267572
rect 435358 267560 435364 267572
rect 409656 267532 435364 267560
rect 409656 267520 409662 267532
rect 435358 267520 435364 267532
rect 435416 267520 435422 267572
rect 445294 267520 445300 267572
rect 445352 267560 445358 267572
rect 485056 267560 485084 267668
rect 492766 267656 492772 267668
rect 492824 267656 492830 267708
rect 492950 267656 492956 267708
rect 493008 267696 493014 267708
rect 558914 267696 558920 267708
rect 493008 267668 558920 267696
rect 493008 267656 493014 267668
rect 558914 267656 558920 267668
rect 558972 267656 558978 267708
rect 445352 267532 485084 267560
rect 445352 267520 445358 267532
rect 485222 267520 485228 267572
rect 485280 267560 485286 267572
rect 502334 267560 502340 267572
rect 485280 267532 502340 267560
rect 485280 267520 485286 267532
rect 502334 267520 502340 267532
rect 502392 267520 502398 267572
rect 502794 267520 502800 267572
rect 502852 267560 502858 267572
rect 506198 267560 506204 267572
rect 502852 267532 506204 267560
rect 502852 267520 502858 267532
rect 506198 267520 506204 267532
rect 506256 267520 506262 267572
rect 506474 267520 506480 267572
rect 506532 267560 506538 267572
rect 507210 267560 507216 267572
rect 506532 267532 507216 267560
rect 506532 267520 506538 267532
rect 507210 267520 507216 267532
rect 507268 267520 507274 267572
rect 507394 267520 507400 267572
rect 507452 267560 507458 267572
rect 578878 267560 578884 267572
rect 507452 267532 578884 267560
rect 507452 267520 507458 267532
rect 578878 267520 578884 267532
rect 578936 267520 578942 267572
rect 107562 267384 107568 267436
rect 107620 267424 107626 267436
rect 167086 267424 167092 267436
rect 107620 267396 167092 267424
rect 107620 267384 107626 267396
rect 167086 267384 167092 267396
rect 167144 267384 167150 267436
rect 167730 267384 167736 267436
rect 167788 267424 167794 267436
rect 204346 267424 204352 267436
rect 167788 267396 204352 267424
rect 167788 267384 167794 267396
rect 204346 267384 204352 267396
rect 204404 267384 204410 267436
rect 211982 267384 211988 267436
rect 212040 267424 212046 267436
rect 222562 267424 222568 267436
rect 212040 267396 222568 267424
rect 212040 267384 212046 267396
rect 222562 267384 222568 267396
rect 222620 267384 222626 267436
rect 224218 267384 224224 267436
rect 224276 267424 224282 267436
rect 231670 267424 231676 267436
rect 224276 267396 231676 267424
rect 224276 267384 224282 267396
rect 231670 267384 231676 267396
rect 231728 267384 231734 267436
rect 233878 267384 233884 267436
rect 233936 267424 233942 267436
rect 246574 267424 246580 267436
rect 233936 267396 246580 267424
rect 233936 267384 233942 267396
rect 246574 267384 246580 267396
rect 246632 267384 246638 267436
rect 313642 267384 313648 267436
rect 313700 267424 313706 267436
rect 317782 267424 317788 267436
rect 313700 267396 317788 267424
rect 313700 267384 313706 267396
rect 317782 267384 317788 267396
rect 317840 267384 317846 267436
rect 334342 267384 334348 267436
rect 334400 267424 334406 267436
rect 342898 267424 342904 267436
rect 334400 267396 342904 267424
rect 334400 267384 334406 267396
rect 342898 267384 342904 267396
rect 342956 267384 342962 267436
rect 350902 267384 350908 267436
rect 350960 267424 350966 267436
rect 361022 267424 361028 267436
rect 350960 267396 361028 267424
rect 350960 267384 350966 267396
rect 361022 267384 361028 267396
rect 361080 267384 361086 267436
rect 365806 267384 365812 267436
rect 365864 267424 365870 267436
rect 382918 267424 382924 267436
rect 365864 267396 382924 267424
rect 365864 267384 365870 267396
rect 382918 267384 382924 267396
rect 382976 267384 382982 267436
rect 397086 267384 397092 267436
rect 397144 267424 397150 267436
rect 422294 267424 422300 267436
rect 397144 267396 422300 267424
rect 397144 267384 397150 267396
rect 422294 267384 422300 267396
rect 422352 267384 422358 267436
rect 440326 267384 440332 267436
rect 440384 267424 440390 267436
rect 494698 267424 494704 267436
rect 440384 267396 494704 267424
rect 440384 267384 440390 267396
rect 494698 267384 494704 267396
rect 494756 267384 494762 267436
rect 497458 267384 497464 267436
rect 497516 267424 497522 267436
rect 552842 267424 552848 267436
rect 497516 267396 552848 267424
rect 497516 267384 497522 267396
rect 552842 267384 552848 267396
rect 552900 267384 552906 267436
rect 553026 267384 553032 267436
rect 553084 267424 553090 267436
rect 570874 267424 570880 267436
rect 553084 267396 570880 267424
rect 553084 267384 553090 267396
rect 570874 267384 570880 267396
rect 570932 267384 570938 267436
rect 100662 267248 100668 267300
rect 100720 267288 100726 267300
rect 162118 267288 162124 267300
rect 100720 267260 162124 267288
rect 100720 267248 100726 267260
rect 162118 267248 162124 267260
rect 162176 267248 162182 267300
rect 166902 267248 166908 267300
rect 166960 267288 166966 267300
rect 174538 267288 174544 267300
rect 166960 267260 174544 267288
rect 166960 267248 166966 267260
rect 174538 267248 174544 267260
rect 174596 267248 174602 267300
rect 175090 267248 175096 267300
rect 175148 267288 175154 267300
rect 214282 267288 214288 267300
rect 175148 267260 214288 267288
rect 175148 267248 175154 267260
rect 214282 267248 214288 267260
rect 214340 267248 214346 267300
rect 220078 267248 220084 267300
rect 220136 267288 220142 267300
rect 239122 267288 239128 267300
rect 220136 267260 239128 267288
rect 220136 267248 220142 267260
rect 239122 267248 239128 267260
rect 239180 267248 239186 267300
rect 254578 267248 254584 267300
rect 254636 267288 254642 267300
rect 262306 267288 262312 267300
rect 254636 267260 262312 267288
rect 254636 267248 254642 267260
rect 262306 267248 262312 267260
rect 262364 267248 262370 267300
rect 312814 267248 312820 267300
rect 312872 267288 312878 267300
rect 316034 267288 316040 267300
rect 312872 267260 316040 267288
rect 312872 267248 312878 267260
rect 316034 267248 316040 267260
rect 316092 267248 316098 267300
rect 343450 267248 343456 267300
rect 343508 267288 343514 267300
rect 353938 267288 353944 267300
rect 343508 267260 353944 267288
rect 343508 267248 343514 267260
rect 353938 267248 353944 267260
rect 353996 267248 354002 267300
rect 359182 267248 359188 267300
rect 359240 267288 359246 267300
rect 373258 267288 373264 267300
rect 359240 267260 373264 267288
rect 359240 267248 359246 267260
rect 373258 267248 373264 267260
rect 373316 267248 373322 267300
rect 375742 267248 375748 267300
rect 375800 267288 375806 267300
rect 393958 267288 393964 267300
rect 375800 267260 393964 267288
rect 375800 267248 375806 267260
rect 393958 267248 393964 267260
rect 394016 267248 394022 267300
rect 399754 267248 399760 267300
rect 399812 267288 399818 267300
rect 418982 267288 418988 267300
rect 399812 267260 418988 267288
rect 399812 267248 399818 267260
rect 418982 267248 418988 267260
rect 419040 267248 419046 267300
rect 421282 267248 421288 267300
rect 421340 267288 421346 267300
rect 464154 267288 464160 267300
rect 421340 267260 464160 267288
rect 421340 267248 421346 267260
rect 464154 267248 464160 267260
rect 464212 267248 464218 267300
rect 465534 267248 465540 267300
rect 465592 267288 465598 267300
rect 471238 267288 471244 267300
rect 465592 267260 471244 267288
rect 465592 267248 465598 267260
rect 471238 267248 471244 267260
rect 471296 267248 471302 267300
rect 471790 267248 471796 267300
rect 471848 267288 471854 267300
rect 475378 267288 475384 267300
rect 471848 267260 475384 267288
rect 471848 267248 471854 267260
rect 475378 267248 475384 267260
rect 475436 267248 475442 267300
rect 475930 267248 475936 267300
rect 475988 267288 475994 267300
rect 518894 267288 518900 267300
rect 475988 267260 518900 267288
rect 475988 267248 475994 267260
rect 518894 267248 518900 267260
rect 518952 267248 518958 267300
rect 519170 267248 519176 267300
rect 519228 267288 519234 267300
rect 521654 267288 521660 267300
rect 519228 267260 521660 267288
rect 519228 267248 519234 267260
rect 521654 267248 521660 267260
rect 521712 267248 521718 267300
rect 522942 267248 522948 267300
rect 523000 267288 523006 267300
rect 523000 267260 523816 267288
rect 523000 267248 523006 267260
rect 73798 267112 73804 267164
rect 73856 267152 73862 267164
rect 141418 267152 141424 267164
rect 73856 267124 141424 267152
rect 73856 267112 73862 267124
rect 141418 267112 141424 267124
rect 141476 267112 141482 267164
rect 144546 267112 144552 267164
rect 144604 267152 144610 267164
rect 147398 267152 147404 267164
rect 144604 267124 147404 267152
rect 144604 267112 144610 267124
rect 147398 267112 147404 267124
rect 147456 267112 147462 267164
rect 147582 267112 147588 267164
rect 147640 267152 147646 267164
rect 149054 267152 149060 267164
rect 147640 267124 149060 267152
rect 147640 267112 147646 267124
rect 149054 267112 149060 267124
rect 149112 267112 149118 267164
rect 149882 267112 149888 267164
rect 149940 267152 149946 267164
rect 194410 267152 194416 267164
rect 149940 267124 194416 267152
rect 149940 267112 149946 267124
rect 194410 267112 194416 267124
rect 194468 267112 194474 267164
rect 199654 267112 199660 267164
rect 199712 267152 199718 267164
rect 218422 267152 218428 267164
rect 199712 267124 218428 267152
rect 199712 267112 199718 267124
rect 218422 267112 218428 267124
rect 218480 267112 218486 267164
rect 221458 267112 221464 267164
rect 221516 267152 221522 267164
rect 241606 267152 241612 267164
rect 221516 267124 241612 267152
rect 221516 267112 221522 267124
rect 241606 267112 241612 267124
rect 241664 267112 241670 267164
rect 246850 267112 246856 267164
rect 246908 267152 246914 267164
rect 263962 267152 263968 267164
rect 246908 267124 263968 267152
rect 246908 267112 246914 267124
rect 263962 267112 263968 267124
rect 264020 267112 264026 267164
rect 342622 267112 342628 267164
rect 342680 267152 342686 267164
rect 356514 267152 356520 267164
rect 342680 267124 356520 267152
rect 342680 267112 342686 267124
rect 356514 267112 356520 267124
rect 356572 267112 356578 267164
rect 363322 267112 363328 267164
rect 363380 267152 363386 267164
rect 370498 267152 370504 267164
rect 363380 267124 370504 267152
rect 363380 267112 363386 267124
rect 370498 267112 370504 267124
rect 370556 267112 370562 267164
rect 373258 267112 373264 267164
rect 373316 267152 373322 267164
rect 392578 267152 392584 267164
rect 373316 267124 392584 267152
rect 373316 267112 373322 267124
rect 392578 267112 392584 267124
rect 392636 267112 392642 267164
rect 404722 267112 404728 267164
rect 404780 267152 404786 267164
rect 431954 267152 431960 267164
rect 404780 267124 431960 267152
rect 404780 267112 404786 267124
rect 431954 267112 431960 267124
rect 432012 267112 432018 267164
rect 449894 267152 449900 267164
rect 441586 267124 449900 267152
rect 71038 266976 71044 267028
rect 71096 267016 71102 267028
rect 138106 267016 138112 267028
rect 71096 266988 138112 267016
rect 71096 266976 71102 266988
rect 138106 266976 138112 266988
rect 138164 266976 138170 267028
rect 141602 266976 141608 267028
rect 141660 267016 141666 267028
rect 184014 267016 184020 267028
rect 141660 266988 184020 267016
rect 141660 266976 141666 266988
rect 184014 266976 184020 266988
rect 184072 266976 184078 267028
rect 184198 266976 184204 267028
rect 184256 267016 184262 267028
rect 184256 266988 190454 267016
rect 184256 266976 184262 266988
rect 132402 266840 132408 266892
rect 132460 266880 132466 266892
rect 184474 266880 184480 266892
rect 132460 266852 184480 266880
rect 132460 266840 132466 266852
rect 184474 266840 184480 266852
rect 184532 266840 184538 266892
rect 190426 266880 190454 266988
rect 193858 266976 193864 267028
rect 193916 267016 193922 267028
rect 201862 267016 201868 267028
rect 193916 266988 201868 267016
rect 193916 266976 193922 266988
rect 201862 266976 201868 266988
rect 201920 266976 201926 267028
rect 206278 266976 206284 267028
rect 206336 267016 206342 267028
rect 228358 267016 228364 267028
rect 206336 266988 228364 267016
rect 206336 266976 206342 266988
rect 228358 266976 228364 266988
rect 228416 266976 228422 267028
rect 237282 266976 237288 267028
rect 237340 267016 237346 267028
rect 254026 267016 254032 267028
rect 237340 266988 254032 267016
rect 237340 266976 237346 266988
rect 254026 266976 254032 266988
rect 254084 266976 254090 267028
rect 271414 267016 271420 267028
rect 258046 266988 271420 267016
rect 258046 266892 258074 266988
rect 271414 266976 271420 266988
rect 271472 266976 271478 267028
rect 276658 266976 276664 267028
rect 276716 267016 276722 267028
rect 278038 267016 278044 267028
rect 276716 266988 278044 267016
rect 276716 266976 276722 266988
rect 278038 266976 278044 266988
rect 278096 266976 278102 267028
rect 286962 266976 286968 267028
rect 287020 267016 287026 267028
rect 291286 267016 291292 267028
rect 287020 266988 291292 267016
rect 287020 266976 287026 266988
rect 291286 266976 291292 266988
rect 291344 266976 291350 267028
rect 295150 266976 295156 267028
rect 295208 267016 295214 267028
rect 297082 267016 297088 267028
rect 295208 266988 297088 267016
rect 295208 266976 295214 266988
rect 297082 266976 297088 266988
rect 297140 266976 297146 267028
rect 324406 266976 324412 267028
rect 324464 267016 324470 267028
rect 332502 267016 332508 267028
rect 324464 266988 332508 267016
rect 324464 266976 324470 266988
rect 332502 266976 332508 266988
rect 332560 266976 332566 267028
rect 353386 266976 353392 267028
rect 353444 267016 353450 267028
rect 355318 267016 355324 267028
rect 353444 266988 355324 267016
rect 353444 266976 353450 266988
rect 355318 266976 355324 266988
rect 355376 266976 355382 267028
rect 355870 266976 355876 267028
rect 355928 267016 355934 267028
rect 369118 267016 369124 267028
rect 355928 266988 369124 267016
rect 355928 266976 355934 266988
rect 369118 266976 369124 266988
rect 369176 266976 369182 267028
rect 378226 266976 378232 267028
rect 378284 267016 378290 267028
rect 409138 267016 409144 267028
rect 378284 266988 409144 267016
rect 378284 266976 378290 266988
rect 409138 266976 409144 266988
rect 409196 266976 409202 267028
rect 422110 266976 422116 267028
rect 422168 267016 422174 267028
rect 441586 267016 441614 267124
rect 449894 267112 449900 267124
rect 449952 267112 449958 267164
rect 450262 267112 450268 267164
rect 450320 267152 450326 267164
rect 499758 267152 499764 267164
rect 450320 267124 499764 267152
rect 450320 267112 450326 267124
rect 499758 267112 499764 267124
rect 499816 267112 499822 267164
rect 499942 267112 499948 267164
rect 500000 267152 500006 267164
rect 500862 267152 500868 267164
rect 500000 267124 500868 267152
rect 500000 267112 500006 267124
rect 500862 267112 500868 267124
rect 500920 267112 500926 267164
rect 501046 267112 501052 267164
rect 501104 267152 501110 267164
rect 506382 267152 506388 267164
rect 501104 267124 506388 267152
rect 501104 267112 501110 267124
rect 506382 267112 506388 267124
rect 506440 267112 506446 267164
rect 506566 267112 506572 267164
rect 506624 267152 506630 267164
rect 507670 267152 507676 267164
rect 506624 267124 507676 267152
rect 506624 267112 506630 267124
rect 507670 267112 507676 267124
rect 507728 267112 507734 267164
rect 507854 267112 507860 267164
rect 507912 267152 507918 267164
rect 523586 267152 523592 267164
rect 507912 267124 523592 267152
rect 507912 267112 507918 267124
rect 523586 267112 523592 267124
rect 523644 267112 523650 267164
rect 523788 267152 523816 267260
rect 523954 267248 523960 267300
rect 524012 267288 524018 267300
rect 543550 267288 543556 267300
rect 524012 267260 543556 267288
rect 524012 267248 524018 267260
rect 543550 267248 543556 267260
rect 543608 267248 543614 267300
rect 543688 267248 543694 267300
rect 543746 267288 543752 267300
rect 621658 267288 621664 267300
rect 543746 267260 621664 267288
rect 543746 267248 543752 267260
rect 621658 267248 621664 267260
rect 621716 267248 621722 267300
rect 585778 267152 585784 267164
rect 523788 267124 585784 267152
rect 585778 267112 585784 267124
rect 585836 267112 585842 267164
rect 422168 266988 441614 267016
rect 422168 266976 422174 266988
rect 446398 266976 446404 267028
rect 446456 267016 446462 267028
rect 451734 267016 451740 267028
rect 446456 266988 451740 267016
rect 446456 266976 446462 266988
rect 451734 266976 451740 266988
rect 451792 266976 451798 267028
rect 451918 266976 451924 267028
rect 451976 267016 451982 267028
rect 460014 267016 460020 267028
rect 451976 266988 460020 267016
rect 451976 266976 451982 266988
rect 460014 266976 460020 266988
rect 460072 266976 460078 267028
rect 465166 266976 465172 267028
rect 465224 267016 465230 267028
rect 519170 267016 519176 267028
rect 465224 266988 519176 267016
rect 465224 266976 465230 266988
rect 519170 266976 519176 266988
rect 519228 266976 519234 267028
rect 519354 266976 519360 267028
rect 519412 267016 519418 267028
rect 520090 267016 520096 267028
rect 519412 266988 520096 267016
rect 519412 266976 519418 266988
rect 520090 266976 520096 266988
rect 520148 266976 520154 267028
rect 520274 266976 520280 267028
rect 520332 267016 520338 267028
rect 522942 267016 522948 267028
rect 520332 266988 522948 267016
rect 520332 266976 520338 266988
rect 522942 266976 522948 266988
rect 523000 266976 523006 267028
rect 523126 266976 523132 267028
rect 523184 267016 523190 267028
rect 524322 267016 524328 267028
rect 523184 266988 524328 267016
rect 523184 266976 523190 266988
rect 524322 266976 524328 266988
rect 524380 266976 524386 267028
rect 524782 266976 524788 267028
rect 524840 267016 524846 267028
rect 525702 267016 525708 267028
rect 524840 266988 525708 267016
rect 524840 266976 524846 266988
rect 525702 266976 525708 266988
rect 525760 266976 525766 267028
rect 525886 266976 525892 267028
rect 525944 267016 525950 267028
rect 533890 267016 533896 267028
rect 525944 266988 533896 267016
rect 525944 266976 525950 266988
rect 533890 266976 533896 266988
rect 533948 266976 533954 267028
rect 534028 266976 534034 267028
rect 534086 267016 534092 267028
rect 622394 267016 622400 267028
rect 534086 266988 622400 267016
rect 534086 266976 534092 266988
rect 622394 266976 622400 266988
rect 622452 266976 622458 267028
rect 209314 266880 209320 266892
rect 190426 266852 209320 266880
rect 209314 266840 209320 266852
rect 209372 266840 209378 266892
rect 216122 266840 216128 266892
rect 216180 266880 216186 266892
rect 223390 266880 223396 266892
rect 216180 266852 223396 266880
rect 216180 266840 216186 266852
rect 223390 266840 223396 266852
rect 223448 266840 223454 266892
rect 249058 266840 249064 266892
rect 249116 266880 249122 266892
rect 251542 266880 251548 266892
rect 249116 266852 251548 266880
rect 249116 266840 249122 266852
rect 251542 266840 251548 266852
rect 251600 266840 251606 266892
rect 257982 266840 257988 266892
rect 258040 266852 258074 266892
rect 258040 266840 258046 266852
rect 316126 266840 316132 266892
rect 316184 266880 316190 266892
rect 320174 266880 320180 266892
rect 316184 266852 320180 266880
rect 316184 266840 316190 266852
rect 320174 266840 320180 266852
rect 320232 266840 320238 266892
rect 331858 266840 331864 266892
rect 331916 266880 331922 266892
rect 335630 266880 335636 266892
rect 331916 266852 335636 266880
rect 331916 266840 331922 266852
rect 335630 266840 335636 266852
rect 335688 266840 335694 266892
rect 335998 266840 336004 266892
rect 336056 266880 336062 266892
rect 347038 266880 347044 266892
rect 336056 266852 347044 266880
rect 336056 266840 336062 266852
rect 347038 266840 347044 266852
rect 347096 266840 347102 266892
rect 393130 266840 393136 266892
rect 393188 266880 393194 266892
rect 401594 266880 401600 266892
rect 393188 266852 401600 266880
rect 393188 266840 393194 266852
rect 401594 266840 401600 266852
rect 401652 266840 401658 266892
rect 405550 266840 405556 266892
rect 405608 266880 405614 266892
rect 425698 266880 425704 266892
rect 405608 266852 425704 266880
rect 405608 266840 405614 266852
rect 425698 266840 425704 266852
rect 425756 266840 425762 266892
rect 451228 266880 451234 266892
rect 431926 266852 451234 266880
rect 265066 266772 265072 266824
rect 265124 266812 265130 266824
rect 268930 266812 268936 266824
rect 265124 266784 268936 266812
rect 265124 266772 265130 266784
rect 268930 266772 268936 266784
rect 268988 266772 268994 266824
rect 120718 266704 120724 266756
rect 120776 266744 120782 266756
rect 156414 266744 156420 266756
rect 120776 266716 156420 266744
rect 120776 266704 120782 266716
rect 156414 266704 156420 266716
rect 156472 266704 156478 266756
rect 156598 266704 156604 266756
rect 156656 266744 156662 266756
rect 159634 266744 159640 266756
rect 156656 266716 159640 266744
rect 156656 266704 156662 266716
rect 159634 266704 159640 266716
rect 159692 266704 159698 266756
rect 169018 266704 169024 266756
rect 169076 266744 169082 266756
rect 172054 266744 172060 266756
rect 169076 266716 172060 266744
rect 169076 266704 169082 266716
rect 172054 266704 172060 266716
rect 172112 266704 172118 266756
rect 184014 266704 184020 266756
rect 184072 266744 184078 266756
rect 189442 266744 189448 266756
rect 184072 266716 189448 266744
rect 184072 266704 184078 266716
rect 189442 266704 189448 266716
rect 189500 266704 189506 266756
rect 245102 266704 245108 266756
rect 245160 266744 245166 266756
rect 249058 266744 249064 266756
rect 245160 266716 249064 266744
rect 245160 266704 245166 266716
rect 249058 266704 249064 266716
rect 249116 266704 249122 266756
rect 320266 266704 320272 266756
rect 320324 266744 320330 266756
rect 327442 266744 327448 266756
rect 320324 266716 327448 266744
rect 320324 266704 320330 266716
rect 327442 266704 327448 266716
rect 327500 266704 327506 266756
rect 358354 266704 358360 266756
rect 358412 266744 358418 266756
rect 360838 266744 360844 266756
rect 358412 266716 360844 266744
rect 358412 266704 358418 266716
rect 360838 266704 360844 266716
rect 360896 266704 360902 266756
rect 388162 266704 388168 266756
rect 388220 266744 388226 266756
rect 396258 266744 396264 266756
rect 388220 266716 396264 266744
rect 388220 266704 388226 266716
rect 396258 266704 396264 266716
rect 396316 266704 396322 266756
rect 412174 266704 412180 266756
rect 412232 266744 412238 266756
rect 412232 266716 412634 266744
rect 412232 266704 412238 266716
rect 330202 266636 330208 266688
rect 330260 266676 330266 266688
rect 334618 266676 334624 266688
rect 330260 266648 334624 266676
rect 330260 266636 330266 266648
rect 334618 266636 334624 266648
rect 334676 266636 334682 266688
rect 138658 266568 138664 266620
rect 138716 266608 138722 266620
rect 138716 266580 145328 266608
rect 138716 266568 138722 266580
rect 119798 266432 119804 266484
rect 119856 266472 119862 266484
rect 144914 266472 144920 266484
rect 119856 266444 144920 266472
rect 119856 266432 119862 266444
rect 144914 266432 144920 266444
rect 144972 266432 144978 266484
rect 145300 266404 145328 266580
rect 149054 266568 149060 266620
rect 149112 266608 149118 266620
rect 179506 266608 179512 266620
rect 149112 266580 179512 266608
rect 149112 266568 149118 266580
rect 179506 266568 179512 266580
rect 179564 266568 179570 266620
rect 208670 266568 208676 266620
rect 208728 266608 208734 266620
rect 210970 266608 210976 266620
rect 208728 266580 210976 266608
rect 208728 266568 208734 266580
rect 210970 266568 210976 266580
rect 211028 266568 211034 266620
rect 213822 266568 213828 266620
rect 213880 266608 213886 266620
rect 220078 266608 220084 266620
rect 213880 266580 220084 266608
rect 213880 266568 213886 266580
rect 220078 266568 220084 266580
rect 220136 266568 220142 266620
rect 360838 266568 360844 266620
rect 360896 266608 360902 266620
rect 362218 266608 362224 266620
rect 360896 266580 362224 266608
rect 360896 266568 360902 266580
rect 362218 266568 362224 266580
rect 362276 266568 362282 266620
rect 412606 266608 412634 266716
rect 417970 266704 417976 266756
rect 418028 266744 418034 266756
rect 428458 266744 428464 266756
rect 418028 266716 428464 266744
rect 418028 266704 418034 266716
rect 428458 266704 428464 266716
rect 428516 266704 428522 266756
rect 430390 266704 430396 266756
rect 430448 266744 430454 266756
rect 431926 266744 431954 266852
rect 451228 266840 451234 266852
rect 451286 266840 451292 266892
rect 456426 266840 456432 266892
rect 456484 266880 456490 266892
rect 469214 266880 469220 266892
rect 456484 266852 469220 266880
rect 456484 266840 456490 266852
rect 469214 266840 469220 266852
rect 469272 266840 469278 266892
rect 470134 266840 470140 266892
rect 470192 266880 470198 266892
rect 470192 266852 519032 266880
rect 470192 266840 470198 266852
rect 453298 266812 453304 266824
rect 451384 266784 453304 266812
rect 430448 266716 431954 266744
rect 430448 266704 430454 266716
rect 432046 266704 432052 266756
rect 432104 266744 432110 266756
rect 446398 266744 446404 266756
rect 432104 266716 446404 266744
rect 432104 266704 432110 266716
rect 446398 266704 446404 266716
rect 446456 266704 446462 266756
rect 449434 266704 449440 266756
rect 449492 266744 449498 266756
rect 449492 266716 451274 266744
rect 449492 266704 449498 266716
rect 451246 266676 451274 266716
rect 451384 266676 451412 266784
rect 453298 266772 453304 266784
rect 453356 266772 453362 266824
rect 455230 266772 455236 266824
rect 455288 266812 455294 266824
rect 455288 266784 456012 266812
rect 455288 266772 455294 266784
rect 455984 266744 456012 266784
rect 512914 266744 512920 266756
rect 455984 266716 512920 266744
rect 512914 266704 512920 266716
rect 512972 266704 512978 266756
rect 513374 266704 513380 266756
rect 513432 266744 513438 266756
rect 515490 266744 515496 266756
rect 513432 266716 515496 266744
rect 513432 266704 513438 266716
rect 515490 266704 515496 266716
rect 515548 266704 515554 266756
rect 516502 266704 516508 266756
rect 516560 266744 516566 266756
rect 518710 266744 518716 266756
rect 516560 266716 518716 266744
rect 516560 266704 516566 266716
rect 518710 266704 518716 266716
rect 518768 266704 518774 266756
rect 519004 266744 519032 266852
rect 519170 266840 519176 266892
rect 519228 266880 519234 266892
rect 533982 266880 533988 266892
rect 519228 266852 533988 266880
rect 519228 266840 519234 266852
rect 533982 266840 533988 266852
rect 534040 266840 534046 266892
rect 534166 266840 534172 266892
rect 534224 266880 534230 266892
rect 537202 266880 537208 266892
rect 534224 266852 537208 266880
rect 534224 266840 534230 266852
rect 537202 266840 537208 266852
rect 537260 266840 537266 266892
rect 537386 266840 537392 266892
rect 537444 266880 537450 266892
rect 539502 266880 539508 266892
rect 537444 266852 539508 266880
rect 537444 266840 537450 266852
rect 539502 266840 539508 266852
rect 539560 266840 539566 266892
rect 539686 266840 539692 266892
rect 539744 266880 539750 266892
rect 580258 266880 580264 266892
rect 539744 266852 580264 266880
rect 539744 266840 539750 266852
rect 580258 266840 580264 266852
rect 580316 266840 580322 266892
rect 524368 266744 524374 266756
rect 519004 266716 524374 266744
rect 524368 266704 524374 266716
rect 524426 266704 524432 266756
rect 524506 266704 524512 266756
rect 524564 266744 524570 266756
rect 613378 266744 613384 266756
rect 524564 266716 613384 266744
rect 524564 266704 524570 266716
rect 613378 266704 613384 266716
rect 613436 266704 613442 266756
rect 451246 266648 451412 266676
rect 452746 266636 452752 266688
rect 452804 266676 452810 266688
rect 455782 266676 455788 266688
rect 452804 266648 455788 266676
rect 452804 266636 452810 266648
rect 455782 266636 455788 266648
rect 455840 266636 455846 266688
rect 421558 266608 421564 266620
rect 412606 266580 421564 266608
rect 421558 266568 421564 266580
rect 421616 266568 421622 266620
rect 422938 266568 422944 266620
rect 422996 266608 423002 266620
rect 439314 266608 439320 266620
rect 422996 266580 439320 266608
rect 422996 266568 423002 266580
rect 439314 266568 439320 266580
rect 439372 266568 439378 266620
rect 439498 266568 439504 266620
rect 439556 266608 439562 266620
rect 439556 266580 443316 266608
rect 439556 266568 439562 266580
rect 145558 266500 145564 266552
rect 145616 266540 145622 266552
rect 148870 266540 148876 266552
rect 145616 266512 148876 266540
rect 145616 266500 145622 266512
rect 148870 266500 148876 266512
rect 148928 266500 148934 266552
rect 240686 266500 240692 266552
rect 240744 266540 240750 266552
rect 245746 266540 245752 266552
rect 240744 266512 245752 266540
rect 240744 266500 240750 266512
rect 245746 266500 245752 266512
rect 245804 266500 245810 266552
rect 308674 266500 308680 266552
rect 308732 266540 308738 266552
rect 310882 266540 310888 266552
rect 308732 266512 310888 266540
rect 308732 266500 308738 266512
rect 310882 266500 310888 266512
rect 310940 266500 310946 266552
rect 311158 266500 311164 266552
rect 311216 266540 311222 266552
rect 313274 266540 313280 266552
rect 311216 266512 313280 266540
rect 311216 266500 311222 266512
rect 313274 266500 313280 266512
rect 313332 266500 313338 266552
rect 327718 266500 327724 266552
rect 327776 266540 327782 266552
rect 332318 266540 332324 266552
rect 327776 266512 332324 266540
rect 327776 266500 327782 266512
rect 332318 266500 332324 266512
rect 332376 266500 332382 266552
rect 346762 266500 346768 266552
rect 346820 266540 346826 266552
rect 351638 266540 351644 266552
rect 346820 266512 351644 266540
rect 346820 266500 346826 266512
rect 351638 266500 351644 266512
rect 351696 266500 351702 266552
rect 355042 266500 355048 266552
rect 355100 266540 355106 266552
rect 358998 266540 359004 266552
rect 355100 266512 359004 266540
rect 355100 266500 355106 266512
rect 358998 266500 359004 266512
rect 359056 266500 359062 266552
rect 394786 266500 394792 266552
rect 394844 266540 394850 266552
rect 398098 266540 398104 266552
rect 394844 266512 398104 266540
rect 394844 266500 394850 266512
rect 398098 266500 398104 266512
rect 398156 266500 398162 266552
rect 151078 266432 151084 266484
rect 151136 266472 151142 266484
rect 172882 266472 172888 266484
rect 151136 266444 172888 266472
rect 151136 266432 151142 266444
rect 172882 266432 172888 266444
rect 172940 266432 172946 266484
rect 361666 266432 361672 266484
rect 361724 266472 361730 266484
rect 362770 266472 362776 266484
rect 361724 266444 362776 266472
rect 361724 266432 361730 266444
rect 362770 266432 362776 266444
rect 362828 266432 362834 266484
rect 427906 266432 427912 266484
rect 427964 266472 427970 266484
rect 427964 266444 431954 266472
rect 427964 266432 427970 266444
rect 147214 266404 147220 266416
rect 145300 266376 147220 266404
rect 147214 266364 147220 266376
rect 147272 266364 147278 266416
rect 148318 266364 148324 266416
rect 148376 266404 148382 266416
rect 149698 266404 149704 266416
rect 148376 266376 149704 266404
rect 148376 266364 148382 266376
rect 149698 266364 149704 266376
rect 149756 266364 149762 266416
rect 182174 266364 182180 266416
rect 182232 266404 182238 266416
rect 186130 266404 186136 266416
rect 182232 266376 186136 266404
rect 182232 266364 182238 266376
rect 186130 266364 186136 266376
rect 186188 266364 186194 266416
rect 202138 266364 202144 266416
rect 202196 266404 202202 266416
rect 206830 266404 206836 266416
rect 202196 266376 206836 266404
rect 202196 266364 202202 266376
rect 206830 266364 206836 266376
rect 206888 266364 206894 266416
rect 222838 266364 222844 266416
rect 222896 266404 222902 266416
rect 224218 266404 224224 266416
rect 222896 266376 224224 266404
rect 222896 266364 222902 266376
rect 224218 266364 224224 266376
rect 224276 266364 224282 266416
rect 230750 266364 230756 266416
rect 230808 266404 230814 266416
rect 236638 266404 236644 266416
rect 230808 266376 236644 266404
rect 230808 266364 230814 266376
rect 236638 266364 236644 266376
rect 236696 266364 236702 266416
rect 242250 266364 242256 266416
rect 242308 266404 242314 266416
rect 243262 266404 243268 266416
rect 242308 266376 243268 266404
rect 242308 266364 242314 266376
rect 243262 266364 243268 266376
rect 243320 266364 243326 266416
rect 252002 266364 252008 266416
rect 252060 266404 252066 266416
rect 257338 266404 257344 266416
rect 252060 266376 257344 266404
rect 252060 266364 252066 266376
rect 257338 266364 257344 266376
rect 257396 266364 257402 266416
rect 263318 266364 263324 266416
rect 263376 266404 263382 266416
rect 265618 266404 265624 266416
rect 263376 266376 265624 266404
rect 263376 266364 263382 266376
rect 265618 266364 265624 266376
rect 265676 266364 265682 266416
rect 269114 266364 269120 266416
rect 269172 266404 269178 266416
rect 276382 266404 276388 266416
rect 269172 266376 276388 266404
rect 269172 266364 269178 266376
rect 276382 266364 276388 266376
rect 276440 266364 276446 266416
rect 278590 266364 278596 266416
rect 278648 266404 278654 266416
rect 286318 266404 286324 266416
rect 278648 266376 286324 266404
rect 278648 266364 278654 266376
rect 286318 266364 286324 266376
rect 286376 266364 286382 266416
rect 290458 266364 290464 266416
rect 290516 266404 290522 266416
rect 292942 266404 292948 266416
rect 290516 266376 292948 266404
rect 290516 266364 290522 266376
rect 292942 266364 292948 266376
rect 293000 266364 293006 266416
rect 297910 266364 297916 266416
rect 297968 266404 297974 266416
rect 299566 266404 299572 266416
rect 297968 266376 299572 266404
rect 297968 266364 297974 266376
rect 299566 266364 299572 266376
rect 299624 266364 299630 266416
rect 301038 266364 301044 266416
rect 301096 266404 301102 266416
rect 302050 266404 302056 266416
rect 301096 266376 302056 266404
rect 301096 266364 301102 266376
rect 302050 266364 302056 266376
rect 302108 266364 302114 266416
rect 307846 266364 307852 266416
rect 307904 266404 307910 266416
rect 309502 266404 309508 266416
rect 307904 266376 309508 266404
rect 307904 266364 307910 266376
rect 309502 266364 309508 266376
rect 309560 266364 309566 266416
rect 310330 266364 310336 266416
rect 310388 266404 310394 266416
rect 311894 266404 311900 266416
rect 310388 266376 311900 266404
rect 310388 266364 310394 266376
rect 311894 266364 311900 266376
rect 311952 266364 311958 266416
rect 312354 266364 312360 266416
rect 312412 266404 312418 266416
rect 314654 266404 314660 266416
rect 312412 266376 314660 266404
rect 312412 266364 312418 266376
rect 314654 266364 314660 266376
rect 314712 266364 314718 266416
rect 317782 266364 317788 266416
rect 317840 266404 317846 266416
rect 323118 266404 323124 266416
rect 317840 266376 323124 266404
rect 317840 266364 317846 266376
rect 323118 266364 323124 266376
rect 323176 266364 323182 266416
rect 328546 266364 328552 266416
rect 328604 266404 328610 266416
rect 329466 266404 329472 266416
rect 328604 266376 329472 266404
rect 328604 266364 328610 266376
rect 329466 266364 329472 266376
rect 329524 266364 329530 266416
rect 332686 266364 332692 266416
rect 332744 266404 332750 266416
rect 333882 266404 333888 266416
rect 332744 266376 333888 266404
rect 332744 266364 332750 266376
rect 333882 266364 333888 266376
rect 333940 266364 333946 266416
rect 340966 266364 340972 266416
rect 341024 266404 341030 266416
rect 342162 266404 342168 266416
rect 341024 266376 342168 266404
rect 341024 266364 341030 266376
rect 342162 266364 342168 266376
rect 342220 266364 342226 266416
rect 345106 266364 345112 266416
rect 345164 266404 345170 266416
rect 346302 266404 346308 266416
rect 345164 266376 346308 266404
rect 345164 266364 345170 266376
rect 346302 266364 346308 266376
rect 346360 266364 346366 266416
rect 349246 266364 349252 266416
rect 349304 266404 349310 266416
rect 350258 266404 350264 266416
rect 349304 266376 350264 266404
rect 349304 266364 349310 266376
rect 350258 266364 350264 266376
rect 350316 266364 350322 266416
rect 357526 266364 357532 266416
rect 357584 266404 357590 266416
rect 358630 266404 358636 266416
rect 357584 266376 358636 266404
rect 357584 266364 357590 266376
rect 358630 266364 358636 266376
rect 358688 266364 358694 266416
rect 367462 266364 367468 266416
rect 367520 266404 367526 266416
rect 368382 266404 368388 266416
rect 367520 266376 368388 266404
rect 367520 266364 367526 266376
rect 368382 266364 368388 266376
rect 368440 266364 368446 266416
rect 371602 266364 371608 266416
rect 371660 266404 371666 266416
rect 372522 266404 372528 266416
rect 371660 266376 372528 266404
rect 371660 266364 371666 266376
rect 372522 266364 372528 266376
rect 372580 266364 372586 266416
rect 374086 266364 374092 266416
rect 374144 266404 374150 266416
rect 375098 266404 375104 266416
rect 374144 266376 375104 266404
rect 374144 266364 374150 266376
rect 375098 266364 375104 266376
rect 375156 266364 375162 266416
rect 379882 266364 379888 266416
rect 379940 266404 379946 266416
rect 380710 266404 380716 266416
rect 379940 266376 380716 266404
rect 379940 266364 379946 266376
rect 380710 266364 380716 266376
rect 380768 266364 380774 266416
rect 386506 266364 386512 266416
rect 386564 266404 386570 266416
rect 387702 266404 387708 266416
rect 386564 266376 387708 266404
rect 386564 266364 386570 266376
rect 387702 266364 387708 266376
rect 387760 266364 387766 266416
rect 396442 266364 396448 266416
rect 396500 266404 396506 266416
rect 397270 266404 397276 266416
rect 396500 266376 397276 266404
rect 396500 266364 396506 266376
rect 397270 266364 397276 266376
rect 397328 266364 397334 266416
rect 398926 266364 398932 266416
rect 398984 266404 398990 266416
rect 400122 266404 400128 266416
rect 398984 266376 400128 266404
rect 398984 266364 398990 266376
rect 400122 266364 400128 266376
rect 400180 266364 400186 266416
rect 408862 266364 408868 266416
rect 408920 266404 408926 266416
rect 409782 266404 409788 266416
rect 408920 266376 409788 266404
rect 408920 266364 408926 266376
rect 409782 266364 409788 266376
rect 409840 266364 409846 266416
rect 411346 266364 411352 266416
rect 411404 266404 411410 266416
rect 412450 266404 412456 266416
rect 411404 266376 412456 266404
rect 411404 266364 411410 266376
rect 412450 266364 412456 266376
rect 412508 266364 412514 266416
rect 415486 266364 415492 266416
rect 415544 266404 415550 266416
rect 416406 266404 416412 266416
rect 415544 266376 416412 266404
rect 415544 266364 415550 266376
rect 416406 266364 416412 266376
rect 416464 266364 416470 266416
rect 423766 266364 423772 266416
rect 423824 266404 423830 266416
rect 424962 266404 424968 266416
rect 423824 266376 424968 266404
rect 423824 266364 423830 266376
rect 424962 266364 424968 266376
rect 425020 266364 425026 266416
rect 425422 266364 425428 266416
rect 425480 266404 425486 266416
rect 426894 266404 426900 266416
rect 425480 266376 426900 266404
rect 425480 266364 425486 266376
rect 426894 266364 426900 266376
rect 426952 266364 426958 266416
rect 431926 266404 431954 266444
rect 432046 266404 432052 266416
rect 431926 266376 432052 266404
rect 432046 266364 432052 266376
rect 432104 266364 432110 266416
rect 432322 266364 432328 266416
rect 432380 266404 432386 266416
rect 433150 266404 433156 266416
rect 432380 266376 433156 266404
rect 432380 266364 432386 266376
rect 433150 266364 433156 266376
rect 433208 266364 433214 266416
rect 433702 266364 433708 266416
rect 433760 266404 433766 266416
rect 434622 266404 434628 266416
rect 433760 266376 434628 266404
rect 433760 266364 433766 266376
rect 434622 266364 434628 266376
rect 434680 266364 434686 266416
rect 437014 266364 437020 266416
rect 437072 266404 437078 266416
rect 440878 266404 440884 266416
rect 437072 266376 440884 266404
rect 437072 266364 437078 266376
rect 440878 266364 440884 266376
rect 440936 266364 440942 266416
rect 441982 266364 441988 266416
rect 442040 266404 442046 266416
rect 442902 266404 442908 266416
rect 442040 266376 442908 266404
rect 442040 266364 442046 266376
rect 442902 266364 442908 266376
rect 442960 266364 442966 266416
rect 443288 266404 443316 266580
rect 459186 266568 459192 266620
rect 459244 266608 459250 266620
rect 464154 266608 464160 266620
rect 459244 266580 464160 266608
rect 459244 266568 459250 266580
rect 464154 266568 464160 266580
rect 464212 266568 464218 266620
rect 464338 266568 464344 266620
rect 464396 266608 464402 266620
rect 465718 266608 465724 266620
rect 464396 266580 465724 266608
rect 464396 266568 464402 266580
rect 465718 266568 465724 266580
rect 465776 266568 465782 266620
rect 469306 266568 469312 266620
rect 469364 266608 469370 266620
rect 473262 266608 473268 266620
rect 469364 266580 473268 266608
rect 469364 266568 469370 266580
rect 473262 266568 473268 266580
rect 473320 266568 473326 266620
rect 473446 266568 473452 266620
rect 473504 266608 473510 266620
rect 474642 266608 474648 266620
rect 473504 266580 474648 266608
rect 473504 266568 473510 266580
rect 474642 266568 474648 266580
rect 474700 266568 474706 266620
rect 474826 266568 474832 266620
rect 474884 266608 474890 266620
rect 478138 266608 478144 266620
rect 474884 266580 478144 266608
rect 474884 266568 474890 266580
rect 478138 266568 478144 266580
rect 478196 266568 478202 266620
rect 481726 266568 481732 266620
rect 481784 266608 481790 266620
rect 485222 266608 485228 266620
rect 481784 266580 485228 266608
rect 481784 266568 481790 266580
rect 485222 266568 485228 266580
rect 485280 266568 485286 266620
rect 485866 266568 485872 266620
rect 485924 266608 485930 266620
rect 487062 266608 487068 266620
rect 485924 266580 487068 266608
rect 485924 266568 485930 266580
rect 487062 266568 487068 266580
rect 487120 266568 487126 266620
rect 490006 266568 490012 266620
rect 490064 266608 490070 266620
rect 490064 266580 536328 266608
rect 490064 266568 490070 266580
rect 444466 266500 444472 266552
rect 444524 266540 444530 266552
rect 447778 266540 447784 266552
rect 444524 266512 447784 266540
rect 444524 266500 444530 266512
rect 447778 266500 447784 266512
rect 447836 266500 447842 266552
rect 454402 266500 454408 266552
rect 454460 266540 454466 266552
rect 457438 266540 457444 266552
rect 454460 266512 457444 266540
rect 454460 266500 454466 266512
rect 457438 266500 457444 266512
rect 457496 266500 457502 266552
rect 536300 266540 536328 266580
rect 543688 266568 543694 266620
rect 543746 266608 543752 266620
rect 553026 266608 553032 266620
rect 543746 266580 553032 266608
rect 543746 266568 543752 266580
rect 553026 266568 553032 266580
rect 553084 266568 553090 266620
rect 536300 266512 543596 266540
rect 460198 266432 460204 266484
rect 460256 266472 460262 266484
rect 460256 266444 512224 266472
rect 460256 266432 460262 266444
rect 445018 266404 445024 266416
rect 443288 266376 445024 266404
rect 445018 266364 445024 266376
rect 445076 266364 445082 266416
rect 447778 266364 447784 266416
rect 447836 266404 447842 266416
rect 449158 266404 449164 266416
rect 447836 266376 449164 266404
rect 447836 266364 447842 266376
rect 449158 266364 449164 266376
rect 449216 266364 449222 266416
rect 451918 266364 451924 266416
rect 451976 266404 451982 266416
rect 454678 266404 454684 266416
rect 451976 266376 454684 266404
rect 451976 266364 451982 266376
rect 454678 266364 454684 266376
rect 454736 266364 454742 266416
rect 456886 266364 456892 266416
rect 456944 266404 456950 266416
rect 458082 266404 458088 266416
rect 456944 266376 458088 266404
rect 456944 266364 456950 266376
rect 458082 266364 458088 266376
rect 458140 266364 458146 266416
rect 458542 266364 458548 266416
rect 458600 266404 458606 266416
rect 459370 266404 459376 266416
rect 458600 266376 459376 266404
rect 458600 266364 458606 266376
rect 459370 266364 459376 266376
rect 459428 266364 459434 266416
rect 498562 266296 498568 266348
rect 498620 266336 498626 266348
rect 501598 266336 501604 266348
rect 498620 266308 501604 266336
rect 498620 266296 498626 266308
rect 501598 266296 501604 266308
rect 501656 266296 501662 266348
rect 512196 266268 512224 266444
rect 517330 266432 517336 266484
rect 517388 266472 517394 266484
rect 543568 266472 543596 266512
rect 549622 266472 549628 266484
rect 517388 266444 534074 266472
rect 543568 266444 549628 266472
rect 517388 266432 517394 266444
rect 512362 266364 512368 266416
rect 512420 266404 512426 266416
rect 512420 266376 514708 266404
rect 512420 266364 512426 266376
rect 513374 266268 513380 266280
rect 512196 266240 513380 266268
rect 513374 266228 513380 266240
rect 513432 266228 513438 266280
rect 514680 266268 514708 266376
rect 514846 266364 514852 266416
rect 514904 266404 514910 266416
rect 516778 266404 516784 266416
rect 514904 266376 516784 266404
rect 514904 266364 514910 266376
rect 516778 266364 516784 266376
rect 516836 266364 516842 266416
rect 534046 266404 534074 266444
rect 549622 266432 549628 266444
rect 549680 266432 549686 266484
rect 534046 266376 543504 266404
rect 520274 266336 520280 266348
rect 518866 266308 520280 266336
rect 518866 266268 518894 266308
rect 520274 266296 520280 266308
rect 520332 266296 520338 266348
rect 522666 266296 522672 266348
rect 522724 266336 522730 266348
rect 524506 266336 524512 266348
rect 522724 266308 524512 266336
rect 522724 266296 522730 266308
rect 524506 266296 524512 266308
rect 524564 266296 524570 266348
rect 543476 266336 543504 266376
rect 546402 266336 546408 266348
rect 543476 266308 546408 266336
rect 546402 266296 546408 266308
rect 546460 266296 546466 266348
rect 514680 266240 518894 266268
rect 475102 266024 475108 266076
rect 475160 266064 475166 266076
rect 547874 266064 547880 266076
rect 475160 266036 547880 266064
rect 475160 266024 475166 266036
rect 547874 266024 547880 266036
rect 547932 266024 547938 266076
rect 485038 265888 485044 265940
rect 485096 265928 485102 265940
rect 561674 265928 561680 265940
rect 485096 265900 561680 265928
rect 485096 265888 485102 265900
rect 561674 265888 561680 265900
rect 561732 265888 561738 265940
rect 494974 265752 494980 265804
rect 495032 265792 495038 265804
rect 575566 265792 575572 265804
rect 495032 265764 575572 265792
rect 495032 265752 495038 265764
rect 575566 265752 575572 265764
rect 575624 265752 575630 265804
rect 187694 265616 187700 265668
rect 187752 265656 187758 265668
rect 188246 265656 188252 265668
rect 187752 265628 188252 265656
rect 187752 265616 187758 265628
rect 188246 265616 188252 265628
rect 188304 265616 188310 265668
rect 247126 265616 247132 265668
rect 247184 265656 247190 265668
rect 247862 265656 247868 265668
rect 247184 265628 247868 265656
rect 247184 265616 247190 265628
rect 247862 265616 247868 265628
rect 247920 265616 247926 265668
rect 259546 265616 259552 265668
rect 259604 265656 259610 265668
rect 260374 265656 260380 265668
rect 259604 265628 260380 265656
rect 259604 265616 259610 265628
rect 260374 265616 260380 265628
rect 260432 265616 260438 265668
rect 284294 265616 284300 265668
rect 284352 265656 284358 265668
rect 285214 265656 285220 265668
rect 284352 265628 285220 265656
rect 284352 265616 284358 265628
rect 285214 265616 285220 265628
rect 285272 265616 285278 265668
rect 480070 265616 480076 265668
rect 480128 265656 480134 265668
rect 554774 265656 554780 265668
rect 480128 265628 554780 265656
rect 480128 265616 480134 265628
rect 554774 265616 554780 265628
rect 554832 265616 554838 265668
rect 558178 265616 558184 265668
rect 558236 265656 558242 265668
rect 647234 265656 647240 265668
rect 558236 265628 647240 265656
rect 558236 265616 558242 265628
rect 647234 265616 647240 265628
rect 647292 265616 647298 265668
rect 570598 261468 570604 261520
rect 570656 261508 570662 261520
rect 645854 261508 645860 261520
rect 570656 261480 645860 261508
rect 570656 261468 570662 261480
rect 645854 261468 645860 261480
rect 645912 261468 645918 261520
rect 554406 260856 554412 260908
rect 554464 260896 554470 260908
rect 568574 260896 568580 260908
rect 554464 260868 568580 260896
rect 554464 260856 554470 260868
rect 568574 260856 568580 260868
rect 568632 260856 568638 260908
rect 554314 259428 554320 259480
rect 554372 259468 554378 259480
rect 567838 259468 567844 259480
rect 554372 259440 567844 259468
rect 554372 259428 554378 259440
rect 567838 259428 567844 259440
rect 567896 259428 567902 259480
rect 35802 256708 35808 256760
rect 35860 256748 35866 256760
rect 40678 256748 40684 256760
rect 35860 256720 40684 256748
rect 35860 256708 35866 256720
rect 40678 256708 40684 256720
rect 40736 256708 40742 256760
rect 553946 256708 553952 256760
rect 554004 256748 554010 256760
rect 562318 256748 562324 256760
rect 554004 256720 562324 256748
rect 554004 256708 554010 256720
rect 562318 256708 562324 256720
rect 562376 256708 562382 256760
rect 554498 253376 554504 253428
rect 554556 253416 554562 253428
rect 559558 253416 559564 253428
rect 554556 253388 559564 253416
rect 554556 253376 554562 253388
rect 559558 253376 559564 253388
rect 559616 253376 559622 253428
rect 35618 252832 35624 252884
rect 35676 252872 35682 252884
rect 41690 252872 41696 252884
rect 35676 252844 41696 252872
rect 35676 252832 35682 252844
rect 41690 252832 41696 252844
rect 41748 252832 41754 252884
rect 35802 252696 35808 252748
rect 35860 252736 35866 252748
rect 40678 252736 40684 252748
rect 35860 252708 40684 252736
rect 35860 252696 35866 252708
rect 40678 252696 40684 252708
rect 40736 252696 40742 252748
rect 35434 252560 35440 252612
rect 35492 252600 35498 252612
rect 41690 252600 41696 252612
rect 35492 252572 41696 252600
rect 35492 252560 35498 252572
rect 41690 252560 41696 252572
rect 41748 252560 41754 252612
rect 675846 252220 675852 252272
rect 675904 252260 675910 252272
rect 678238 252260 678244 252272
rect 675904 252232 678244 252260
rect 675904 252220 675910 252232
rect 678238 252220 678244 252232
rect 678296 252220 678302 252272
rect 675846 251540 675852 251592
rect 675904 251580 675910 251592
rect 678422 251580 678428 251592
rect 675904 251552 678428 251580
rect 675904 251540 675910 251552
rect 678422 251540 678428 251552
rect 678480 251540 678486 251592
rect 35802 251200 35808 251252
rect 35860 251240 35866 251252
rect 36538 251240 36544 251252
rect 35860 251212 36544 251240
rect 35860 251200 35866 251212
rect 36538 251200 36544 251212
rect 36596 251200 36602 251252
rect 553486 251200 553492 251252
rect 553544 251240 553550 251252
rect 555418 251240 555424 251252
rect 553544 251212 555424 251240
rect 553544 251200 553550 251212
rect 555418 251200 555424 251212
rect 555476 251200 555482 251252
rect 553670 249024 553676 249076
rect 553728 249064 553734 249076
rect 571334 249064 571340 249076
rect 553728 249036 571340 249064
rect 553728 249024 553734 249036
rect 571334 249024 571340 249036
rect 571392 249024 571398 249076
rect 553854 246304 553860 246356
rect 553912 246344 553918 246356
rect 632698 246344 632704 246356
rect 553912 246316 632704 246344
rect 553912 246304 553918 246316
rect 632698 246304 632704 246316
rect 632756 246304 632762 246356
rect 554406 245624 554412 245676
rect 554464 245664 554470 245676
rect 591298 245664 591304 245676
rect 554464 245636 591304 245664
rect 554464 245624 554470 245636
rect 591298 245624 591304 245636
rect 591356 245624 591362 245676
rect 554498 244264 554504 244316
rect 554556 244304 554562 244316
rect 624418 244304 624424 244316
rect 554556 244276 624424 244304
rect 554556 244264 554562 244276
rect 624418 244264 624424 244276
rect 624476 244264 624482 244316
rect 36538 242836 36544 242888
rect 36596 242876 36602 242888
rect 41690 242876 41696 242888
rect 36596 242848 41696 242876
rect 36596 242836 36602 242848
rect 41690 242836 41696 242848
rect 41748 242836 41754 242888
rect 576118 242156 576124 242208
rect 576176 242196 576182 242208
rect 648614 242196 648620 242208
rect 576176 242168 648620 242196
rect 576176 242156 576182 242168
rect 648614 242156 648620 242168
rect 648672 242156 648678 242208
rect 553946 241476 553952 241528
rect 554004 241516 554010 241528
rect 628558 241516 628564 241528
rect 554004 241488 628564 241516
rect 554004 241476 554010 241488
rect 628558 241476 628564 241488
rect 628616 241476 628622 241528
rect 553854 240116 553860 240168
rect 553912 240156 553918 240168
rect 577498 240156 577504 240168
rect 553912 240128 577504 240156
rect 553912 240116 553918 240128
rect 577498 240116 577504 240128
rect 577556 240116 577562 240168
rect 554314 238688 554320 238740
rect 554372 238728 554378 238740
rect 576118 238728 576124 238740
rect 554372 238700 576124 238728
rect 554372 238688 554378 238700
rect 576118 238688 576124 238700
rect 576176 238688 576182 238740
rect 672166 238008 672172 238060
rect 672224 238048 672230 238060
rect 672756 238048 672784 238102
rect 672224 238020 672784 238048
rect 672224 238008 672230 238020
rect 672874 237776 672902 237898
rect 672756 237748 672902 237776
rect 671246 237600 671252 237652
rect 671304 237640 671310 237652
rect 672756 237640 672784 237748
rect 672966 237640 672994 237694
rect 671304 237612 672784 237640
rect 672874 237612 672994 237640
rect 671304 237600 671310 237612
rect 672874 237572 672902 237612
rect 672828 237544 672902 237572
rect 668762 237396 668768 237448
rect 668820 237436 668826 237448
rect 672828 237436 672856 237544
rect 668820 237408 672856 237436
rect 668820 237396 668826 237408
rect 671430 237124 671436 237176
rect 671488 237164 671494 237176
rect 673104 237164 673132 237490
rect 671488 237136 673132 237164
rect 671488 237124 671494 237136
rect 673196 237028 673224 237286
rect 673304 237108 673356 237114
rect 673304 237050 673356 237056
rect 673104 237000 673224 237028
rect 671614 236920 671620 236972
rect 671672 236960 671678 236972
rect 673104 236960 673132 237000
rect 671672 236932 673132 236960
rect 671672 236920 671678 236932
rect 673414 236904 673466 236910
rect 673414 236846 673466 236852
rect 673528 236700 673580 236706
rect 673528 236642 673580 236648
rect 673408 236444 673414 236496
rect 673466 236484 673472 236496
rect 673466 236456 673670 236484
rect 673466 236444 673472 236456
rect 673752 236292 673804 236298
rect 673752 236234 673804 236240
rect 672626 236104 672632 236156
rect 672684 236144 672690 236156
rect 672684 236116 673900 236144
rect 672684 236104 672690 236116
rect 554498 236036 554504 236088
rect 554556 236076 554562 236088
rect 558178 236076 558184 236088
rect 554556 236048 558184 236076
rect 554556 236036 554562 236048
rect 558178 236036 558184 236048
rect 558236 236036 558242 236088
rect 673886 235912 673992 235940
rect 671062 235832 671068 235884
rect 671120 235872 671126 235884
rect 673886 235872 673914 235912
rect 671120 235844 673914 235872
rect 671120 235832 671126 235844
rect 672994 235696 673000 235748
rect 673052 235736 673058 235748
rect 673052 235708 674114 235736
rect 673052 235696 673058 235708
rect 669774 235492 669780 235544
rect 669832 235532 669838 235544
rect 669832 235504 674222 235532
rect 669832 235492 669838 235504
rect 668118 235288 668124 235340
rect 668176 235328 668182 235340
rect 668176 235300 674338 235328
rect 668176 235288 668182 235300
rect 591298 235220 591304 235272
rect 591356 235260 591362 235272
rect 633618 235260 633624 235272
rect 591356 235232 633624 235260
rect 591356 235220 591362 235232
rect 633618 235220 633624 235232
rect 633676 235220 633682 235272
rect 674438 234796 674466 235110
rect 674420 234744 674426 234796
rect 674478 234744 674484 234796
rect 672534 234608 672540 234660
rect 672592 234648 672598 234660
rect 674548 234648 674576 234906
rect 672592 234620 674576 234648
rect 672592 234608 672598 234620
rect 554406 234540 554412 234592
rect 554464 234580 554470 234592
rect 570598 234580 570604 234592
rect 554464 234552 570604 234580
rect 554464 234540 554470 234552
rect 570598 234540 570604 234552
rect 570656 234540 570662 234592
rect 674668 234444 674696 234702
rect 675846 234540 675852 234592
rect 675904 234580 675910 234592
rect 679618 234580 679624 234592
rect 675904 234552 679624 234580
rect 675904 234540 675910 234552
rect 679618 234540 679624 234552
rect 679676 234540 679682 234592
rect 673960 234416 674696 234444
rect 669590 234200 669596 234252
rect 669648 234240 669654 234252
rect 673960 234240 673988 234416
rect 669648 234212 673988 234240
rect 669648 234200 669654 234212
rect 674558 234200 674564 234252
rect 674616 234240 674622 234252
rect 674760 234240 674788 234498
rect 675846 234336 675852 234388
rect 675904 234376 675910 234388
rect 679986 234376 679992 234388
rect 675904 234348 679992 234376
rect 675904 234336 675910 234348
rect 679986 234336 679992 234348
rect 680044 234336 680050 234388
rect 674886 234320 674938 234326
rect 674886 234262 674938 234268
rect 674616 234212 674788 234240
rect 674616 234200 674622 234212
rect 675846 234200 675852 234252
rect 675904 234240 675910 234252
rect 679802 234240 679808 234252
rect 675904 234212 679808 234240
rect 675904 234200 675910 234212
rect 679802 234200 679808 234212
rect 679860 234200 679866 234252
rect 674978 234116 675030 234122
rect 674978 234058 675030 234064
rect 670786 233996 670792 234048
rect 670844 234036 670850 234048
rect 671798 234036 671804 234048
rect 670844 234008 671804 234036
rect 670844 233996 670850 234008
rect 671798 233996 671804 234008
rect 671856 233996 671862 234048
rect 675096 233912 675148 233918
rect 675096 233854 675148 233860
rect 669130 233588 669136 233640
rect 669188 233628 669194 233640
rect 675248 233628 675276 233682
rect 675846 233656 675852 233708
rect 675904 233696 675910 233708
rect 677778 233696 677784 233708
rect 675904 233668 677784 233696
rect 675904 233656 675910 233668
rect 677778 233656 677784 233668
rect 677836 233656 677842 233708
rect 669188 233600 675276 233628
rect 669188 233588 669194 233600
rect 671798 233316 671804 233368
rect 671856 233356 671862 233368
rect 671856 233328 674788 233356
rect 671856 233316 671862 233328
rect 674760 233220 674788 233328
rect 675358 233220 675386 233478
rect 676030 233384 676036 233436
rect 676088 233424 676094 233436
rect 683482 233424 683488 233436
rect 676088 233396 683488 233424
rect 676088 233384 676094 233396
rect 683482 233384 683488 233396
rect 683540 233384 683546 233436
rect 674760 233192 675386 233220
rect 671154 232976 671160 233028
rect 671212 233016 671218 233028
rect 674742 233016 674748 233028
rect 671212 232988 674748 233016
rect 671212 232976 671218 232988
rect 674742 232976 674748 232988
rect 674800 232976 674806 233028
rect 670878 232772 670884 232824
rect 670936 232812 670942 232824
rect 675018 232812 675024 232824
rect 670936 232784 675024 232812
rect 670936 232772 670942 232784
rect 675018 232772 675024 232784
rect 675076 232772 675082 232824
rect 652018 232500 652024 232552
rect 652076 232540 652082 232552
rect 675478 232540 675484 232552
rect 652076 232512 675484 232540
rect 652076 232500 652082 232512
rect 675478 232500 675484 232512
rect 675536 232500 675542 232552
rect 675846 232500 675852 232552
rect 675904 232540 675910 232552
rect 680170 232540 680176 232552
rect 675904 232512 680176 232540
rect 675904 232500 675910 232512
rect 680170 232500 680176 232512
rect 680228 232500 680234 232552
rect 662322 232364 662328 232416
rect 662380 232404 662386 232416
rect 662380 232376 663794 232404
rect 662380 232364 662386 232376
rect 663766 232336 663794 232376
rect 675340 232336 675346 232348
rect 663766 232308 675346 232336
rect 675340 232296 675346 232308
rect 675398 232296 675404 232348
rect 665082 232160 665088 232212
rect 665140 232200 665146 232212
rect 665140 232172 675556 232200
rect 665140 232160 665146 232172
rect 675346 232076 675398 232082
rect 673914 232024 673920 232076
rect 673972 232064 673978 232076
rect 674558 232064 674564 232076
rect 673972 232036 674564 232064
rect 673972 232024 673978 232036
rect 674558 232024 674564 232036
rect 674616 232024 674622 232076
rect 675346 232018 675398 232024
rect 675180 231804 675232 231810
rect 675180 231746 675232 231752
rect 675070 231600 675122 231606
rect 675070 231542 675122 231548
rect 674956 231328 675008 231334
rect 674956 231270 675008 231276
rect 675846 231208 675852 231260
rect 675904 231248 675910 231260
rect 677594 231248 677600 231260
rect 675904 231220 677600 231248
rect 675904 231208 675910 231220
rect 677594 231208 677600 231220
rect 677652 231208 677658 231260
rect 674840 231192 674892 231198
rect 674840 231134 674892 231140
rect 673546 231004 673552 231056
rect 673604 231044 673610 231056
rect 674558 231044 674564 231056
rect 673604 231016 674564 231044
rect 673604 231004 673610 231016
rect 674558 231004 674564 231016
rect 674616 231004 674622 231056
rect 674732 230920 674784 230926
rect 674732 230862 674784 230868
rect 673454 230800 673460 230852
rect 673512 230840 673518 230852
rect 673512 230812 674636 230840
rect 673512 230800 673518 230812
rect 158254 230704 158260 230716
rect 157306 230676 158260 230704
rect 144638 230528 144644 230580
rect 144696 230568 144702 230580
rect 150526 230568 150532 230580
rect 144696 230540 150532 230568
rect 144696 230528 144702 230540
rect 150526 230528 150532 230540
rect 150584 230528 150590 230580
rect 150894 230528 150900 230580
rect 150952 230568 150958 230580
rect 157306 230568 157334 230676
rect 158254 230664 158260 230676
rect 158312 230664 158318 230716
rect 150952 230540 157334 230568
rect 157536 230540 158760 230568
rect 150952 230528 150958 230540
rect 90358 230392 90364 230444
rect 90416 230432 90422 230444
rect 157536 230432 157564 230540
rect 90416 230404 157564 230432
rect 158732 230432 158760 230540
rect 165430 230528 165436 230580
rect 165488 230568 165494 230580
rect 172054 230568 172060 230580
rect 165488 230540 172060 230568
rect 165488 230528 165494 230540
rect 172054 230528 172060 230540
rect 172112 230528 172118 230580
rect 176102 230528 176108 230580
rect 176160 230568 176166 230580
rect 181070 230568 181076 230580
rect 176160 230540 181076 230568
rect 176160 230528 176166 230540
rect 181070 230528 181076 230540
rect 181128 230528 181134 230580
rect 439314 230528 439320 230580
rect 439372 230568 439378 230580
rect 439372 230540 439544 230568
rect 439372 230528 439378 230540
rect 161106 230432 161112 230444
rect 158732 230404 161112 230432
rect 90416 230392 90422 230404
rect 161106 230392 161112 230404
rect 161164 230392 161170 230444
rect 161290 230392 161296 230444
rect 161348 230432 161354 230444
rect 215202 230432 215208 230444
rect 161348 230404 215208 230432
rect 161348 230392 161354 230404
rect 215202 230392 215208 230404
rect 215260 230392 215266 230444
rect 223390 230392 223396 230444
rect 223448 230432 223454 230444
rect 271874 230432 271880 230444
rect 223448 230404 271880 230432
rect 223448 230392 223454 230404
rect 271874 230392 271880 230404
rect 271932 230392 271938 230444
rect 274174 230392 274180 230444
rect 274232 230432 274238 230444
rect 307938 230432 307944 230444
rect 274232 230404 307944 230432
rect 274232 230392 274238 230404
rect 307938 230392 307944 230404
rect 307996 230392 308002 230444
rect 312538 230392 312544 230444
rect 312596 230432 312602 230444
rect 315666 230432 315672 230444
rect 312596 230404 315672 230432
rect 312596 230392 312602 230404
rect 315666 230392 315672 230404
rect 315724 230392 315730 230444
rect 377398 230392 377404 230444
rect 377456 230432 377462 230444
rect 378778 230432 378784 230444
rect 377456 230404 378784 230432
rect 377456 230392 377462 230404
rect 378778 230392 378784 230404
rect 378836 230392 378842 230444
rect 439516 230432 439544 230540
rect 674006 230528 674012 230580
rect 674064 230568 674070 230580
rect 674064 230528 674098 230568
rect 440694 230432 440700 230444
rect 439516 230404 440700 230432
rect 440694 230392 440700 230404
rect 440752 230392 440758 230444
rect 441890 230392 441896 230444
rect 441948 230432 441954 230444
rect 443454 230432 443460 230444
rect 441948 230404 443460 230432
rect 441948 230392 441954 230404
rect 443454 230392 443460 230404
rect 443512 230392 443518 230444
rect 468294 230392 468300 230444
rect 468352 230432 468358 230444
rect 469030 230432 469036 230444
rect 468352 230404 469036 230432
rect 468352 230392 468358 230404
rect 469030 230392 469036 230404
rect 469088 230392 469094 230444
rect 534626 230392 534632 230444
rect 534684 230432 534690 230444
rect 544194 230432 544200 230444
rect 534684 230404 544200 230432
rect 534684 230392 534690 230404
rect 544194 230392 544200 230404
rect 544252 230392 544258 230444
rect 669314 230392 669320 230444
rect 669372 230432 669378 230444
rect 673914 230432 673920 230444
rect 669372 230404 673920 230432
rect 669372 230392 669378 230404
rect 673914 230392 673920 230404
rect 673972 230392 673978 230444
rect 674070 230432 674098 230528
rect 674518 230512 674570 230518
rect 674518 230454 674570 230460
rect 674070 230404 674422 230432
rect 404262 230324 404268 230376
rect 404320 230364 404326 230376
rect 412266 230364 412272 230376
rect 404320 230336 412272 230364
rect 404320 230324 404326 230336
rect 412266 230324 412272 230336
rect 412324 230324 412330 230376
rect 436094 230324 436100 230376
rect 436152 230364 436158 230376
rect 436738 230364 436744 230376
rect 436152 230336 436744 230364
rect 436152 230324 436158 230336
rect 436738 230324 436744 230336
rect 436796 230324 436802 230376
rect 438670 230324 438676 230376
rect 438728 230364 438734 230376
rect 439314 230364 439320 230376
rect 438728 230336 439320 230364
rect 438728 230324 438734 230336
rect 439314 230324 439320 230336
rect 439372 230324 439378 230376
rect 443822 230324 443828 230376
rect 443880 230364 443886 230376
rect 444834 230364 444840 230376
rect 443880 230336 444840 230364
rect 443880 230324 443886 230336
rect 444834 230324 444840 230336
rect 444892 230324 444898 230376
rect 446398 230324 446404 230376
rect 446456 230364 446462 230376
rect 449158 230364 449164 230376
rect 446456 230336 449164 230364
rect 446456 230324 446462 230336
rect 449158 230324 449164 230336
rect 449216 230324 449222 230376
rect 449618 230324 449624 230376
rect 449676 230364 449682 230376
rect 450538 230364 450544 230376
rect 449676 230336 450544 230364
rect 449676 230324 449682 230336
rect 450538 230324 450544 230336
rect 450596 230324 450602 230376
rect 452838 230324 452844 230376
rect 452896 230364 452902 230376
rect 454310 230364 454316 230376
rect 452896 230336 454316 230364
rect 452896 230324 452902 230336
rect 454310 230324 454316 230336
rect 454368 230324 454374 230376
rect 455414 230324 455420 230376
rect 455472 230364 455478 230376
rect 457162 230364 457168 230376
rect 455472 230336 457168 230364
rect 455472 230324 455478 230336
rect 457162 230324 457168 230336
rect 457220 230324 457226 230376
rect 463786 230324 463792 230376
rect 463844 230364 463850 230376
rect 465718 230364 465724 230376
rect 463844 230336 465724 230364
rect 463844 230324 463850 230336
rect 465718 230324 465724 230336
rect 465776 230324 465782 230376
rect 475378 230324 475384 230376
rect 475436 230364 475442 230376
rect 478322 230364 478328 230376
rect 475436 230336 478328 230364
rect 475436 230324 475442 230336
rect 478322 230324 478328 230336
rect 478380 230324 478386 230376
rect 480530 230324 480536 230376
rect 480588 230364 480594 230376
rect 481542 230364 481548 230376
rect 480588 230336 481548 230364
rect 480588 230324 480594 230336
rect 481542 230324 481548 230336
rect 481600 230324 481606 230376
rect 492766 230324 492772 230376
rect 492824 230364 492830 230376
rect 493962 230364 493968 230376
rect 492824 230336 493968 230364
rect 492824 230324 492830 230336
rect 493962 230324 493968 230336
rect 494020 230324 494026 230376
rect 494698 230324 494704 230376
rect 494756 230364 494762 230376
rect 496354 230364 496360 230376
rect 494756 230336 496360 230364
rect 494756 230324 494762 230336
rect 496354 230324 496360 230336
rect 496412 230324 496418 230376
rect 499850 230324 499856 230376
rect 499908 230364 499914 230376
rect 501138 230364 501144 230376
rect 499908 230336 501144 230364
rect 499908 230324 499914 230336
rect 501138 230324 501144 230336
rect 501196 230324 501202 230376
rect 503714 230324 503720 230376
rect 503772 230364 503778 230376
rect 506934 230364 506940 230376
rect 503772 230336 506940 230364
rect 503772 230324 503778 230336
rect 506934 230324 506940 230336
rect 506992 230324 506998 230376
rect 516594 230324 516600 230376
rect 516652 230364 516658 230376
rect 517422 230364 517428 230376
rect 516652 230336 517428 230364
rect 516652 230324 516658 230336
rect 517422 230324 517428 230336
rect 517480 230324 517486 230376
rect 520458 230324 520464 230376
rect 520516 230364 520522 230376
rect 521562 230364 521568 230376
rect 520516 230336 521568 230364
rect 520516 230324 520522 230336
rect 521562 230324 521568 230336
rect 521620 230324 521626 230376
rect 526898 230324 526904 230376
rect 526956 230364 526962 230376
rect 527818 230364 527824 230376
rect 526956 230336 527824 230364
rect 526956 230324 526962 230336
rect 527818 230324 527824 230336
rect 527876 230324 527882 230376
rect 118418 230256 118424 230308
rect 118476 230296 118482 230308
rect 189442 230296 189448 230308
rect 118476 230268 189448 230296
rect 118476 230256 118482 230268
rect 189442 230256 189448 230268
rect 189500 230256 189506 230308
rect 190914 230256 190920 230308
rect 190972 230296 190978 230308
rect 202322 230296 202328 230308
rect 190972 230268 202328 230296
rect 190972 230256 190978 230268
rect 202322 230256 202328 230268
rect 202380 230256 202386 230308
rect 203702 230256 203708 230308
rect 203760 230296 203766 230308
rect 256418 230296 256424 230308
rect 203760 230268 256424 230296
rect 203760 230256 203766 230268
rect 256418 230256 256424 230268
rect 256476 230256 256482 230308
rect 261386 230256 261392 230308
rect 261444 230296 261450 230308
rect 297634 230296 297640 230308
rect 261444 230268 297640 230296
rect 261444 230256 261450 230268
rect 297634 230256 297640 230268
rect 297692 230256 297698 230308
rect 302878 230256 302884 230308
rect 302936 230296 302942 230308
rect 305362 230296 305368 230308
rect 302936 230268 305368 230296
rect 302936 230256 302942 230268
rect 305362 230256 305368 230268
rect 305420 230256 305426 230308
rect 307846 230256 307852 230308
rect 307904 230296 307910 230308
rect 323394 230296 323400 230308
rect 307904 230268 323400 230296
rect 307904 230256 307910 230268
rect 323394 230256 323400 230268
rect 323452 230256 323458 230308
rect 497918 230256 497924 230308
rect 497976 230296 497982 230308
rect 499666 230296 499672 230308
rect 497976 230268 499672 230296
rect 497976 230256 497982 230268
rect 499666 230256 499672 230268
rect 499724 230256 499730 230308
rect 518728 230268 519032 230296
rect 408862 230188 408868 230240
rect 408920 230228 408926 230240
rect 410978 230228 410984 230240
rect 408920 230200 410984 230228
rect 408920 230188 408926 230200
rect 410978 230188 410984 230200
rect 411036 230188 411042 230240
rect 447042 230188 447048 230240
rect 447100 230228 447106 230240
rect 449894 230228 449900 230240
rect 447100 230200 449900 230228
rect 447100 230188 447106 230200
rect 449894 230188 449900 230200
rect 449952 230188 449958 230240
rect 451550 230188 451556 230240
rect 451608 230228 451614 230240
rect 453298 230228 453304 230240
rect 451608 230200 453304 230228
rect 451608 230188 451614 230200
rect 453298 230188 453304 230200
rect 453356 230188 453362 230240
rect 454126 230188 454132 230240
rect 454184 230228 454190 230240
rect 455230 230228 455236 230240
rect 454184 230200 455236 230228
rect 454184 230188 454190 230200
rect 455230 230188 455236 230200
rect 455288 230188 455294 230240
rect 470870 230188 470876 230240
rect 470928 230228 470934 230240
rect 471882 230228 471888 230240
rect 470928 230200 471888 230228
rect 470928 230188 470934 230200
rect 471882 230188 471888 230200
rect 471940 230188 471946 230240
rect 493410 230188 493416 230240
rect 493468 230228 493474 230240
rect 495158 230228 495164 230240
rect 493468 230200 495164 230228
rect 493468 230188 493474 230200
rect 495158 230188 495164 230200
rect 495216 230188 495222 230240
rect 513374 230188 513380 230240
rect 513432 230228 513438 230240
rect 515398 230228 515404 230240
rect 513432 230200 515404 230228
rect 513432 230188 513438 230200
rect 515398 230188 515404 230200
rect 515456 230188 515462 230240
rect 517238 230188 517244 230240
rect 517296 230228 517302 230240
rect 518728 230228 518756 230268
rect 517296 230200 518756 230228
rect 519004 230228 519032 230268
rect 529198 230256 529204 230308
rect 529256 230296 529262 230308
rect 541618 230296 541624 230308
rect 529256 230268 541624 230296
rect 529256 230256 529262 230268
rect 541618 230256 541624 230268
rect 541676 230256 541682 230308
rect 667934 230256 667940 230308
rect 667992 230296 667998 230308
rect 673822 230296 673828 230308
rect 667992 230268 673828 230296
rect 667992 230256 667998 230268
rect 673822 230256 673828 230268
rect 673880 230256 673886 230308
rect 522298 230228 522304 230240
rect 519004 230200 522304 230228
rect 517296 230188 517302 230200
rect 522298 230188 522304 230200
rect 522356 230188 522362 230240
rect 529014 230228 529020 230240
rect 522868 230200 529020 230228
rect 111058 230120 111064 230172
rect 111116 230160 111122 230172
rect 184290 230160 184296 230172
rect 111116 230132 184296 230160
rect 111116 230120 111122 230132
rect 184290 230120 184296 230132
rect 184348 230120 184354 230172
rect 191558 230160 191564 230172
rect 186286 230132 191564 230160
rect 88242 229984 88248 230036
rect 88300 230024 88306 230036
rect 166258 230024 166264 230036
rect 88300 229996 166264 230024
rect 88300 229984 88306 229996
rect 166258 229984 166264 229996
rect 166316 229984 166322 230036
rect 166442 229984 166448 230036
rect 166500 230024 166506 230036
rect 181714 230024 181720 230036
rect 166500 229996 181720 230024
rect 166500 229984 166506 229996
rect 181714 229984 181720 229996
rect 181772 229984 181778 230036
rect 184198 229984 184204 230036
rect 184256 230024 184262 230036
rect 186286 230024 186314 230132
rect 191558 230120 191564 230132
rect 191616 230120 191622 230172
rect 196986 230120 196992 230172
rect 197044 230160 197050 230172
rect 251266 230160 251272 230172
rect 197044 230132 251272 230160
rect 197044 230120 197050 230132
rect 251266 230120 251272 230132
rect 251324 230120 251330 230172
rect 276842 230120 276848 230172
rect 276900 230160 276906 230172
rect 313090 230160 313096 230172
rect 276900 230132 313096 230160
rect 276900 230120 276906 230132
rect 313090 230120 313096 230132
rect 313148 230120 313154 230172
rect 315298 230120 315304 230172
rect 315356 230160 315362 230172
rect 340138 230160 340144 230172
rect 315356 230132 340144 230160
rect 315356 230120 315362 230132
rect 340138 230120 340144 230132
rect 340196 230120 340202 230172
rect 476666 230120 476672 230172
rect 476724 230160 476730 230172
rect 479702 230160 479708 230172
rect 476724 230132 479708 230160
rect 476724 230120 476730 230132
rect 479702 230120 479708 230132
rect 479760 230120 479766 230172
rect 503254 230160 503260 230172
rect 499546 230132 503260 230160
rect 345658 230052 345664 230104
rect 345716 230092 345722 230104
rect 353018 230092 353024 230104
rect 345716 230064 353024 230092
rect 345716 230052 345722 230064
rect 353018 230052 353024 230064
rect 353076 230052 353082 230104
rect 444466 230052 444472 230104
rect 444524 230092 444530 230104
rect 447594 230092 447600 230104
rect 444524 230064 447600 230092
rect 444524 230052 444530 230064
rect 447594 230052 447600 230064
rect 447652 230052 447658 230104
rect 490834 230052 490840 230104
rect 490892 230092 490898 230104
rect 493778 230092 493784 230104
rect 490892 230064 493784 230092
rect 490892 230052 490898 230064
rect 493778 230052 493784 230064
rect 493836 230052 493842 230104
rect 494330 230052 494336 230104
rect 494388 230092 494394 230104
rect 499546 230092 499574 230132
rect 503254 230120 503260 230132
rect 503312 230120 503318 230172
rect 518820 230132 518940 230160
rect 494388 230064 499574 230092
rect 494388 230052 494394 230064
rect 515674 230052 515680 230104
rect 515732 230092 515738 230104
rect 518820 230092 518848 230132
rect 515732 230064 518848 230092
rect 518912 230092 518940 230132
rect 518912 230064 519032 230092
rect 515732 230052 515738 230064
rect 184256 229996 186314 230024
rect 184256 229984 184262 229996
rect 189718 229984 189724 230036
rect 189776 230024 189782 230036
rect 246114 230024 246120 230036
rect 189776 229996 246120 230024
rect 189776 229984 189782 229996
rect 246114 229984 246120 229996
rect 246172 229984 246178 230036
rect 251726 229984 251732 230036
rect 251784 230024 251790 230036
rect 292482 230024 292488 230036
rect 251784 229996 292488 230024
rect 251784 229984 251790 229996
rect 292482 229984 292488 229996
rect 292540 229984 292546 230036
rect 296898 229984 296904 230036
rect 296956 230024 296962 230036
rect 302510 230024 302516 230036
rect 296956 229996 302516 230024
rect 296956 229984 296962 229996
rect 302510 229984 302516 229996
rect 302568 229984 302574 230036
rect 305638 229984 305644 230036
rect 305696 230024 305702 230036
rect 334986 230024 334992 230036
rect 305696 229996 334992 230024
rect 305696 229984 305702 229996
rect 334986 229984 334992 229996
rect 335044 229984 335050 230036
rect 380434 229984 380440 230036
rect 380492 230024 380498 230036
rect 389082 230024 389088 230036
rect 380492 229996 389088 230024
rect 380492 229984 380498 229996
rect 389082 229984 389088 229996
rect 389140 229984 389146 230036
rect 468846 229984 468852 230036
rect 468904 230024 468910 230036
rect 475378 230024 475384 230036
rect 468904 229996 475384 230024
rect 468904 229984 468910 229996
rect 475378 229984 475384 229996
rect 475436 229984 475442 230036
rect 476022 229984 476028 230036
rect 476080 230024 476086 230036
rect 479518 230024 479524 230036
rect 476080 229996 479524 230024
rect 476080 229984 476086 229996
rect 479518 229984 479524 229996
rect 479576 229984 479582 230036
rect 483106 229984 483112 230036
rect 483164 230024 483170 230036
rect 484302 230024 484308 230036
rect 483164 229996 484308 230024
rect 483164 229984 483170 229996
rect 484302 229984 484308 229996
rect 484360 229984 484366 230036
rect 484762 229984 484768 230036
rect 484820 230024 484826 230036
rect 490650 230024 490656 230036
rect 484820 229996 490656 230024
rect 484820 229984 484826 229996
rect 490650 229984 490656 229996
rect 490708 229984 490714 230036
rect 499666 229984 499672 230036
rect 499724 230024 499730 230036
rect 504358 230024 504364 230036
rect 499724 229996 504364 230024
rect 499724 229984 499730 229996
rect 504358 229984 504364 229996
rect 504416 229984 504422 230036
rect 511442 229916 511448 229968
rect 511500 229956 511506 229968
rect 516778 229956 516784 229968
rect 511500 229928 516784 229956
rect 511500 229916 511506 229928
rect 516778 229916 516784 229928
rect 516836 229916 516842 229968
rect 74442 229848 74448 229900
rect 74500 229888 74506 229900
rect 155954 229888 155960 229900
rect 74500 229860 155960 229888
rect 74500 229848 74506 229860
rect 155954 229848 155960 229860
rect 156012 229848 156018 229900
rect 156322 229848 156328 229900
rect 156380 229888 156386 229900
rect 176562 229888 176568 229900
rect 156380 229860 176568 229888
rect 156380 229848 156386 229860
rect 176562 229848 176568 229860
rect 176620 229848 176626 229900
rect 177574 229848 177580 229900
rect 177632 229888 177638 229900
rect 177632 229860 191144 229888
rect 177632 229848 177638 229860
rect 67542 229712 67548 229764
rect 67600 229752 67606 229764
rect 144638 229752 144644 229764
rect 67600 229724 144644 229752
rect 67600 229712 67606 229724
rect 144638 229712 144644 229724
rect 144696 229712 144702 229764
rect 144822 229712 144828 229764
rect 144880 229752 144886 229764
rect 144880 229724 147168 229752
rect 144880 229712 144886 229724
rect 140038 229576 140044 229628
rect 140096 229616 140102 229628
rect 146938 229616 146944 229628
rect 140096 229588 146944 229616
rect 140096 229576 140102 229588
rect 146938 229576 146944 229588
rect 146996 229576 147002 229628
rect 147140 229616 147168 229724
rect 148594 229712 148600 229764
rect 148652 229752 148658 229764
rect 150894 229752 150900 229764
rect 148652 229724 150900 229752
rect 148652 229712 148658 229724
rect 150894 229712 150900 229724
rect 150952 229712 150958 229764
rect 151354 229712 151360 229764
rect 151412 229752 151418 229764
rect 190914 229752 190920 229764
rect 151412 229724 190920 229752
rect 151412 229712 151418 229724
rect 190914 229712 190920 229724
rect 190972 229712 190978 229764
rect 191116 229752 191144 229860
rect 191558 229848 191564 229900
rect 191616 229888 191622 229900
rect 240962 229888 240968 229900
rect 191616 229860 240968 229888
rect 191616 229848 191622 229860
rect 240962 229848 240968 229860
rect 241020 229848 241026 229900
rect 245654 229848 245660 229900
rect 245712 229888 245718 229900
rect 287330 229888 287336 229900
rect 245712 229860 287336 229888
rect 245712 229848 245718 229860
rect 287330 229848 287336 229860
rect 287388 229848 287394 229900
rect 300118 229848 300124 229900
rect 300176 229888 300182 229900
rect 329834 229888 329840 229900
rect 300176 229860 329840 229888
rect 300176 229848 300182 229860
rect 329834 229848 329840 229860
rect 329892 229848 329898 229900
rect 334250 229848 334256 229900
rect 334308 229888 334314 229900
rect 345290 229888 345296 229900
rect 334308 229860 345296 229888
rect 334308 229848 334314 229860
rect 345290 229848 345296 229860
rect 345348 229848 345354 229900
rect 352558 229848 352564 229900
rect 352616 229888 352622 229900
rect 358170 229888 358176 229900
rect 352616 229860 358176 229888
rect 352616 229848 352622 229860
rect 358170 229848 358176 229860
rect 358228 229848 358234 229900
rect 364150 229848 364156 229900
rect 364208 229888 364214 229900
rect 381354 229888 381360 229900
rect 364208 229860 381360 229888
rect 364208 229848 364214 229860
rect 381354 229848 381360 229860
rect 381412 229848 381418 229900
rect 384298 229848 384304 229900
rect 384356 229888 384362 229900
rect 394234 229888 394240 229900
rect 384356 229860 394240 229888
rect 384356 229848 384362 229860
rect 394234 229848 394240 229860
rect 394292 229848 394298 229900
rect 412450 229848 412456 229900
rect 412508 229888 412514 229900
rect 419350 229888 419356 229900
rect 412508 229860 419356 229888
rect 412508 229848 412514 229860
rect 419350 229848 419356 229860
rect 419408 229848 419414 229900
rect 467006 229848 467012 229900
rect 467064 229888 467070 229900
rect 473998 229888 474004 229900
rect 467064 229860 474004 229888
rect 467064 229848 467070 229860
rect 473998 229848 474004 229860
rect 474056 229848 474062 229900
rect 481818 229848 481824 229900
rect 481876 229888 481882 229900
rect 489914 229888 489920 229900
rect 481876 229860 489920 229888
rect 481876 229848 481882 229860
rect 489914 229848 489920 229860
rect 489972 229848 489978 229900
rect 495986 229848 495992 229900
rect 496044 229888 496050 229900
rect 509234 229888 509240 229900
rect 496044 229860 509240 229888
rect 496044 229848 496050 229860
rect 509234 229848 509240 229860
rect 509292 229848 509298 229900
rect 519004 229888 519032 230064
rect 519170 230052 519176 230104
rect 519228 230092 519234 230104
rect 522868 230092 522896 230200
rect 529014 230188 529020 230200
rect 529072 230188 529078 230240
rect 674052 230188 674058 230240
rect 674110 230228 674116 230240
rect 674110 230200 674314 230228
rect 674110 230188 674116 230200
rect 530762 230120 530768 230172
rect 530820 230160 530826 230172
rect 530820 230132 534948 230160
rect 530820 230120 530826 230132
rect 519228 230064 522896 230092
rect 519228 230052 519234 230064
rect 523034 229984 523040 230036
rect 523092 230024 523098 230036
rect 534718 230024 534724 230036
rect 523092 229996 534724 230024
rect 523092 229984 523098 229996
rect 534718 229984 534724 229996
rect 534776 229984 534782 230036
rect 534920 230024 534948 230132
rect 536558 230120 536564 230172
rect 536616 230160 536622 230172
rect 549254 230160 549260 230172
rect 536616 230132 549260 230160
rect 536616 230120 536622 230132
rect 549254 230120 549260 230132
rect 549312 230120 549318 230172
rect 673638 230052 673644 230104
rect 673696 230092 673702 230104
rect 673696 230064 674198 230092
rect 673696 230052 673702 230064
rect 547138 230024 547144 230036
rect 534920 229996 547144 230024
rect 547138 229984 547144 229996
rect 547196 229984 547202 230036
rect 555418 229984 555424 230036
rect 555476 230024 555482 230036
rect 569954 230024 569960 230036
rect 555476 229996 569960 230024
rect 555476 229984 555482 229996
rect 569954 229984 569960 229996
rect 570012 229984 570018 230036
rect 673942 229916 673948 229968
rect 674000 229916 674006 229968
rect 525518 229888 525524 229900
rect 519004 229860 525524 229888
rect 525518 229848 525524 229860
rect 525576 229848 525582 229900
rect 538490 229848 538496 229900
rect 538548 229888 538554 229900
rect 556798 229888 556804 229900
rect 538548 229860 556804 229888
rect 538548 229848 538554 229860
rect 556798 229848 556804 229860
rect 556856 229848 556862 229900
rect 433518 229780 433524 229832
rect 433576 229820 433582 229832
rect 434162 229820 434168 229832
rect 433576 229792 434168 229820
rect 433576 229780 433582 229792
rect 434162 229780 434168 229792
rect 434220 229780 434226 229832
rect 673960 229820 673988 229916
rect 675846 229848 675852 229900
rect 675904 229888 675910 229900
rect 676950 229888 676956 229900
rect 675904 229860 676956 229888
rect 675904 229848 675910 229860
rect 676950 229848 676956 229860
rect 677008 229848 677014 229900
rect 673960 229792 674084 229820
rect 235810 229752 235816 229764
rect 191116 229724 235816 229752
rect 235810 229712 235816 229724
rect 235868 229712 235874 229764
rect 236914 229712 236920 229764
rect 236972 229752 236978 229764
rect 282178 229752 282184 229764
rect 236972 229724 282184 229752
rect 236972 229712 236978 229724
rect 282178 229712 282184 229724
rect 282236 229712 282242 229764
rect 285306 229712 285312 229764
rect 285364 229752 285370 229764
rect 318242 229752 318248 229764
rect 285364 229724 318248 229752
rect 285364 229712 285370 229724
rect 318242 229712 318248 229724
rect 318300 229712 318306 229764
rect 324038 229712 324044 229764
rect 324096 229752 324102 229764
rect 350442 229752 350448 229764
rect 324096 229724 350448 229752
rect 324096 229712 324102 229724
rect 350442 229712 350448 229724
rect 350500 229712 350506 229764
rect 371050 229752 371056 229764
rect 354646 229724 371056 229752
rect 210050 229616 210056 229628
rect 147140 229588 210056 229616
rect 210050 229576 210056 229588
rect 210108 229576 210114 229628
rect 210234 229576 210240 229628
rect 210292 229616 210298 229628
rect 261570 229616 261576 229628
rect 210292 229588 261576 229616
rect 210292 229576 210298 229588
rect 261570 229576 261576 229588
rect 261628 229576 261634 229628
rect 350534 229576 350540 229628
rect 350592 229616 350598 229628
rect 354646 229616 354674 229724
rect 371050 229712 371056 229724
rect 371108 229712 371114 229764
rect 386506 229752 386512 229764
rect 373966 229724 386512 229752
rect 350592 229588 354674 229616
rect 350592 229576 350598 229588
rect 370958 229576 370964 229628
rect 371016 229616 371022 229628
rect 373966 229616 373994 229724
rect 386506 229712 386512 229724
rect 386564 229712 386570 229764
rect 386966 229712 386972 229764
rect 387024 229752 387030 229764
rect 396810 229752 396816 229764
rect 387024 229724 396816 229752
rect 387024 229712 387030 229724
rect 396810 229712 396816 229724
rect 396868 229712 396874 229764
rect 399846 229712 399852 229764
rect 399904 229752 399910 229764
rect 409690 229752 409696 229764
rect 399904 229724 409696 229752
rect 399904 229712 399910 229724
rect 409690 229712 409696 229724
rect 409748 229712 409754 229764
rect 411162 229712 411168 229764
rect 411220 229752 411226 229764
rect 417418 229752 417424 229764
rect 411220 229724 417424 229752
rect 411220 229712 411226 229724
rect 417418 229712 417424 229724
rect 417476 229712 417482 229764
rect 457346 229712 457352 229764
rect 457404 229752 457410 229764
rect 463878 229752 463884 229764
rect 457404 229724 463884 229752
rect 457404 229712 457410 229724
rect 463878 229712 463884 229724
rect 463936 229712 463942 229764
rect 465442 229712 465448 229764
rect 465500 229752 465506 229764
rect 467466 229752 467472 229764
rect 465500 229724 467472 229752
rect 465500 229712 465506 229724
rect 467466 229712 467472 229724
rect 467524 229712 467530 229764
rect 469582 229712 469588 229764
rect 469640 229752 469646 229764
rect 476758 229752 476764 229764
rect 469640 229724 476764 229752
rect 469640 229712 469646 229724
rect 476758 229712 476764 229724
rect 476816 229712 476822 229764
rect 479242 229712 479248 229764
rect 479300 229752 479306 229764
rect 484118 229752 484124 229764
rect 479300 229724 484124 229752
rect 479300 229712 479306 229724
rect 484118 229712 484124 229724
rect 484176 229712 484182 229764
rect 486326 229712 486332 229764
rect 486384 229752 486390 229764
rect 500218 229752 500224 229764
rect 486384 229724 500224 229752
rect 486384 229712 486390 229724
rect 500218 229712 500224 229724
rect 500276 229712 500282 229764
rect 505646 229712 505652 229764
rect 505704 229752 505710 229764
rect 516042 229752 516048 229764
rect 505704 229724 516048 229752
rect 505704 229712 505710 229724
rect 516042 229712 516048 229724
rect 516100 229712 516106 229764
rect 518894 229752 518900 229764
rect 518866 229712 518900 229752
rect 518952 229712 518958 229764
rect 521102 229712 521108 229764
rect 521160 229752 521166 229764
rect 529934 229752 529940 229764
rect 521160 229724 529940 229752
rect 521160 229712 521166 229724
rect 529934 229712 529940 229724
rect 529992 229712 529998 229764
rect 532694 229712 532700 229764
rect 532752 229752 532758 229764
rect 555602 229752 555608 229764
rect 532752 229724 555608 229752
rect 532752 229712 532758 229724
rect 555602 229712 555608 229724
rect 555660 229712 555666 229764
rect 371016 229588 373994 229616
rect 371016 229576 371022 229588
rect 490650 229576 490656 229628
rect 490708 229616 490714 229628
rect 497458 229616 497464 229628
rect 490708 229588 497464 229616
rect 490708 229576 490714 229588
rect 497458 229576 497464 229588
rect 497516 229576 497522 229628
rect 509510 229576 509516 229628
rect 509568 229616 509574 229628
rect 518866 229616 518894 229712
rect 666830 229644 666836 229696
rect 666888 229684 666894 229696
rect 666888 229656 673974 229684
rect 666888 229644 666894 229656
rect 509568 229588 518894 229616
rect 509568 229576 509574 229588
rect 524966 229576 524972 229628
rect 525024 229616 525030 229628
rect 532418 229616 532424 229628
rect 525024 229588 532424 229616
rect 525024 229576 525030 229588
rect 532418 229576 532424 229588
rect 532476 229576 532482 229628
rect 675846 229576 675852 229628
rect 675904 229616 675910 229628
rect 677134 229616 677140 229628
rect 675904 229588 677140 229616
rect 675904 229576 675910 229588
rect 677134 229576 677140 229588
rect 677192 229576 677198 229628
rect 673828 229492 673880 229498
rect 131114 229440 131120 229492
rect 131172 229480 131178 229492
rect 197170 229480 197176 229492
rect 131172 229452 197176 229480
rect 131172 229440 131178 229452
rect 197170 229440 197176 229452
rect 197228 229440 197234 229492
rect 200206 229440 200212 229492
rect 200264 229480 200270 229492
rect 200758 229480 200764 229492
rect 200264 229452 200764 229480
rect 200264 229440 200270 229452
rect 200758 229440 200764 229452
rect 200816 229440 200822 229492
rect 231118 229440 231124 229492
rect 231176 229480 231182 229492
rect 277026 229480 277032 229492
rect 231176 229452 277032 229480
rect 231176 229440 231182 229452
rect 277026 229440 277032 229452
rect 277084 229440 277090 229492
rect 673828 229434 673880 229440
rect 448974 229372 448980 229424
rect 449032 229412 449038 229424
rect 451366 229412 451372 229424
rect 449032 229384 451372 229412
rect 449032 229372 449038 229384
rect 451366 229372 451372 229384
rect 451424 229372 451430 229424
rect 122926 229304 122932 229356
rect 122984 229344 122990 229356
rect 179138 229344 179144 229356
rect 122984 229316 179144 229344
rect 122984 229304 122990 229316
rect 179138 229304 179144 229316
rect 179196 229304 179202 229356
rect 181346 229304 181352 229356
rect 181404 229344 181410 229356
rect 230658 229344 230664 229356
rect 181404 229316 230664 229344
rect 181404 229304 181410 229316
rect 230658 229304 230664 229316
rect 230716 229304 230722 229356
rect 453482 229304 453488 229356
rect 453540 229344 453546 229356
rect 455782 229344 455788 229356
rect 453540 229316 455788 229344
rect 453540 229304 453546 229316
rect 455782 229304 455788 229316
rect 455840 229304 455846 229356
rect 673454 229304 673460 229356
rect 673512 229344 673518 229356
rect 673512 229316 673638 229344
rect 673512 229304 673518 229316
rect 358078 229236 358084 229288
rect 358136 229276 358142 229288
rect 360746 229276 360752 229288
rect 358136 229248 360752 229276
rect 358136 229236 358142 229248
rect 360746 229236 360752 229248
rect 360804 229236 360810 229288
rect 360930 229236 360936 229288
rect 360988 229276 360994 229288
rect 363322 229276 363328 229288
rect 360988 229248 363328 229276
rect 360988 229236 360994 229248
rect 363322 229236 363328 229248
rect 363380 229236 363386 229288
rect 419442 229236 419448 229288
rect 419500 229276 419506 229288
rect 424502 229276 424508 229288
rect 419500 229248 424508 229276
rect 419500 229236 419506 229248
rect 424502 229236 424508 229248
rect 424560 229236 424566 229288
rect 450262 229236 450268 229288
rect 450320 229276 450326 229288
rect 451826 229276 451832 229288
rect 450320 229248 451832 229276
rect 450320 229236 450326 229248
rect 451826 229236 451832 229248
rect 451884 229236 451890 229288
rect 479886 229236 479892 229288
rect 479944 229276 479950 229288
rect 482278 229276 482284 229288
rect 479944 229248 482284 229276
rect 479944 229236 479950 229248
rect 482278 229236 482284 229248
rect 482336 229236 482342 229288
rect 483750 229236 483756 229288
rect 483808 229276 483814 229288
rect 486786 229276 486792 229288
rect 483808 229248 486792 229276
rect 483808 229236 483814 229248
rect 486786 229236 486792 229248
rect 486844 229236 486850 229288
rect 501782 229236 501788 229288
rect 501840 229276 501846 229288
rect 507118 229276 507124 229288
rect 501840 229248 507124 229276
rect 501840 229236 501846 229248
rect 507118 229236 507124 229248
rect 507176 229236 507182 229288
rect 673610 229276 673638 229316
rect 675846 229304 675852 229356
rect 675904 229344 675910 229356
rect 677318 229344 677324 229356
rect 675904 229316 677324 229344
rect 675904 229304 675910 229316
rect 677318 229304 677324 229316
rect 677376 229304 677382 229356
rect 673610 229248 673762 229276
rect 92474 229168 92480 229220
rect 92532 229208 92538 229220
rect 146294 229208 146300 229220
rect 92532 229180 146300 229208
rect 92532 229168 92538 229180
rect 146294 229168 146300 229180
rect 146352 229168 146358 229220
rect 146938 229168 146944 229220
rect 146996 229208 147002 229220
rect 153378 229208 153384 229220
rect 146996 229180 153384 229208
rect 146996 229168 147002 229180
rect 153378 229168 153384 229180
rect 153436 229168 153442 229220
rect 153838 229168 153844 229220
rect 153896 229208 153902 229220
rect 163682 229208 163688 229220
rect 153896 229180 163688 229208
rect 153896 229168 153902 229180
rect 163682 229168 163688 229180
rect 163740 229168 163746 229220
rect 163866 229168 163872 229220
rect 163924 229208 163930 229220
rect 166442 229208 166448 229220
rect 163924 229180 166448 229208
rect 163924 229168 163930 229180
rect 166442 229168 166448 229180
rect 166500 229168 166506 229220
rect 166902 229168 166908 229220
rect 166960 229208 166966 229220
rect 172238 229208 172244 229220
rect 166960 229180 172244 229208
rect 166960 229168 166966 229180
rect 172238 229168 172244 229180
rect 172296 229168 172302 229220
rect 172422 229168 172428 229220
rect 172480 229208 172486 229220
rect 220354 229208 220360 229220
rect 172480 229180 220360 229208
rect 172480 229168 172486 229180
rect 220354 229168 220360 229180
rect 220412 229168 220418 229220
rect 378962 229100 378968 229152
rect 379020 229140 379026 229152
rect 383930 229140 383936 229152
rect 379020 229112 383936 229140
rect 379020 229100 379026 229112
rect 383930 229100 383936 229112
rect 383988 229100 383994 229152
rect 419994 229140 420000 229152
rect 418126 229112 420000 229140
rect 97902 229032 97908 229084
rect 97960 229072 97966 229084
rect 107286 229072 107292 229084
rect 97960 229044 107292 229072
rect 97960 229032 97966 229044
rect 107286 229032 107292 229044
rect 107344 229032 107350 229084
rect 107470 229032 107476 229084
rect 107528 229072 107534 229084
rect 107528 229044 167868 229072
rect 107528 229032 107534 229044
rect 102042 228896 102048 228948
rect 102100 228936 102106 228948
rect 166902 228936 166908 228948
rect 102100 228908 166908 228936
rect 102100 228896 102106 228908
rect 166902 228896 166908 228908
rect 166960 228896 166966 228948
rect 107102 228800 107108 228812
rect 84166 228772 107108 228800
rect 82078 228624 82084 228676
rect 82136 228664 82142 228676
rect 84166 228664 84194 228772
rect 107102 228760 107108 228772
rect 107160 228760 107166 228812
rect 107286 228760 107292 228812
rect 107344 228800 107350 228812
rect 166442 228800 166448 228812
rect 107344 228772 166448 228800
rect 107344 228760 107350 228772
rect 166442 228760 166448 228772
rect 166500 228760 166506 228812
rect 82136 228636 84194 228664
rect 82136 228624 82142 228636
rect 96246 228624 96252 228676
rect 96304 228664 96310 228676
rect 165430 228664 165436 228676
rect 96304 228636 165436 228664
rect 96304 228624 96310 228636
rect 165430 228624 165436 228636
rect 165488 228624 165494 228676
rect 167840 228664 167868 229044
rect 168190 229032 168196 229084
rect 168248 229072 168254 229084
rect 173986 229072 173992 229084
rect 168248 229044 173992 229072
rect 168248 229032 168254 229044
rect 173986 229032 173992 229044
rect 174044 229032 174050 229084
rect 174814 229032 174820 229084
rect 174872 229072 174878 229084
rect 174872 229044 181576 229072
rect 174872 229032 174878 229044
rect 172238 228896 172244 228948
rect 172296 228936 172302 228948
rect 175274 228936 175280 228948
rect 172296 228908 175280 228936
rect 172296 228896 172302 228908
rect 175274 228896 175280 228908
rect 175332 228896 175338 228948
rect 175642 228896 175648 228948
rect 175700 228936 175706 228948
rect 175700 228908 181484 228936
rect 175700 228896 175706 228908
rect 168006 228760 168012 228812
rect 168064 228800 168070 228812
rect 168064 228772 180012 228800
rect 168064 228760 168070 228772
rect 179984 228732 180012 228772
rect 181254 228732 181260 228744
rect 179984 228704 181260 228732
rect 181254 228692 181260 228704
rect 181312 228692 181318 228744
rect 179782 228664 179788 228676
rect 167840 228636 179788 228664
rect 179782 228624 179788 228636
rect 179840 228624 179846 228676
rect 181456 228664 181484 228908
rect 181548 228800 181576 229044
rect 181714 229032 181720 229084
rect 181772 229072 181778 229084
rect 192662 229072 192668 229084
rect 181772 229044 192668 229072
rect 181772 229032 181778 229044
rect 192662 229032 192668 229044
rect 192720 229032 192726 229084
rect 192846 229032 192852 229084
rect 192904 229072 192910 229084
rect 194594 229072 194600 229084
rect 192904 229044 194600 229072
rect 192904 229032 192910 229044
rect 194594 229032 194600 229044
rect 194652 229032 194658 229084
rect 195606 229032 195612 229084
rect 195664 229072 195670 229084
rect 250622 229072 250628 229084
rect 195664 229044 250628 229072
rect 195664 229032 195670 229044
rect 250622 229032 250628 229044
rect 250680 229032 250686 229084
rect 259270 229032 259276 229084
rect 259328 229072 259334 229084
rect 298278 229072 298284 229084
rect 259328 229044 298284 229072
rect 259328 229032 259334 229044
rect 298278 229032 298284 229044
rect 298336 229032 298342 229084
rect 413830 229032 413836 229084
rect 413888 229072 413894 229084
rect 418126 229072 418154 229112
rect 419994 229100 420000 229112
rect 420052 229100 420058 229152
rect 420178 229100 420184 229152
rect 420236 229140 420242 229152
rect 421926 229140 421932 229152
rect 420236 229112 421932 229140
rect 420236 229100 420242 229112
rect 421926 229100 421932 229112
rect 421984 229100 421990 229152
rect 424318 229100 424324 229152
rect 424376 229140 424382 229152
rect 427722 229140 427728 229152
rect 424376 229112 427728 229140
rect 424376 229100 424382 229112
rect 427722 229100 427728 229112
rect 427780 229100 427786 229152
rect 441246 229100 441252 229152
rect 441304 229140 441310 229152
rect 442074 229140 442080 229152
rect 441304 229112 442080 229140
rect 441304 229100 441310 229112
rect 442074 229100 442080 229112
rect 442132 229100 442138 229152
rect 450906 229100 450912 229152
rect 450964 229140 450970 229152
rect 452746 229140 452752 229152
rect 450964 229112 452752 229140
rect 450964 229100 450970 229112
rect 452746 229100 452752 229112
rect 452804 229100 452810 229152
rect 507578 229100 507584 229152
rect 507636 229140 507642 229152
rect 511258 229140 511264 229152
rect 507636 229112 511264 229140
rect 507636 229100 507642 229112
rect 511258 229100 511264 229112
rect 511316 229100 511322 229152
rect 673598 229084 673650 229090
rect 413888 229044 418154 229072
rect 413888 229032 413894 229044
rect 517882 229032 517888 229084
rect 517940 229072 517946 229084
rect 540514 229072 540520 229084
rect 517940 229044 540520 229072
rect 517940 229032 517946 229044
rect 540514 229032 540520 229044
rect 540572 229032 540578 229084
rect 675846 229032 675852 229084
rect 675904 229072 675910 229084
rect 676398 229072 676404 229084
rect 675904 229044 676404 229072
rect 675904 229032 675910 229044
rect 676398 229032 676404 229044
rect 676456 229032 676462 229084
rect 673598 229026 673650 229032
rect 181898 228896 181904 228948
rect 181956 228936 181962 228948
rect 237098 228936 237104 228948
rect 181956 228908 237104 228936
rect 181956 228896 181962 228908
rect 237098 228896 237104 228908
rect 237156 228896 237162 228948
rect 251082 228896 251088 228948
rect 251140 228936 251146 228948
rect 291194 228936 291200 228948
rect 251140 228908 291200 228936
rect 251140 228896 251146 228908
rect 291194 228896 291200 228908
rect 291252 228896 291258 228948
rect 319806 228896 319812 228948
rect 319864 228936 319870 228948
rect 345934 228936 345940 228948
rect 319864 228908 345940 228936
rect 319864 228896 319870 228908
rect 345934 228896 345940 228908
rect 345992 228896 345998 228948
rect 350166 228896 350172 228948
rect 350224 228936 350230 228948
rect 369118 228936 369124 228948
rect 350224 228908 369124 228936
rect 350224 228896 350230 228908
rect 369118 228896 369124 228908
rect 369176 228896 369182 228948
rect 507118 228896 507124 228948
rect 507176 228936 507182 228948
rect 520090 228936 520096 228948
rect 507176 228908 520096 228936
rect 507176 228896 507182 228908
rect 520090 228896 520096 228908
rect 520148 228896 520154 228948
rect 526254 228896 526260 228948
rect 526312 228936 526318 228948
rect 551554 228936 551560 228948
rect 526312 228908 551560 228936
rect 526312 228896 526318 228908
rect 551554 228896 551560 228908
rect 551612 228896 551618 228948
rect 673506 228880 673558 228886
rect 673506 228822 673558 228828
rect 190546 228800 190552 228812
rect 181548 228772 190552 228800
rect 190546 228760 190552 228772
rect 190604 228760 190610 228812
rect 190730 228760 190736 228812
rect 190788 228800 190794 228812
rect 241606 228800 241612 228812
rect 190788 228772 241612 228800
rect 190788 228760 190794 228772
rect 241606 228760 241612 228772
rect 241664 228760 241670 228812
rect 246298 228760 246304 228812
rect 246356 228800 246362 228812
rect 253842 228800 253848 228812
rect 246356 228772 253848 228800
rect 246356 228760 246362 228772
rect 253842 228760 253848 228772
rect 253900 228760 253906 228812
rect 255130 228760 255136 228812
rect 255188 228800 255194 228812
rect 295702 228800 295708 228812
rect 255188 228772 295708 228800
rect 255188 228760 255194 228772
rect 295702 228760 295708 228772
rect 295760 228760 295766 228812
rect 317966 228760 317972 228812
rect 318024 228800 318030 228812
rect 344646 228800 344652 228812
rect 318024 228772 344652 228800
rect 318024 228760 318030 228772
rect 344646 228760 344652 228772
rect 344704 228760 344710 228812
rect 346210 228760 346216 228812
rect 346268 228800 346274 228812
rect 366542 228800 366548 228812
rect 346268 228772 366548 228800
rect 346268 228760 346274 228772
rect 366542 228760 366548 228772
rect 366600 228760 366606 228812
rect 376570 228760 376576 228812
rect 376628 228800 376634 228812
rect 389726 228800 389732 228812
rect 376628 228772 389732 228800
rect 376628 228760 376634 228772
rect 389726 228760 389732 228772
rect 389784 228760 389790 228812
rect 401410 228760 401416 228812
rect 401468 228800 401474 228812
rect 408402 228800 408408 228812
rect 401468 228772 408408 228800
rect 401468 228760 401474 228772
rect 408402 228760 408408 228772
rect 408460 228760 408466 228812
rect 493778 228760 493784 228812
rect 493836 228800 493842 228812
rect 506014 228800 506020 228812
rect 493836 228772 506020 228800
rect 493836 228760 493842 228772
rect 506014 228760 506020 228772
rect 506072 228760 506078 228812
rect 519814 228760 519820 228812
rect 519872 228800 519878 228812
rect 543182 228800 543188 228812
rect 519872 228772 543188 228800
rect 519872 228760 519878 228772
rect 543182 228760 543188 228772
rect 543240 228760 543246 228812
rect 675846 228760 675852 228812
rect 675904 228800 675910 228812
rect 676214 228800 676220 228812
rect 675904 228772 676220 228800
rect 675904 228760 675910 228772
rect 676214 228760 676220 228772
rect 676272 228760 676278 228812
rect 231302 228664 231308 228676
rect 181456 228636 231308 228664
rect 231302 228624 231308 228636
rect 231360 228624 231366 228676
rect 239398 228624 239404 228676
rect 239456 228664 239462 228676
rect 284110 228664 284116 228676
rect 239456 228636 284116 228664
rect 239456 228624 239462 228636
rect 284110 228624 284116 228636
rect 284168 228624 284174 228676
rect 292390 228624 292396 228676
rect 292448 228664 292454 228676
rect 326614 228664 326620 228676
rect 292448 228636 326620 228664
rect 292448 228624 292454 228636
rect 326614 228624 326620 228636
rect 326672 228624 326678 228676
rect 333238 228624 333244 228676
rect 333296 228664 333302 228676
rect 355594 228664 355600 228676
rect 333296 228636 355600 228664
rect 333296 228624 333302 228636
rect 355594 228624 355600 228636
rect 355652 228624 355658 228676
rect 369762 228664 369768 228676
rect 359016 228636 369768 228664
rect 62758 228488 62764 228540
rect 62816 228528 62822 228540
rect 140774 228528 140780 228540
rect 62816 228500 140780 228528
rect 62816 228488 62822 228500
rect 140774 228488 140780 228500
rect 140832 228488 140838 228540
rect 140958 228488 140964 228540
rect 141016 228528 141022 228540
rect 141016 228500 149744 228528
rect 141016 228488 141022 228500
rect 66162 228352 66168 228404
rect 66220 228392 66226 228404
rect 147628 228392 147634 228404
rect 66220 228364 147634 228392
rect 66220 228352 66226 228364
rect 147628 228352 147634 228364
rect 147686 228352 147692 228404
rect 149716 228392 149744 228500
rect 153286 228488 153292 228540
rect 153344 228528 153350 228540
rect 200574 228528 200580 228540
rect 153344 228500 200580 228528
rect 153344 228488 153350 228500
rect 200574 228488 200580 228500
rect 200632 228488 200638 228540
rect 200758 228488 200764 228540
rect 200816 228528 200822 228540
rect 200816 228500 212672 228528
rect 200816 228488 200822 228500
rect 212644 228460 212672 228500
rect 219342 228488 219348 228540
rect 219400 228528 219406 228540
rect 267366 228528 267372 228540
rect 219400 228500 267372 228528
rect 219400 228488 219406 228500
rect 267366 228488 267372 228500
rect 267424 228488 267430 228540
rect 267550 228488 267556 228540
rect 267608 228528 267614 228540
rect 307294 228528 307300 228540
rect 267608 228500 307300 228528
rect 267608 228488 267614 228500
rect 307294 228488 307300 228500
rect 307352 228488 307358 228540
rect 307662 228488 307668 228540
rect 307720 228528 307726 228540
rect 335630 228528 335636 228540
rect 307720 228500 335636 228528
rect 307720 228488 307726 228500
rect 335630 228488 335636 228500
rect 335688 228488 335694 228540
rect 336642 228488 336648 228540
rect 336700 228528 336706 228540
rect 358814 228528 358820 228540
rect 336700 228500 358820 228528
rect 336700 228488 336706 228500
rect 358814 228488 358820 228500
rect 358872 228488 358878 228540
rect 212644 228432 214236 228460
rect 157426 228392 157432 228404
rect 149716 228364 157432 228392
rect 157426 228352 157432 228364
rect 157484 228352 157490 228404
rect 157794 228352 157800 228404
rect 157852 228392 157858 228404
rect 212166 228392 212172 228404
rect 157852 228364 212172 228392
rect 157852 228352 157858 228364
rect 212166 228352 212172 228364
rect 212224 228352 212230 228404
rect 214208 228392 214236 228432
rect 226150 228392 226156 228404
rect 214208 228364 226156 228392
rect 226150 228352 226156 228364
rect 226208 228352 226214 228404
rect 226334 228352 226340 228404
rect 226392 228392 226398 228404
rect 273806 228392 273812 228404
rect 226392 228364 273812 228392
rect 226392 228352 226398 228364
rect 273806 228352 273812 228364
rect 273864 228352 273870 228404
rect 284110 228352 284116 228404
rect 284168 228392 284174 228404
rect 320174 228392 320180 228404
rect 284168 228364 320180 228392
rect 284168 228352 284174 228364
rect 320174 228352 320180 228364
rect 320232 228352 320238 228404
rect 326890 228352 326896 228404
rect 326948 228392 326954 228404
rect 351086 228392 351092 228404
rect 326948 228364 351092 228392
rect 326948 228352 326954 228364
rect 351086 228352 351092 228364
rect 351144 228352 351150 228404
rect 355226 228352 355232 228404
rect 355284 228392 355290 228404
rect 359016 228392 359044 228636
rect 369762 228624 369768 228636
rect 369820 228624 369826 228676
rect 373810 228624 373816 228676
rect 373868 228664 373874 228676
rect 387242 228664 387248 228676
rect 373868 228636 387248 228664
rect 373868 228624 373874 228636
rect 387242 228624 387248 228636
rect 387300 228624 387306 228676
rect 390278 228624 390284 228676
rect 390336 228664 390342 228676
rect 400030 228664 400036 228676
rect 390336 228636 400036 228664
rect 390336 228624 390342 228636
rect 400030 228624 400036 228636
rect 400088 228624 400094 228676
rect 410886 228624 410892 228676
rect 410944 228664 410950 228676
rect 416130 228664 416136 228676
rect 410944 228636 416136 228664
rect 410944 228624 410950 228636
rect 416130 228624 416136 228636
rect 416188 228624 416194 228676
rect 478782 228624 478788 228676
rect 478840 228664 478846 228676
rect 483566 228664 483572 228676
rect 478840 228636 483572 228664
rect 478840 228624 478846 228636
rect 483566 228624 483572 228636
rect 483624 228624 483630 228676
rect 484118 228624 484124 228676
rect 484176 228664 484182 228676
rect 490558 228664 490564 228676
rect 484176 228636 490564 228664
rect 484176 228624 484182 228636
rect 490558 228624 490564 228636
rect 490616 228624 490622 228676
rect 495342 228624 495348 228676
rect 495400 228664 495406 228676
rect 511810 228664 511816 228676
rect 495400 228636 511816 228664
rect 495400 228624 495406 228636
rect 511810 228624 511816 228636
rect 511868 228624 511874 228676
rect 512086 228624 512092 228676
rect 512144 228664 512150 228676
rect 533522 228664 533528 228676
rect 512144 228636 533528 228664
rect 512144 228624 512150 228636
rect 533522 228624 533528 228636
rect 533580 228624 533586 228676
rect 533982 228624 533988 228676
rect 534040 228664 534046 228676
rect 561582 228664 561588 228676
rect 534040 228636 561588 228664
rect 534040 228624 534046 228636
rect 561582 228624 561588 228636
rect 561640 228624 561646 228676
rect 673388 228540 673440 228546
rect 366910 228488 366916 228540
rect 366968 228528 366974 228540
rect 381998 228528 382004 228540
rect 366968 228500 382004 228528
rect 366968 228488 366974 228500
rect 381998 228488 382004 228500
rect 382056 228488 382062 228540
rect 392946 228528 392952 228540
rect 383626 228500 392952 228528
rect 355284 228364 359044 228392
rect 355284 228352 355290 228364
rect 362862 228352 362868 228404
rect 362920 228392 362926 228404
rect 379422 228392 379428 228404
rect 362920 228364 379428 228392
rect 362920 228352 362926 228364
rect 379422 228352 379428 228364
rect 379480 228352 379486 228404
rect 381722 228352 381728 228404
rect 381780 228392 381786 228404
rect 383626 228392 383654 228500
rect 392946 228488 392952 228500
rect 393004 228488 393010 228540
rect 393222 228488 393228 228540
rect 393280 228528 393286 228540
rect 393280 228500 397960 228528
rect 393280 228488 393286 228500
rect 381780 228364 383654 228392
rect 381780 228352 381786 228364
rect 391842 228352 391848 228404
rect 391900 228392 391906 228404
rect 397932 228392 397960 228500
rect 400122 228488 400128 228540
rect 400180 228528 400186 228540
rect 407758 228528 407764 228540
rect 400180 228500 407764 228528
rect 400180 228488 400186 228500
rect 407758 228488 407764 228500
rect 407816 228488 407822 228540
rect 482462 228488 482468 228540
rect 482520 228528 482526 228540
rect 494606 228528 494612 228540
rect 482520 228500 494612 228528
rect 482520 228488 482526 228500
rect 494606 228488 494612 228500
rect 494664 228488 494670 228540
rect 502426 228488 502432 228540
rect 502484 228528 502490 228540
rect 520918 228528 520924 228540
rect 502484 228500 520924 228528
rect 502484 228488 502490 228500
rect 520918 228488 520924 228500
rect 520976 228488 520982 228540
rect 531406 228488 531412 228540
rect 531464 228528 531470 228540
rect 558178 228528 558184 228540
rect 531464 228500 558184 228528
rect 531464 228488 531470 228500
rect 558178 228488 558184 228500
rect 558236 228488 558242 228540
rect 673388 228482 673440 228488
rect 671798 228420 671804 228472
rect 671856 228460 671862 228472
rect 671856 228432 673302 228460
rect 671856 228420 671862 228432
rect 402606 228392 402612 228404
rect 391900 228364 393314 228392
rect 397932 228364 402612 228392
rect 391900 228352 391906 228364
rect 107102 228216 107108 228268
rect 107160 228256 107166 228268
rect 140958 228256 140964 228268
rect 107160 228228 140964 228256
rect 107160 228216 107166 228228
rect 140958 228216 140964 228228
rect 141016 228216 141022 228268
rect 141142 228216 141148 228268
rect 141200 228256 141206 228268
rect 190914 228256 190920 228268
rect 141200 228228 190920 228256
rect 141200 228216 141206 228228
rect 190914 228216 190920 228228
rect 190972 228216 190978 228268
rect 200758 228256 200764 228268
rect 191116 228228 200764 228256
rect 106182 228080 106188 228132
rect 106240 228120 106246 228132
rect 107470 228120 107476 228132
rect 106240 228092 107476 228120
rect 106240 228080 106246 228092
rect 107470 228080 107476 228092
rect 107528 228080 107534 228132
rect 112990 228080 112996 228132
rect 113048 228120 113054 228132
rect 113048 228092 181300 228120
rect 113048 228080 113054 228092
rect 122742 227944 122748 227996
rect 122800 227984 122806 227996
rect 181070 227984 181076 227996
rect 122800 227956 181076 227984
rect 122800 227944 122806 227956
rect 181070 227944 181076 227956
rect 181128 227944 181134 227996
rect 181272 227984 181300 228092
rect 181898 228080 181904 228132
rect 181956 228120 181962 228132
rect 191116 228120 191144 228228
rect 200758 228216 200764 228228
rect 200816 228216 200822 228268
rect 201402 228216 201408 228268
rect 201460 228256 201466 228268
rect 252554 228256 252560 228268
rect 201460 228228 252560 228256
rect 201460 228216 201466 228228
rect 252554 228216 252560 228228
rect 252612 228216 252618 228268
rect 277210 228216 277216 228268
rect 277268 228256 277274 228268
rect 311802 228256 311808 228268
rect 277268 228228 311808 228256
rect 277268 228216 277274 228228
rect 311802 228216 311808 228228
rect 311860 228216 311866 228268
rect 393286 228256 393314 228364
rect 402606 228352 402612 228364
rect 402664 228352 402670 228404
rect 409782 228352 409788 228404
rect 409840 228392 409846 228404
rect 415486 228392 415492 228404
rect 409840 228364 415492 228392
rect 409840 228352 409846 228364
rect 415486 228352 415492 228364
rect 415544 228352 415550 228404
rect 487614 228352 487620 228404
rect 487672 228392 487678 228404
rect 501506 228392 501512 228404
rect 487672 228364 501512 228392
rect 487672 228352 487678 228364
rect 501506 228352 501512 228364
rect 501564 228352 501570 228404
rect 506290 228352 506296 228404
rect 506348 228392 506354 228404
rect 525886 228392 525892 228404
rect 506348 228364 525892 228392
rect 506348 228352 506354 228364
rect 525886 228352 525892 228364
rect 525944 228352 525950 228404
rect 537846 228352 537852 228404
rect 537904 228392 537910 228404
rect 566366 228392 566372 228404
rect 537904 228364 566372 228392
rect 537904 228352 537910 228364
rect 566366 228352 566372 228364
rect 566424 228352 566430 228404
rect 403894 228256 403900 228268
rect 393286 228228 403900 228256
rect 403894 228216 403900 228228
rect 403952 228216 403958 228268
rect 479702 228216 479708 228268
rect 479760 228256 479766 228268
rect 487798 228256 487804 228268
rect 479760 228228 487804 228256
rect 479760 228216 479766 228228
rect 487798 228216 487804 228228
rect 487856 228216 487862 228268
rect 671062 228216 671068 228268
rect 671120 228256 671126 228268
rect 671120 228228 673190 228256
rect 671120 228216 671126 228228
rect 181956 228092 191144 228120
rect 181956 228080 181962 228092
rect 197906 228080 197912 228132
rect 197964 228120 197970 228132
rect 204898 228120 204904 228132
rect 197964 228092 204904 228120
rect 197964 228080 197970 228092
rect 204898 228080 204904 228092
rect 204956 228080 204962 228132
rect 205358 228080 205364 228132
rect 205416 228120 205422 228132
rect 257062 228120 257068 228132
rect 205416 228092 257068 228120
rect 205416 228080 205422 228092
rect 257062 228080 257068 228092
rect 257120 228080 257126 228132
rect 288158 228080 288164 228132
rect 288216 228120 288222 228132
rect 321462 228120 321468 228132
rect 288216 228092 321468 228120
rect 288216 228080 288222 228092
rect 321462 228080 321468 228092
rect 321520 228080 321526 228132
rect 184934 227984 184940 227996
rect 181272 227956 184940 227984
rect 184934 227944 184940 227956
rect 184992 227944 184998 227996
rect 186130 227944 186136 227996
rect 186188 227984 186194 227996
rect 190730 227984 190736 227996
rect 186188 227956 190736 227984
rect 186188 227944 186194 227956
rect 190730 227944 190736 227956
rect 190788 227944 190794 227996
rect 190914 227944 190920 227996
rect 190972 227984 190978 227996
rect 200206 227984 200212 227996
rect 190972 227956 200212 227984
rect 190972 227944 190978 227956
rect 200206 227944 200212 227956
rect 200264 227944 200270 227996
rect 200574 227944 200580 227996
rect 200632 227984 200638 227996
rect 210694 227984 210700 227996
rect 200632 227956 210700 227984
rect 200632 227944 200638 227956
rect 210694 227944 210700 227956
rect 210752 227944 210758 227996
rect 212166 227944 212172 227996
rect 212224 227984 212230 227996
rect 218422 227984 218428 227996
rect 212224 227956 218428 227984
rect 212224 227944 212230 227956
rect 218422 227944 218428 227956
rect 218480 227944 218486 227996
rect 226150 227944 226156 227996
rect 226208 227984 226214 227996
rect 272518 227984 272524 227996
rect 226208 227956 272524 227984
rect 226208 227944 226214 227956
rect 272518 227944 272524 227956
rect 272576 227944 272582 227996
rect 673046 227928 673098 227934
rect 369118 227876 369124 227928
rect 369176 227916 369182 227928
rect 375558 227916 375564 227928
rect 369176 227888 375564 227916
rect 369176 227876 369182 227888
rect 375558 227876 375564 227888
rect 375616 227876 375622 227928
rect 407758 227876 407764 227928
rect 407816 227916 407822 227928
rect 411622 227916 411628 227928
rect 407816 227888 411628 227916
rect 407816 227876 407822 227888
rect 411622 227876 411628 227888
rect 411680 227876 411686 227928
rect 471514 227876 471520 227928
rect 471572 227916 471578 227928
rect 479334 227916 479340 227928
rect 471572 227888 479340 227916
rect 471572 227876 471578 227888
rect 479334 227876 479340 227888
rect 479392 227876 479398 227928
rect 673046 227870 673098 227876
rect 133782 227808 133788 227860
rect 133840 227848 133846 227860
rect 200390 227848 200396 227860
rect 133840 227820 200396 227848
rect 133840 227808 133846 227820
rect 200390 227808 200396 227820
rect 200448 227808 200454 227860
rect 225690 227808 225696 227860
rect 225748 227848 225754 227860
rect 226334 227848 226340 227860
rect 225748 227820 226340 227848
rect 225748 227808 225754 227820
rect 226334 227808 226340 227820
rect 226392 227808 226398 227860
rect 671798 227808 671804 227860
rect 671856 227848 671862 227860
rect 671856 227820 672980 227848
rect 671856 227808 671862 227820
rect 242710 227740 242716 227792
rect 242768 227780 242774 227792
rect 245654 227780 245660 227792
rect 242768 227752 245660 227780
rect 242768 227740 242774 227752
rect 245654 227740 245660 227752
rect 245712 227740 245718 227792
rect 255958 227740 255964 227792
rect 256016 227780 256022 227792
rect 258994 227780 259000 227792
rect 256016 227752 259000 227780
rect 256016 227740 256022 227752
rect 258994 227740 259000 227752
rect 259052 227740 259058 227792
rect 366358 227740 366364 227792
rect 366416 227780 366422 227792
rect 372982 227780 372988 227792
rect 366416 227752 372988 227780
rect 366416 227740 366422 227752
rect 372982 227740 372988 227752
rect 373040 227740 373046 227792
rect 393958 227740 393964 227792
rect 394016 227780 394022 227792
rect 395522 227780 395528 227792
rect 394016 227752 395528 227780
rect 394016 227740 394022 227752
rect 395522 227740 395528 227752
rect 395580 227740 395586 227792
rect 396626 227740 396632 227792
rect 396684 227780 396690 227792
rect 397454 227780 397460 227792
rect 396684 227752 397460 227780
rect 396684 227740 396690 227752
rect 397454 227740 397460 227752
rect 397512 227740 397518 227792
rect 402238 227740 402244 227792
rect 402296 227780 402302 227792
rect 403250 227780 403256 227792
rect 402296 227752 403256 227780
rect 402296 227740 402302 227752
rect 403250 227740 403256 227752
rect 403308 227740 403314 227792
rect 404078 227740 404084 227792
rect 404136 227780 404142 227792
rect 408862 227780 408868 227792
rect 404136 227752 408868 227780
rect 404136 227740 404142 227752
rect 408862 227740 408868 227752
rect 408920 227740 408926 227792
rect 409046 227740 409052 227792
rect 409104 227780 409110 227792
rect 410334 227780 410340 227792
rect 409104 227752 410340 227780
rect 409104 227740 409110 227752
rect 410334 227740 410340 227752
rect 410392 227740 410398 227792
rect 411898 227740 411904 227792
rect 411956 227780 411962 227792
rect 413554 227780 413560 227792
rect 411956 227752 413560 227780
rect 411956 227740 411962 227752
rect 413554 227740 413560 227752
rect 413612 227740 413618 227792
rect 416682 227740 416688 227792
rect 416740 227780 416746 227792
rect 420638 227780 420644 227792
rect 416740 227752 420644 227780
rect 416740 227740 416746 227752
rect 420638 227740 420644 227752
rect 420696 227740 420702 227792
rect 475010 227740 475016 227792
rect 475068 227780 475074 227792
rect 482922 227780 482928 227792
rect 475068 227752 482928 227780
rect 475068 227740 475074 227752
rect 482922 227740 482928 227752
rect 482980 227740 482986 227792
rect 110138 227672 110144 227724
rect 110196 227712 110202 227724
rect 182358 227712 182364 227724
rect 110196 227684 182364 227712
rect 110196 227672 110202 227684
rect 182358 227672 182364 227684
rect 182416 227672 182422 227724
rect 185486 227672 185492 227724
rect 185544 227712 185550 227724
rect 187510 227712 187516 227724
rect 185544 227684 187516 227712
rect 185544 227672 185550 227684
rect 187510 227672 187516 227684
rect 187568 227672 187574 227724
rect 191558 227672 191564 227724
rect 191616 227712 191622 227724
rect 191616 227684 238754 227712
rect 191616 227672 191622 227684
rect 238726 227644 238754 227684
rect 270126 227672 270132 227724
rect 270184 227712 270190 227724
rect 306650 227712 306656 227724
rect 270184 227684 306656 227712
rect 270184 227672 270190 227684
rect 306650 227672 306656 227684
rect 306708 227672 306714 227724
rect 321370 227672 321376 227724
rect 321428 227712 321434 227724
rect 346578 227712 346584 227724
rect 321428 227684 346584 227712
rect 321428 227672 321434 227684
rect 346578 227672 346584 227684
rect 346636 227672 346642 227724
rect 525518 227672 525524 227724
rect 525576 227712 525582 227724
rect 537478 227712 537484 227724
rect 525576 227684 537484 227712
rect 525576 227672 525582 227684
rect 537478 227672 537484 227684
rect 537536 227672 537542 227724
rect 248046 227644 248052 227656
rect 238726 227616 248052 227644
rect 248046 227604 248052 227616
rect 248104 227604 248110 227656
rect 465902 227604 465908 227656
rect 465960 227644 465966 227656
rect 469858 227644 469864 227656
rect 465960 227616 469864 227644
rect 465960 227604 465966 227616
rect 469858 227604 469864 227616
rect 469916 227604 469922 227656
rect 672598 227604 672604 227656
rect 672656 227644 672662 227656
rect 672656 227616 672842 227644
rect 672656 227604 672662 227616
rect 100662 227536 100668 227588
rect 100720 227576 100726 227588
rect 174630 227576 174636 227588
rect 100720 227548 174636 227576
rect 100720 227536 100726 227548
rect 174630 227536 174636 227548
rect 174688 227536 174694 227588
rect 179046 227536 179052 227588
rect 179104 227576 179110 227588
rect 236454 227576 236460 227588
rect 179104 227548 236460 227576
rect 179104 227536 179110 227548
rect 236454 227536 236460 227548
rect 236512 227536 236518 227588
rect 252462 227536 252468 227588
rect 252520 227576 252526 227588
rect 293126 227576 293132 227588
rect 252520 227548 293132 227576
rect 252520 227536 252526 227548
rect 293126 227536 293132 227548
rect 293184 227536 293190 227588
rect 299290 227536 299296 227588
rect 299348 227576 299354 227588
rect 328546 227576 328552 227588
rect 299348 227548 328552 227576
rect 299348 227536 299354 227548
rect 328546 227536 328552 227548
rect 328604 227536 328610 227588
rect 359366 227536 359372 227588
rect 359424 227576 359430 227588
rect 374914 227576 374920 227588
rect 359424 227548 374920 227576
rect 359424 227536 359430 227548
rect 374914 227536 374920 227548
rect 374972 227536 374978 227588
rect 515858 227536 515864 227588
rect 515916 227576 515922 227588
rect 538950 227576 538956 227588
rect 515916 227548 538956 227576
rect 515916 227536 515922 227548
rect 538950 227536 538956 227548
rect 539008 227536 539014 227588
rect 89622 227400 89628 227452
rect 89680 227440 89686 227452
rect 159634 227440 159640 227452
rect 89680 227412 159640 227440
rect 89680 227400 89686 227412
rect 159634 227400 159640 227412
rect 159692 227400 159698 227452
rect 160002 227400 160008 227452
rect 160060 227440 160066 227452
rect 166810 227440 166816 227452
rect 160060 227412 166816 227440
rect 160060 227400 160066 227412
rect 166810 227400 166816 227412
rect 166868 227400 166874 227452
rect 175182 227400 175188 227452
rect 175240 227440 175246 227452
rect 231946 227440 231952 227452
rect 175240 227412 231952 227440
rect 175240 227400 175246 227412
rect 231946 227400 231952 227412
rect 232004 227400 232010 227452
rect 248230 227400 248236 227452
rect 248288 227440 248294 227452
rect 291838 227440 291844 227452
rect 248288 227412 291844 227440
rect 248288 227400 248294 227412
rect 291838 227400 291844 227412
rect 291896 227400 291902 227452
rect 293770 227400 293776 227452
rect 293828 227440 293834 227452
rect 325326 227440 325332 227452
rect 293828 227412 325332 227440
rect 293828 227400 293834 227412
rect 325326 227400 325332 227412
rect 325384 227400 325390 227452
rect 340598 227400 340604 227452
rect 340656 227440 340662 227452
rect 361390 227440 361396 227452
rect 340656 227412 361396 227440
rect 340656 227400 340662 227412
rect 361390 227400 361396 227412
rect 361448 227400 361454 227452
rect 369762 227400 369768 227452
rect 369820 227440 369826 227452
rect 385862 227440 385868 227452
rect 369820 227412 385868 227440
rect 369820 227400 369826 227412
rect 385862 227400 385868 227412
rect 385920 227400 385926 227452
rect 524322 227400 524328 227452
rect 524380 227440 524386 227452
rect 547874 227440 547880 227452
rect 524380 227412 547880 227440
rect 524380 227400 524386 227412
rect 547874 227400 547880 227412
rect 547932 227400 547938 227452
rect 672442 227400 672448 227452
rect 672500 227440 672506 227452
rect 672500 227412 672750 227440
rect 672500 227400 672506 227412
rect 676398 227332 676404 227384
rect 676456 227372 676462 227384
rect 677042 227372 677048 227384
rect 676456 227344 677048 227372
rect 676456 227332 676462 227344
rect 677042 227332 677048 227344
rect 677100 227332 677106 227384
rect 86862 227264 86868 227316
rect 86920 227304 86926 227316
rect 151906 227304 151912 227316
rect 86920 227276 151912 227304
rect 86920 227264 86926 227276
rect 151906 227264 151912 227276
rect 151964 227264 151970 227316
rect 152918 227264 152924 227316
rect 152976 227304 152982 227316
rect 164326 227304 164332 227316
rect 152976 227276 164332 227304
rect 152976 227264 152982 227276
rect 164326 227264 164332 227276
rect 164384 227264 164390 227316
rect 165430 227264 165436 227316
rect 165488 227304 165494 227316
rect 227438 227304 227444 227316
rect 165488 227276 227444 227304
rect 165488 227264 165494 227276
rect 227438 227264 227444 227276
rect 227496 227264 227502 227316
rect 233234 227304 233240 227316
rect 228928 227276 233240 227304
rect 75822 227128 75828 227180
rect 75880 227168 75886 227180
rect 150158 227168 150164 227180
rect 75880 227140 150164 227168
rect 75880 227128 75886 227140
rect 150158 227128 150164 227140
rect 150216 227128 150222 227180
rect 150342 227128 150348 227180
rect 150400 227168 150406 227180
rect 150400 227140 152136 227168
rect 150400 227128 150406 227140
rect 57882 226992 57888 227044
rect 57940 227032 57946 227044
rect 134978 227032 134984 227044
rect 57940 227004 134984 227032
rect 57940 226992 57946 227004
rect 134978 226992 134984 227004
rect 135036 226992 135042 227044
rect 135438 226992 135444 227044
rect 135496 227032 135502 227044
rect 151906 227032 151912 227044
rect 135496 227004 151912 227032
rect 135496 226992 135502 227004
rect 151906 226992 151912 227004
rect 151964 226992 151970 227044
rect 152108 227032 152136 227140
rect 152274 227128 152280 227180
rect 152332 227168 152338 227180
rect 168834 227168 168840 227180
rect 152332 227140 168840 227168
rect 152332 227128 152338 227140
rect 168834 227128 168840 227140
rect 168892 227128 168898 227180
rect 169570 227128 169576 227180
rect 169628 227168 169634 227180
rect 228726 227168 228732 227180
rect 169628 227140 228732 227168
rect 169628 227128 169634 227140
rect 228726 227128 228732 227140
rect 228784 227128 228790 227180
rect 213270 227032 213276 227044
rect 152108 227004 213276 227032
rect 213270 226992 213276 227004
rect 213328 226992 213334 227044
rect 226886 226992 226892 227044
rect 226944 227032 226950 227044
rect 228928 227032 228956 227276
rect 233234 227264 233240 227276
rect 233292 227264 233298 227316
rect 234522 227264 234528 227316
rect 234580 227304 234586 227316
rect 278314 227304 278320 227316
rect 234580 227276 278320 227304
rect 234580 227264 234586 227276
rect 278314 227264 278320 227276
rect 278372 227264 278378 227316
rect 280706 227264 280712 227316
rect 280764 227304 280770 227316
rect 312078 227304 312084 227316
rect 280764 227276 312084 227304
rect 280764 227264 280770 227276
rect 312078 227264 312084 227276
rect 312136 227264 312142 227316
rect 326338 227264 326344 227316
rect 326396 227304 326402 227316
rect 352374 227304 352380 227316
rect 326396 227276 352380 227304
rect 326396 227264 326402 227276
rect 352374 227264 352380 227276
rect 352432 227264 352438 227316
rect 355502 227264 355508 227316
rect 355560 227304 355566 227316
rect 372338 227304 372344 227316
rect 355560 227276 372344 227304
rect 355560 227264 355566 227276
rect 372338 227264 372344 227276
rect 372396 227264 372402 227316
rect 373626 227304 373632 227316
rect 372540 227276 373632 227304
rect 235902 227128 235908 227180
rect 235960 227168 235966 227180
rect 280246 227168 280252 227180
rect 235960 227140 280252 227168
rect 235960 227128 235966 227140
rect 280246 227128 280252 227140
rect 280304 227128 280310 227180
rect 296438 227128 296444 227180
rect 296496 227168 296502 227180
rect 329190 227168 329196 227180
rect 296496 227140 329196 227168
rect 296496 227128 296502 227140
rect 329190 227128 329196 227140
rect 329248 227128 329254 227180
rect 329742 227128 329748 227180
rect 329800 227168 329806 227180
rect 353662 227168 353668 227180
rect 329800 227140 353668 227168
rect 329800 227128 329806 227140
rect 353662 227128 353668 227140
rect 353720 227128 353726 227180
rect 354582 227128 354588 227180
rect 354640 227168 354646 227180
rect 372540 227168 372568 227276
rect 373626 227264 373632 227276
rect 373684 227264 373690 227316
rect 382918 227264 382924 227316
rect 382976 227304 382982 227316
rect 391658 227304 391664 227316
rect 382976 227276 391664 227304
rect 382976 227264 382982 227276
rect 391658 227264 391664 227276
rect 391716 227264 391722 227316
rect 395982 227264 395988 227316
rect 396040 227304 396046 227316
rect 406470 227304 406476 227316
rect 396040 227276 406476 227304
rect 396040 227264 396046 227276
rect 406470 227264 406476 227276
rect 406528 227264 406534 227316
rect 485038 227264 485044 227316
rect 485096 227304 485102 227316
rect 498746 227304 498752 227316
rect 485096 227276 498752 227304
rect 485096 227264 485102 227276
rect 498746 227264 498752 227276
rect 498804 227264 498810 227316
rect 501138 227264 501144 227316
rect 501196 227304 501202 227316
rect 517790 227304 517796 227316
rect 501196 227276 517796 227304
rect 501196 227264 501202 227276
rect 517790 227264 517796 227276
rect 517848 227264 517854 227316
rect 521746 227264 521752 227316
rect 521804 227304 521810 227316
rect 545114 227304 545120 227316
rect 521804 227276 545120 227304
rect 521804 227264 521810 227276
rect 545114 227264 545120 227276
rect 545172 227264 545178 227316
rect 354640 227140 372568 227168
rect 354640 227128 354646 227140
rect 373258 227128 373264 227180
rect 373316 227168 373322 227180
rect 383286 227168 383292 227180
rect 373316 227140 383292 227168
rect 373316 227128 373322 227140
rect 383286 227128 383292 227140
rect 383344 227128 383350 227180
rect 386322 227128 386328 227180
rect 386380 227168 386386 227180
rect 398742 227168 398748 227180
rect 386380 227140 398748 227168
rect 386380 227128 386386 227140
rect 398742 227128 398748 227140
rect 398800 227128 398806 227180
rect 481174 227128 481180 227180
rect 481232 227168 481238 227180
rect 492950 227168 492956 227180
rect 481232 227140 492956 227168
rect 481232 227128 481238 227140
rect 492950 227128 492956 227140
rect 493008 227128 493014 227180
rect 498562 227128 498568 227180
rect 498620 227168 498626 227180
rect 515858 227168 515864 227180
rect 498620 227140 515864 227168
rect 498620 227128 498626 227140
rect 515858 227128 515864 227140
rect 515916 227128 515922 227180
rect 516042 227128 516048 227180
rect 516100 227168 516106 227180
rect 525058 227168 525064 227180
rect 516100 227140 525064 227168
rect 516100 227128 516106 227140
rect 525058 227128 525064 227140
rect 525116 227128 525122 227180
rect 535914 227128 535920 227180
rect 535972 227168 535978 227180
rect 563882 227168 563888 227180
rect 535972 227140 563888 227168
rect 535972 227128 535978 227140
rect 563882 227128 563888 227140
rect 563940 227128 563946 227180
rect 672604 227112 672656 227118
rect 672604 227054 672656 227060
rect 226944 227004 228956 227032
rect 226944 226992 226950 227004
rect 229048 226992 229054 227044
rect 229106 227032 229112 227044
rect 271230 227032 271236 227044
rect 229106 227004 271236 227032
rect 229106 226992 229112 227004
rect 271230 226992 271236 227004
rect 271288 226992 271294 227044
rect 271782 226992 271788 227044
rect 271840 227032 271846 227044
rect 308582 227032 308588 227044
rect 271840 227004 308588 227032
rect 271840 226992 271846 227004
rect 308582 226992 308588 227004
rect 308640 226992 308646 227044
rect 308766 226992 308772 227044
rect 308824 227032 308830 227044
rect 336274 227032 336280 227044
rect 308824 227004 336280 227032
rect 308824 226992 308830 227004
rect 336274 226992 336280 227004
rect 336332 226992 336338 227044
rect 336458 226992 336464 227044
rect 336516 227032 336522 227044
rect 360102 227032 360108 227044
rect 336516 227004 360108 227032
rect 336516 226992 336522 227004
rect 360102 226992 360108 227004
rect 360160 226992 360166 227044
rect 361206 226992 361212 227044
rect 361264 227032 361270 227044
rect 377214 227032 377220 227044
rect 361264 227004 377220 227032
rect 361264 226992 361270 227004
rect 377214 226992 377220 227004
rect 377272 226992 377278 227044
rect 381906 226992 381912 227044
rect 381964 227032 381970 227044
rect 396166 227032 396172 227044
rect 381964 227004 396172 227032
rect 381964 226992 381970 227004
rect 396166 226992 396172 227004
rect 396224 226992 396230 227044
rect 398466 226992 398472 227044
rect 398524 227032 398530 227044
rect 408678 227032 408684 227044
rect 398524 227004 408684 227032
rect 398524 226992 398530 227004
rect 408678 226992 408684 227004
rect 408736 226992 408742 227044
rect 472158 226992 472164 227044
rect 472216 227032 472222 227044
rect 481174 227032 481180 227044
rect 472216 227004 481180 227032
rect 472216 226992 472222 227004
rect 481174 226992 481180 227004
rect 481232 226992 481238 227044
rect 497274 226992 497280 227044
rect 497332 227032 497338 227044
rect 497332 227004 509234 227032
rect 497332 226992 497338 227004
rect 106918 226856 106924 226908
rect 106976 226896 106982 226908
rect 125778 226896 125784 226908
rect 106976 226868 125784 226896
rect 106976 226856 106982 226868
rect 125778 226856 125784 226868
rect 125836 226856 125842 226908
rect 191098 226896 191104 226908
rect 125980 226868 191104 226896
rect 121086 226720 121092 226772
rect 121144 226760 121150 226772
rect 125980 226760 126008 226868
rect 191098 226856 191104 226868
rect 191156 226856 191162 226908
rect 200022 226856 200028 226908
rect 200080 226896 200086 226908
rect 251910 226896 251916 226908
rect 200080 226868 251916 226896
rect 200080 226856 200086 226868
rect 251910 226856 251916 226868
rect 251968 226856 251974 226908
rect 272426 226856 272432 226908
rect 272484 226896 272490 226908
rect 284754 226896 284760 226908
rect 272484 226868 284760 226896
rect 272484 226856 272490 226868
rect 284754 226856 284760 226868
rect 284812 226856 284818 226908
rect 509206 226896 509234 227004
rect 514018 226992 514024 227044
rect 514076 227032 514082 227044
rect 535638 227032 535644 227044
rect 514076 227004 535644 227032
rect 514076 226992 514082 227004
rect 535638 226992 535644 227004
rect 535696 226992 535702 227044
rect 537202 226992 537208 227044
rect 537260 227032 537266 227044
rect 565630 227032 565636 227044
rect 537260 227004 565636 227032
rect 537260 226992 537266 227004
rect 565630 226992 565636 227004
rect 565688 226992 565694 227044
rect 672494 226908 672546 226914
rect 514294 226896 514300 226908
rect 509206 226868 514300 226896
rect 514294 226856 514300 226868
rect 514352 226856 514358 226908
rect 672494 226850 672546 226856
rect 672380 226772 672432 226778
rect 190086 226760 190092 226772
rect 121144 226732 126008 226760
rect 126072 226732 190092 226760
rect 121144 226720 121150 226732
rect 119982 226584 119988 226636
rect 120040 226624 120046 226636
rect 126072 226624 126100 226732
rect 190086 226720 190092 226732
rect 190144 226720 190150 226772
rect 195790 226720 195796 226772
rect 195848 226760 195854 226772
rect 199470 226760 199476 226772
rect 195848 226732 199476 226760
rect 195848 226720 195854 226732
rect 199470 226720 199476 226732
rect 199528 226720 199534 226772
rect 212166 226720 212172 226772
rect 212224 226760 212230 226772
rect 262214 226760 262220 226772
rect 212224 226732 262220 226760
rect 212224 226720 212230 226732
rect 262214 226720 262220 226732
rect 262272 226720 262278 226772
rect 672380 226714 672432 226720
rect 135438 226624 135444 226636
rect 120040 226596 126100 226624
rect 126164 226596 135444 226624
rect 120040 226584 120046 226596
rect 125778 226448 125784 226500
rect 125836 226488 125842 226500
rect 126164 226488 126192 226596
rect 135438 226584 135444 226596
rect 135496 226584 135502 226636
rect 135622 226584 135628 226636
rect 135680 226624 135686 226636
rect 135680 226596 137416 226624
rect 135680 226584 135686 226596
rect 125836 226460 126192 226488
rect 125836 226448 125842 226460
rect 129366 226448 129372 226500
rect 129424 226488 129430 226500
rect 137186 226488 137192 226500
rect 129424 226460 137192 226488
rect 129424 226448 129430 226460
rect 137186 226448 137192 226460
rect 137244 226448 137250 226500
rect 137388 226488 137416 226596
rect 137554 226584 137560 226636
rect 137612 226624 137618 226636
rect 197446 226624 197452 226636
rect 137612 226596 197452 226624
rect 137612 226584 137618 226596
rect 197446 226584 197452 226596
rect 197504 226584 197510 226636
rect 222010 226584 222016 226636
rect 222068 226624 222074 226636
rect 269942 226624 269948 226636
rect 222068 226596 269948 226624
rect 222068 226584 222074 226596
rect 269942 226584 269948 226596
rect 270000 226584 270006 226636
rect 668302 226584 668308 226636
rect 668360 226624 668366 226636
rect 668360 226596 672290 226624
rect 668360 226584 668366 226596
rect 142108 226488 142114 226500
rect 137388 226460 142114 226488
rect 142108 226448 142114 226460
rect 142166 226448 142172 226500
rect 142246 226448 142252 226500
rect 142304 226488 142310 226500
rect 205542 226488 205548 226500
rect 142304 226460 205548 226488
rect 142304 226448 142310 226460
rect 205542 226448 205548 226460
rect 205600 226448 205606 226500
rect 213178 226448 213184 226500
rect 213236 226488 213242 226500
rect 217778 226488 217784 226500
rect 213236 226460 217784 226488
rect 213236 226448 213242 226460
rect 217778 226448 217784 226460
rect 217836 226448 217842 226500
rect 221826 226448 221832 226500
rect 221884 226488 221890 226500
rect 229002 226488 229008 226500
rect 221884 226460 229008 226488
rect 221884 226448 221890 226460
rect 229002 226448 229008 226460
rect 229060 226448 229066 226500
rect 232498 226448 232504 226500
rect 232556 226488 232562 226500
rect 266722 226488 266728 226500
rect 232556 226460 266728 226488
rect 232556 226448 232562 226460
rect 266722 226448 266728 226460
rect 266780 226448 266786 226500
rect 666646 226448 666652 226500
rect 666704 226488 666710 226500
rect 666704 226460 672182 226488
rect 666704 226448 666710 226460
rect 291838 226380 291844 226432
rect 291896 226420 291902 226432
rect 295058 226420 295064 226432
rect 291896 226392 295064 226420
rect 291896 226380 291902 226392
rect 295058 226380 295064 226392
rect 295116 226380 295122 226432
rect 152200 226324 152688 226352
rect 83458 226244 83464 226296
rect 83516 226284 83522 226296
rect 152200 226284 152228 226324
rect 83516 226256 152228 226284
rect 83516 226244 83522 226256
rect 69566 226108 69572 226160
rect 69624 226148 69630 226160
rect 137462 226148 137468 226160
rect 69624 226120 137468 226148
rect 69624 226108 69630 226120
rect 137462 226108 137468 226120
rect 137520 226108 137526 226160
rect 137646 226108 137652 226160
rect 137704 226148 137710 226160
rect 141510 226148 141516 226160
rect 137704 226120 141516 226148
rect 137704 226108 137710 226120
rect 141510 226108 141516 226120
rect 141568 226108 141574 226160
rect 141694 226108 141700 226160
rect 141752 226148 141758 226160
rect 146754 226148 146760 226160
rect 141752 226120 146760 226148
rect 141752 226108 141758 226120
rect 146754 226108 146760 226120
rect 146812 226108 146818 226160
rect 152660 226148 152688 226324
rect 166810 226312 166816 226364
rect 166868 226352 166874 226364
rect 220998 226352 221004 226364
rect 166868 226324 221004 226352
rect 166868 226312 166874 226324
rect 220998 226312 221004 226324
rect 221056 226312 221062 226364
rect 672034 226296 672086 226302
rect 152826 226244 152832 226296
rect 152884 226284 152890 226296
rect 161934 226284 161940 226296
rect 152884 226256 161940 226284
rect 152884 226244 152890 226256
rect 161934 226244 161940 226256
rect 161992 226244 161998 226296
rect 162302 226244 162308 226296
rect 162360 226284 162366 226296
rect 166626 226284 166632 226296
rect 162360 226256 166632 226284
rect 162360 226244 162366 226256
rect 166626 226244 166632 226256
rect 166684 226244 166690 226296
rect 222470 226244 222476 226296
rect 222528 226284 222534 226296
rect 225506 226284 225512 226296
rect 222528 226256 225512 226284
rect 222528 226244 222534 226256
rect 225506 226244 225512 226256
rect 225564 226244 225570 226296
rect 228726 226244 228732 226296
rect 228784 226284 228790 226296
rect 275094 226284 275100 226296
rect 228784 226256 275100 226284
rect 228784 226244 228790 226256
rect 275094 226244 275100 226256
rect 275152 226244 275158 226296
rect 278498 226244 278504 226296
rect 278556 226284 278562 226296
rect 315022 226284 315028 226296
rect 278556 226256 315028 226284
rect 278556 226244 278562 226256
rect 315022 226244 315028 226256
rect 315080 226244 315086 226296
rect 317322 226244 317328 226296
rect 317380 226284 317386 226296
rect 334250 226284 334256 226296
rect 317380 226256 334256 226284
rect 317380 226244 317386 226256
rect 334250 226244 334256 226256
rect 334308 226244 334314 226296
rect 503254 226244 503260 226296
rect 503312 226284 503318 226296
rect 510154 226284 510160 226296
rect 503312 226256 510160 226284
rect 503312 226244 503318 226256
rect 510154 226244 510160 226256
rect 510212 226244 510218 226296
rect 529934 226244 529940 226296
rect 529992 226284 529998 226296
rect 544930 226284 544936 226296
rect 529992 226256 544936 226284
rect 529992 226244 529998 226256
rect 544930 226244 544936 226256
rect 544988 226244 544994 226296
rect 562318 226244 562324 226296
rect 562376 226284 562382 226296
rect 567562 226284 567568 226296
rect 562376 226256 567568 226284
rect 562376 226244 562382 226256
rect 567562 226244 567568 226256
rect 567620 226244 567626 226296
rect 672034 226238 672086 226244
rect 157426 226148 157432 226160
rect 152660 226120 157432 226148
rect 157426 226108 157432 226120
rect 157484 226108 157490 226160
rect 157610 226108 157616 226160
rect 157668 226148 157674 226160
rect 215846 226148 215852 226160
rect 157668 226120 215852 226148
rect 157668 226108 157674 226120
rect 215846 226108 215852 226120
rect 215904 226108 215910 226160
rect 216490 226108 216496 226160
rect 216548 226148 216554 226160
rect 264790 226148 264796 226160
rect 216548 226120 264796 226148
rect 216548 226108 216554 226120
rect 264790 226108 264796 226120
rect 264848 226108 264854 226160
rect 266262 226108 266268 226160
rect 266320 226148 266326 226160
rect 303430 226148 303436 226160
rect 266320 226120 303436 226148
rect 266320 226108 266326 226120
rect 303430 226108 303436 226120
rect 303488 226108 303494 226160
rect 325418 226108 325424 226160
rect 325476 226148 325482 226160
rect 349154 226148 349160 226160
rect 325476 226120 349160 226148
rect 325476 226108 325482 226120
rect 349154 226108 349160 226120
rect 349212 226108 349218 226160
rect 510798 226108 510804 226160
rect 510856 226148 510862 226160
rect 531682 226148 531688 226160
rect 510856 226120 531688 226148
rect 510856 226108 510862 226120
rect 531682 226108 531688 226120
rect 531740 226108 531746 226160
rect 666002 226040 666008 226092
rect 666060 226080 666066 226092
rect 666060 226052 671968 226080
rect 666060 226040 666066 226052
rect 93762 225972 93768 226024
rect 93820 226012 93826 226024
rect 166810 226012 166816 226024
rect 93820 225984 166816 226012
rect 93820 225972 93826 225984
rect 166810 225972 166816 225984
rect 166868 225972 166874 226024
rect 166948 225972 166954 226024
rect 167006 226012 167012 226024
rect 176470 226012 176476 226024
rect 167006 225984 176476 226012
rect 167006 225972 167012 225984
rect 176470 225972 176476 225984
rect 176528 225972 176534 226024
rect 178678 225972 178684 226024
rect 178736 226012 178742 226024
rect 187142 226012 187148 226024
rect 178736 225984 187148 226012
rect 178736 225972 178742 225984
rect 187142 225972 187148 225984
rect 187200 225972 187206 226024
rect 187326 225972 187332 226024
rect 187384 226012 187390 226024
rect 224218 226012 224224 226024
rect 187384 225984 224224 226012
rect 187384 225972 187390 225984
rect 224218 225972 224224 225984
rect 224276 225972 224282 226024
rect 233878 226012 233884 226024
rect 229066 225984 233884 226012
rect 95142 225836 95148 225888
rect 95200 225876 95206 225888
rect 161198 225876 161204 225888
rect 95200 225848 161204 225876
rect 95200 225836 95206 225848
rect 161198 225836 161204 225848
rect 161256 225836 161262 225888
rect 161934 225836 161940 225888
rect 161992 225876 161998 225888
rect 176102 225876 176108 225888
rect 161992 225848 176108 225876
rect 161992 225836 161998 225848
rect 176102 225836 176108 225848
rect 176160 225836 176166 225888
rect 177206 225836 177212 225888
rect 177264 225876 177270 225888
rect 229066 225876 229094 225984
rect 233878 225972 233884 225984
rect 233936 225972 233942 226024
rect 243446 225972 243452 226024
rect 243504 226012 243510 226024
rect 248690 226012 248696 226024
rect 243504 225984 248696 226012
rect 243504 225972 243510 225984
rect 248690 225972 248696 225984
rect 248748 225972 248754 226024
rect 267688 225972 267694 226024
rect 267746 226012 267752 226024
rect 304074 226012 304080 226024
rect 267746 225984 304080 226012
rect 267746 225972 267752 225984
rect 304074 225972 304080 225984
rect 304132 225972 304138 226024
rect 313090 225972 313096 226024
rect 313148 226012 313154 226024
rect 340782 226012 340788 226024
rect 313148 225984 340788 226012
rect 313148 225972 313154 225984
rect 340782 225972 340788 225984
rect 340840 225972 340846 226024
rect 347866 226012 347872 226024
rect 344986 225984 347872 226012
rect 239030 225876 239036 225888
rect 177264 225848 229094 225876
rect 232700 225848 239036 225876
rect 177264 225836 177270 225848
rect 64782 225700 64788 225752
rect 64840 225740 64846 225752
rect 92474 225740 92480 225752
rect 64840 225712 92480 225740
rect 64840 225700 64846 225712
rect 92474 225700 92480 225712
rect 92532 225700 92538 225752
rect 108298 225700 108304 225752
rect 108356 225740 108362 225752
rect 176470 225740 176476 225752
rect 108356 225712 176476 225740
rect 108356 225700 108362 225712
rect 176470 225700 176476 225712
rect 176528 225700 176534 225752
rect 176654 225700 176660 225752
rect 176712 225740 176718 225752
rect 185670 225740 185676 225752
rect 176712 225712 185676 225740
rect 176712 225700 176718 225712
rect 185670 225700 185676 225712
rect 185728 225700 185734 225752
rect 187510 225700 187516 225752
rect 187568 225740 187574 225752
rect 232700 225740 232728 225848
rect 239030 225836 239036 225848
rect 239088 225836 239094 225888
rect 249702 225836 249708 225888
rect 249760 225876 249766 225888
rect 290550 225876 290556 225888
rect 249760 225848 290556 225876
rect 249760 225836 249766 225848
rect 290550 225836 290556 225848
rect 290608 225836 290614 225888
rect 294966 225836 294972 225888
rect 295024 225876 295030 225888
rect 325970 225876 325976 225888
rect 295024 225848 325976 225876
rect 295024 225836 295030 225848
rect 325970 225836 325976 225848
rect 326028 225836 326034 225888
rect 340138 225836 340144 225888
rect 340196 225876 340202 225888
rect 344986 225876 345014 225984
rect 347866 225972 347872 225984
rect 347924 225972 347930 226024
rect 349062 225972 349068 226024
rect 349120 226012 349126 226024
rect 367186 226012 367192 226024
rect 349120 225984 367192 226012
rect 349120 225972 349126 225984
rect 367186 225972 367192 225984
rect 367244 225972 367250 226024
rect 518526 225972 518532 226024
rect 518584 226012 518590 226024
rect 541434 226012 541440 226024
rect 518584 225984 541440 226012
rect 518584 225972 518590 225984
rect 541434 225972 541440 225984
rect 541492 225972 541498 226024
rect 544194 225972 544200 226024
rect 544252 226012 544258 226024
rect 562686 226012 562692 226024
rect 544252 225984 562692 226012
rect 544252 225972 544258 225984
rect 562686 225972 562692 225984
rect 562744 225972 562750 226024
rect 340196 225848 345014 225876
rect 340196 225836 340202 225848
rect 347038 225836 347044 225888
rect 347096 225876 347102 225888
rect 365898 225876 365904 225888
rect 347096 225848 365904 225876
rect 347096 225836 347102 225848
rect 365898 225836 365904 225848
rect 365956 225836 365962 225888
rect 367646 225836 367652 225888
rect 367704 225876 367710 225888
rect 380066 225876 380072 225888
rect 367704 225848 380072 225876
rect 367704 225836 367710 225848
rect 380066 225836 380072 225848
rect 380124 225836 380130 225888
rect 488902 225836 488908 225888
rect 488960 225876 488966 225888
rect 502978 225876 502984 225888
rect 488960 225848 502984 225876
rect 488960 225836 488966 225848
rect 502978 225836 502984 225848
rect 503036 225836 503042 225888
rect 528186 225836 528192 225888
rect 528244 225876 528250 225888
rect 554038 225876 554044 225888
rect 528244 225848 554044 225876
rect 528244 225836 528250 225848
rect 554038 225836 554044 225848
rect 554096 225836 554102 225888
rect 458634 225768 458640 225820
rect 458692 225808 458698 225820
rect 462958 225808 462964 225820
rect 458692 225780 462964 225808
rect 458692 225768 458698 225780
rect 462958 225768 462964 225780
rect 463016 225768 463022 225820
rect 671820 225752 671872 225758
rect 242894 225740 242900 225752
rect 187568 225712 232728 225740
rect 232792 225712 242900 225740
rect 187568 225700 187574 225712
rect 186608 225644 186820 225672
rect 61286 225564 61292 225616
rect 61344 225604 61350 225616
rect 136818 225604 136824 225616
rect 61344 225576 136824 225604
rect 61344 225564 61350 225576
rect 136818 225564 136824 225576
rect 136876 225564 136882 225616
rect 137002 225564 137008 225616
rect 137060 225604 137066 225616
rect 146938 225604 146944 225616
rect 137060 225576 146944 225604
rect 137060 225564 137066 225576
rect 146938 225564 146944 225576
rect 146996 225564 147002 225616
rect 147122 225564 147128 225616
rect 147180 225604 147186 225616
rect 186608 225604 186636 225644
rect 147180 225576 186636 225604
rect 186792 225604 186820 225644
rect 186792 225576 200804 225604
rect 147180 225564 147186 225576
rect 200776 225536 200804 225576
rect 201034 225564 201040 225616
rect 201092 225604 201098 225616
rect 222470 225604 222476 225616
rect 201092 225576 222476 225604
rect 201092 225564 201098 225576
rect 222470 225564 222476 225576
rect 222528 225564 222534 225616
rect 224218 225564 224224 225616
rect 224276 225604 224282 225616
rect 232792 225604 232820 225712
rect 242894 225700 242900 225712
rect 242952 225700 242958 225752
rect 257706 225700 257712 225752
rect 257764 225740 257770 225752
rect 299566 225740 299572 225752
rect 257764 225712 299572 225740
rect 257764 225700 257770 225712
rect 299566 225700 299572 225712
rect 299624 225700 299630 225752
rect 304902 225700 304908 225752
rect 304960 225740 304966 225752
rect 333698 225740 333704 225752
rect 304960 225712 333704 225740
rect 304960 225700 304966 225712
rect 333698 225700 333704 225712
rect 333756 225700 333762 225752
rect 335262 225700 335268 225752
rect 335320 225740 335326 225752
rect 356882 225740 356888 225752
rect 335320 225712 356888 225740
rect 335320 225700 335326 225712
rect 356882 225700 356888 225712
rect 356940 225700 356946 225752
rect 379330 225700 379336 225752
rect 379388 225740 379394 225752
rect 393590 225740 393596 225752
rect 379388 225712 393596 225740
rect 379388 225700 379394 225712
rect 393590 225700 393596 225712
rect 393648 225700 393654 225752
rect 394602 225700 394608 225752
rect 394660 225740 394666 225752
rect 404538 225740 404544 225752
rect 394660 225712 404544 225740
rect 394660 225700 394666 225712
rect 404538 225700 404544 225712
rect 404596 225700 404602 225752
rect 491478 225700 491484 225752
rect 491536 225740 491542 225752
rect 506842 225740 506848 225752
rect 491536 225712 506848 225740
rect 491536 225700 491542 225712
rect 506842 225700 506848 225712
rect 506900 225700 506906 225752
rect 507302 225700 507308 225752
rect 507360 225740 507366 225752
rect 526714 225740 526720 225752
rect 507360 225712 526720 225740
rect 507360 225700 507366 225712
rect 526714 225700 526720 225712
rect 526772 225700 526778 225752
rect 527542 225700 527548 225752
rect 527600 225740 527606 225752
rect 553210 225740 553216 225752
rect 527600 225712 553216 225740
rect 527600 225700 527606 225712
rect 553210 225700 553216 225712
rect 553268 225700 553274 225752
rect 671820 225694 671872 225700
rect 224276 225576 232820 225604
rect 224276 225564 224282 225576
rect 234338 225564 234344 225616
rect 234396 225604 234402 225616
rect 281534 225604 281540 225616
rect 234396 225576 281540 225604
rect 234396 225564 234402 225576
rect 281534 225564 281540 225576
rect 281592 225564 281598 225616
rect 285490 225564 285496 225616
rect 285548 225604 285554 225616
rect 318886 225604 318892 225616
rect 285548 225576 318892 225604
rect 285548 225564 285554 225576
rect 318886 225564 318892 225576
rect 318944 225564 318950 225616
rect 322842 225564 322848 225616
rect 322900 225604 322906 225616
rect 349798 225604 349804 225616
rect 322900 225576 349804 225604
rect 322900 225564 322906 225576
rect 349798 225564 349804 225576
rect 349856 225564 349862 225616
rect 351178 225564 351184 225616
rect 351236 225604 351242 225616
rect 370406 225604 370412 225616
rect 351236 225576 370412 225604
rect 351236 225564 351242 225576
rect 370406 225564 370412 225576
rect 370464 225564 370470 225616
rect 372522 225564 372528 225616
rect 372580 225604 372586 225616
rect 388070 225604 388076 225616
rect 372580 225576 388076 225604
rect 372580 225564 372586 225576
rect 388070 225564 388076 225576
rect 388128 225564 388134 225616
rect 388438 225564 388444 225616
rect 388496 225604 388502 225616
rect 399386 225604 399392 225616
rect 388496 225576 399392 225604
rect 388496 225564 388502 225576
rect 399386 225564 399392 225576
rect 399444 225564 399450 225616
rect 467650 225564 467656 225616
rect 467708 225604 467714 225616
rect 476574 225604 476580 225616
rect 467708 225576 476580 225604
rect 467708 225564 467714 225576
rect 476574 225564 476580 225576
rect 476632 225564 476638 225616
rect 477310 225564 477316 225616
rect 477368 225604 477374 225616
rect 489178 225604 489184 225616
rect 477368 225576 489184 225604
rect 477368 225564 477374 225576
rect 489178 225564 489184 225576
rect 489236 225564 489242 225616
rect 495158 225564 495164 225616
rect 495216 225604 495222 225616
rect 509694 225604 509700 225616
rect 495216 225576 509700 225604
rect 495216 225564 495222 225576
rect 509694 225564 509700 225576
rect 509752 225564 509758 225616
rect 510338 225564 510344 225616
rect 510396 225604 510402 225616
rect 530486 225604 530492 225616
rect 510396 225576 530492 225604
rect 510396 225564 510402 225576
rect 530486 225564 530492 225576
rect 530544 225564 530550 225616
rect 532050 225564 532056 225616
rect 532108 225604 532114 225616
rect 559006 225604 559012 225616
rect 532108 225576 559012 225604
rect 532108 225564 532114 225576
rect 559006 225564 559012 225576
rect 559064 225564 559070 225616
rect 671712 225548 671764 225554
rect 200776 225508 200896 225536
rect 103422 225428 103428 225480
rect 103480 225468 103486 225480
rect 108298 225468 108304 225480
rect 103480 225440 108304 225468
rect 103480 225428 103486 225440
rect 108298 225428 108304 225440
rect 108356 225428 108362 225480
rect 127434 225468 127440 225480
rect 113146 225440 127440 225468
rect 105998 225292 106004 225344
rect 106056 225332 106062 225344
rect 113146 225332 113174 225440
rect 127434 225428 127440 225440
rect 127492 225428 127498 225480
rect 185486 225468 185492 225480
rect 127636 225440 185492 225468
rect 106056 225304 113174 225332
rect 106056 225292 106062 225304
rect 117222 225292 117228 225344
rect 117280 225332 117286 225344
rect 127636 225332 127664 225440
rect 185486 225428 185492 225440
rect 185544 225428 185550 225480
rect 187326 225428 187332 225480
rect 187384 225468 187390 225480
rect 195790 225468 195796 225480
rect 187384 225440 195796 225468
rect 187384 225428 187390 225440
rect 195790 225428 195796 225440
rect 195848 225428 195854 225480
rect 199378 225428 199384 225480
rect 199436 225468 199442 225480
rect 200482 225468 200488 225480
rect 199436 225440 200488 225468
rect 199436 225428 199442 225440
rect 200482 225428 200488 225440
rect 200540 225428 200546 225480
rect 137002 225332 137008 225344
rect 117280 225304 127664 225332
rect 127728 225304 137008 225332
rect 117280 225292 117286 225304
rect 127434 225156 127440 225208
rect 127492 225196 127498 225208
rect 127728 225196 127756 225304
rect 137002 225292 137008 225304
rect 137060 225292 137066 225344
rect 146938 225332 146944 225344
rect 137204 225304 146944 225332
rect 127492 225168 127756 225196
rect 127492 225156 127498 225168
rect 128262 225156 128268 225208
rect 128320 225196 128326 225208
rect 137204 225196 137232 225304
rect 146938 225292 146944 225304
rect 146996 225292 147002 225344
rect 147122 225292 147128 225344
rect 147180 225332 147186 225344
rect 200868 225332 200896 225508
rect 671712 225490 671764 225496
rect 201034 225428 201040 225480
rect 201092 225468 201098 225480
rect 242250 225468 242256 225480
rect 201092 225440 242256 225468
rect 201092 225428 201098 225440
rect 242250 225428 242256 225440
rect 242308 225428 242314 225480
rect 669406 225428 669412 225480
rect 669464 225468 669470 225480
rect 669464 225440 671622 225468
rect 669464 225428 669470 225440
rect 463142 225360 463148 225412
rect 463200 225400 463206 225412
rect 467282 225400 467288 225412
rect 463200 225372 467288 225400
rect 463200 225360 463206 225372
rect 467282 225360 467288 225372
rect 467340 225360 467346 225412
rect 207750 225332 207756 225344
rect 147180 225304 186268 225332
rect 147180 225292 147186 225304
rect 186240 225264 186268 225304
rect 186608 225304 200804 225332
rect 200868 225304 207756 225332
rect 186608 225264 186636 225304
rect 186240 225236 186636 225264
rect 185670 225196 185676 225208
rect 128320 225168 137232 225196
rect 137296 225168 185676 225196
rect 128320 225156 128326 225168
rect 126882 225020 126888 225072
rect 126940 225060 126946 225072
rect 137296 225060 137324 225168
rect 185670 225156 185676 225168
rect 185728 225156 185734 225208
rect 187326 225156 187332 225208
rect 187384 225196 187390 225208
rect 200574 225196 200580 225208
rect 187384 225168 200580 225196
rect 187384 225156 187390 225168
rect 200574 225156 200580 225168
rect 200632 225156 200638 225208
rect 200776 225196 200804 225304
rect 207750 225292 207756 225304
rect 207808 225292 207814 225344
rect 208026 225292 208032 225344
rect 208084 225332 208090 225344
rect 260926 225332 260932 225344
rect 208084 225304 260932 225332
rect 208084 225292 208090 225304
rect 260926 225292 260932 225304
rect 260984 225292 260990 225344
rect 671062 225224 671068 225276
rect 671120 225264 671126 225276
rect 671120 225236 671508 225264
rect 671120 225224 671126 225236
rect 202506 225196 202512 225208
rect 200776 225168 202512 225196
rect 202506 225156 202512 225168
rect 202564 225156 202570 225208
rect 202690 225156 202696 225208
rect 202748 225196 202754 225208
rect 254486 225196 254492 225208
rect 202748 225168 254492 225196
rect 202748 225156 202754 225168
rect 254486 225156 254492 225168
rect 254544 225156 254550 225208
rect 126940 225032 137324 225060
rect 126940 225020 126946 225032
rect 137462 225020 137468 225072
rect 137520 225060 137526 225072
rect 143534 225060 143540 225072
rect 137520 225032 143540 225060
rect 137520 225020 137526 225032
rect 143534 225020 143540 225032
rect 143592 225020 143598 225072
rect 146938 225020 146944 225072
rect 146996 225060 147002 225072
rect 162302 225060 162308 225072
rect 146996 225032 162308 225060
rect 146996 225020 147002 225032
rect 162302 225020 162308 225032
rect 162360 225020 162366 225072
rect 162486 225020 162492 225072
rect 162544 225060 162550 225072
rect 166442 225060 166448 225072
rect 162544 225032 166448 225060
rect 162544 225020 162550 225032
rect 166442 225020 166448 225032
rect 166500 225020 166506 225072
rect 166810 225020 166816 225072
rect 166868 225060 166874 225072
rect 166994 225060 167000 225072
rect 166868 225032 167000 225060
rect 166868 225020 166874 225032
rect 166994 225020 167000 225032
rect 167052 225020 167058 225072
rect 167362 225020 167368 225072
rect 167420 225060 167426 225072
rect 185670 225060 185676 225072
rect 167420 225032 185676 225060
rect 167420 225020 167426 225032
rect 185670 225020 185676 225032
rect 185728 225020 185734 225072
rect 187050 225020 187056 225072
rect 187108 225060 187114 225072
rect 223574 225060 223580 225072
rect 187108 225032 223580 225060
rect 187108 225020 187114 225032
rect 223574 225020 223580 225032
rect 223632 225020 223638 225072
rect 224862 225020 224868 225072
rect 224920 225060 224926 225072
rect 270586 225060 270592 225072
rect 224920 225032 270592 225060
rect 224920 225020 224926 225032
rect 270586 225020 270592 225032
rect 270644 225020 270650 225072
rect 668302 225020 668308 225072
rect 668360 225060 668366 225072
rect 668360 225032 671398 225060
rect 668360 225020 668366 225032
rect 275830 224952 275836 225004
rect 275888 224992 275894 225004
rect 276842 224992 276848 225004
rect 275888 224964 276848 224992
rect 275888 224952 275894 224964
rect 276842 224952 276848 224964
rect 276900 224952 276906 225004
rect 282730 224952 282736 225004
rect 282788 224992 282794 225004
rect 285306 224992 285312 225004
rect 282788 224964 285312 224992
rect 282788 224952 282794 224964
rect 285306 224952 285312 224964
rect 285364 224952 285370 225004
rect 489914 224952 489920 225004
rect 489972 224992 489978 225004
rect 494790 224992 494796 225004
rect 489972 224964 494796 224992
rect 489972 224952 489978 224964
rect 494790 224952 494796 224964
rect 494848 224952 494854 225004
rect 509234 224952 509240 225004
rect 509292 224992 509298 225004
rect 512638 224992 512644 225004
rect 509292 224964 512644 224992
rect 509292 224952 509298 224964
rect 512638 224952 512644 224964
rect 512696 224952 512702 225004
rect 122558 224884 122564 224936
rect 122616 224924 122622 224936
rect 193950 224924 193956 224936
rect 122616 224896 193956 224924
rect 122616 224884 122622 224896
rect 193950 224884 193956 224896
rect 194008 224884 194014 224936
rect 194502 224884 194508 224936
rect 194560 224924 194566 224936
rect 247402 224924 247408 224936
rect 194560 224896 247408 224924
rect 194560 224884 194566 224896
rect 247402 224884 247408 224896
rect 247460 224884 247466 224936
rect 264146 224884 264152 224936
rect 264204 224924 264210 224936
rect 269298 224924 269304 224936
rect 264204 224896 269304 224924
rect 264204 224884 264210 224896
rect 269298 224884 269304 224896
rect 269356 224884 269362 224936
rect 285674 224884 285680 224936
rect 285732 224924 285738 224936
rect 316310 224924 316316 224936
rect 285732 224896 316316 224924
rect 285732 224884 285738 224896
rect 316310 224884 316316 224896
rect 316368 224884 316374 224936
rect 406746 224884 406752 224936
rect 406804 224924 406810 224936
rect 414842 224924 414848 224936
rect 406804 224896 414848 224924
rect 406804 224884 406810 224896
rect 414842 224884 414848 224896
rect 414900 224884 414906 224936
rect 516778 224884 516784 224936
rect 516836 224924 516842 224936
rect 531314 224924 531320 224936
rect 516836 224896 531320 224924
rect 516836 224884 516842 224896
rect 531314 224884 531320 224896
rect 531372 224884 531378 224936
rect 667934 224884 667940 224936
rect 667992 224924 667998 224936
rect 668302 224924 668308 224936
rect 667992 224896 668308 224924
rect 667992 224884 667998 224896
rect 668302 224884 668308 224896
rect 668360 224884 668366 224936
rect 671062 224884 671068 224936
rect 671120 224924 671126 224936
rect 671120 224896 671278 224924
rect 671120 224884 671126 224896
rect 115842 224748 115848 224800
rect 115900 224788 115906 224800
rect 115900 224760 118372 224788
rect 115900 224748 115906 224760
rect 116762 224612 116768 224664
rect 116820 224652 116826 224664
rect 118142 224652 118148 224664
rect 116820 224624 118148 224652
rect 116820 224612 116826 224624
rect 118142 224612 118148 224624
rect 118200 224612 118206 224664
rect 118344 224652 118372 224760
rect 118786 224748 118792 224800
rect 118844 224788 118850 224800
rect 191374 224788 191380 224800
rect 118844 224760 191380 224788
rect 118844 224748 118850 224760
rect 191374 224748 191380 224760
rect 191432 224748 191438 224800
rect 192478 224748 192484 224800
rect 192536 224788 192542 224800
rect 246758 224788 246764 224800
rect 192536 224760 246764 224788
rect 192536 224748 192542 224760
rect 246758 224748 246764 224760
rect 246816 224748 246822 224800
rect 247586 224748 247592 224800
rect 247644 224788 247650 224800
rect 289262 224788 289268 224800
rect 247644 224760 289268 224788
rect 247644 224748 247650 224760
rect 289262 224748 289268 224760
rect 289320 224748 289326 224800
rect 315850 224748 315856 224800
rect 315908 224788 315914 224800
rect 341426 224788 341432 224800
rect 315908 224760 341432 224788
rect 315908 224748 315914 224760
rect 341426 224748 341432 224760
rect 341484 224748 341490 224800
rect 532418 224748 532424 224800
rect 532476 224788 532482 224800
rect 549898 224788 549904 224800
rect 532476 224760 549904 224788
rect 532476 224748 532482 224760
rect 549898 224748 549904 224760
rect 549956 224748 549962 224800
rect 460566 224680 460572 224732
rect 460624 224720 460630 224732
rect 463142 224720 463148 224732
rect 460624 224692 463148 224720
rect 460624 224680 460630 224692
rect 463142 224680 463148 224692
rect 463200 224680 463206 224732
rect 188798 224652 188804 224664
rect 118344 224624 188804 224652
rect 188798 224612 188804 224624
rect 188856 224612 188862 224664
rect 195606 224612 195612 224664
rect 195664 224652 195670 224664
rect 248874 224652 248880 224664
rect 195664 224624 248880 224652
rect 195664 224612 195670 224624
rect 248874 224612 248880 224624
rect 248932 224612 248938 224664
rect 249058 224612 249064 224664
rect 249116 224652 249122 224664
rect 263870 224652 263876 224664
rect 249116 224624 263876 224652
rect 249116 224612 249122 224624
rect 263870 224612 263876 224624
rect 263928 224612 263934 224664
rect 271598 224612 271604 224664
rect 271656 224652 271662 224664
rect 309870 224652 309876 224664
rect 271656 224624 309876 224652
rect 271656 224612 271662 224624
rect 309870 224612 309876 224624
rect 309928 224612 309934 224664
rect 319990 224612 319996 224664
rect 320048 224652 320054 224664
rect 347222 224652 347228 224664
rect 320048 224624 347228 224652
rect 320048 224612 320054 224624
rect 347222 224612 347228 224624
rect 347280 224612 347286 224664
rect 514662 224612 514668 224664
rect 514720 224652 514726 224664
rect 536650 224652 536656 224664
rect 514720 224624 536656 224652
rect 514720 224612 514726 224624
rect 536650 224612 536656 224624
rect 536708 224612 536714 224664
rect 667934 224612 667940 224664
rect 667992 224652 667998 224664
rect 667992 224624 671186 224652
rect 667992 224612 667998 224624
rect 456058 224544 456064 224596
rect 456116 224584 456122 224596
rect 459646 224584 459652 224596
rect 456116 224556 459652 224584
rect 456116 224544 456122 224556
rect 459646 224544 459652 224556
rect 459704 224544 459710 224596
rect 60642 224476 60648 224528
rect 60700 224516 60706 224528
rect 103606 224516 103612 224528
rect 60700 224488 103612 224516
rect 60700 224476 60706 224488
rect 103606 224476 103612 224488
rect 103664 224476 103670 224528
rect 108666 224476 108672 224528
rect 108724 224516 108730 224528
rect 118602 224516 118608 224528
rect 108724 224488 118608 224516
rect 108724 224476 108730 224488
rect 118602 224476 118608 224488
rect 118660 224476 118666 224528
rect 126698 224476 126704 224528
rect 126756 224516 126762 224528
rect 131114 224516 131120 224528
rect 126756 224488 131120 224516
rect 126756 224476 126762 224488
rect 131114 224476 131120 224488
rect 131172 224476 131178 224528
rect 131298 224476 131304 224528
rect 131356 224516 131362 224528
rect 196526 224516 196532 224528
rect 131356 224488 196532 224516
rect 131356 224476 131362 224488
rect 196526 224476 196532 224488
rect 196584 224476 196590 224528
rect 201218 224476 201224 224528
rect 201276 224516 201282 224528
rect 255774 224516 255780 224528
rect 201276 224488 255780 224516
rect 201276 224476 201282 224488
rect 255774 224476 255780 224488
rect 255832 224476 255838 224528
rect 261846 224476 261852 224528
rect 261904 224516 261910 224528
rect 300854 224516 300860 224528
rect 261904 224488 300860 224516
rect 261904 224476 261910 224488
rect 300854 224476 300860 224488
rect 300912 224476 300918 224528
rect 303246 224476 303252 224528
rect 303304 224516 303310 224528
rect 333054 224516 333060 224528
rect 303304 224488 333060 224516
rect 303304 224476 303310 224488
rect 333054 224476 333060 224488
rect 333112 224476 333118 224528
rect 333882 224476 333888 224528
rect 333940 224516 333946 224528
rect 356238 224516 356244 224528
rect 333940 224488 356244 224516
rect 333940 224476 333946 224488
rect 356238 224476 356244 224488
rect 356296 224476 356302 224528
rect 357342 224476 357348 224528
rect 357400 224516 357406 224528
rect 374270 224516 374276 224528
rect 357400 224488 374276 224516
rect 357400 224476 357406 224488
rect 374270 224476 374276 224488
rect 374328 224476 374334 224528
rect 479518 224476 479524 224528
rect 479576 224516 479582 224528
rect 486602 224516 486608 224528
rect 479576 224488 486608 224516
rect 479576 224476 479582 224488
rect 486602 224476 486608 224488
rect 486660 224476 486666 224528
rect 508222 224476 508228 224528
rect 508280 224516 508286 224528
rect 528370 224516 528376 224528
rect 508280 224488 528376 224516
rect 508280 224476 508286 224488
rect 528370 224476 528376 224488
rect 528428 224476 528434 224528
rect 530118 224476 530124 224528
rect 530176 224516 530182 224528
rect 556522 224516 556528 224528
rect 530176 224488 556528 224516
rect 530176 224476 530182 224488
rect 556522 224476 556528 224488
rect 556580 224476 556586 224528
rect 671022 224460 671074 224466
rect 671022 224402 671074 224408
rect 82722 224340 82728 224392
rect 82780 224380 82786 224392
rect 157288 224380 157294 224392
rect 82780 224352 157294 224380
rect 82780 224340 82786 224352
rect 157288 224340 157294 224352
rect 157346 224340 157352 224392
rect 157426 224340 157432 224392
rect 157484 224380 157490 224392
rect 170950 224380 170956 224392
rect 157484 224352 170956 224380
rect 157484 224340 157490 224352
rect 170950 224340 170956 224352
rect 171008 224340 171014 224392
rect 171088 224340 171094 224392
rect 171146 224380 171152 224392
rect 186866 224380 186872 224392
rect 171146 224352 186872 224380
rect 171146 224340 171152 224352
rect 186866 224340 186872 224352
rect 186924 224340 186930 224392
rect 188982 224340 188988 224392
rect 189040 224380 189046 224392
rect 243814 224380 243820 224392
rect 189040 224352 243820 224380
rect 189040 224340 189046 224352
rect 243814 224340 243820 224352
rect 243872 224340 243878 224392
rect 246942 224340 246948 224392
rect 247000 224380 247006 224392
rect 288618 224380 288624 224392
rect 247000 224352 288624 224380
rect 247000 224340 247006 224352
rect 288618 224340 288624 224352
rect 288676 224340 288682 224392
rect 289630 224340 289636 224392
rect 289688 224380 289694 224392
rect 307846 224380 307852 224392
rect 289688 224352 307852 224380
rect 289688 224340 289694 224352
rect 307846 224340 307852 224352
rect 307904 224340 307910 224392
rect 308950 224340 308956 224392
rect 309008 224380 309014 224392
rect 339494 224380 339500 224392
rect 309008 224352 339500 224380
rect 309008 224340 309014 224352
rect 339494 224340 339500 224352
rect 339552 224340 339558 224392
rect 344646 224340 344652 224392
rect 344704 224380 344710 224392
rect 364610 224380 364616 224392
rect 344704 224352 364616 224380
rect 344704 224340 344710 224352
rect 364610 224340 364616 224352
rect 364668 224340 364674 224392
rect 375282 224340 375288 224392
rect 375340 224380 375346 224392
rect 387794 224380 387800 224392
rect 375340 224352 387800 224380
rect 375340 224340 375346 224352
rect 387794 224340 387800 224352
rect 387852 224340 387858 224392
rect 462498 224340 462504 224392
rect 462556 224380 462562 224392
rect 469306 224380 469312 224392
rect 462556 224352 469312 224380
rect 462556 224340 462562 224352
rect 469306 224340 469312 224352
rect 469364 224340 469370 224392
rect 470226 224340 470232 224392
rect 470284 224380 470290 224392
rect 479702 224380 479708 224392
rect 470284 224352 479708 224380
rect 470284 224340 470290 224352
rect 479702 224340 479708 224352
rect 479760 224340 479766 224392
rect 486786 224340 486792 224392
rect 486844 224380 486850 224392
rect 496906 224380 496912 224392
rect 486844 224352 496912 224380
rect 486844 224340 486850 224352
rect 496906 224340 496912 224352
rect 496964 224340 496970 224392
rect 499206 224340 499212 224392
rect 499264 224380 499270 224392
rect 516778 224380 516784 224392
rect 499264 224352 516784 224380
rect 499264 224340 499270 224352
rect 516778 224340 516784 224352
rect 516836 224340 516842 224392
rect 525702 224340 525708 224392
rect 525760 224380 525766 224392
rect 550634 224380 550640 224392
rect 525760 224352 550640 224380
rect 525760 224340 525766 224352
rect 550634 224340 550640 224352
rect 550692 224340 550698 224392
rect 58986 224204 58992 224256
rect 59044 224244 59050 224256
rect 116762 224244 116768 224256
rect 59044 224216 116768 224244
rect 59044 224204 59050 224216
rect 116762 224204 116768 224216
rect 116820 224204 116826 224256
rect 116946 224204 116952 224256
rect 117004 224244 117010 224256
rect 118418 224244 118424 224256
rect 117004 224216 118424 224244
rect 117004 224204 117010 224216
rect 118418 224204 118424 224216
rect 118476 224204 118482 224256
rect 118602 224204 118608 224256
rect 118660 224244 118666 224256
rect 183830 224244 183836 224256
rect 118660 224216 183836 224244
rect 118660 224204 118666 224216
rect 183830 224204 183836 224216
rect 183888 224204 183894 224256
rect 184658 224204 184664 224256
rect 184716 224244 184722 224256
rect 239674 224244 239680 224256
rect 184716 224216 239680 224244
rect 184716 224204 184722 224216
rect 239674 224204 239680 224216
rect 239732 224204 239738 224256
rect 241974 224204 241980 224256
rect 242032 224244 242038 224256
rect 242032 224216 277394 224244
rect 242032 224204 242038 224216
rect 104802 224068 104808 224120
rect 104860 224108 104866 224120
rect 117958 224108 117964 224120
rect 104860 224080 117964 224108
rect 104860 224068 104866 224080
rect 117958 224068 117964 224080
rect 118016 224068 118022 224120
rect 118142 224068 118148 224120
rect 118200 224108 118206 224120
rect 118200 224080 142476 224108
rect 118200 224068 118206 224080
rect 76558 223932 76564 223984
rect 76616 223972 76622 223984
rect 142154 223972 142160 223984
rect 76616 223944 142160 223972
rect 76616 223932 76622 223944
rect 142154 223932 142160 223944
rect 142212 223932 142218 223984
rect 142448 223972 142476 224080
rect 142614 224068 142620 224120
rect 142672 224108 142678 224120
rect 209406 224108 209412 224120
rect 142672 224080 209412 224108
rect 142672 224068 142678 224080
rect 209406 224068 209412 224080
rect 209464 224068 209470 224120
rect 209682 224068 209688 224120
rect 209740 224108 209746 224120
rect 259638 224108 259644 224120
rect 209740 224080 259644 224108
rect 209740 224068 209746 224080
rect 259638 224068 259644 224080
rect 259696 224068 259702 224120
rect 277366 224108 277394 224216
rect 282546 224204 282552 224256
rect 282604 224244 282610 224256
rect 285674 224244 285680 224256
rect 282604 224216 285680 224244
rect 282604 224204 282610 224216
rect 285674 224204 285680 224216
rect 285732 224204 285738 224256
rect 288342 224204 288348 224256
rect 288400 224244 288406 224256
rect 322382 224244 322388 224256
rect 288400 224216 322388 224244
rect 288400 224204 288406 224216
rect 322382 224204 322388 224216
rect 322440 224204 322446 224256
rect 342070 224204 342076 224256
rect 342128 224244 342134 224256
rect 364794 224244 364800 224256
rect 342128 224216 364800 224244
rect 342128 224204 342134 224216
rect 364794 224204 364800 224216
rect 364852 224204 364858 224256
rect 364978 224204 364984 224256
rect 365036 224244 365042 224256
rect 378134 224244 378140 224256
rect 365036 224216 378140 224244
rect 365036 224204 365042 224216
rect 378134 224204 378140 224216
rect 378192 224204 378198 224256
rect 389082 224204 389088 224256
rect 389140 224244 389146 224256
rect 400950 224244 400956 224256
rect 389140 224216 400956 224244
rect 389140 224204 389146 224216
rect 400950 224204 400956 224216
rect 401008 224204 401014 224256
rect 416498 224204 416504 224256
rect 416556 224244 416562 224256
rect 422202 224244 422208 224256
rect 416556 224216 422208 224244
rect 416556 224204 416562 224216
rect 422202 224204 422208 224216
rect 422260 224204 422266 224256
rect 423306 224204 423312 224256
rect 423364 224244 423370 224256
rect 424318 224244 424324 224256
rect 423364 224216 424324 224244
rect 423364 224204 423370 224216
rect 424318 224204 424324 224216
rect 424376 224204 424382 224256
rect 451366 224204 451372 224256
rect 451424 224244 451430 224256
rect 452194 224244 452200 224256
rect 451424 224216 452200 224244
rect 451424 224204 451430 224216
rect 452194 224204 452200 224216
rect 452252 224204 452258 224256
rect 474734 224204 474740 224256
rect 474792 224244 474798 224256
rect 484578 224244 484584 224256
rect 474792 224216 484584 224244
rect 474792 224204 474798 224216
rect 484578 224204 484584 224216
rect 484636 224204 484642 224256
rect 485682 224204 485688 224256
rect 485740 224244 485746 224256
rect 499390 224244 499396 224256
rect 485740 224216 499396 224244
rect 485740 224204 485746 224216
rect 499390 224204 499396 224216
rect 499448 224204 499454 224256
rect 508866 224204 508872 224256
rect 508924 224244 508930 224256
rect 529382 224244 529388 224256
rect 508924 224216 529388 224244
rect 508924 224204 508930 224216
rect 529382 224204 529388 224216
rect 529440 224204 529446 224256
rect 535270 224204 535276 224256
rect 535328 224244 535334 224256
rect 563790 224244 563796 224256
rect 535328 224216 563796 224244
rect 535328 224204 535334 224216
rect 563790 224204 563796 224216
rect 563848 224204 563854 224256
rect 567838 224204 567844 224256
rect 567896 224244 567902 224256
rect 568942 224244 568948 224256
rect 567896 224216 568948 224244
rect 567896 224204 567902 224216
rect 568942 224204 568948 224216
rect 569000 224204 569006 224256
rect 669406 224136 669412 224188
rect 669464 224176 669470 224188
rect 669464 224148 670956 224176
rect 669464 224136 669470 224148
rect 285030 224108 285036 224120
rect 277366 224080 285036 224108
rect 285030 224068 285036 224080
rect 285088 224068 285094 224120
rect 286686 224068 286692 224120
rect 286744 224108 286750 224120
rect 319530 224108 319536 224120
rect 286744 224080 319536 224108
rect 286744 224068 286750 224080
rect 319530 224068 319536 224080
rect 319588 224068 319594 224120
rect 145190 223972 145196 223984
rect 142448 223944 145196 223972
rect 145190 223932 145196 223944
rect 145248 223932 145254 223984
rect 147674 223932 147680 223984
rect 147732 223972 147738 223984
rect 154574 223972 154580 223984
rect 147732 223944 154580 223972
rect 147732 223932 147738 223944
rect 154574 223932 154580 223944
rect 154632 223932 154638 223984
rect 156874 223932 156880 223984
rect 156932 223972 156938 223984
rect 217134 223972 217140 223984
rect 156932 223944 217140 223972
rect 156932 223932 156938 223944
rect 217134 223932 217140 223944
rect 217192 223932 217198 223984
rect 217318 223932 217324 223984
rect 217376 223972 217382 223984
rect 228082 223972 228088 223984
rect 217376 223944 228088 223972
rect 217376 223932 217382 223944
rect 228082 223932 228088 223944
rect 228140 223932 228146 223984
rect 231302 223932 231308 223984
rect 231360 223972 231366 223984
rect 278958 223972 278964 223984
rect 231360 223944 278964 223972
rect 231360 223932 231366 223944
rect 278958 223932 278964 223944
rect 279016 223932 279022 223984
rect 117958 223796 117964 223848
rect 118016 223836 118022 223848
rect 122926 223836 122932 223848
rect 118016 223808 122932 223836
rect 118016 223796 118022 223808
rect 122926 223796 122932 223808
rect 122984 223796 122990 223848
rect 125226 223796 125232 223848
rect 125284 223836 125290 223848
rect 131298 223836 131304 223848
rect 125284 223808 131304 223836
rect 125284 223796 125290 223808
rect 131298 223796 131304 223808
rect 131356 223796 131362 223848
rect 134978 223796 134984 223848
rect 135036 223836 135042 223848
rect 204254 223836 204260 223848
rect 135036 223808 204260 223836
rect 135036 223796 135042 223808
rect 204254 223796 204260 223808
rect 204312 223796 204318 223848
rect 205266 223796 205272 223848
rect 205324 223836 205330 223848
rect 212626 223836 212632 223848
rect 205324 223808 212632 223836
rect 205324 223796 205330 223808
rect 212626 223796 212632 223808
rect 212684 223796 212690 223848
rect 215938 223796 215944 223848
rect 215996 223836 216002 223848
rect 222930 223836 222936 223848
rect 215996 223808 222936 223836
rect 215996 223796 216002 223808
rect 222930 223796 222936 223808
rect 222988 223796 222994 223848
rect 238662 223796 238668 223848
rect 238720 223836 238726 223848
rect 282362 223836 282368 223848
rect 238720 223808 282368 223836
rect 238720 223796 238726 223808
rect 282362 223796 282368 223808
rect 282420 223796 282426 223848
rect 132402 223660 132408 223712
rect 132460 223700 132466 223712
rect 201678 223700 201684 223712
rect 132460 223672 201684 223700
rect 132460 223660 132466 223672
rect 201678 223660 201684 223672
rect 201736 223660 201742 223712
rect 297836 223672 300348 223700
rect 85482 223524 85488 223576
rect 85540 223564 85546 223576
rect 161934 223564 161940 223576
rect 85540 223536 161940 223564
rect 85540 223524 85546 223536
rect 161934 223524 161940 223536
rect 161992 223524 161998 223576
rect 162118 223524 162124 223576
rect 162176 223564 162182 223576
rect 167822 223564 167828 223576
rect 162176 223536 167828 223564
rect 162176 223524 162182 223536
rect 167822 223524 167828 223536
rect 167880 223524 167886 223576
rect 168282 223524 168288 223576
rect 168340 223564 168346 223576
rect 226702 223564 226708 223576
rect 168340 223536 226708 223564
rect 168340 223524 168346 223536
rect 226702 223524 226708 223536
rect 226760 223524 226766 223576
rect 269022 223524 269028 223576
rect 269080 223564 269086 223576
rect 297836 223564 297864 223672
rect 269080 223536 297864 223564
rect 269080 223524 269086 223536
rect 298002 223524 298008 223576
rect 298060 223564 298066 223576
rect 300118 223564 300124 223576
rect 298060 223536 300124 223564
rect 298060 223524 298066 223536
rect 300118 223524 300124 223536
rect 300176 223524 300182 223576
rect 300320 223564 300348 223672
rect 426434 223592 426440 223644
rect 426492 223632 426498 223644
rect 426986 223632 426992 223644
rect 426492 223604 426992 223632
rect 426492 223592 426498 223604
rect 426986 223592 426992 223604
rect 427044 223592 427050 223644
rect 306006 223564 306012 223576
rect 300320 223536 306012 223564
rect 306006 223524 306012 223536
rect 306064 223524 306070 223576
rect 329098 223524 329104 223576
rect 329156 223564 329162 223576
rect 342714 223564 342720 223576
rect 329156 223536 342720 223564
rect 329156 223524 329162 223536
rect 342714 223524 342720 223536
rect 342772 223524 342778 223576
rect 457990 223524 457996 223576
rect 458048 223564 458054 223576
rect 460198 223564 460204 223576
rect 458048 223536 460204 223564
rect 458048 223524 458054 223536
rect 460198 223524 460204 223536
rect 460256 223524 460262 223576
rect 473446 223524 473452 223576
rect 473504 223564 473510 223576
rect 475562 223564 475568 223576
rect 473504 223536 475568 223564
rect 473504 223524 473510 223536
rect 475562 223524 475568 223536
rect 475620 223524 475626 223576
rect 679250 223524 679256 223576
rect 679308 223564 679314 223576
rect 680170 223564 680176 223576
rect 679308 223536 680176 223564
rect 679308 223524 679314 223536
rect 680170 223524 680176 223536
rect 680228 223524 680234 223576
rect 112806 223388 112812 223440
rect 112864 223428 112870 223440
rect 185854 223428 185860 223440
rect 112864 223400 185860 223428
rect 112864 223388 112870 223400
rect 185854 223388 185860 223400
rect 185912 223388 185918 223440
rect 203886 223388 203892 223440
rect 203944 223428 203950 223440
rect 254854 223428 254860 223440
rect 203944 223400 254860 223428
rect 203944 223388 203950 223400
rect 254854 223388 254860 223400
rect 254912 223388 254918 223440
rect 260098 223388 260104 223440
rect 260156 223428 260162 223440
rect 298922 223428 298928 223440
rect 260156 223400 298928 223428
rect 260156 223388 260162 223400
rect 298922 223388 298928 223400
rect 298980 223388 298986 223440
rect 302142 223388 302148 223440
rect 302200 223428 302206 223440
rect 331122 223428 331128 223440
rect 302200 223400 331128 223428
rect 302200 223388 302206 223400
rect 331122 223388 331128 223400
rect 331180 223388 331186 223440
rect 518894 223388 518900 223440
rect 518952 223428 518958 223440
rect 530026 223428 530032 223440
rect 518952 223400 530032 223428
rect 518952 223388 518958 223400
rect 530026 223388 530032 223400
rect 530084 223388 530090 223440
rect 81342 223252 81348 223304
rect 81400 223292 81406 223304
rect 156874 223292 156880 223304
rect 81400 223264 156880 223292
rect 81400 223252 81406 223264
rect 156874 223252 156880 223264
rect 156932 223252 156938 223304
rect 157426 223252 157432 223304
rect 157484 223292 157490 223304
rect 159818 223292 159824 223304
rect 157484 223264 159824 223292
rect 157484 223252 157490 223264
rect 159818 223252 159824 223264
rect 159876 223252 159882 223304
rect 160922 223252 160928 223304
rect 160980 223292 160986 223304
rect 164510 223292 164516 223304
rect 160980 223264 164516 223292
rect 160980 223252 160986 223264
rect 164510 223252 164516 223264
rect 164568 223252 164574 223304
rect 224034 223292 224040 223304
rect 164942 223264 224040 223292
rect 78582 223116 78588 223168
rect 78640 223156 78646 223168
rect 157058 223156 157064 223168
rect 78640 223128 157064 223156
rect 78640 223116 78646 223128
rect 157058 223116 157064 223128
rect 157116 223116 157122 223168
rect 157242 223116 157248 223168
rect 157300 223156 157306 223168
rect 161198 223156 161204 223168
rect 157300 223128 161204 223156
rect 157300 223116 157306 223128
rect 161198 223116 161204 223128
rect 161256 223116 161262 223168
rect 161382 223116 161388 223168
rect 161440 223156 161446 223168
rect 161440 223128 162348 223156
rect 161440 223116 161446 223128
rect 89438 222980 89444 223032
rect 89496 223020 89502 223032
rect 162118 223020 162124 223032
rect 89496 222992 162124 223020
rect 89496 222980 89502 222992
rect 162118 222980 162124 222992
rect 162176 222980 162182 223032
rect 162320 223020 162348 223128
rect 164142 223116 164148 223168
rect 164200 223156 164206 223168
rect 164942 223156 164970 223264
rect 224034 223252 224040 223264
rect 224092 223252 224098 223304
rect 264790 223252 264796 223304
rect 264848 223292 264854 223304
rect 304718 223292 304724 223304
rect 264848 223264 304724 223292
rect 264848 223252 264854 223264
rect 304718 223252 304724 223264
rect 304776 223252 304782 223304
rect 306282 223252 306288 223304
rect 306340 223292 306346 223304
rect 336918 223292 336924 223304
rect 306340 223264 336924 223292
rect 306340 223252 306346 223264
rect 336918 223252 336924 223264
rect 336976 223252 336982 223304
rect 343542 223252 343548 223304
rect 343600 223292 343606 223304
rect 363966 223292 363972 223304
rect 343600 223264 363972 223292
rect 343600 223252 343606 223264
rect 363966 223252 363972 223264
rect 364024 223252 364030 223304
rect 489546 223252 489552 223304
rect 489604 223292 489610 223304
rect 504358 223292 504364 223304
rect 489604 223264 504364 223292
rect 489604 223252 489610 223264
rect 504358 223252 504364 223264
rect 504416 223252 504422 223304
rect 505094 223252 505100 223304
rect 505152 223292 505158 223304
rect 523954 223292 523960 223304
rect 505152 223264 523960 223292
rect 505152 223252 505158 223264
rect 523954 223252 523960 223264
rect 524012 223252 524018 223304
rect 529014 223252 529020 223304
rect 529072 223292 529078 223304
rect 543642 223292 543648 223304
rect 529072 223264 543648 223292
rect 529072 223252 529078 223264
rect 543642 223252 543648 223264
rect 543700 223252 543706 223304
rect 164200 223128 164970 223156
rect 164200 223116 164206 223128
rect 165062 223116 165068 223168
rect 165120 223156 165126 223168
rect 222286 223156 222292 223168
rect 165120 223128 222292 223156
rect 165120 223116 165126 223128
rect 222286 223116 222292 223128
rect 222344 223116 222350 223168
rect 224218 223116 224224 223168
rect 224276 223156 224282 223168
rect 238386 223156 238392 223168
rect 224276 223128 238392 223156
rect 224276 223116 224282 223128
rect 238386 223116 238392 223128
rect 238444 223116 238450 223168
rect 245286 223116 245292 223168
rect 245344 223156 245350 223168
rect 287606 223156 287612 223168
rect 245344 223128 287612 223156
rect 245344 223116 245350 223128
rect 287606 223116 287612 223128
rect 287664 223116 287670 223168
rect 290826 223116 290832 223168
rect 290884 223156 290890 223168
rect 323670 223156 323676 223168
rect 290884 223128 323676 223156
rect 290884 223116 290890 223128
rect 323670 223116 323676 223128
rect 323728 223116 323734 223168
rect 330478 223116 330484 223168
rect 330536 223156 330542 223168
rect 354950 223156 354956 223168
rect 330536 223128 354956 223156
rect 330536 223116 330542 223128
rect 354950 223116 354956 223128
rect 355008 223116 355014 223168
rect 357066 223116 357072 223168
rect 357124 223156 357130 223168
rect 376202 223156 376208 223168
rect 357124 223128 376208 223156
rect 357124 223116 357130 223128
rect 376202 223116 376208 223128
rect 376260 223116 376266 223168
rect 490190 223116 490196 223168
rect 490248 223156 490254 223168
rect 505646 223156 505652 223168
rect 490248 223128 505652 223156
rect 490248 223116 490254 223128
rect 505646 223116 505652 223128
rect 505704 223116 505710 223168
rect 513098 223116 513104 223168
rect 513156 223156 513162 223168
rect 534442 223156 534448 223168
rect 513156 223128 534448 223156
rect 513156 223116 513162 223128
rect 534442 223116 534448 223128
rect 534500 223116 534506 223168
rect 534718 223116 534724 223168
rect 534776 223156 534782 223168
rect 547414 223156 547420 223168
rect 534776 223128 547420 223156
rect 534776 223116 534782 223128
rect 547414 223116 547420 223128
rect 547472 223116 547478 223168
rect 162320 222992 166626 223020
rect 92106 222844 92112 222896
rect 92164 222884 92170 222896
rect 166442 222884 166448 222896
rect 92164 222856 166448 222884
rect 92164 222844 92170 222856
rect 166442 222844 166448 222856
rect 166500 222844 166506 222896
rect 166598 222884 166626 222992
rect 166948 222980 166954 223032
rect 167006 223020 167012 223032
rect 176102 223020 176108 223032
rect 167006 222992 176108 223020
rect 167006 222980 167012 222992
rect 176102 222980 176108 222992
rect 176160 222980 176166 223032
rect 176286 222980 176292 223032
rect 176344 223020 176350 223032
rect 234798 223020 234804 223032
rect 176344 222992 234804 223020
rect 176344 222980 176350 222992
rect 234798 222980 234804 222992
rect 234856 222980 234862 223032
rect 235166 222980 235172 223032
rect 235224 223020 235230 223032
rect 243262 223020 243268 223032
rect 235224 222992 243268 223020
rect 235224 222980 235230 222992
rect 243262 222980 243268 222992
rect 243320 222980 243326 223032
rect 250898 222980 250904 223032
rect 250956 223020 250962 223032
rect 294414 223020 294420 223032
rect 250956 222992 294420 223020
rect 250956 222980 250962 222992
rect 294414 222980 294420 222992
rect 294472 222980 294478 223032
rect 300302 222980 300308 223032
rect 300360 223020 300366 223032
rect 331306 223020 331312 223032
rect 300360 222992 331312 223020
rect 300360 222980 300366 222992
rect 331306 222980 331312 222992
rect 331364 222980 331370 223032
rect 337930 222980 337936 223032
rect 337988 223020 337994 223032
rect 359182 223020 359188 223032
rect 337988 222992 359188 223020
rect 337988 222980 337994 222992
rect 359182 222980 359188 222992
rect 359240 222980 359246 223032
rect 370498 222980 370504 223032
rect 370556 223020 370562 223032
rect 384574 223020 384580 223032
rect 370556 222992 384580 223020
rect 370556 222980 370562 222992
rect 384574 222980 384580 222992
rect 384632 222980 384638 223032
rect 387702 222980 387708 223032
rect 387760 223020 387766 223032
rect 398098 223020 398104 223032
rect 387760 222992 398104 223020
rect 387760 222980 387766 222992
rect 398098 222980 398104 222992
rect 398156 222980 398162 223032
rect 501782 222980 501788 223032
rect 501840 223020 501846 223032
rect 519262 223020 519268 223032
rect 501840 222992 519268 223020
rect 501840 222980 501846 222992
rect 519262 222980 519268 222992
rect 519320 222980 519326 223032
rect 523678 222980 523684 223032
rect 523736 223020 523742 223032
rect 548058 223020 548064 223032
rect 523736 222992 548064 223020
rect 523736 222980 523742 222992
rect 548058 222980 548064 222992
rect 548116 222980 548122 223032
rect 549254 222980 549260 223032
rect 549312 223020 549318 223032
rect 564802 223020 564808 223032
rect 549312 222992 564808 223020
rect 549312 222980 549318 222992
rect 564802 222980 564808 222992
rect 564860 222980 564866 223032
rect 566826 222912 566832 222964
rect 566884 222952 566890 222964
rect 576394 222952 576400 222964
rect 566884 222924 576400 222952
rect 566884 222912 566890 222924
rect 576394 222912 576400 222924
rect 576452 222912 576458 222964
rect 221642 222884 221648 222896
rect 166598 222856 221648 222884
rect 221642 222844 221648 222856
rect 221700 222844 221706 222896
rect 231946 222844 231952 222896
rect 232004 222884 232010 222896
rect 277670 222884 277676 222896
rect 232004 222856 277676 222884
rect 232004 222844 232010 222856
rect 277670 222844 277676 222856
rect 277728 222844 277734 222896
rect 283374 222844 283380 222896
rect 283432 222884 283438 222896
rect 316954 222884 316960 222896
rect 283432 222856 316960 222884
rect 283432 222844 283438 222856
rect 316954 222844 316960 222856
rect 317012 222844 317018 222896
rect 317138 222844 317144 222896
rect 317196 222884 317202 222896
rect 343358 222884 343364 222896
rect 317196 222856 343364 222884
rect 317196 222844 317202 222856
rect 343358 222844 343364 222856
rect 343416 222844 343422 222896
rect 347590 222844 347596 222896
rect 347648 222884 347654 222896
rect 368474 222884 368480 222896
rect 347648 222856 368480 222884
rect 347648 222844 347654 222856
rect 368474 222844 368480 222856
rect 368532 222844 368538 222896
rect 375098 222844 375104 222896
rect 375156 222884 375162 222896
rect 391014 222884 391020 222896
rect 375156 222856 391020 222884
rect 375156 222844 375162 222856
rect 391014 222844 391020 222856
rect 391072 222844 391078 222896
rect 397362 222844 397368 222896
rect 397420 222884 397426 222896
rect 407114 222884 407120 222896
rect 397420 222856 407120 222884
rect 397420 222844 397426 222856
rect 407114 222844 407120 222856
rect 407172 222844 407178 222896
rect 408402 222844 408408 222896
rect 408460 222884 408466 222896
rect 416866 222884 416872 222896
rect 408460 222856 416872 222884
rect 408460 222844 408466 222856
rect 416866 222844 416872 222856
rect 416924 222844 416930 222896
rect 420822 222844 420828 222896
rect 420880 222884 420886 222896
rect 425146 222884 425152 222896
rect 420880 222856 425152 222884
rect 420880 222844 420886 222856
rect 425146 222844 425152 222856
rect 425204 222844 425210 222896
rect 459922 222844 459928 222896
rect 459980 222884 459986 222896
rect 467098 222884 467104 222896
rect 459980 222856 467104 222884
rect 459980 222844 459986 222856
rect 467098 222844 467104 222856
rect 467156 222844 467162 222896
rect 467466 222844 467472 222896
rect 467524 222884 467530 222896
rect 473722 222884 473728 222896
rect 467524 222856 473728 222884
rect 467524 222844 467530 222856
rect 473722 222844 473728 222856
rect 473780 222844 473786 222896
rect 478322 222844 478328 222896
rect 478380 222884 478386 222896
rect 486142 222884 486148 222896
rect 478380 222856 486148 222884
rect 478380 222844 478386 222856
rect 486142 222844 486148 222856
rect 486200 222844 486206 222896
rect 486970 222844 486976 222896
rect 487028 222884 487034 222896
rect 501046 222884 501052 222896
rect 487028 222856 501052 222884
rect 487028 222844 487034 222856
rect 501046 222844 501052 222856
rect 501104 222844 501110 222896
rect 504634 222844 504640 222896
rect 504692 222884 504698 222896
rect 523770 222884 523776 222896
rect 504692 222856 523776 222884
rect 504692 222844 504698 222856
rect 523770 222844 523776 222856
rect 523828 222844 523834 222896
rect 533706 222844 533712 222896
rect 533764 222884 533770 222896
rect 560662 222884 560668 222896
rect 533764 222856 560668 222884
rect 533764 222844 533770 222856
rect 560662 222844 560668 222856
rect 560720 222844 560726 222896
rect 563790 222776 563796 222828
rect 563848 222816 563854 222828
rect 569954 222816 569960 222828
rect 563848 222788 569960 222816
rect 563848 222776 563854 222788
rect 569954 222776 569960 222788
rect 570012 222776 570018 222828
rect 87966 222708 87972 222760
rect 88024 222748 88030 222760
rect 160922 222748 160928 222760
rect 88024 222720 160928 222748
rect 88024 222708 88030 222720
rect 160922 222708 160928 222720
rect 160980 222708 160986 222760
rect 161198 222708 161204 222760
rect 161256 222748 161262 222760
rect 161256 222720 175964 222748
rect 161256 222708 161262 222720
rect 99282 222572 99288 222624
rect 99340 222612 99346 222624
rect 175458 222612 175464 222624
rect 99340 222584 175464 222612
rect 99340 222572 99346 222584
rect 175458 222572 175464 222584
rect 175516 222572 175522 222624
rect 175936 222612 175964 222720
rect 176102 222708 176108 222760
rect 176160 222748 176166 222760
rect 192018 222748 192024 222760
rect 176160 222720 192024 222748
rect 176160 222708 176166 222720
rect 192018 222708 192024 222720
rect 192076 222708 192082 222760
rect 192294 222708 192300 222760
rect 192352 222748 192358 222760
rect 207474 222748 207480 222760
rect 192352 222720 207480 222748
rect 192352 222708 192358 222720
rect 207474 222708 207480 222720
rect 207532 222708 207538 222760
rect 209498 222708 209504 222760
rect 209556 222748 209562 222760
rect 210234 222748 210240 222760
rect 209556 222720 210240 222748
rect 209556 222708 209562 222720
rect 210234 222708 210240 222720
rect 210292 222708 210298 222760
rect 213822 222708 213828 222760
rect 213880 222748 213886 222760
rect 262858 222748 262864 222760
rect 213880 222720 262864 222748
rect 213880 222708 213886 222720
rect 262858 222708 262864 222720
rect 262916 222708 262922 222760
rect 263502 222708 263508 222760
rect 263560 222748 263566 222760
rect 296898 222748 296904 222760
rect 263560 222720 296904 222748
rect 263560 222708 263566 222720
rect 296898 222708 296904 222720
rect 296956 222708 296962 222760
rect 562502 222640 562508 222692
rect 562560 222680 562566 222692
rect 564618 222680 564624 222692
rect 562560 222652 564624 222680
rect 562560 222640 562566 222652
rect 564618 222640 564624 222652
rect 564676 222640 564682 222692
rect 564802 222640 564808 222692
rect 564860 222680 564866 222692
rect 574094 222680 574100 222692
rect 564860 222652 574100 222680
rect 564860 222640 564866 222652
rect 574094 222640 574100 222652
rect 574152 222640 574158 222692
rect 175936 222584 214604 222612
rect 56502 222436 56508 222488
rect 56560 222476 56566 222488
rect 56560 222448 122834 222476
rect 56560 222436 56566 222448
rect 122806 222340 122834 222448
rect 133506 222436 133512 222488
rect 133564 222476 133570 222488
rect 142982 222476 142988 222488
rect 133564 222448 142988 222476
rect 133564 222436 133570 222448
rect 142982 222436 142988 222448
rect 143040 222436 143046 222488
rect 143350 222436 143356 222488
rect 143408 222476 143414 222488
rect 144822 222476 144828 222488
rect 143408 222448 144828 222476
rect 143408 222436 143414 222448
rect 144822 222436 144828 222448
rect 144880 222436 144886 222488
rect 145006 222436 145012 222488
rect 145064 222476 145070 222488
rect 151354 222476 151360 222488
rect 145064 222448 151360 222476
rect 145064 222436 145070 222448
rect 151354 222436 151360 222448
rect 151412 222436 151418 222488
rect 154206 222436 154212 222488
rect 154264 222476 154270 222488
rect 214374 222476 214380 222488
rect 154264 222448 214380 222476
rect 154264 222436 154270 222448
rect 214374 222436 214380 222448
rect 214432 222436 214438 222488
rect 214576 222476 214604 222584
rect 214742 222572 214748 222624
rect 214800 222612 214806 222624
rect 260282 222612 260288 222624
rect 214800 222584 260288 222612
rect 214800 222572 214806 222584
rect 260282 222572 260288 222584
rect 260340 222572 260346 222624
rect 571702 222544 571708 222556
rect 563440 222516 571708 222544
rect 219710 222476 219716 222488
rect 214576 222448 219716 222476
rect 219710 222436 219716 222448
rect 219768 222436 219774 222488
rect 220078 222436 220084 222488
rect 220136 222476 220142 222488
rect 268654 222476 268660 222488
rect 220136 222448 268660 222476
rect 220136 222436 220142 222448
rect 268654 222436 268660 222448
rect 268712 222436 268718 222488
rect 142338 222340 142344 222352
rect 122806 222312 142344 222340
rect 142338 222300 142344 222312
rect 142396 222300 142402 222352
rect 144270 222300 144276 222352
rect 144328 222340 144334 222352
rect 208762 222340 208768 222352
rect 144328 222312 208768 222340
rect 144328 222300 144334 222312
rect 208762 222300 208768 222312
rect 208820 222300 208826 222352
rect 210970 222300 210976 222352
rect 211028 222340 211034 222352
rect 214742 222340 214748 222352
rect 211028 222312 214748 222340
rect 211028 222300 211034 222312
rect 214742 222300 214748 222312
rect 214800 222300 214806 222352
rect 220446 222300 220452 222352
rect 220504 222340 220510 222352
rect 268010 222340 268016 222352
rect 220504 222312 268016 222340
rect 220504 222300 220510 222312
rect 268010 222300 268016 222312
rect 268068 222300 268074 222352
rect 214926 222232 214932 222284
rect 214984 222272 214990 222284
rect 216214 222272 216220 222284
rect 214984 222244 216220 222272
rect 214984 222232 214990 222244
rect 216214 222232 216220 222244
rect 216272 222232 216278 222284
rect 562502 222272 562508 222284
rect 543706 222244 562508 222272
rect 171244 222176 171456 222204
rect 107838 222096 107844 222148
rect 107896 222136 107902 222148
rect 171042 222136 171048 222148
rect 107896 222108 171048 222136
rect 107896 222096 107902 222108
rect 171042 222096 171048 222108
rect 171100 222096 171106 222148
rect 104526 221960 104532 222012
rect 104584 222000 104590 222012
rect 171244 222000 171272 222176
rect 171428 222136 171456 222176
rect 173084 222176 173204 222204
rect 173084 222136 173112 222176
rect 171428 222108 173112 222136
rect 173176 222068 173204 222176
rect 174906 222164 174912 222216
rect 174964 222204 174970 222216
rect 176286 222204 176292 222216
rect 174964 222176 176292 222204
rect 174964 222164 174970 222176
rect 176286 222164 176292 222176
rect 176344 222164 176350 222216
rect 482922 222164 482928 222216
rect 482980 222204 482986 222216
rect 543706 222204 543734 222244
rect 562502 222232 562508 222244
rect 562560 222232 562566 222284
rect 563440 222204 563468 222516
rect 571702 222504 571708 222516
rect 571760 222504 571766 222556
rect 572806 222544 572812 222556
rect 572686 222516 572812 222544
rect 567378 222368 567384 222420
rect 567436 222408 567442 222420
rect 572686 222408 572714 222516
rect 572806 222504 572812 222516
rect 572864 222504 572870 222556
rect 593966 222408 593972 222420
rect 567436 222380 572714 222408
rect 582346 222380 593972 222408
rect 567436 222368 567442 222380
rect 564618 222232 564624 222284
rect 564676 222272 564682 222284
rect 582346 222272 582374 222380
rect 593966 222368 593972 222380
rect 594024 222368 594030 222420
rect 597554 222272 597560 222284
rect 564676 222244 582374 222272
rect 593064 222244 597560 222272
rect 564676 222232 564682 222244
rect 482980 222176 543734 222204
rect 563348 222194 563468 222204
rect 563256 222176 563468 222194
rect 482980 222164 482986 222176
rect 563256 222166 563376 222176
rect 178218 222096 178224 222148
rect 178276 222136 178282 222148
rect 178276 222108 180794 222136
rect 178276 222096 178282 222108
rect 176102 222068 176108 222080
rect 173176 222040 176108 222068
rect 176102 222028 176108 222040
rect 176160 222028 176166 222080
rect 172974 222000 172980 222012
rect 104584 221972 171272 222000
rect 171336 221972 172980 222000
rect 104584 221960 104590 221972
rect 71406 221824 71412 221876
rect 71464 221864 71470 221876
rect 71464 221836 147812 221864
rect 71464 221824 71470 221836
rect 68094 221688 68100 221740
rect 68152 221728 68158 221740
rect 142108 221728 142114 221740
rect 68152 221700 142114 221728
rect 68152 221688 68158 221700
rect 142108 221688 142114 221700
rect 142166 221688 142172 221740
rect 142338 221688 142344 221740
rect 142396 221728 142402 221740
rect 144454 221728 144460 221740
rect 142396 221700 144460 221728
rect 142396 221688 142402 221700
rect 144454 221688 144460 221700
rect 144512 221688 144518 221740
rect 146202 221688 146208 221740
rect 146260 221728 146266 221740
rect 147784 221728 147812 221836
rect 149238 221824 149244 221876
rect 149296 221864 149302 221876
rect 149296 221836 157334 221864
rect 149296 221824 149302 221836
rect 152090 221728 152096 221740
rect 146260 221700 147674 221728
rect 147784 221700 152096 221728
rect 146260 221688 146266 221700
rect 61470 221552 61476 221604
rect 61528 221592 61534 221604
rect 137278 221592 137284 221604
rect 61528 221564 137284 221592
rect 61528 221552 61534 221564
rect 137278 221552 137284 221564
rect 137336 221552 137342 221604
rect 137462 221552 137468 221604
rect 137520 221592 137526 221604
rect 147646 221592 147674 221700
rect 152090 221688 152096 221700
rect 152148 221688 152154 221740
rect 157306 221728 157334 221836
rect 162118 221824 162124 221876
rect 162176 221864 162182 221876
rect 171336 221864 171364 221972
rect 172974 221960 172980 221972
rect 173032 221960 173038 222012
rect 176286 221960 176292 222012
rect 176344 222000 176350 222012
rect 180610 222000 180616 222012
rect 176344 221972 180616 222000
rect 176344 221960 176350 221972
rect 180610 221960 180616 221972
rect 180668 221960 180674 222012
rect 180766 222000 180794 222108
rect 181622 222096 181628 222148
rect 181680 222136 181686 222148
rect 240134 222136 240140 222148
rect 181680 222108 240140 222136
rect 181680 222096 181686 222108
rect 240134 222096 240140 222108
rect 240192 222096 240198 222148
rect 261018 222096 261024 222148
rect 261076 222136 261082 222148
rect 301682 222136 301688 222148
rect 261076 222108 301688 222136
rect 261076 222096 261082 222108
rect 301682 222096 301688 222108
rect 301740 222096 301746 222148
rect 331398 222096 331404 222148
rect 331456 222136 331462 222148
rect 353938 222136 353944 222148
rect 331456 222108 353944 222136
rect 331456 222096 331462 222108
rect 353938 222096 353944 222108
rect 353996 222096 354002 222148
rect 424962 222096 424968 222148
rect 425020 222136 425026 222148
rect 429286 222136 429292 222148
rect 425020 222108 429292 222136
rect 425020 222096 425026 222108
rect 429286 222096 429292 222108
rect 429344 222096 429350 222148
rect 462130 222096 462136 222148
rect 462188 222136 462194 222148
rect 468754 222136 468760 222148
rect 462188 222108 468760 222136
rect 462188 222096 462194 222108
rect 468754 222096 468760 222108
rect 468812 222096 468818 222148
rect 471882 222096 471888 222148
rect 471940 222136 471946 222148
rect 477862 222136 477868 222148
rect 471940 222108 477868 222136
rect 471940 222096 471946 222108
rect 477862 222096 477868 222108
rect 477920 222096 477926 222148
rect 553578 222096 553584 222148
rect 553636 222136 553642 222148
rect 553636 222108 562916 222136
rect 553636 222096 553642 222108
rect 562888 222068 562916 222108
rect 563256 222068 563284 222166
rect 563698 222096 563704 222148
rect 563756 222136 563762 222148
rect 593064 222136 593092 222244
rect 597554 222232 597560 222244
rect 597612 222232 597618 222284
rect 563756 222108 593092 222136
rect 563756 222096 563762 222108
rect 593230 222096 593236 222148
rect 593288 222136 593294 222148
rect 607490 222136 607496 222148
rect 593288 222108 607496 222136
rect 593288 222096 593294 222108
rect 607490 222096 607496 222108
rect 607548 222096 607554 222148
rect 562888 222040 563284 222068
rect 237558 222000 237564 222012
rect 180766 221972 237564 222000
rect 237558 221960 237564 221972
rect 237616 221960 237622 222012
rect 243630 221960 243636 222012
rect 243688 222000 243694 222012
rect 285858 222000 285864 222012
rect 243688 221972 285864 222000
rect 243688 221960 243694 221972
rect 285858 221960 285864 221972
rect 285916 221960 285922 222012
rect 309870 221960 309876 222012
rect 309928 222000 309934 222012
rect 338390 222000 338396 222012
rect 309928 221972 338396 222000
rect 309928 221960 309934 221972
rect 338390 221960 338396 221972
rect 338448 221960 338454 222012
rect 529750 221960 529756 222012
rect 529808 222000 529814 222012
rect 555786 222000 555792 222012
rect 529808 221972 555792 222000
rect 529808 221960 529814 221972
rect 555786 221960 555792 221972
rect 555844 221960 555850 222012
rect 556798 221960 556804 222012
rect 556856 222000 556862 222012
rect 562686 222000 562692 222012
rect 556856 221972 562692 222000
rect 556856 221960 556862 221972
rect 562686 221960 562692 221972
rect 562744 221960 562750 222012
rect 563422 221960 563428 222012
rect 563480 222000 563486 222012
rect 569310 222000 569316 222012
rect 563480 221972 569316 222000
rect 563480 221960 563486 221972
rect 569310 221960 569316 221972
rect 569368 221960 569374 222012
rect 569586 221960 569592 222012
rect 569644 222000 569650 222012
rect 596450 222000 596456 222012
rect 569644 221972 596456 222000
rect 569644 221960 569650 221972
rect 596450 221960 596456 221972
rect 596508 221960 596514 222012
rect 596634 221960 596640 222012
rect 596692 222000 596698 222012
rect 596692 221972 597048 222000
rect 596692 221960 596698 221972
rect 162176 221836 171364 221864
rect 162176 221824 162182 221836
rect 171502 221824 171508 221876
rect 171560 221864 171566 221876
rect 229646 221864 229652 221876
rect 171560 221836 229652 221864
rect 171560 221824 171566 221836
rect 229646 221824 229652 221836
rect 229704 221824 229710 221876
rect 230382 221824 230388 221876
rect 230440 221864 230446 221876
rect 258718 221864 258724 221876
rect 230440 221836 258724 221864
rect 230440 221824 230446 221836
rect 258718 221824 258724 221836
rect 258776 221824 258782 221876
rect 267826 221824 267832 221876
rect 267884 221864 267890 221876
rect 273990 221864 273996 221876
rect 267884 221836 273996 221864
rect 267884 221824 267890 221836
rect 273990 221824 273996 221836
rect 274048 221824 274054 221876
rect 303706 221824 303712 221876
rect 303764 221864 303770 221876
rect 334066 221864 334072 221876
rect 303764 221836 334072 221864
rect 303764 221824 303770 221836
rect 334066 221824 334072 221836
rect 334124 221824 334130 221876
rect 496170 221824 496176 221876
rect 496228 221864 496234 221876
rect 513374 221864 513380 221876
rect 496228 221836 513380 221864
rect 496228 221824 496234 221836
rect 513374 221824 513380 221836
rect 513432 221824 513438 221876
rect 515398 221824 515404 221876
rect 515456 221864 515462 221876
rect 534994 221864 535000 221876
rect 515456 221836 535000 221864
rect 515456 221824 515462 221836
rect 534994 221824 535000 221836
rect 535052 221824 535058 221876
rect 545114 221824 545120 221876
rect 545172 221864 545178 221876
rect 596818 221864 596824 221876
rect 545172 221836 596824 221864
rect 545172 221824 545178 221836
rect 596818 221824 596824 221836
rect 596876 221824 596882 221876
rect 597020 221864 597048 221972
rect 597186 221960 597192 222012
rect 597244 222000 597250 222012
rect 607306 222000 607312 222012
rect 597244 221972 607312 222000
rect 597244 221960 597250 221972
rect 607306 221960 607312 221972
rect 607364 221960 607370 222012
rect 606018 221864 606024 221876
rect 597020 221836 606024 221864
rect 606018 221824 606024 221836
rect 606076 221824 606082 221876
rect 162302 221728 162308 221740
rect 157306 221700 162308 221728
rect 162302 221688 162308 221700
rect 162360 221688 162366 221740
rect 162670 221688 162676 221740
rect 162728 221728 162734 221740
rect 224494 221728 224500 221740
rect 162728 221700 224500 221728
rect 162728 221688 162734 221700
rect 224494 221688 224500 221700
rect 224552 221688 224558 221740
rect 227070 221688 227076 221740
rect 227128 221728 227134 221740
rect 272702 221728 272708 221740
rect 227128 221700 272708 221728
rect 227128 221688 227134 221700
rect 272702 221688 272708 221700
rect 272760 221688 272766 221740
rect 275094 221688 275100 221740
rect 275152 221728 275158 221740
rect 310882 221728 310888 221740
rect 275152 221700 310888 221728
rect 275152 221688 275158 221700
rect 310882 221688 310888 221700
rect 310940 221688 310946 221740
rect 311526 221688 311532 221740
rect 311584 221728 311590 221740
rect 338574 221728 338580 221740
rect 311584 221700 338580 221728
rect 311584 221688 311590 221700
rect 338574 221688 338580 221700
rect 338632 221688 338638 221740
rect 341610 221728 341616 221740
rect 338776 221700 341616 221728
rect 204898 221592 204904 221604
rect 137520 221564 146984 221592
rect 147646 221564 204904 221592
rect 137520 221552 137526 221564
rect 64598 221416 64604 221468
rect 64656 221456 64662 221468
rect 142108 221456 142114 221468
rect 64656 221428 142114 221456
rect 64656 221416 64662 221428
rect 142108 221416 142114 221428
rect 142166 221416 142172 221468
rect 142246 221416 142252 221468
rect 142304 221456 142310 221468
rect 143994 221456 144000 221468
rect 142304 221428 144000 221456
rect 142304 221416 142310 221428
rect 143994 221416 144000 221428
rect 144052 221416 144058 221468
rect 144454 221416 144460 221468
rect 144512 221456 144518 221468
rect 146662 221456 146668 221468
rect 144512 221428 146668 221456
rect 144512 221416 144518 221428
rect 146662 221416 146668 221428
rect 146720 221416 146726 221468
rect 146956 221456 146984 221564
rect 204898 221552 204904 221564
rect 204956 221552 204962 221604
rect 205082 221552 205088 221604
rect 205140 221592 205146 221604
rect 214190 221592 214196 221604
rect 205140 221564 214196 221592
rect 205140 221552 205146 221564
rect 214190 221552 214196 221564
rect 214248 221552 214254 221604
rect 214650 221552 214656 221604
rect 214708 221592 214714 221604
rect 258534 221592 258540 221604
rect 214708 221564 258540 221592
rect 214708 221552 214714 221564
rect 258534 221552 258540 221564
rect 258592 221552 258598 221604
rect 258718 221552 258724 221604
rect 258776 221592 258782 221604
rect 275278 221592 275284 221604
rect 258776 221564 275284 221592
rect 258776 221552 258782 221564
rect 275278 221552 275284 221564
rect 275336 221552 275342 221604
rect 278314 221552 278320 221604
rect 278372 221592 278378 221604
rect 313274 221592 313280 221604
rect 278372 221564 313280 221592
rect 278372 221552 278378 221564
rect 313274 221552 313280 221564
rect 313332 221552 313338 221604
rect 314470 221552 314476 221604
rect 314528 221592 314534 221604
rect 338776 221592 338804 221700
rect 341610 221688 341616 221700
rect 341668 221688 341674 221740
rect 359550 221688 359556 221740
rect 359608 221728 359614 221740
rect 376846 221728 376852 221740
rect 359608 221700 376852 221728
rect 359608 221688 359614 221700
rect 376846 221688 376852 221700
rect 376904 221688 376910 221740
rect 500034 221688 500040 221740
rect 500092 221728 500098 221740
rect 518434 221728 518440 221740
rect 500092 221700 518440 221728
rect 500092 221688 500098 221700
rect 518434 221688 518440 221700
rect 518492 221688 518498 221740
rect 522850 221688 522856 221740
rect 522908 221728 522914 221740
rect 546586 221728 546592 221740
rect 522908 221700 546592 221728
rect 522908 221688 522914 221700
rect 546586 221688 546592 221700
rect 546644 221688 546650 221740
rect 547138 221688 547144 221740
rect 547196 221728 547202 221740
rect 556706 221728 556712 221740
rect 547196 221700 556712 221728
rect 547196 221688 547202 221700
rect 556706 221688 556712 221700
rect 556764 221688 556770 221740
rect 557810 221688 557816 221740
rect 557868 221728 557874 221740
rect 558270 221728 558276 221740
rect 557868 221700 558276 221728
rect 557868 221688 557874 221700
rect 558270 221688 558276 221700
rect 558328 221728 558334 221740
rect 562870 221728 562876 221740
rect 558328 221700 562876 221728
rect 558328 221688 558334 221700
rect 562870 221688 562876 221700
rect 562928 221688 562934 221740
rect 563054 221688 563060 221740
rect 563112 221728 563118 221740
rect 566642 221728 566648 221740
rect 563112 221700 566648 221728
rect 563112 221688 563118 221700
rect 566642 221688 566648 221700
rect 566700 221728 566706 221740
rect 567378 221728 567384 221740
rect 566700 221700 567384 221728
rect 566700 221688 566706 221700
rect 567378 221688 567384 221700
rect 567436 221688 567442 221740
rect 567746 221688 567752 221740
rect 567804 221728 567810 221740
rect 569586 221728 569592 221740
rect 567804 221700 569592 221728
rect 567804 221688 567810 221700
rect 569586 221688 569592 221700
rect 569644 221688 569650 221740
rect 569954 221688 569960 221740
rect 570012 221728 570018 221740
rect 610526 221728 610532 221740
rect 570012 221700 610532 221728
rect 570012 221688 570018 221700
rect 610526 221688 610532 221700
rect 610584 221688 610590 221740
rect 314528 221564 338804 221592
rect 314528 221552 314534 221564
rect 341334 221552 341340 221604
rect 341392 221592 341398 221604
rect 361574 221592 361580 221604
rect 341392 221564 361580 221592
rect 341392 221552 341398 221564
rect 361574 221552 361580 221564
rect 361632 221552 361638 221604
rect 362218 221592 362224 221604
rect 361776 221564 362224 221592
rect 162118 221456 162124 221468
rect 146956 221428 162124 221456
rect 162118 221416 162124 221428
rect 162176 221416 162182 221468
rect 162302 221416 162308 221468
rect 162360 221456 162366 221468
rect 162360 221428 185624 221456
rect 162360 221416 162366 221428
rect 95418 221280 95424 221332
rect 95476 221320 95482 221332
rect 95476 221292 103514 221320
rect 95476 221280 95482 221292
rect 103486 221184 103514 221292
rect 114462 221280 114468 221332
rect 114520 221320 114526 221332
rect 185118 221320 185124 221332
rect 114520 221292 185124 221320
rect 114520 221280 114526 221292
rect 185118 221280 185124 221292
rect 185176 221280 185182 221332
rect 185596 221320 185624 221428
rect 185762 221416 185768 221468
rect 185820 221456 185826 221468
rect 232130 221456 232136 221468
rect 185820 221428 232136 221456
rect 185820 221416 185826 221428
rect 232130 221416 232136 221428
rect 232188 221416 232194 221468
rect 241146 221416 241152 221468
rect 241204 221456 241210 221468
rect 285858 221456 285864 221468
rect 241204 221428 285864 221456
rect 241204 221416 241210 221428
rect 285858 221416 285864 221428
rect 285916 221416 285922 221468
rect 286042 221416 286048 221468
rect 286100 221456 286106 221468
rect 289814 221456 289820 221468
rect 286100 221428 289820 221456
rect 286100 221416 286106 221428
rect 289814 221416 289820 221428
rect 289872 221416 289878 221468
rect 289998 221416 290004 221468
rect 290056 221456 290062 221468
rect 321738 221456 321744 221468
rect 290056 221428 321744 221456
rect 290056 221416 290062 221428
rect 321738 221416 321744 221428
rect 321796 221416 321802 221468
rect 338850 221416 338856 221468
rect 338908 221456 338914 221468
rect 361776 221456 361804 221564
rect 362218 221552 362224 221564
rect 362276 221552 362282 221604
rect 377766 221552 377772 221604
rect 377824 221592 377830 221604
rect 390002 221592 390008 221604
rect 377824 221564 390008 221592
rect 377824 221552 377830 221564
rect 390002 221552 390008 221564
rect 390060 221552 390066 221604
rect 456702 221552 456708 221604
rect 456760 221592 456766 221604
rect 462130 221592 462136 221604
rect 456760 221564 462136 221592
rect 456760 221552 456766 221564
rect 462130 221552 462136 221564
rect 462188 221552 462194 221604
rect 484302 221552 484308 221604
rect 484360 221592 484366 221604
rect 496078 221592 496084 221604
rect 484360 221564 496084 221592
rect 484360 221552 484366 221564
rect 496078 221552 496084 221564
rect 496136 221552 496142 221604
rect 503438 221552 503444 221604
rect 503496 221592 503502 221604
rect 521746 221592 521752 221604
rect 503496 221564 521752 221592
rect 503496 221552 503502 221564
rect 521746 221552 521752 221564
rect 521804 221552 521810 221604
rect 525886 221552 525892 221604
rect 525944 221592 525950 221604
rect 601510 221592 601516 221604
rect 525944 221564 601516 221592
rect 525944 221552 525950 221564
rect 601510 221552 601516 221564
rect 601568 221552 601574 221604
rect 606662 221592 606668 221604
rect 601666 221564 606668 221592
rect 338908 221428 361804 221456
rect 338908 221416 338914 221428
rect 362034 221416 362040 221468
rect 362092 221456 362098 221468
rect 379882 221456 379888 221468
rect 362092 221428 379888 221456
rect 362092 221416 362098 221428
rect 379882 221416 379888 221428
rect 379940 221416 379946 221468
rect 391014 221416 391020 221468
rect 391072 221456 391078 221468
rect 400398 221456 400404 221468
rect 391072 221428 400404 221456
rect 391072 221416 391078 221428
rect 400398 221416 400404 221428
rect 400456 221416 400462 221468
rect 405090 221416 405096 221468
rect 405148 221456 405154 221468
rect 414198 221456 414204 221468
rect 405148 221428 414204 221456
rect 405148 221416 405154 221428
rect 414198 221416 414204 221428
rect 414256 221416 414262 221468
rect 452562 221416 452568 221468
rect 452620 221456 452626 221468
rect 456702 221456 456708 221468
rect 452620 221428 456708 221456
rect 452620 221416 452626 221428
rect 456702 221416 456708 221428
rect 456760 221416 456766 221468
rect 483750 221416 483756 221468
rect 483808 221456 483814 221468
rect 538674 221456 538680 221468
rect 483808 221428 538680 221456
rect 483808 221416 483814 221428
rect 538674 221416 538680 221428
rect 538732 221416 538738 221468
rect 543274 221416 543280 221468
rect 543332 221456 543338 221468
rect 596634 221456 596640 221468
rect 543332 221428 596640 221456
rect 543332 221416 543338 221428
rect 596634 221416 596640 221428
rect 596692 221416 596698 221468
rect 596818 221416 596824 221468
rect 596876 221456 596882 221468
rect 601666 221456 601694 221564
rect 606662 221552 606668 221564
rect 606720 221552 606726 221604
rect 655698 221552 655704 221604
rect 655756 221592 655762 221604
rect 659286 221592 659292 221604
rect 655756 221564 659292 221592
rect 655756 221552 655762 221564
rect 659286 221552 659292 221564
rect 659344 221552 659350 221604
rect 596876 221428 601694 221456
rect 596876 221416 596882 221428
rect 654226 221416 654232 221468
rect 654284 221456 654290 221468
rect 655514 221456 655520 221468
rect 654284 221428 655520 221456
rect 654284 221416 654290 221428
rect 655514 221416 655520 221428
rect 655572 221416 655578 221468
rect 195238 221320 195244 221332
rect 185596 221292 195244 221320
rect 195238 221280 195244 221292
rect 195296 221280 195302 221332
rect 195422 221280 195428 221332
rect 195480 221320 195486 221332
rect 245102 221320 245108 221332
rect 195480 221292 245108 221320
rect 195480 221280 195486 221292
rect 245102 221280 245108 221292
rect 245160 221280 245166 221332
rect 258534 221280 258540 221332
rect 258592 221320 258598 221332
rect 265710 221320 265716 221332
rect 258592 221292 265716 221320
rect 258592 221280 258598 221292
rect 265710 221280 265716 221292
rect 265768 221280 265774 221332
rect 273438 221280 273444 221332
rect 273496 221320 273502 221332
rect 309226 221320 309232 221332
rect 273496 221292 309232 221320
rect 273496 221280 273502 221292
rect 309226 221280 309232 221292
rect 309284 221280 309290 221332
rect 542906 221212 542912 221264
rect 542964 221252 542970 221264
rect 550358 221252 550364 221264
rect 542964 221224 550364 221252
rect 542964 221212 542970 221224
rect 550358 221212 550364 221224
rect 550416 221212 550422 221264
rect 550634 221212 550640 221264
rect 550692 221252 550698 221264
rect 551278 221252 551284 221264
rect 550692 221224 551284 221252
rect 550692 221212 550698 221224
rect 551278 221212 551284 221224
rect 551336 221252 551342 221264
rect 569126 221252 569132 221264
rect 551336 221224 569132 221252
rect 551336 221212 551342 221224
rect 569126 221212 569132 221224
rect 569184 221212 569190 221264
rect 569310 221212 569316 221264
rect 569368 221252 569374 221264
rect 610066 221252 610072 221264
rect 569368 221224 610072 221252
rect 569368 221212 569374 221224
rect 610066 221212 610072 221224
rect 610124 221212 610130 221264
rect 137094 221184 137100 221196
rect 103486 221156 137100 221184
rect 137094 221144 137100 221156
rect 137152 221144 137158 221196
rect 137278 221144 137284 221196
rect 137336 221184 137342 221196
rect 142108 221184 142114 221196
rect 137336 221156 142114 221184
rect 137336 221144 137342 221156
rect 142108 221144 142114 221156
rect 142166 221144 142172 221196
rect 142246 221144 142252 221196
rect 142304 221184 142310 221196
rect 203242 221184 203248 221196
rect 142304 221156 203248 221184
rect 142304 221144 142310 221156
rect 203242 221144 203248 221156
rect 203300 221144 203306 221196
rect 205082 221184 205088 221196
rect 204732 221156 205088 221184
rect 117774 221008 117780 221060
rect 117832 221048 117838 221060
rect 180748 221048 180754 221060
rect 117832 221020 180754 221048
rect 117832 221008 117838 221020
rect 180748 221008 180754 221020
rect 180806 221008 180812 221060
rect 180886 221008 180892 221060
rect 180944 221048 180950 221060
rect 185762 221048 185768 221060
rect 180944 221020 185768 221048
rect 180944 221008 180950 221020
rect 185762 221008 185768 221020
rect 185820 221008 185826 221060
rect 185946 221008 185952 221060
rect 186004 221048 186010 221060
rect 187878 221048 187884 221060
rect 186004 221020 187884 221048
rect 186004 221008 186010 221020
rect 187878 221008 187884 221020
rect 187936 221008 187942 221060
rect 188154 221008 188160 221060
rect 188212 221048 188218 221060
rect 188212 221020 195100 221048
rect 188212 221008 188218 221020
rect 128538 220872 128544 220924
rect 128596 220912 128602 220924
rect 195072 220912 195100 221020
rect 195238 221008 195244 221060
rect 195296 221048 195302 221060
rect 204732 221048 204760 221156
rect 205082 221144 205088 221156
rect 205140 221144 205146 221196
rect 206002 221144 206008 221196
rect 206060 221184 206066 221196
rect 258350 221184 258356 221196
rect 206060 221156 258356 221184
rect 206060 221144 206066 221156
rect 258350 221144 258356 221156
rect 258408 221144 258414 221196
rect 548058 221076 548064 221128
rect 548116 221116 548122 221128
rect 593230 221116 593236 221128
rect 548116 221088 593236 221116
rect 548116 221076 548122 221088
rect 593230 221076 593236 221088
rect 593288 221076 593294 221128
rect 596450 221076 596456 221128
rect 596508 221116 596514 221128
rect 596508 221088 597416 221116
rect 596508 221076 596514 221088
rect 195296 221020 204760 221048
rect 195296 221008 195302 221020
rect 204898 221008 204904 221060
rect 204956 221048 204962 221060
rect 211614 221048 211620 221060
rect 204956 221020 211620 221048
rect 204956 221008 204962 221020
rect 211614 221008 211620 221020
rect 211672 221008 211678 221060
rect 237098 221008 237104 221060
rect 237156 221048 237162 221060
rect 280430 221048 280436 221060
rect 237156 221020 280436 221048
rect 237156 221008 237162 221020
rect 280430 221008 280436 221020
rect 280488 221008 280494 221060
rect 415026 221008 415032 221060
rect 415084 221048 415090 221060
rect 420178 221048 420184 221060
rect 415084 221020 420184 221048
rect 415084 221008 415090 221020
rect 420178 221008 420184 221020
rect 420236 221008 420242 221060
rect 545114 221008 545120 221060
rect 545172 221048 545178 221060
rect 545758 221048 545764 221060
rect 545172 221020 545764 221048
rect 545172 221008 545178 221020
rect 545758 221008 545764 221020
rect 545816 221008 545822 221060
rect 552842 220940 552848 220992
rect 552900 220980 552906 220992
rect 553210 220980 553216 220992
rect 552900 220952 553216 220980
rect 552900 220940 552906 220952
rect 553210 220940 553216 220952
rect 553268 220980 553274 220992
rect 567746 220980 567752 220992
rect 553268 220952 567752 220980
rect 553268 220940 553274 220952
rect 567746 220940 567752 220952
rect 567804 220940 567810 220992
rect 569126 220940 569132 220992
rect 569184 220980 569190 220992
rect 597186 220980 597192 220992
rect 569184 220952 597192 220980
rect 569184 220940 569190 220952
rect 597186 220940 597192 220952
rect 597244 220940 597250 220992
rect 597388 220980 597416 221088
rect 597554 221076 597560 221128
rect 597612 221116 597618 221128
rect 608686 221116 608692 221128
rect 597612 221088 608692 221116
rect 597612 221076 597618 221088
rect 608686 221076 608692 221088
rect 608744 221076 608750 221128
rect 608870 220980 608876 220992
rect 597388 220952 608876 220980
rect 608870 220940 608876 220952
rect 608928 220940 608934 220992
rect 195422 220912 195428 220924
rect 128596 220884 195008 220912
rect 195072 220884 195428 220912
rect 128596 220872 128602 220884
rect 91278 220736 91284 220788
rect 91336 220776 91342 220788
rect 91336 220748 162164 220776
rect 91336 220736 91342 220748
rect 97718 220600 97724 220652
rect 97776 220640 97782 220652
rect 162136 220640 162164 220748
rect 162302 220736 162308 220788
rect 162360 220776 162366 220788
rect 172698 220776 172704 220788
rect 162360 220748 172704 220776
rect 162360 220736 162366 220748
rect 172698 220736 172704 220748
rect 172756 220736 172762 220788
rect 173342 220736 173348 220788
rect 173400 220776 173406 220788
rect 182634 220776 182640 220788
rect 173400 220748 182640 220776
rect 173400 220736 173406 220748
rect 182634 220736 182640 220748
rect 182692 220736 182698 220788
rect 183094 220736 183100 220788
rect 183152 220776 183158 220788
rect 184198 220776 184204 220788
rect 183152 220748 184204 220776
rect 183152 220736 183158 220748
rect 184198 220736 184204 220748
rect 184256 220736 184262 220788
rect 190454 220736 190460 220788
rect 190512 220776 190518 220788
rect 194778 220776 194784 220788
rect 190512 220748 194784 220776
rect 190512 220736 190518 220748
rect 194778 220736 194784 220748
rect 194836 220736 194842 220788
rect 194980 220776 195008 220884
rect 195422 220872 195428 220884
rect 195480 220872 195486 220924
rect 198918 220912 198924 220924
rect 195624 220884 198924 220912
rect 195624 220776 195652 220884
rect 198918 220872 198924 220884
rect 198976 220872 198982 220924
rect 203242 220872 203248 220924
rect 203300 220912 203306 220924
rect 206370 220912 206376 220924
rect 203300 220884 206376 220912
rect 203300 220872 203306 220884
rect 206370 220872 206376 220884
rect 206428 220872 206434 220924
rect 256050 220872 256056 220924
rect 256108 220912 256114 220924
rect 261386 220912 261392 220924
rect 256108 220884 261392 220912
rect 256108 220872 256114 220884
rect 261386 220872 261392 220884
rect 261444 220872 261450 220924
rect 420638 220804 420644 220856
rect 420696 220844 420702 220856
rect 423766 220844 423772 220856
rect 420696 220816 423772 220844
rect 420696 220804 420702 220816
rect 423766 220804 423772 220816
rect 423824 220804 423830 220856
rect 466086 220804 466092 220856
rect 466144 220844 466150 220856
rect 470594 220844 470600 220856
rect 466144 220816 470600 220844
rect 466144 220804 466150 220816
rect 470594 220804 470600 220816
rect 470652 220804 470658 220856
rect 518434 220804 518440 220856
rect 518492 220844 518498 220856
rect 591942 220844 591948 220856
rect 518492 220816 591948 220844
rect 518492 220804 518498 220816
rect 591942 220804 591948 220816
rect 592000 220804 592006 220856
rect 194980 220748 195652 220776
rect 196066 220736 196072 220788
rect 196124 220776 196130 220788
rect 197722 220776 197728 220788
rect 196124 220748 197728 220776
rect 196124 220736 196130 220748
rect 197722 220736 197728 220748
rect 197780 220736 197786 220788
rect 198090 220736 198096 220788
rect 198148 220776 198154 220788
rect 252738 220776 252744 220788
rect 198148 220748 252744 220776
rect 198148 220736 198154 220748
rect 252738 220736 252744 220748
rect 252796 220736 252802 220788
rect 253566 220736 253572 220788
rect 253624 220776 253630 220788
rect 293310 220776 293316 220788
rect 253624 220748 293316 220776
rect 253624 220736 253630 220748
rect 293310 220736 293316 220748
rect 293368 220736 293374 220788
rect 293586 220736 293592 220788
rect 293644 220776 293650 220788
rect 299934 220776 299940 220788
rect 293644 220748 299940 220776
rect 293644 220736 293650 220748
rect 299934 220736 299940 220748
rect 299992 220736 299998 220788
rect 306742 220736 306748 220788
rect 306800 220776 306806 220788
rect 320358 220776 320364 220788
rect 306800 220748 320364 220776
rect 306800 220736 306806 220748
rect 320358 220736 320364 220748
rect 320416 220736 320422 220788
rect 329558 220736 329564 220788
rect 329616 220776 329622 220788
rect 331950 220776 331956 220788
rect 329616 220748 331956 220776
rect 329616 220736 329622 220748
rect 331950 220736 331956 220748
rect 332008 220736 332014 220788
rect 414198 220736 414204 220788
rect 414256 220776 414262 220788
rect 418246 220776 418252 220788
rect 414256 220748 418252 220776
rect 414256 220736 414262 220748
rect 418246 220736 418252 220748
rect 418304 220736 418310 220788
rect 455230 220736 455236 220788
rect 455288 220776 455294 220788
rect 458818 220776 458824 220788
rect 455288 220748 458824 220776
rect 455288 220736 455294 220748
rect 458818 220736 458824 220748
rect 458876 220736 458882 220788
rect 475378 220736 475384 220788
rect 475436 220776 475442 220788
rect 476206 220776 476212 220788
rect 475436 220748 476212 220776
rect 475436 220736 475442 220748
rect 476206 220736 476212 220748
rect 476264 220736 476270 220788
rect 476758 220736 476764 220788
rect 476816 220776 476822 220788
rect 478690 220776 478696 220788
rect 476816 220748 478696 220776
rect 476816 220736 476822 220748
rect 478690 220736 478696 220748
rect 478748 220736 478754 220788
rect 504174 220736 504180 220788
rect 504232 220776 504238 220788
rect 515766 220776 515772 220788
rect 504232 220748 515772 220776
rect 504232 220736 504238 220748
rect 515766 220736 515772 220748
rect 515824 220736 515830 220788
rect 592126 220736 592132 220788
rect 592184 220776 592190 220788
rect 620278 220776 620284 220788
rect 592184 220748 620284 220776
rect 592184 220736 592190 220748
rect 620278 220736 620284 220748
rect 620336 220736 620342 220788
rect 465718 220668 465724 220720
rect 465776 220708 465782 220720
rect 469582 220708 469588 220720
rect 465776 220680 469588 220708
rect 465776 220668 465782 220680
rect 469582 220668 469588 220680
rect 469640 220668 469646 220720
rect 676030 220668 676036 220720
rect 676088 220708 676094 220720
rect 677410 220708 677416 220720
rect 676088 220680 677416 220708
rect 676088 220668 676094 220680
rect 677410 220668 677416 220680
rect 677468 220668 677474 220720
rect 167178 220640 167184 220652
rect 97776 220612 162072 220640
rect 162136 220612 167184 220640
rect 97776 220600 97782 220612
rect 82998 220464 83004 220516
rect 83056 220504 83062 220516
rect 157334 220504 157340 220516
rect 83056 220476 157340 220504
rect 83056 220464 83062 220476
rect 157334 220464 157340 220476
rect 157392 220464 157398 220516
rect 157518 220464 157524 220516
rect 157576 220504 157582 220516
rect 162044 220504 162072 220612
rect 167178 220600 167184 220612
rect 167236 220600 167242 220652
rect 170766 220600 170772 220652
rect 170824 220640 170830 220652
rect 170824 220612 173756 220640
rect 170824 220600 170830 220612
rect 162302 220504 162308 220516
rect 157576 220476 161980 220504
rect 162044 220476 162308 220504
rect 157576 220464 157582 220476
rect 76374 220328 76380 220380
rect 76432 220368 76438 220380
rect 150710 220368 150716 220380
rect 76432 220340 150716 220368
rect 76432 220328 76438 220340
rect 150710 220328 150716 220340
rect 150768 220328 150774 220380
rect 150894 220328 150900 220380
rect 150952 220368 150958 220380
rect 161750 220368 161756 220380
rect 150952 220340 161756 220368
rect 150952 220328 150958 220340
rect 161750 220328 161756 220340
rect 161808 220328 161814 220380
rect 161952 220368 161980 220476
rect 162302 220464 162308 220476
rect 162360 220464 162366 220516
rect 162854 220464 162860 220516
rect 162912 220504 162918 220516
rect 173526 220504 173532 220516
rect 162912 220476 173532 220504
rect 162912 220464 162918 220476
rect 173526 220464 173532 220476
rect 173584 220464 173590 220516
rect 173728 220504 173756 220612
rect 177390 220600 177396 220652
rect 177448 220640 177454 220652
rect 234062 220640 234068 220652
rect 177448 220612 234068 220640
rect 177448 220600 177454 220612
rect 234062 220600 234068 220612
rect 234120 220600 234126 220652
rect 254394 220600 254400 220652
rect 254452 220640 254458 220652
rect 296714 220640 296720 220652
rect 254452 220612 296720 220640
rect 254452 220600 254458 220612
rect 296714 220600 296720 220612
rect 296772 220600 296778 220652
rect 299934 220600 299940 220652
rect 299992 220640 299998 220652
rect 330018 220640 330024 220652
rect 299992 220612 330024 220640
rect 299992 220600 299998 220612
rect 330018 220600 330024 220612
rect 330076 220600 330082 220652
rect 473998 220600 474004 220652
rect 474056 220640 474062 220652
rect 475378 220640 475384 220652
rect 474056 220612 475384 220640
rect 474056 220600 474062 220612
rect 475378 220600 475384 220612
rect 475436 220600 475442 220652
rect 511258 220600 511264 220652
rect 511316 220640 511322 220652
rect 527542 220640 527548 220652
rect 511316 220612 527548 220640
rect 511316 220600 511322 220612
rect 527542 220600 527548 220612
rect 527600 220600 527606 220652
rect 542722 220600 542728 220652
rect 542780 220640 542786 220652
rect 543642 220640 543648 220652
rect 542780 220612 543648 220640
rect 542780 220600 542786 220612
rect 543642 220600 543648 220612
rect 543700 220640 543706 220652
rect 545942 220640 545948 220652
rect 543700 220612 545948 220640
rect 543700 220600 543706 220612
rect 545942 220600 545948 220612
rect 546000 220600 546006 220652
rect 546126 220600 546132 220652
rect 546184 220640 546190 220652
rect 550266 220640 550272 220652
rect 546184 220612 550272 220640
rect 546184 220600 546190 220612
rect 550266 220600 550272 220612
rect 550324 220600 550330 220652
rect 550542 220600 550548 220652
rect 550600 220640 550606 220652
rect 553762 220640 553768 220652
rect 550600 220612 553768 220640
rect 550600 220600 550606 220612
rect 553762 220600 553768 220612
rect 553820 220600 553826 220652
rect 555602 220600 555608 220652
rect 555660 220640 555666 220652
rect 559834 220640 559840 220652
rect 555660 220612 559840 220640
rect 555660 220600 555666 220612
rect 559834 220600 559840 220612
rect 559892 220640 559898 220652
rect 626626 220640 626632 220652
rect 559892 220612 626632 220640
rect 559892 220600 559898 220612
rect 626626 220600 626632 220612
rect 626684 220600 626690 220652
rect 229278 220504 229284 220516
rect 173728 220476 229284 220504
rect 229278 220464 229284 220476
rect 229336 220464 229342 220516
rect 240318 220464 240324 220516
rect 240376 220504 240382 220516
rect 283006 220504 283012 220516
rect 240376 220476 283012 220504
rect 240376 220464 240382 220476
rect 283006 220464 283012 220476
rect 283064 220464 283070 220516
rect 296622 220464 296628 220516
rect 296680 220504 296686 220516
rect 327534 220504 327540 220516
rect 296680 220476 327540 220504
rect 296680 220464 296686 220476
rect 327534 220464 327540 220476
rect 327592 220464 327598 220516
rect 328086 220464 328092 220516
rect 328144 220504 328150 220516
rect 351362 220504 351368 220516
rect 328144 220476 351368 220504
rect 328144 220464 328150 220476
rect 351362 220464 351368 220476
rect 351420 220464 351426 220516
rect 371142 220464 371148 220516
rect 371200 220504 371206 220516
rect 385218 220504 385224 220516
rect 371200 220476 385224 220504
rect 371200 220464 371206 220476
rect 385218 220464 385224 220476
rect 385276 220464 385282 220516
rect 482278 220464 482284 220516
rect 482336 220504 482342 220516
rect 491938 220504 491944 220516
rect 482336 220476 491944 220504
rect 482336 220464 482342 220476
rect 491938 220464 491944 220476
rect 491996 220464 492002 220516
rect 493962 220464 493968 220516
rect 494020 220504 494026 220516
rect 508498 220504 508504 220516
rect 494020 220476 508504 220504
rect 494020 220464 494026 220476
rect 508498 220464 508504 220476
rect 508556 220464 508562 220516
rect 522298 220464 522304 220516
rect 522356 220504 522362 220516
rect 540054 220504 540060 220516
rect 522356 220476 540060 220504
rect 522356 220464 522362 220476
rect 540054 220464 540060 220476
rect 540112 220504 540118 220516
rect 622670 220504 622676 220516
rect 540112 220476 622676 220504
rect 540112 220464 540118 220476
rect 622670 220464 622676 220476
rect 622728 220464 622734 220516
rect 218606 220368 218612 220380
rect 161952 220340 218612 220368
rect 218606 220328 218612 220340
rect 218664 220328 218670 220380
rect 229738 220328 229744 220380
rect 229796 220368 229802 220380
rect 276106 220368 276112 220380
rect 229796 220340 276112 220368
rect 229796 220328 229802 220340
rect 276106 220328 276112 220340
rect 276164 220328 276170 220380
rect 280062 220328 280068 220380
rect 280120 220368 280126 220380
rect 313918 220368 313924 220380
rect 280120 220340 313924 220368
rect 280120 220328 280126 220340
rect 313918 220328 313924 220340
rect 313976 220328 313982 220380
rect 323118 220328 323124 220380
rect 323176 220368 323182 220380
rect 348142 220368 348148 220380
rect 323176 220340 348148 220368
rect 323176 220328 323182 220340
rect 348142 220328 348148 220340
rect 348200 220328 348206 220380
rect 352926 220328 352932 220380
rect 352984 220368 352990 220380
rect 371418 220368 371424 220380
rect 352984 220340 371424 220368
rect 352984 220328 352990 220340
rect 371418 220328 371424 220340
rect 371476 220328 371482 220380
rect 481542 220328 481548 220380
rect 481600 220368 481606 220380
rect 492766 220368 492772 220380
rect 481600 220340 492772 220368
rect 481600 220328 481606 220340
rect 492766 220328 492772 220340
rect 492824 220328 492830 220380
rect 496354 220328 496360 220380
rect 496412 220368 496418 220380
rect 510982 220368 510988 220380
rect 496412 220340 510988 220368
rect 496412 220328 496418 220340
rect 510982 220328 510988 220340
rect 511040 220328 511046 220380
rect 517422 220328 517428 220380
rect 517480 220368 517486 220380
rect 539134 220368 539140 220380
rect 517480 220340 539140 220368
rect 517480 220328 517486 220340
rect 539134 220328 539140 220340
rect 539192 220328 539198 220380
rect 541710 220328 541716 220380
rect 541768 220368 541774 220380
rect 554958 220368 554964 220380
rect 541768 220340 554964 220368
rect 541768 220328 541774 220340
rect 554958 220328 554964 220340
rect 555016 220368 555022 220380
rect 555016 220340 558316 220368
rect 555016 220328 555022 220340
rect 66438 220192 66444 220244
rect 66496 220232 66502 220244
rect 142108 220232 142114 220244
rect 66496 220204 142114 220232
rect 66496 220192 66502 220204
rect 142108 220192 142114 220204
rect 142166 220192 142172 220244
rect 142246 220192 142252 220244
rect 142304 220232 142310 220244
rect 205726 220232 205732 220244
rect 142304 220204 205732 220232
rect 142304 220192 142310 220204
rect 205726 220192 205732 220204
rect 205784 220192 205790 220244
rect 211338 220192 211344 220244
rect 211396 220232 211402 220244
rect 263042 220232 263048 220244
rect 211396 220204 263048 220232
rect 211396 220192 211402 220204
rect 263042 220192 263048 220204
rect 263100 220192 263106 220244
rect 263318 220192 263324 220244
rect 263376 220232 263382 220244
rect 301038 220232 301044 220244
rect 263376 220204 301044 220232
rect 263376 220192 263382 220204
rect 301038 220192 301044 220204
rect 301096 220192 301102 220244
rect 311802 220192 311808 220244
rect 311860 220232 311866 220244
rect 327258 220232 327264 220244
rect 311860 220204 327264 220232
rect 311860 220192 311866 220204
rect 327258 220192 327264 220204
rect 327316 220192 327322 220244
rect 332226 220192 332232 220244
rect 332284 220232 332290 220244
rect 357526 220232 357532 220244
rect 332284 220204 357532 220232
rect 332284 220192 332290 220204
rect 357526 220192 357532 220204
rect 357584 220192 357590 220244
rect 360378 220192 360384 220244
rect 360436 220232 360442 220244
rect 377398 220232 377404 220244
rect 360436 220204 377404 220232
rect 360436 220192 360442 220204
rect 377398 220192 377404 220204
rect 377456 220192 377462 220244
rect 390094 220192 390100 220244
rect 390152 220232 390158 220244
rect 401686 220232 401692 220244
rect 390152 220204 401692 220232
rect 390152 220192 390158 220204
rect 401686 220192 401692 220204
rect 401744 220192 401750 220244
rect 432230 220192 432236 220244
rect 432288 220232 432294 220244
rect 434806 220232 434812 220244
rect 432288 220204 434812 220232
rect 432288 220192 432294 220204
rect 434806 220192 434812 220204
rect 434864 220192 434870 220244
rect 459462 220192 459468 220244
rect 459520 220232 459526 220244
rect 465442 220232 465448 220244
rect 459520 220204 465448 220232
rect 459520 220192 459526 220204
rect 465442 220192 465448 220204
rect 465500 220192 465506 220244
rect 469030 220192 469036 220244
rect 469088 220232 469094 220244
rect 474550 220232 474556 220244
rect 469088 220204 474556 220232
rect 469088 220192 469094 220204
rect 474550 220192 474556 220204
rect 474608 220192 474614 220244
rect 478506 220192 478512 220244
rect 478564 220232 478570 220244
rect 489454 220232 489460 220244
rect 478564 220204 489460 220232
rect 478564 220192 478570 220204
rect 489454 220192 489460 220204
rect 489512 220192 489518 220244
rect 492306 220192 492312 220244
rect 492364 220232 492370 220244
rect 507670 220232 507676 220244
rect 492364 220204 507676 220232
rect 492364 220192 492370 220204
rect 507670 220192 507676 220204
rect 507728 220192 507734 220244
rect 521562 220192 521568 220244
rect 521620 220232 521626 220244
rect 544194 220232 544200 220244
rect 521620 220204 544200 220232
rect 521620 220192 521626 220204
rect 544194 220192 544200 220204
rect 544252 220192 544258 220244
rect 552474 220232 552480 220244
rect 549824 220204 552480 220232
rect 63126 220056 63132 220108
rect 63184 220096 63190 220108
rect 146478 220096 146484 220108
rect 63184 220068 146484 220096
rect 63184 220056 63190 220068
rect 146478 220056 146484 220068
rect 146536 220056 146542 220108
rect 147582 220056 147588 220108
rect 147640 220096 147646 220108
rect 204530 220096 204536 220108
rect 147640 220068 204536 220096
rect 147640 220056 147646 220068
rect 204530 220056 204536 220068
rect 204588 220056 204594 220108
rect 204714 220056 204720 220108
rect 204772 220096 204778 220108
rect 214006 220096 214012 220108
rect 204772 220068 214012 220096
rect 204772 220056 204778 220068
rect 214006 220056 214012 220068
rect 214064 220056 214070 220108
rect 217134 220056 217140 220108
rect 217192 220096 217198 220108
rect 265158 220096 265164 220108
rect 217192 220068 265164 220096
rect 217192 220056 217198 220068
rect 265158 220056 265164 220068
rect 265216 220056 265222 220108
rect 280890 220056 280896 220108
rect 280948 220096 280954 220108
rect 317506 220096 317512 220108
rect 280948 220068 317512 220096
rect 280948 220056 280954 220068
rect 317506 220056 317512 220068
rect 317564 220056 317570 220108
rect 318150 220056 318156 220108
rect 318208 220096 318214 220108
rect 343726 220096 343732 220108
rect 318208 220068 343732 220096
rect 318208 220056 318214 220068
rect 343726 220056 343732 220068
rect 343784 220056 343790 220108
rect 345474 220056 345480 220108
rect 345532 220096 345538 220108
rect 367370 220096 367376 220108
rect 345532 220068 367376 220096
rect 345532 220056 345538 220068
rect 367370 220056 367376 220068
rect 367428 220056 367434 220108
rect 367830 220056 367836 220108
rect 367888 220096 367894 220108
rect 382458 220096 382464 220108
rect 367888 220068 382464 220096
rect 367888 220056 367894 220068
rect 382458 220056 382464 220068
rect 382516 220056 382522 220108
rect 382734 220056 382740 220108
rect 382792 220096 382798 220108
rect 394786 220096 394792 220108
rect 382792 220068 394792 220096
rect 382792 220056 382798 220068
rect 394786 220056 394792 220068
rect 394844 220056 394850 220108
rect 397638 220056 397644 220108
rect 397696 220096 397702 220108
rect 405826 220096 405832 220108
rect 397696 220068 405832 220096
rect 397696 220056 397702 220068
rect 405826 220056 405832 220068
rect 405884 220056 405890 220108
rect 421650 220056 421656 220108
rect 421708 220096 421714 220108
rect 426802 220096 426808 220108
rect 421708 220068 426808 220096
rect 421708 220056 421714 220068
rect 426802 220056 426808 220068
rect 426860 220056 426866 220108
rect 427906 220056 427912 220108
rect 427964 220096 427970 220108
rect 428734 220096 428740 220108
rect 427964 220068 428740 220096
rect 427964 220056 427970 220068
rect 428734 220056 428740 220068
rect 428792 220056 428798 220108
rect 472986 220056 472992 220108
rect 473044 220096 473050 220108
rect 482002 220096 482008 220108
rect 473044 220068 482008 220096
rect 473044 220056 473050 220068
rect 482002 220056 482008 220068
rect 482060 220056 482066 220108
rect 488258 220056 488264 220108
rect 488316 220096 488322 220108
rect 502702 220096 502708 220108
rect 488316 220068 502708 220096
rect 488316 220056 488322 220068
rect 502702 220056 502708 220068
rect 502760 220056 502766 220108
rect 507026 220056 507032 220108
rect 507084 220096 507090 220108
rect 522574 220096 522580 220108
rect 507084 220068 522580 220096
rect 507084 220056 507090 220068
rect 522574 220056 522580 220068
rect 522632 220056 522638 220108
rect 527818 220056 527824 220108
rect 527876 220096 527882 220108
rect 527876 220068 543734 220096
rect 527876 220056 527882 220068
rect 543706 220028 543734 220068
rect 549824 220028 549852 220204
rect 552474 220192 552480 220204
rect 552532 220232 552538 220244
rect 558288 220232 558316 220340
rect 559558 220328 559564 220380
rect 559616 220368 559622 220380
rect 567194 220368 567200 220380
rect 559616 220340 567200 220368
rect 559616 220328 559622 220340
rect 567194 220328 567200 220340
rect 567252 220328 567258 220380
rect 567378 220328 567384 220380
rect 567436 220368 567442 220380
rect 572346 220368 572352 220380
rect 567436 220340 572352 220368
rect 567436 220328 567442 220340
rect 572346 220328 572352 220340
rect 572404 220328 572410 220380
rect 572806 220328 572812 220380
rect 572864 220368 572870 220380
rect 582190 220368 582196 220380
rect 572864 220340 582196 220368
rect 572864 220328 572870 220340
rect 582190 220328 582196 220340
rect 582248 220328 582254 220380
rect 582374 220328 582380 220380
rect 582432 220368 582438 220380
rect 591850 220368 591856 220380
rect 582432 220340 591856 220368
rect 582432 220328 582438 220340
rect 591850 220328 591856 220340
rect 591908 220328 591914 220380
rect 591988 220328 591994 220380
rect 592046 220368 592052 220380
rect 628190 220368 628196 220380
rect 592046 220340 628196 220368
rect 592046 220328 592052 220340
rect 628190 220328 628196 220340
rect 628248 220328 628254 220380
rect 562686 220232 562692 220244
rect 552532 220204 553394 220232
rect 558288 220204 562692 220232
rect 552532 220192 552538 220204
rect 553366 220164 553394 220204
rect 562686 220192 562692 220204
rect 562744 220192 562750 220244
rect 563054 220192 563060 220244
rect 563112 220232 563118 220244
rect 620094 220232 620100 220244
rect 563112 220204 620100 220232
rect 563112 220192 563118 220204
rect 620094 220192 620100 220204
rect 620152 220192 620158 220244
rect 620278 220192 620284 220244
rect 620336 220232 620342 220244
rect 628006 220232 628012 220244
rect 620336 220204 628012 220232
rect 620336 220192 620342 220204
rect 628006 220192 628012 220204
rect 628064 220192 628070 220244
rect 553366 220136 558224 220164
rect 558196 220096 558224 220136
rect 625522 220096 625528 220108
rect 558196 220068 625528 220096
rect 625522 220056 625528 220068
rect 625580 220056 625586 220108
rect 647234 220056 647240 220108
rect 647292 220096 647298 220108
rect 652754 220096 652760 220108
rect 647292 220068 652760 220096
rect 647292 220056 647298 220068
rect 652754 220056 652760 220068
rect 652812 220056 652818 220108
rect 543706 220000 549852 220028
rect 553210 219988 553216 220040
rect 553268 220028 553274 220040
rect 553578 220028 553584 220040
rect 553268 220000 553584 220028
rect 553268 219988 553274 220000
rect 553578 219988 553584 220000
rect 553636 219988 553642 220040
rect 553762 219988 553768 220040
rect 553820 220028 553826 220040
rect 557994 220028 558000 220040
rect 553820 220000 558000 220028
rect 553820 219988 553826 220000
rect 557994 219988 558000 220000
rect 558052 219988 558058 220040
rect 111242 219920 111248 219972
rect 111300 219960 111306 219972
rect 173342 219960 173348 219972
rect 111300 219932 173348 219960
rect 111300 219920 111306 219932
rect 173342 219920 173348 219932
rect 173400 219920 173406 219972
rect 173526 219920 173532 219972
rect 173584 219960 173590 219972
rect 173584 219932 195284 219960
rect 173584 219920 173590 219932
rect 124398 219784 124404 219836
rect 124456 219824 124462 219836
rect 193306 219824 193312 219836
rect 124456 219796 193312 219824
rect 124456 219784 124462 219796
rect 193306 219784 193312 219796
rect 193364 219784 193370 219836
rect 195256 219824 195284 219932
rect 195422 219920 195428 219972
rect 195480 219960 195486 219972
rect 244458 219960 244464 219972
rect 195480 219932 244464 219960
rect 195480 219920 195486 219932
rect 244458 219920 244464 219932
rect 244516 219920 244522 219972
rect 256878 219920 256884 219972
rect 256936 219960 256942 219972
rect 295886 219960 295892 219972
rect 256936 219932 295892 219960
rect 256936 219920 256942 219932
rect 295886 219920 295892 219932
rect 295944 219920 295950 219972
rect 296806 219920 296812 219972
rect 296864 219960 296870 219972
rect 310698 219960 310704 219972
rect 296864 219932 310704 219960
rect 296864 219920 296870 219932
rect 310698 219920 310704 219932
rect 310756 219920 310762 219972
rect 540790 219852 540796 219904
rect 540848 219892 540854 219904
rect 548886 219892 548892 219904
rect 540848 219864 548892 219892
rect 540848 219852 540854 219864
rect 548886 219852 548892 219864
rect 548944 219852 548950 219904
rect 550082 219852 550088 219904
rect 550140 219892 550146 219904
rect 625338 219892 625344 219904
rect 550140 219864 625344 219892
rect 550140 219852 550146 219864
rect 625338 219852 625344 219864
rect 625396 219852 625402 219904
rect 204714 219824 204720 219836
rect 195256 219796 204720 219824
rect 204714 219784 204720 219796
rect 204772 219784 204778 219836
rect 249886 219824 249892 219836
rect 204916 219796 249892 219824
rect 131022 219648 131028 219700
rect 131080 219688 131086 219700
rect 190454 219688 190460 219700
rect 131080 219660 190460 219688
rect 131080 219648 131086 219660
rect 190454 219648 190460 219660
rect 190512 219648 190518 219700
rect 190638 219648 190644 219700
rect 190696 219688 190702 219700
rect 195422 219688 195428 219700
rect 190696 219660 195428 219688
rect 190696 219648 190702 219660
rect 195422 219648 195428 219660
rect 195480 219648 195486 219700
rect 197262 219648 197268 219700
rect 197320 219688 197326 219700
rect 204916 219688 204944 219796
rect 249886 219784 249892 219796
rect 249944 219784 249950 219836
rect 531314 219716 531320 219768
rect 531372 219756 531378 219768
rect 532602 219756 532608 219768
rect 531372 219728 532608 219756
rect 531372 219716 531378 219728
rect 532602 219716 532608 219728
rect 532660 219756 532666 219768
rect 621014 219756 621020 219768
rect 532660 219728 621020 219756
rect 532660 219716 532666 219728
rect 621014 219716 621020 219728
rect 621072 219716 621078 219768
rect 197320 219660 204944 219688
rect 197320 219648 197326 219660
rect 207198 219648 207204 219700
rect 207256 219688 207262 219700
rect 257246 219688 257252 219700
rect 207256 219660 257252 219688
rect 207256 219648 207262 219660
rect 257246 219648 257252 219660
rect 257304 219648 257310 219700
rect 520090 219648 520096 219700
rect 520148 219688 520154 219700
rect 520148 219660 524414 219688
rect 520148 219648 520154 219660
rect 464982 219580 464988 219632
rect 465040 219620 465046 219632
rect 472066 219620 472072 219632
rect 465040 219592 472072 219620
rect 465040 219580 465046 219592
rect 472066 219580 472072 219592
rect 472124 219580 472130 219632
rect 524386 219620 524414 219660
rect 618254 219620 618260 219632
rect 524386 219592 618260 219620
rect 618254 219580 618260 219592
rect 618312 219580 618318 219632
rect 620094 219580 620100 219632
rect 620152 219620 620158 219632
rect 626810 219620 626816 219632
rect 620152 219592 626816 219620
rect 620152 219580 620158 219592
rect 626810 219580 626816 219592
rect 626868 219580 626874 219632
rect 137646 219512 137652 219564
rect 137704 219552 137710 219564
rect 140774 219552 140780 219564
rect 137704 219524 140780 219552
rect 137704 219512 137710 219524
rect 140774 219512 140780 219524
rect 140832 219512 140838 219564
rect 140958 219512 140964 219564
rect 141016 219552 141022 219564
rect 141970 219552 141976 219564
rect 141016 219524 141976 219552
rect 141016 219512 141022 219524
rect 141970 219512 141976 219524
rect 142028 219512 142034 219564
rect 142154 219512 142160 219564
rect 142212 219552 142218 219564
rect 203426 219552 203432 219564
rect 142212 219524 203432 219552
rect 142212 219512 142218 219524
rect 203426 219512 203432 219524
rect 203484 219512 203490 219564
rect 204530 219512 204536 219564
rect 204588 219552 204594 219564
rect 211154 219552 211160 219564
rect 204588 219524 211160 219552
rect 204588 219512 204594 219524
rect 211154 219512 211160 219524
rect 211212 219512 211218 219564
rect 432046 219552 432052 219564
rect 431926 219524 432052 219552
rect 105814 219444 105820 219496
rect 105872 219484 105878 219496
rect 279234 219484 279240 219496
rect 105872 219456 107148 219484
rect 105872 219444 105878 219456
rect 63954 219376 63960 219428
rect 64012 219416 64018 219428
rect 64874 219416 64880 219428
rect 64012 219388 64880 219416
rect 64012 219376 64018 219388
rect 64874 219376 64880 219388
rect 64932 219376 64938 219428
rect 72234 219376 72240 219428
rect 72292 219416 72298 219428
rect 73154 219416 73160 219428
rect 72292 219388 73160 219416
rect 72292 219376 72298 219388
rect 73154 219376 73160 219388
rect 73212 219376 73218 219428
rect 80514 219376 80520 219428
rect 80572 219416 80578 219428
rect 90266 219416 90272 219428
rect 80572 219388 90272 219416
rect 80572 219376 80578 219388
rect 90266 219376 90272 219388
rect 90324 219376 90330 219428
rect 90450 219376 90456 219428
rect 90508 219416 90514 219428
rect 90508 219388 103514 219416
rect 90508 219376 90514 219388
rect 103486 219280 103514 219388
rect 106918 219280 106924 219292
rect 103486 219252 106924 219280
rect 106918 219240 106924 219252
rect 106976 219240 106982 219292
rect 107120 219280 107148 219456
rect 224420 219456 224954 219484
rect 117958 219376 117964 219428
rect 118016 219416 118022 219428
rect 123478 219416 123484 219428
rect 118016 219388 123484 219416
rect 118016 219376 118022 219388
rect 123478 219376 123484 219388
rect 123536 219376 123542 219428
rect 126054 219376 126060 219428
rect 126112 219416 126118 219428
rect 126974 219416 126980 219428
rect 126112 219388 126980 219416
rect 126112 219376 126118 219388
rect 126974 219376 126980 219388
rect 127032 219376 127038 219428
rect 130194 219376 130200 219428
rect 130252 219416 130258 219428
rect 134150 219416 134156 219428
rect 130252 219388 134156 219416
rect 130252 219376 130258 219388
rect 134150 219376 134156 219388
rect 134208 219376 134214 219428
rect 134334 219376 134340 219428
rect 134392 219416 134398 219428
rect 135254 219416 135260 219428
rect 134392 219388 135260 219416
rect 134392 219376 134398 219388
rect 135254 219376 135260 219388
rect 135312 219376 135318 219428
rect 135806 219376 135812 219428
rect 135864 219416 135870 219428
rect 139946 219416 139952 219428
rect 135864 219388 139952 219416
rect 135864 219376 135870 219388
rect 139946 219376 139952 219388
rect 140004 219376 140010 219428
rect 140130 219376 140136 219428
rect 140188 219416 140194 219428
rect 145742 219416 145748 219428
rect 140188 219388 145748 219416
rect 140188 219376 140194 219388
rect 145742 219376 145748 219388
rect 145800 219376 145806 219428
rect 146478 219376 146484 219428
rect 146536 219416 146542 219428
rect 197906 219416 197912 219428
rect 146536 219388 197912 219416
rect 146536 219376 146542 219388
rect 197906 219376 197912 219388
rect 197964 219376 197970 219428
rect 199746 219376 199752 219428
rect 199804 219416 199810 219428
rect 203334 219416 203340 219428
rect 199804 219388 203340 219416
rect 199804 219376 199810 219388
rect 203334 219376 203340 219388
rect 203392 219376 203398 219428
rect 208854 219376 208860 219428
rect 208912 219416 208918 219428
rect 209774 219416 209780 219428
rect 208912 219388 209780 219416
rect 208912 219376 208918 219388
rect 209774 219376 209780 219388
rect 209832 219376 209838 219428
rect 148364 219280 148370 219292
rect 107120 219252 148370 219280
rect 148364 219240 148370 219252
rect 148422 219240 148428 219292
rect 149238 219240 149244 219292
rect 149296 219280 149302 219292
rect 150342 219280 150348 219292
rect 149296 219252 150348 219280
rect 149296 219240 149302 219252
rect 150342 219240 150348 219252
rect 150400 219240 150406 219292
rect 152550 219240 152556 219292
rect 152608 219280 152614 219292
rect 153102 219280 153108 219292
rect 152608 219252 153108 219280
rect 152608 219240 152614 219252
rect 153102 219240 153108 219252
rect 153160 219240 153166 219292
rect 153378 219240 153384 219292
rect 153436 219280 153442 219292
rect 162302 219280 162308 219292
rect 153436 219252 162308 219280
rect 153436 219240 153442 219252
rect 162302 219240 162308 219252
rect 162360 219240 162366 219292
rect 162854 219240 162860 219292
rect 162912 219280 162918 219292
rect 163958 219280 163964 219292
rect 162912 219252 163964 219280
rect 162912 219240 162918 219252
rect 163958 219240 163964 219252
rect 164016 219240 164022 219292
rect 164970 219240 164976 219292
rect 165028 219280 165034 219292
rect 165430 219280 165436 219292
rect 165028 219252 165436 219280
rect 165028 219240 165034 219252
rect 165430 219240 165436 219252
rect 165488 219240 165494 219292
rect 165798 219240 165804 219292
rect 165856 219280 165862 219292
rect 166442 219280 166448 219292
rect 165856 219252 166448 219280
rect 165856 219240 165862 219252
rect 166442 219240 166448 219252
rect 166500 219240 166506 219292
rect 168926 219280 168932 219292
rect 166644 219252 168932 219280
rect 85298 219104 85304 219156
rect 85356 219144 85362 219156
rect 117958 219144 117964 219156
rect 85356 219116 117964 219144
rect 85356 219104 85362 219116
rect 117958 219104 117964 219116
rect 118016 219104 118022 219156
rect 123570 219104 123576 219156
rect 123628 219144 123634 219156
rect 128722 219144 128728 219156
rect 123628 219116 128728 219144
rect 123628 219104 123634 219116
rect 128722 219104 128728 219116
rect 128780 219104 128786 219156
rect 131850 219104 131856 219156
rect 131908 219144 131914 219156
rect 132402 219144 132408 219156
rect 131908 219116 132408 219144
rect 131908 219104 131914 219116
rect 132402 219104 132408 219116
rect 132460 219104 132466 219156
rect 132604 219116 134012 219144
rect 70578 218968 70584 219020
rect 70636 219008 70642 219020
rect 132604 219008 132632 219116
rect 70636 218980 132632 219008
rect 70636 218968 70642 218980
rect 132770 218968 132776 219020
rect 132828 219008 132834 219020
rect 133782 219008 133788 219020
rect 132828 218980 133788 219008
rect 132828 218968 132834 218980
rect 133782 218968 133788 218980
rect 133840 218968 133846 219020
rect 133984 219008 134012 219116
rect 134150 219104 134156 219156
rect 134208 219144 134214 219156
rect 134208 219116 136772 219144
rect 134208 219104 134214 219116
rect 135806 219008 135812 219020
rect 133984 218980 135812 219008
rect 135806 218968 135812 218980
rect 135864 218968 135870 219020
rect 135990 218968 135996 219020
rect 136048 219008 136054 219020
rect 136542 219008 136548 219020
rect 136048 218980 136548 219008
rect 136048 218968 136054 218980
rect 136542 218968 136548 218980
rect 136600 218968 136606 219020
rect 136744 219008 136772 219116
rect 136910 219104 136916 219156
rect 136968 219144 136974 219156
rect 146478 219144 146484 219156
rect 136968 219116 146484 219144
rect 136968 219104 136974 219116
rect 146478 219104 146484 219116
rect 146536 219104 146542 219156
rect 146938 219104 146944 219156
rect 146996 219144 147002 219156
rect 152274 219144 152280 219156
rect 146996 219116 152280 219144
rect 146996 219104 147002 219116
rect 152274 219104 152280 219116
rect 152332 219104 152338 219156
rect 166644 219144 166672 219252
rect 168926 219240 168932 219252
rect 168984 219240 168990 219292
rect 169110 219240 169116 219292
rect 169168 219280 169174 219292
rect 169168 219252 190454 219280
rect 169168 219240 169174 219252
rect 152476 219116 166672 219144
rect 152476 219008 152504 219116
rect 167086 219104 167092 219156
rect 167144 219144 167150 219156
rect 185762 219144 185768 219156
rect 167144 219116 185768 219144
rect 167144 219104 167150 219116
rect 185762 219104 185768 219116
rect 185820 219104 185826 219156
rect 190426 219144 190454 219252
rect 193122 219240 193128 219292
rect 193180 219280 193186 219292
rect 195422 219280 195428 219292
rect 193180 219252 195428 219280
rect 193180 219240 193186 219252
rect 195422 219240 195428 219252
rect 195480 219240 195486 219292
rect 196066 219240 196072 219292
rect 196124 219280 196130 219292
rect 199378 219280 199384 219292
rect 196124 219252 199384 219280
rect 196124 219240 196130 219252
rect 199378 219240 199384 219252
rect 199436 219240 199442 219292
rect 224420 219280 224448 219456
rect 200086 219252 224448 219280
rect 224926 219280 224954 219456
rect 270788 219456 279240 219484
rect 225414 219376 225420 219428
rect 225472 219416 225478 219428
rect 226150 219416 226156 219428
rect 225472 219388 226156 219416
rect 225472 219376 225478 219388
rect 226150 219376 226156 219388
rect 226208 219376 226214 219428
rect 228542 219376 228548 219428
rect 228600 219416 228606 219428
rect 232498 219416 232504 219428
rect 228600 219388 232504 219416
rect 228600 219376 228606 219388
rect 232498 219376 232504 219388
rect 232556 219376 232562 219428
rect 233694 219376 233700 219428
rect 233752 219416 233758 219428
rect 234614 219416 234620 219428
rect 233752 219388 234620 219416
rect 233752 219376 233758 219388
rect 234614 219376 234620 219388
rect 234672 219376 234678 219428
rect 234798 219376 234804 219428
rect 234856 219416 234862 219428
rect 270788 219416 270816 219456
rect 279234 219444 279240 219456
rect 279292 219444 279298 219496
rect 405918 219444 405924 219496
rect 405976 219484 405982 219496
rect 412726 219484 412732 219496
rect 405976 219456 412732 219484
rect 405976 219444 405982 219456
rect 412726 219444 412732 219456
rect 412784 219444 412790 219496
rect 421006 219484 421012 219496
rect 418172 219456 421012 219484
rect 234856 219388 270816 219416
rect 234856 219376 234862 219388
rect 285858 219376 285864 219428
rect 285916 219416 285922 219428
rect 301498 219416 301504 219428
rect 285916 219388 301504 219416
rect 285916 219376 285922 219388
rect 301498 219376 301504 219388
rect 301556 219376 301562 219428
rect 325602 219376 325608 219428
rect 325660 219416 325666 219428
rect 326338 219416 326344 219428
rect 325660 219388 326344 219416
rect 325660 219376 325666 219388
rect 326338 219376 326344 219388
rect 326396 219376 326402 219428
rect 343818 219376 343824 219428
rect 343876 219416 343882 219428
rect 347038 219416 347044 219428
rect 343876 219388 347044 219416
rect 343876 219376 343882 219388
rect 347038 219376 347044 219388
rect 347096 219376 347102 219428
rect 352098 219376 352104 219428
rect 352156 219416 352162 219428
rect 366358 219416 366364 219428
rect 352156 219388 366364 219416
rect 352156 219376 352162 219388
rect 366358 219376 366364 219388
rect 366416 219376 366422 219428
rect 374454 219376 374460 219428
rect 374512 219416 374518 219428
rect 375374 219416 375380 219428
rect 374512 219388 375380 219416
rect 374512 219376 374518 219388
rect 375374 219376 375380 219388
rect 375432 219376 375438 219428
rect 380250 219376 380256 219428
rect 380308 219416 380314 219428
rect 384298 219416 384304 219428
rect 380308 219388 384304 219416
rect 380308 219376 380314 219388
rect 384298 219376 384304 219388
rect 384356 219376 384362 219428
rect 399294 219376 399300 219428
rect 399352 219416 399358 219428
rect 400214 219416 400220 219428
rect 399352 219388 400220 219416
rect 399352 219376 399358 219388
rect 400214 219376 400220 219388
rect 400272 219376 400278 219428
rect 403434 219376 403440 219428
rect 403492 219416 403498 219428
rect 404354 219416 404360 219428
rect 403492 219388 404360 219416
rect 403492 219376 403498 219388
rect 404354 219376 404360 219388
rect 404412 219376 404418 219428
rect 415854 219376 415860 219428
rect 415912 219416 415918 219428
rect 416774 219416 416780 219428
rect 415912 219388 416780 219416
rect 415912 219376 415918 219388
rect 416774 219376 416780 219388
rect 416832 219376 416838 219428
rect 417510 219376 417516 219428
rect 417568 219416 417574 219428
rect 418172 219416 418200 219456
rect 421006 219444 421012 219456
rect 421064 219444 421070 219496
rect 431926 219484 431954 219524
rect 432046 219512 432052 219524
rect 432104 219512 432110 219564
rect 515214 219512 515220 219564
rect 515272 219552 515278 219564
rect 515766 219552 515772 219564
rect 515272 219524 515772 219552
rect 515272 219512 515278 219524
rect 515766 219512 515772 219524
rect 515824 219552 515830 219564
rect 515824 219524 520044 219552
rect 515824 219512 515830 219524
rect 429212 219456 431954 219484
rect 520016 219484 520044 219524
rect 667934 219512 667940 219564
rect 667992 219552 667998 219564
rect 669314 219552 669320 219564
rect 667992 219524 669320 219552
rect 667992 219512 667998 219524
rect 669314 219512 669320 219524
rect 669372 219512 669378 219564
rect 617242 219484 617248 219496
rect 520016 219456 560294 219484
rect 417568 219388 418200 219416
rect 417568 219376 417574 219388
rect 428274 219376 428280 219428
rect 428332 219416 428338 219428
rect 429212 219416 429240 219456
rect 428332 219388 429240 219416
rect 428332 219376 428338 219388
rect 488718 219376 488724 219428
rect 488776 219416 488782 219428
rect 489178 219416 489184 219428
rect 488776 219388 489184 219416
rect 488776 219376 488782 219388
rect 489178 219376 489184 219388
rect 489236 219376 489242 219428
rect 518802 219376 518808 219428
rect 518860 219416 518866 219428
rect 519814 219416 519820 219428
rect 518860 219388 519820 219416
rect 518860 219376 518866 219388
rect 519814 219376 519820 219388
rect 519872 219376 519878 219428
rect 560266 219416 560294 219456
rect 569926 219456 617248 219484
rect 567838 219416 567844 219428
rect 560266 219388 567844 219416
rect 567838 219376 567844 219388
rect 567896 219376 567902 219428
rect 568114 219376 568120 219428
rect 568172 219416 568178 219428
rect 569926 219416 569954 219456
rect 617242 219444 617248 219456
rect 617300 219444 617306 219496
rect 568172 219388 569954 219416
rect 568172 219376 568178 219388
rect 504634 219308 504640 219360
rect 504692 219348 504698 219360
rect 505278 219348 505284 219360
rect 504692 219320 505284 219348
rect 504692 219308 504698 219320
rect 505278 219308 505284 219320
rect 505336 219308 505342 219360
rect 516594 219348 516600 219360
rect 511966 219320 516600 219348
rect 226886 219280 226892 219292
rect 224926 219252 226892 219280
rect 195054 219144 195060 219156
rect 190426 219116 195060 219144
rect 195054 219104 195060 219116
rect 195112 219104 195118 219156
rect 195238 219104 195244 219156
rect 195296 219144 195302 219156
rect 200086 219144 200114 219252
rect 226886 219240 226892 219252
rect 226944 219240 226950 219292
rect 229370 219240 229376 219292
rect 229428 219280 229434 219292
rect 235166 219280 235172 219292
rect 229428 219252 235172 219280
rect 229428 219240 229434 219252
rect 235166 219240 235172 219252
rect 235224 219240 235230 219292
rect 237834 219240 237840 219292
rect 237892 219280 237898 219292
rect 239398 219280 239404 219292
rect 237892 219252 239404 219280
rect 237892 219240 237898 219252
rect 239398 219240 239404 219252
rect 239456 219240 239462 219292
rect 246114 219240 246120 219292
rect 246172 219280 246178 219292
rect 286042 219280 286048 219292
rect 246172 219252 286048 219280
rect 246172 219240 246178 219252
rect 286042 219240 286048 219252
rect 286100 219240 286106 219292
rect 327258 219240 327264 219292
rect 327316 219280 327322 219292
rect 327316 219252 345014 219280
rect 327316 219240 327322 219252
rect 195296 219116 200114 219144
rect 200408 219116 201724 219144
rect 195296 219104 195302 219116
rect 166736 219048 166948 219076
rect 136744 218980 152504 219008
rect 152734 218968 152740 219020
rect 152792 219008 152798 219020
rect 166736 219008 166764 219048
rect 152792 218980 166764 219008
rect 166920 219008 166948 219048
rect 200408 219008 200436 219116
rect 166920 218980 200436 219008
rect 152792 218968 152798 218980
rect 200574 218968 200580 219020
rect 200632 219008 200638 219020
rect 201494 219008 201500 219020
rect 200632 218980 201500 219008
rect 200632 218968 200638 218980
rect 201494 218968 201500 218980
rect 201552 218968 201558 219020
rect 201696 219008 201724 219116
rect 203334 219104 203340 219156
rect 203392 219144 203398 219156
rect 246298 219144 246304 219156
rect 203392 219116 246304 219144
rect 203392 219104 203398 219116
rect 246298 219104 246304 219116
rect 246356 219104 246362 219156
rect 258534 219104 258540 219156
rect 258592 219144 258598 219156
rect 259270 219144 259276 219156
rect 258592 219116 259276 219144
rect 258592 219104 258598 219116
rect 259270 219104 259276 219116
rect 259328 219104 259334 219156
rect 259454 219104 259460 219156
rect 259512 219144 259518 219156
rect 291838 219144 291844 219156
rect 259512 219116 291844 219144
rect 259512 219104 259518 219116
rect 291838 219104 291844 219116
rect 291896 219104 291902 219156
rect 294138 219104 294144 219156
rect 294196 219144 294202 219156
rect 311802 219144 311808 219156
rect 294196 219116 311808 219144
rect 294196 219104 294202 219116
rect 311802 219104 311808 219116
rect 311860 219104 311866 219156
rect 315666 219104 315672 219156
rect 315724 219144 315730 219156
rect 317966 219144 317972 219156
rect 315724 219116 317972 219144
rect 315724 219104 315730 219116
rect 317966 219104 317972 219116
rect 318024 219104 318030 219156
rect 320634 219104 320640 219156
rect 320692 219144 320698 219156
rect 340138 219144 340144 219156
rect 320692 219116 340144 219144
rect 320692 219104 320698 219116
rect 340138 219104 340144 219116
rect 340196 219104 340202 219156
rect 344986 219144 345014 219252
rect 383562 219240 383568 219292
rect 383620 219280 383626 219292
rect 387058 219280 387064 219292
rect 383620 219252 387064 219280
rect 383620 219240 383626 219252
rect 387058 219240 387064 219252
rect 387116 219240 387122 219292
rect 419166 219240 419172 219292
rect 419224 219280 419230 219292
rect 422662 219280 422668 219292
rect 419224 219252 422668 219280
rect 419224 219240 419230 219252
rect 422662 219240 422668 219252
rect 422720 219240 422726 219292
rect 450722 219240 450728 219292
rect 450780 219280 450786 219292
rect 453850 219280 453856 219292
rect 450780 219252 453856 219280
rect 450780 219240 450786 219252
rect 453850 219240 453856 219252
rect 453908 219240 453914 219292
rect 479702 219240 479708 219292
rect 479760 219280 479766 219292
rect 480346 219280 480352 219292
rect 479760 219252 480352 219280
rect 479760 219240 479766 219252
rect 480346 219240 480352 219252
rect 480404 219240 480410 219292
rect 507118 219172 507124 219224
rect 507176 219212 507182 219224
rect 511966 219212 511994 219320
rect 516594 219308 516600 219320
rect 516652 219308 516658 219360
rect 534994 219308 535000 219360
rect 535052 219348 535058 219360
rect 543826 219348 543832 219360
rect 535052 219320 543832 219348
rect 535052 219308 535058 219320
rect 543826 219308 543832 219320
rect 543884 219308 543890 219360
rect 544010 219308 544016 219360
rect 544068 219348 544074 219360
rect 544068 219320 550634 219348
rect 544068 219308 544074 219320
rect 550606 219280 550634 219320
rect 553210 219280 553216 219292
rect 550606 219252 553216 219280
rect 553210 219240 553216 219252
rect 553268 219240 553274 219292
rect 568022 219280 568028 219292
rect 553366 219252 568028 219280
rect 507176 219184 511994 219212
rect 507176 219172 507182 219184
rect 345658 219144 345664 219156
rect 344986 219116 345664 219144
rect 345658 219104 345664 219116
rect 345716 219104 345722 219156
rect 352558 219144 352564 219156
rect 348758 219116 352564 219144
rect 204898 219008 204904 219020
rect 201696 218980 204904 219008
rect 204898 218968 204904 218980
rect 204956 218968 204962 219020
rect 206370 218968 206376 219020
rect 206428 219008 206434 219020
rect 255866 219008 255872 219020
rect 206428 218980 255872 219008
rect 206428 218968 206434 218980
rect 255866 218968 255872 218980
rect 255924 218968 255930 219020
rect 259270 218968 259276 219020
rect 259328 219008 259334 219020
rect 293586 219008 293592 219020
rect 259328 218980 293592 219008
rect 259328 218968 259334 218980
rect 293586 218968 293592 218980
rect 293644 218968 293650 219020
rect 301498 218968 301504 219020
rect 301556 219008 301562 219020
rect 306742 219008 306748 219020
rect 301556 218980 306748 219008
rect 301556 218968 301562 218980
rect 306742 218968 306748 218980
rect 306800 218968 306806 219020
rect 329558 219008 329564 219020
rect 312740 218980 329564 219008
rect 62298 218832 62304 218884
rect 62356 218872 62362 218884
rect 76558 218872 76564 218884
rect 62356 218844 76564 218872
rect 62356 218832 62362 218844
rect 76558 218832 76564 218844
rect 76616 218832 76622 218884
rect 83826 218832 83832 218884
rect 83884 218872 83890 218884
rect 148226 218872 148232 218884
rect 83884 218844 148232 218872
rect 83884 218832 83890 218844
rect 148226 218832 148232 218844
rect 148284 218832 148290 218884
rect 148410 218832 148416 218884
rect 148468 218872 148474 218884
rect 148962 218872 148968 218884
rect 148468 218844 148968 218872
rect 148468 218832 148474 218844
rect 148962 218832 148968 218844
rect 149020 218832 149026 218884
rect 149882 218832 149888 218884
rect 149940 218872 149946 218884
rect 152090 218872 152096 218884
rect 149940 218844 152096 218872
rect 149940 218832 149946 218844
rect 152090 218832 152096 218844
rect 152148 218832 152154 218884
rect 152274 218832 152280 218884
rect 152332 218872 152338 218884
rect 166074 218872 166080 218884
rect 152332 218844 166080 218872
rect 152332 218832 152338 218844
rect 166074 218832 166080 218844
rect 166132 218832 166138 218884
rect 166948 218832 166954 218884
rect 167006 218872 167012 218884
rect 215938 218872 215944 218884
rect 167006 218844 215944 218872
rect 167006 218832 167012 218844
rect 215938 218832 215944 218844
rect 215996 218832 216002 218884
rect 217962 218832 217968 218884
rect 218020 218872 218026 218884
rect 220078 218872 220084 218884
rect 218020 218844 220084 218872
rect 218020 218832 218026 218844
rect 220078 218832 220084 218844
rect 220136 218832 220142 218884
rect 220280 218844 229784 218872
rect 77202 218696 77208 218748
rect 77260 218736 77266 218748
rect 142246 218736 142252 218748
rect 77260 218708 142252 218736
rect 77260 218696 77266 218708
rect 142246 218696 142252 218708
rect 142304 218696 142310 218748
rect 145558 218736 145564 218748
rect 142448 218708 145564 218736
rect 59814 218560 59820 218612
rect 59872 218600 59878 218612
rect 69566 218600 69572 218612
rect 59872 218572 69572 218600
rect 59872 218560 59878 218572
rect 69566 218560 69572 218572
rect 69624 218560 69630 218612
rect 92934 218560 92940 218612
rect 92992 218600 92998 218612
rect 93762 218600 93768 218612
rect 92992 218572 93768 218600
rect 92992 218560 92998 218572
rect 93762 218560 93768 218572
rect 93820 218560 93826 218612
rect 142448 218600 142476 218708
rect 145558 218696 145564 218708
rect 145616 218696 145622 218748
rect 145742 218696 145748 218748
rect 145800 218736 145806 218748
rect 146938 218736 146944 218748
rect 145800 218708 146944 218736
rect 145800 218696 145806 218708
rect 146938 218696 146944 218708
rect 146996 218696 147002 218748
rect 152734 218736 152740 218748
rect 147140 218708 152740 218736
rect 103486 218572 142476 218600
rect 93762 218424 93768 218476
rect 93820 218464 93826 218476
rect 103486 218464 103514 218572
rect 142614 218560 142620 218612
rect 142672 218600 142678 218612
rect 143166 218600 143172 218612
rect 142672 218572 143172 218600
rect 142672 218560 142678 218572
rect 143166 218560 143172 218572
rect 143224 218560 143230 218612
rect 145098 218560 145104 218612
rect 145156 218600 145162 218612
rect 146202 218600 146208 218612
rect 145156 218572 146208 218600
rect 145156 218560 145162 218572
rect 146202 218560 146208 218572
rect 146260 218560 146266 218612
rect 146754 218560 146760 218612
rect 146812 218600 146818 218612
rect 147140 218600 147168 218708
rect 152734 218696 152740 218708
rect 152792 218696 152798 218748
rect 152918 218696 152924 218748
rect 152976 218736 152982 218748
rect 156322 218736 156328 218748
rect 152976 218708 156328 218736
rect 152976 218696 152982 218708
rect 156322 218696 156328 218708
rect 156380 218696 156386 218748
rect 156690 218696 156696 218748
rect 156748 218736 156754 218748
rect 156748 218708 162164 218736
rect 156748 218696 156754 218708
rect 157978 218600 157984 218612
rect 146812 218572 147168 218600
rect 147646 218572 157984 218600
rect 146812 218560 146818 218572
rect 93820 218436 103514 218464
rect 93820 218424 93826 218436
rect 107010 218424 107016 218476
rect 107068 218464 107074 218476
rect 147646 218464 147674 218572
rect 157978 218560 157984 218572
rect 158036 218560 158042 218612
rect 159174 218560 159180 218612
rect 159232 218600 159238 218612
rect 160002 218600 160008 218612
rect 159232 218572 160008 218600
rect 159232 218560 159238 218572
rect 160002 218560 160008 218572
rect 160060 218560 160066 218612
rect 160830 218560 160836 218612
rect 160888 218600 160894 218612
rect 161382 218600 161388 218612
rect 160888 218572 161388 218600
rect 160888 218560 160894 218572
rect 161382 218560 161388 218572
rect 161440 218560 161446 218612
rect 162136 218600 162164 218708
rect 162302 218696 162308 218748
rect 162360 218736 162366 218748
rect 213178 218736 213184 218748
rect 162360 218708 213184 218736
rect 162360 218696 162366 218708
rect 213178 218696 213184 218708
rect 213236 218696 213242 218748
rect 213546 218696 213552 218748
rect 213604 218736 213610 218748
rect 217318 218736 217324 218748
rect 213604 218708 217324 218736
rect 213604 218696 213610 218708
rect 217318 218696 217324 218708
rect 217376 218696 217382 218748
rect 218790 218696 218796 218748
rect 218848 218736 218854 218748
rect 219342 218736 219348 218748
rect 218848 218708 219348 218736
rect 218848 218696 218854 218708
rect 219342 218696 219348 218708
rect 219400 218696 219406 218748
rect 219618 218696 219624 218748
rect 219676 218736 219682 218748
rect 220280 218736 220308 218844
rect 219676 218708 220308 218736
rect 219676 218696 219682 218708
rect 220906 218696 220912 218748
rect 220964 218736 220970 218748
rect 228542 218736 228548 218748
rect 220964 218708 228548 218736
rect 220964 218696 220970 218708
rect 228542 218696 228548 218708
rect 228600 218696 228606 218748
rect 229756 218736 229784 218844
rect 229922 218832 229928 218884
rect 229980 218872 229986 218884
rect 229980 218844 264330 218872
rect 229980 218832 229986 218844
rect 264146 218736 264152 218748
rect 229756 218708 264152 218736
rect 264146 218696 264152 218708
rect 264204 218696 264210 218748
rect 167270 218600 167276 218612
rect 162136 218572 167276 218600
rect 167270 218560 167276 218572
rect 167328 218560 167334 218612
rect 169938 218560 169944 218612
rect 169996 218600 170002 218612
rect 177574 218600 177580 218612
rect 169996 218572 177580 218600
rect 169996 218560 170002 218572
rect 177574 218560 177580 218572
rect 177632 218560 177638 218612
rect 185578 218560 185584 218612
rect 185636 218600 185642 218612
rect 195238 218600 195244 218612
rect 185636 218572 195244 218600
rect 185636 218560 185642 218572
rect 195238 218560 195244 218572
rect 195296 218560 195302 218612
rect 195422 218560 195428 218612
rect 195480 218600 195486 218612
rect 243446 218600 243452 218612
rect 195480 218572 243452 218600
rect 195480 218560 195486 218572
rect 243446 218560 243452 218572
rect 243504 218560 243510 218612
rect 252738 218560 252744 218612
rect 252796 218600 252802 218612
rect 259454 218600 259460 218612
rect 252796 218572 259460 218600
rect 252796 218560 252802 218572
rect 259454 218560 259460 218572
rect 259512 218560 259518 218612
rect 264302 218600 264330 218844
rect 274266 218832 274272 218884
rect 274324 218872 274330 218884
rect 280706 218872 280712 218884
rect 274324 218844 280712 218872
rect 274324 218832 274330 218844
rect 280706 218832 280712 218844
rect 280764 218832 280770 218884
rect 281074 218832 281080 218884
rect 281132 218872 281138 218884
rect 312538 218872 312544 218884
rect 281132 218844 312544 218872
rect 281132 218832 281138 218844
rect 312538 218832 312544 218844
rect 312596 218832 312602 218884
rect 265986 218696 265992 218748
rect 266044 218736 266050 218748
rect 266044 218708 299796 218736
rect 266044 218696 266050 218708
rect 267826 218600 267832 218612
rect 264302 218572 267832 218600
rect 267826 218560 267832 218572
rect 267884 218560 267890 218612
rect 272610 218560 272616 218612
rect 272668 218600 272674 218612
rect 296806 218600 296812 218612
rect 272668 218572 296812 218600
rect 272668 218560 272674 218572
rect 296806 218560 296812 218572
rect 296864 218560 296870 218612
rect 299768 218600 299796 218708
rect 300762 218696 300768 218748
rect 300820 218736 300826 218748
rect 312740 218736 312768 218980
rect 329558 218968 329564 218980
rect 329616 218968 329622 219020
rect 333698 218968 333704 219020
rect 333756 219008 333762 219020
rect 348758 219008 348786 219116
rect 352558 219104 352564 219116
rect 352616 219104 352622 219156
rect 354398 219104 354404 219156
rect 354456 219144 354462 219156
rect 355502 219144 355508 219156
rect 354456 219116 355508 219144
rect 354456 219104 354462 219116
rect 355502 219104 355508 219116
rect 355560 219104 355566 219156
rect 358722 219104 358728 219156
rect 358780 219144 358786 219156
rect 364978 219144 364984 219156
rect 358780 219116 364984 219144
rect 358780 219104 358786 219116
rect 364978 219104 364984 219116
rect 365036 219104 365042 219156
rect 483566 219104 483572 219156
rect 483624 219144 483630 219156
rect 490282 219144 490288 219156
rect 483624 219116 490288 219144
rect 483624 219104 483630 219116
rect 490282 219104 490288 219116
rect 490340 219104 490346 219156
rect 502978 219104 502984 219156
rect 503036 219144 503042 219156
rect 503530 219144 503536 219156
rect 503036 219116 503536 219144
rect 503036 219104 503042 219116
rect 503530 219104 503536 219116
rect 503588 219104 503594 219156
rect 524414 219104 524420 219156
rect 524472 219144 524478 219156
rect 533890 219144 533896 219156
rect 524472 219116 533896 219144
rect 524472 219104 524478 219116
rect 533890 219104 533896 219116
rect 533948 219104 533954 219156
rect 538858 219104 538864 219156
rect 538916 219144 538922 219156
rect 544010 219144 544016 219156
rect 538916 219116 543320 219144
rect 538916 219104 538922 219116
rect 543292 219076 543320 219116
rect 543476 219116 544016 219144
rect 543476 219076 543504 219116
rect 544010 219104 544016 219116
rect 544068 219104 544074 219156
rect 553366 219144 553394 219252
rect 568022 219240 568028 219252
rect 568080 219240 568086 219292
rect 572162 219280 572168 219292
rect 568178 219252 572168 219280
rect 545040 219116 553394 219144
rect 543292 219048 543504 219076
rect 333756 218980 348786 219008
rect 333756 218968 333762 218980
rect 351362 218968 351368 219020
rect 351420 219008 351426 219020
rect 355226 219008 355232 219020
rect 351420 218980 355232 219008
rect 351420 218968 351426 218980
rect 355226 218968 355232 218980
rect 355284 218968 355290 219020
rect 355410 218968 355416 219020
rect 355468 219008 355474 219020
rect 369118 219008 369124 219020
rect 355468 218980 369124 219008
rect 355468 218968 355474 218980
rect 369118 218968 369124 218980
rect 369176 218968 369182 219020
rect 373626 218968 373632 219020
rect 373684 219008 373690 219020
rect 380066 219008 380072 219020
rect 373684 218980 380072 219008
rect 373684 218968 373690 218980
rect 380066 218968 380072 218980
rect 380124 218968 380130 219020
rect 384390 218968 384396 219020
rect 384448 219008 384454 219020
rect 393958 219008 393964 219020
rect 384448 218980 393964 219008
rect 384448 218968 384454 218980
rect 393958 218968 393964 218980
rect 394016 218968 394022 219020
rect 401778 218968 401784 219020
rect 401836 219008 401842 219020
rect 407758 219008 407764 219020
rect 401836 218980 407764 219008
rect 401836 218968 401842 218980
rect 407758 218968 407764 218980
rect 407816 218968 407822 219020
rect 502518 218968 502524 219020
rect 502576 219008 502582 219020
rect 507302 219008 507308 219020
rect 502576 218980 507308 219008
rect 502576 218968 502582 218980
rect 507302 218968 507308 218980
rect 507360 218968 507366 219020
rect 515030 218968 515036 219020
rect 515088 219008 515094 219020
rect 542538 219008 542544 219020
rect 515088 218980 542544 219008
rect 515088 218968 515094 218980
rect 542538 218968 542544 218980
rect 542596 218968 542602 219020
rect 543826 218968 543832 219020
rect 543884 219008 543890 219020
rect 545040 219008 545068 219116
rect 553486 219104 553492 219156
rect 553544 219144 553550 219156
rect 558546 219144 558552 219156
rect 553544 219116 558552 219144
rect 553544 219104 553550 219116
rect 558546 219104 558552 219116
rect 558604 219104 558610 219156
rect 558730 219104 558736 219156
rect 558788 219144 558794 219156
rect 563008 219144 563014 219156
rect 558788 219116 563014 219144
rect 558788 219104 558794 219116
rect 563008 219104 563014 219116
rect 563066 219104 563072 219156
rect 568178 219144 568206 219252
rect 572162 219240 572168 219252
rect 572220 219240 572226 219292
rect 572346 219240 572352 219292
rect 572404 219280 572410 219292
rect 573726 219280 573732 219292
rect 572404 219252 573732 219280
rect 572404 219240 572410 219252
rect 573726 219240 573732 219252
rect 573784 219240 573790 219292
rect 574094 219240 574100 219292
rect 574152 219280 574158 219292
rect 577866 219280 577872 219292
rect 574152 219252 577872 219280
rect 574152 219240 574158 219252
rect 577866 219240 577872 219252
rect 577924 219240 577930 219292
rect 563164 219116 568206 219144
rect 563164 219020 563192 219116
rect 568390 219104 568396 219156
rect 568448 219144 568454 219156
rect 572346 219144 572352 219156
rect 568448 219116 572352 219144
rect 568448 219104 568454 219116
rect 572346 219104 572352 219116
rect 572404 219104 572410 219156
rect 576026 219144 576032 219156
rect 572548 219116 576032 219144
rect 562870 219008 562876 219020
rect 543884 218980 545068 219008
rect 548628 218980 562876 219008
rect 543884 218968 543890 218980
rect 314010 218832 314016 218884
rect 314068 218872 314074 218884
rect 329098 218872 329104 218884
rect 314068 218844 329104 218872
rect 314068 218832 314074 218844
rect 329098 218832 329104 218844
rect 329156 218832 329162 218884
rect 337194 218832 337200 218884
rect 337252 218872 337258 218884
rect 357710 218872 357716 218884
rect 337252 218844 357716 218872
rect 337252 218832 337258 218844
rect 357710 218832 357716 218844
rect 357768 218832 357774 218884
rect 366726 218832 366732 218884
rect 366784 218872 366790 218884
rect 378778 218872 378784 218884
rect 366784 218844 378784 218872
rect 366784 218832 366790 218844
rect 378778 218832 378784 218844
rect 378836 218832 378842 218884
rect 386046 218832 386052 218884
rect 386104 218872 386110 218884
rect 396626 218872 396632 218884
rect 386104 218844 396632 218872
rect 386104 218832 386110 218844
rect 396626 218832 396632 218844
rect 396684 218832 396690 218884
rect 402606 218832 402612 218884
rect 402664 218872 402670 218884
rect 409046 218872 409052 218884
rect 402664 218844 409052 218872
rect 402664 218832 402670 218844
rect 409046 218832 409052 218844
rect 409104 218832 409110 218884
rect 411714 218832 411720 218884
rect 411772 218872 411778 218884
rect 412450 218872 412456 218884
rect 411772 218844 412456 218872
rect 411772 218832 411778 218844
rect 412450 218832 412456 218844
rect 412508 218832 412514 218884
rect 510154 218832 510160 218884
rect 510212 218872 510218 218884
rect 514754 218872 514760 218884
rect 510212 218844 514760 218872
rect 510212 218832 510218 218844
rect 514754 218832 514760 218844
rect 514812 218832 514818 218884
rect 524138 218832 524144 218884
rect 524196 218872 524202 218884
rect 524598 218872 524604 218884
rect 524196 218844 524604 218872
rect 524196 218832 524202 218844
rect 524598 218832 524604 218844
rect 524656 218832 524662 218884
rect 525058 218832 525064 218884
rect 525116 218872 525122 218884
rect 529566 218872 529572 218884
rect 525116 218844 529572 218872
rect 525116 218832 525122 218844
rect 529566 218832 529572 218844
rect 529624 218832 529630 218884
rect 534258 218832 534264 218884
rect 534316 218872 534322 218884
rect 545298 218872 545304 218884
rect 534316 218844 545304 218872
rect 534316 218832 534322 218844
rect 545298 218832 545304 218844
rect 545356 218832 545362 218884
rect 547414 218832 547420 218884
rect 547472 218872 547478 218884
rect 548242 218872 548248 218884
rect 547472 218844 548248 218872
rect 547472 218832 547478 218844
rect 548242 218832 548248 218844
rect 548300 218832 548306 218884
rect 548628 218872 548656 218980
rect 562870 218968 562876 218980
rect 562928 218968 562934 219020
rect 563146 218968 563152 219020
rect 563204 218968 563210 219020
rect 563330 218968 563336 219020
rect 563388 219008 563394 219020
rect 566918 219008 566924 219020
rect 563388 218980 566924 219008
rect 563388 218968 563394 218980
rect 566918 218968 566924 218980
rect 566976 218968 566982 219020
rect 567194 218968 567200 219020
rect 567252 219008 567258 219020
rect 570966 219008 570972 219020
rect 567252 218980 570972 219008
rect 567252 218968 567258 218980
rect 570966 218968 570972 218980
rect 571024 218968 571030 219020
rect 571150 218968 571156 219020
rect 571208 219008 571214 219020
rect 572548 219008 572576 219116
rect 576026 219104 576032 219116
rect 576084 219104 576090 219156
rect 592126 219104 592132 219156
rect 592184 219144 592190 219156
rect 599210 219144 599216 219156
rect 592184 219116 599216 219144
rect 592184 219104 592190 219116
rect 599210 219104 599216 219116
rect 599268 219104 599274 219156
rect 576210 219008 576216 219020
rect 571208 218980 572576 219008
rect 572640 218980 576216 219008
rect 571208 218968 571214 218980
rect 548444 218844 548656 218872
rect 337010 218736 337016 218748
rect 300820 218708 312768 218736
rect 316006 218708 337016 218736
rect 300820 218696 300826 218708
rect 302878 218600 302884 218612
rect 299768 218572 302884 218600
rect 302878 218560 302884 218572
rect 302936 218560 302942 218612
rect 307386 218560 307392 218612
rect 307444 218600 307450 218612
rect 316006 218600 316034 218708
rect 337010 218696 337016 218708
rect 337068 218696 337074 218748
rect 340506 218696 340512 218748
rect 340564 218736 340570 218748
rect 360838 218736 360844 218748
rect 340564 218708 360844 218736
rect 340564 218696 340570 218708
rect 360838 218696 360844 218708
rect 360896 218696 360902 218748
rect 379146 218696 379152 218748
rect 379204 218736 379210 218748
rect 392118 218736 392124 218748
rect 379204 218708 392124 218736
rect 379204 218696 379210 218708
rect 392118 218696 392124 218708
rect 392176 218696 392182 218748
rect 395798 218696 395804 218748
rect 395856 218736 395862 218748
rect 404538 218736 404544 218748
rect 395856 218708 404544 218736
rect 395856 218696 395862 218708
rect 404538 218696 404544 218708
rect 404596 218696 404602 218748
rect 412542 218696 412548 218748
rect 412600 218736 412606 218748
rect 417142 218736 417148 218748
rect 412600 218708 417148 218736
rect 412600 218696 412606 218708
rect 417142 218696 417148 218708
rect 417200 218696 417206 218748
rect 429930 218696 429936 218748
rect 429988 218736 429994 218748
rect 432690 218736 432696 218748
rect 429988 218708 432696 218736
rect 429988 218696 429994 218708
rect 432690 218696 432696 218708
rect 432748 218696 432754 218748
rect 460198 218696 460204 218748
rect 460256 218736 460262 218748
rect 461302 218736 461308 218748
rect 460256 218708 461308 218736
rect 460256 218696 460262 218708
rect 461302 218696 461308 218708
rect 461360 218696 461366 218748
rect 482922 218696 482928 218748
rect 482980 218736 482986 218748
rect 485314 218736 485320 218748
rect 482980 218708 485320 218736
rect 482980 218696 482986 218708
rect 485314 218696 485320 218708
rect 485372 218696 485378 218748
rect 519722 218696 519728 218748
rect 519780 218736 519786 218748
rect 530302 218736 530308 218748
rect 519780 218708 530308 218736
rect 519780 218696 519786 218708
rect 530302 218696 530308 218708
rect 530360 218696 530366 218748
rect 534074 218696 534080 218748
rect 534132 218736 534138 218748
rect 534626 218736 534632 218748
rect 534132 218708 534632 218736
rect 534132 218696 534138 218708
rect 534626 218696 534632 218708
rect 534684 218696 534690 218748
rect 537478 218696 537484 218748
rect 537536 218736 537542 218748
rect 548444 218736 548472 218844
rect 548886 218832 548892 218884
rect 548944 218872 548950 218884
rect 553578 218872 553584 218884
rect 548944 218844 553584 218872
rect 548944 218832 548950 218844
rect 553578 218832 553584 218844
rect 553636 218832 553642 218884
rect 567194 218872 567200 218884
rect 557092 218844 567200 218872
rect 557092 218736 557120 218844
rect 567194 218832 567200 218844
rect 567252 218832 567258 218884
rect 572640 218872 572668 218980
rect 576210 218968 576216 218980
rect 576268 218968 576274 219020
rect 567488 218844 572668 218872
rect 537536 218708 548472 218736
rect 548536 218708 557120 218736
rect 537536 218696 537542 218708
rect 518802 218668 518808 218680
rect 514726 218640 518808 218668
rect 307444 218572 316034 218600
rect 307444 218560 307450 218572
rect 469858 218560 469864 218612
rect 469916 218600 469922 218612
rect 471238 218600 471244 218612
rect 469916 218572 471244 218600
rect 469916 218560 469922 218572
rect 471238 218560 471244 218572
rect 471296 218560 471302 218612
rect 475562 218560 475568 218612
rect 475620 218600 475626 218612
rect 482830 218600 482836 218612
rect 475620 218572 482836 218600
rect 475620 218560 475626 218572
rect 482830 218560 482836 218572
rect 482888 218560 482894 218612
rect 514726 218600 514754 218640
rect 518802 218628 518808 218640
rect 518860 218628 518866 218680
rect 509896 218572 514754 218600
rect 107068 218436 147674 218464
rect 107068 218424 107074 218436
rect 148226 218424 148232 218476
rect 148284 218464 148290 218476
rect 149882 218464 149888 218476
rect 148284 218436 149888 218464
rect 148284 218424 148290 218436
rect 149882 218424 149888 218436
rect 149940 218424 149946 218476
rect 150066 218424 150072 218476
rect 150124 218464 150130 218476
rect 157242 218464 157248 218476
rect 150124 218436 157248 218464
rect 150124 218424 150130 218436
rect 157242 218424 157248 218436
rect 157300 218424 157306 218476
rect 157702 218424 157708 218476
rect 157760 218464 157766 218476
rect 160646 218464 160652 218476
rect 157760 218436 160652 218464
rect 157760 218424 157766 218436
rect 160646 218424 160652 218436
rect 160704 218424 160710 218476
rect 161658 218424 161664 218476
rect 161716 218464 161722 218476
rect 162670 218464 162676 218476
rect 161716 218436 162676 218464
rect 161716 218424 161722 218436
rect 162670 218424 162676 218436
rect 162728 218424 162734 218476
rect 163314 218424 163320 218476
rect 163372 218464 163378 218476
rect 166258 218464 166264 218476
rect 163372 218436 166264 218464
rect 163372 218424 163378 218436
rect 166258 218424 166264 218436
rect 166316 218424 166322 218476
rect 166994 218424 167000 218476
rect 167052 218464 167058 218476
rect 213546 218464 213552 218476
rect 167052 218436 213552 218464
rect 167052 218424 167058 218436
rect 213546 218424 213552 218436
rect 213604 218424 213610 218476
rect 216306 218424 216312 218476
rect 216364 218464 216370 218476
rect 220906 218464 220912 218476
rect 216364 218436 220912 218464
rect 216364 218424 216370 218436
rect 220906 218424 220912 218436
rect 220964 218424 220970 218476
rect 221090 218424 221096 218476
rect 221148 218464 221154 218476
rect 224218 218464 224224 218476
rect 221148 218436 224224 218464
rect 221148 218424 221154 218436
rect 224218 218424 224224 218436
rect 224276 218424 224282 218476
rect 224586 218424 224592 218476
rect 224644 218464 224650 218476
rect 225690 218464 225696 218476
rect 224644 218436 225696 218464
rect 224644 218424 224650 218436
rect 225690 218424 225696 218436
rect 225748 218424 225754 218476
rect 226242 218424 226248 218476
rect 226300 218464 226306 218476
rect 229922 218464 229928 218476
rect 226300 218436 229928 218464
rect 226300 218424 226306 218436
rect 229922 218424 229928 218436
rect 229980 218424 229986 218476
rect 239490 218424 239496 218476
rect 239548 218464 239554 218476
rect 272426 218464 272432 218476
rect 239548 218436 272432 218464
rect 239548 218424 239554 218436
rect 272426 218424 272432 218436
rect 272484 218424 272490 218476
rect 279234 218424 279240 218476
rect 279292 218464 279298 218476
rect 281074 218464 281080 218476
rect 279292 218436 281080 218464
rect 279292 218424 279298 218436
rect 281074 218424 281080 218436
rect 281132 218424 281138 218476
rect 291654 218424 291660 218476
rect 291712 218464 291718 218476
rect 324590 218464 324596 218476
rect 291712 218436 324596 218464
rect 291712 218424 291718 218436
rect 324590 218424 324596 218436
rect 324648 218424 324654 218476
rect 501046 218424 501052 218476
rect 501104 218464 501110 218476
rect 509896 218464 509924 218572
rect 529198 218560 529204 218612
rect 529256 218600 529262 218612
rect 548536 218600 548564 218708
rect 557258 218696 557264 218748
rect 557316 218736 557322 218748
rect 562870 218736 562876 218748
rect 557316 218708 562876 218736
rect 557316 218696 557322 218708
rect 562870 218696 562876 218708
rect 562928 218696 562934 218748
rect 563330 218696 563336 218748
rect 563388 218736 563394 218748
rect 567488 218736 567516 218844
rect 573082 218832 573088 218884
rect 573140 218872 573146 218884
rect 575428 218872 575434 218884
rect 573140 218844 575434 218872
rect 573140 218832 573146 218844
rect 575428 218832 575434 218844
rect 575486 218832 575492 218884
rect 575566 218832 575572 218884
rect 575624 218872 575630 218884
rect 575624 218844 583754 218872
rect 575624 218832 575630 218844
rect 563388 218708 567516 218736
rect 563388 218696 563394 218708
rect 567654 218696 567660 218748
rect 567712 218736 567718 218748
rect 568114 218736 568120 218748
rect 567712 218708 568120 218736
rect 567712 218696 567718 218708
rect 568114 218696 568120 218708
rect 568172 218696 568178 218748
rect 572714 218736 572720 218748
rect 570616 218708 572720 218736
rect 570616 218600 570644 218708
rect 572714 218696 572720 218708
rect 572772 218696 572778 218748
rect 572898 218696 572904 218748
rect 572956 218736 572962 218748
rect 575566 218736 575572 218748
rect 572956 218708 575244 218736
rect 572956 218696 572962 218708
rect 575216 218668 575244 218708
rect 575446 218708 575572 218736
rect 575446 218668 575474 218708
rect 575566 218696 575572 218708
rect 575624 218696 575630 218748
rect 575842 218696 575848 218748
rect 575900 218736 575906 218748
rect 582926 218736 582932 218748
rect 575900 218708 582932 218736
rect 575900 218696 575906 218708
rect 582926 218696 582932 218708
rect 582984 218696 582990 218748
rect 575216 218640 575474 218668
rect 529256 218572 548564 218600
rect 548628 218572 570644 218600
rect 529256 218560 529262 218572
rect 501104 218436 509924 218464
rect 501104 218424 501110 218436
rect 514754 218424 514760 218476
rect 514812 218464 514818 218476
rect 538858 218464 538864 218476
rect 514812 218436 538864 218464
rect 514812 218424 514818 218436
rect 538858 218424 538864 218436
rect 538916 218424 538922 218476
rect 542354 218424 542360 218476
rect 542412 218464 542418 218476
rect 543642 218464 543648 218476
rect 542412 218436 543648 218464
rect 542412 218424 542418 218436
rect 543642 218424 543648 218436
rect 543700 218424 543706 218476
rect 545942 218424 545948 218476
rect 546000 218464 546006 218476
rect 548628 218464 548656 218572
rect 571150 218560 571156 218612
rect 571208 218600 571214 218612
rect 571978 218600 571984 218612
rect 571208 218572 571984 218600
rect 571208 218560 571214 218572
rect 571978 218560 571984 218572
rect 572036 218560 572042 218612
rect 572530 218560 572536 218612
rect 572588 218600 572594 218612
rect 583726 218600 583754 218844
rect 591942 218696 591948 218748
rect 592000 218736 592006 218748
rect 592126 218736 592132 218748
rect 592000 218708 592132 218736
rect 592000 218696 592006 218708
rect 592126 218696 592132 218708
rect 592184 218696 592190 218748
rect 675846 218628 675852 218680
rect 675904 218668 675910 218680
rect 677042 218668 677048 218680
rect 675904 218640 677048 218668
rect 675904 218628 675910 218640
rect 677042 218628 677048 218640
rect 677100 218628 677106 218680
rect 596818 218600 596824 218612
rect 572588 218572 575152 218600
rect 583726 218572 596824 218600
rect 572588 218560 572594 218572
rect 546000 218436 548656 218464
rect 546000 218424 546006 218436
rect 548794 218424 548800 218476
rect 548852 218464 548858 218476
rect 567378 218464 567384 218476
rect 548852 218436 567384 218464
rect 548852 218424 548858 218436
rect 567378 218424 567384 218436
rect 567436 218424 567442 218476
rect 567562 218424 567568 218476
rect 567620 218464 567626 218476
rect 575124 218464 575152 218572
rect 596818 218560 596824 218572
rect 596876 218560 596882 218612
rect 575750 218464 575756 218476
rect 567620 218436 575060 218464
rect 575124 218436 575756 218464
rect 567620 218424 567626 218436
rect 75546 218288 75552 218340
rect 75604 218328 75610 218340
rect 83458 218328 83464 218340
rect 75604 218300 83464 218328
rect 75604 218288 75610 218300
rect 83458 218288 83464 218300
rect 83516 218288 83522 218340
rect 100386 218288 100392 218340
rect 100444 218328 100450 218340
rect 105814 218328 105820 218340
rect 100444 218300 105820 218328
rect 100444 218288 100450 218300
rect 105814 218288 105820 218300
rect 105872 218288 105878 218340
rect 113634 218288 113640 218340
rect 113692 218328 113698 218340
rect 113692 218300 128492 218328
rect 113692 218288 113698 218300
rect 56318 218152 56324 218204
rect 56376 218192 56382 218204
rect 62758 218192 62764 218204
rect 56376 218164 62764 218192
rect 56376 218152 56382 218164
rect 62758 218152 62764 218164
rect 62816 218152 62822 218204
rect 79686 218152 79692 218204
rect 79744 218192 79750 218204
rect 82078 218192 82084 218204
rect 79744 218164 82084 218192
rect 79744 218152 79750 218164
rect 82078 218152 82084 218164
rect 82136 218152 82142 218204
rect 120258 218152 120264 218204
rect 120316 218192 120322 218204
rect 120316 218164 122742 218192
rect 120316 218152 120322 218164
rect 55674 218016 55680 218068
rect 55732 218056 55738 218068
rect 56502 218056 56508 218068
rect 55732 218028 56508 218056
rect 55732 218016 55738 218028
rect 56502 218016 56508 218028
rect 56560 218016 56566 218068
rect 57330 218016 57336 218068
rect 57388 218056 57394 218068
rect 57882 218056 57888 218068
rect 57388 218028 57888 218056
rect 57388 218016 57394 218028
rect 57882 218016 57888 218028
rect 57940 218016 57946 218068
rect 58158 218016 58164 218068
rect 58216 218056 58222 218068
rect 61286 218056 61292 218068
rect 58216 218028 61292 218056
rect 58216 218016 58222 218028
rect 61286 218016 61292 218028
rect 61344 218016 61350 218068
rect 65610 218016 65616 218068
rect 65668 218056 65674 218068
rect 66162 218056 66168 218068
rect 65668 218028 66168 218056
rect 65668 218016 65674 218028
rect 66162 218016 66168 218028
rect 66220 218016 66226 218068
rect 73890 218016 73896 218068
rect 73948 218056 73954 218068
rect 74442 218056 74448 218068
rect 73948 218028 74448 218056
rect 73948 218016 73954 218028
rect 74442 218016 74448 218028
rect 74500 218016 74506 218068
rect 74718 218016 74724 218068
rect 74776 218056 74782 218068
rect 75822 218056 75828 218068
rect 74776 218028 75828 218056
rect 74776 218016 74782 218028
rect 75822 218016 75828 218028
rect 75880 218016 75886 218068
rect 78030 218016 78036 218068
rect 78088 218056 78094 218068
rect 78582 218056 78588 218068
rect 78088 218028 78588 218056
rect 78088 218016 78094 218028
rect 78582 218016 78588 218028
rect 78640 218016 78646 218068
rect 78858 218016 78864 218068
rect 78916 218056 78922 218068
rect 79962 218056 79968 218068
rect 78916 218028 79968 218056
rect 78916 218016 78922 218028
rect 79962 218016 79968 218028
rect 80020 218016 80026 218068
rect 82170 218016 82176 218068
rect 82228 218056 82234 218068
rect 82722 218056 82728 218068
rect 82228 218028 82728 218056
rect 82228 218016 82234 218028
rect 82722 218016 82728 218028
rect 82780 218016 82786 218068
rect 84654 218016 84660 218068
rect 84712 218056 84718 218068
rect 85482 218056 85488 218068
rect 84712 218028 85488 218056
rect 84712 218016 84718 218028
rect 85482 218016 85488 218028
rect 85540 218016 85546 218068
rect 86310 218016 86316 218068
rect 86368 218056 86374 218068
rect 86862 218056 86868 218068
rect 86368 218028 86868 218056
rect 86368 218016 86374 218028
rect 86862 218016 86868 218028
rect 86920 218016 86926 218068
rect 87138 218016 87144 218068
rect 87196 218056 87202 218068
rect 88242 218056 88248 218068
rect 87196 218028 88248 218056
rect 87196 218016 87202 218028
rect 88242 218016 88248 218028
rect 88300 218016 88306 218068
rect 88794 218016 88800 218068
rect 88852 218056 88858 218068
rect 89438 218056 89444 218068
rect 88852 218028 89444 218056
rect 88852 218016 88858 218028
rect 89438 218016 89444 218028
rect 89496 218016 89502 218068
rect 94590 218016 94596 218068
rect 94648 218056 94654 218068
rect 95142 218056 95148 218068
rect 94648 218028 95148 218056
rect 94648 218016 94654 218028
rect 95142 218016 95148 218028
rect 95200 218016 95206 218068
rect 97074 218016 97080 218068
rect 97132 218056 97138 218068
rect 97994 218056 98000 218068
rect 97132 218028 98000 218056
rect 97132 218016 97138 218028
rect 97994 218016 98000 218028
rect 98052 218016 98058 218068
rect 98730 218016 98736 218068
rect 98788 218056 98794 218068
rect 99282 218056 99288 218068
rect 98788 218028 99288 218056
rect 98788 218016 98794 218028
rect 99282 218016 99288 218028
rect 99340 218016 99346 218068
rect 99558 218016 99564 218068
rect 99616 218056 99622 218068
rect 100662 218056 100668 218068
rect 99616 218028 100668 218056
rect 99616 218016 99622 218028
rect 100662 218016 100668 218028
rect 100720 218016 100726 218068
rect 101214 218016 101220 218068
rect 101272 218056 101278 218068
rect 102134 218056 102140 218068
rect 101272 218028 102140 218056
rect 101272 218016 101278 218028
rect 102134 218016 102140 218028
rect 102192 218016 102198 218068
rect 102870 218016 102876 218068
rect 102928 218056 102934 218068
rect 103422 218056 103428 218068
rect 102928 218028 103428 218056
rect 102928 218016 102934 218028
rect 103422 218016 103428 218028
rect 103480 218016 103486 218068
rect 103698 218016 103704 218068
rect 103756 218056 103762 218068
rect 104802 218056 104808 218068
rect 103756 218028 104808 218056
rect 103756 218016 103762 218028
rect 104802 218016 104808 218028
rect 104860 218016 104866 218068
rect 105354 218016 105360 218068
rect 105412 218056 105418 218068
rect 105998 218056 106004 218068
rect 105412 218028 106004 218056
rect 105412 218016 105418 218028
rect 105998 218016 106004 218028
rect 106056 218016 106062 218068
rect 109494 218016 109500 218068
rect 109552 218056 109558 218068
rect 110138 218056 110144 218068
rect 109552 218028 110144 218056
rect 109552 218016 109558 218028
rect 110138 218016 110144 218028
rect 110196 218016 110202 218068
rect 110322 218016 110328 218068
rect 110380 218056 110386 218068
rect 110966 218056 110972 218068
rect 110380 218028 110972 218056
rect 110380 218016 110386 218028
rect 110966 218016 110972 218028
rect 111024 218016 111030 218068
rect 111978 218016 111984 218068
rect 112036 218056 112042 218068
rect 112806 218056 112812 218068
rect 112036 218028 112812 218056
rect 112036 218016 112042 218028
rect 112806 218016 112812 218028
rect 112864 218016 112870 218068
rect 115290 218016 115296 218068
rect 115348 218056 115354 218068
rect 115842 218056 115848 218068
rect 115348 218028 115848 218056
rect 115348 218016 115354 218028
rect 115842 218016 115848 218028
rect 115900 218016 115906 218068
rect 116118 218016 116124 218068
rect 116176 218056 116182 218068
rect 117222 218056 117228 218068
rect 116176 218028 117228 218056
rect 116176 218016 116182 218028
rect 117222 218016 117228 218028
rect 117280 218016 117286 218068
rect 119430 218016 119436 218068
rect 119488 218056 119494 218068
rect 119982 218056 119988 218068
rect 119488 218028 119988 218056
rect 119488 218016 119494 218028
rect 119982 218016 119988 218028
rect 120040 218016 120046 218068
rect 121914 218016 121920 218068
rect 121972 218056 121978 218068
rect 122558 218056 122564 218068
rect 121972 218028 122564 218056
rect 121972 218016 121978 218028
rect 122558 218016 122564 218028
rect 122616 218016 122622 218068
rect 122714 218056 122742 218164
rect 127710 218152 127716 218204
rect 127768 218192 127774 218204
rect 128262 218192 128268 218204
rect 127768 218164 128268 218192
rect 127768 218152 127774 218164
rect 128262 218152 128268 218164
rect 128320 218152 128326 218204
rect 128464 218192 128492 218300
rect 128722 218288 128728 218340
rect 128780 218328 128786 218340
rect 174538 218328 174544 218340
rect 128780 218300 174544 218328
rect 128780 218288 128786 218300
rect 174538 218288 174544 218300
rect 174596 218288 174602 218340
rect 176286 218328 176292 218340
rect 174740 218300 176292 218328
rect 159634 218192 159640 218204
rect 128464 218164 159640 218192
rect 159634 218152 159640 218164
rect 159692 218152 159698 218204
rect 166442 218192 166448 218204
rect 159836 218164 166448 218192
rect 159836 218056 159864 218164
rect 166442 218152 166448 218164
rect 166500 218152 166506 218204
rect 166626 218152 166632 218204
rect 166684 218192 166690 218204
rect 166994 218192 167000 218204
rect 166684 218164 167000 218192
rect 166684 218152 166690 218164
rect 166994 218152 167000 218164
rect 167052 218152 167058 218204
rect 168098 218152 168104 218204
rect 168156 218192 168162 218204
rect 171042 218192 171048 218204
rect 168156 218164 171048 218192
rect 168156 218152 168162 218164
rect 171042 218152 171048 218164
rect 171100 218152 171106 218204
rect 171594 218152 171600 218204
rect 171652 218192 171658 218204
rect 174740 218192 174768 218300
rect 176286 218288 176292 218300
rect 176344 218288 176350 218340
rect 185578 218328 185584 218340
rect 177362 218300 185584 218328
rect 171652 218164 174768 218192
rect 171652 218152 171658 218164
rect 175734 218152 175740 218204
rect 175792 218192 175798 218204
rect 176470 218192 176476 218204
rect 175792 218164 176476 218192
rect 175792 218152 175798 218164
rect 176470 218152 176476 218164
rect 176528 218152 176534 218204
rect 122714 218028 159864 218056
rect 160002 218016 160008 218068
rect 160060 218056 160066 218068
rect 166810 218056 166816 218068
rect 160060 218028 166816 218056
rect 160060 218016 160066 218028
rect 166810 218016 166816 218028
rect 166868 218016 166874 218068
rect 167454 218016 167460 218068
rect 167512 218056 167518 218068
rect 168282 218056 168288 218068
rect 167512 218028 168288 218056
rect 167512 218016 167518 218028
rect 168282 218016 168288 218028
rect 168340 218016 168346 218068
rect 169110 218016 169116 218068
rect 169168 218056 169174 218068
rect 169570 218056 169576 218068
rect 169168 218028 169576 218056
rect 169168 218016 169174 218028
rect 169570 218016 169576 218028
rect 169628 218016 169634 218068
rect 173250 218016 173256 218068
rect 173308 218056 173314 218068
rect 173308 218028 173940 218056
rect 173308 218016 173314 218028
rect 173912 217920 173940 218028
rect 174078 218016 174084 218068
rect 174136 218056 174142 218068
rect 175182 218056 175188 218068
rect 174136 218028 175188 218056
rect 174136 218016 174142 218028
rect 175182 218016 175188 218028
rect 175240 218016 175246 218068
rect 176562 218016 176568 218068
rect 176620 218056 176626 218068
rect 177206 218056 177212 218068
rect 176620 218028 177212 218056
rect 176620 218016 176626 218028
rect 177206 218016 177212 218028
rect 177264 218016 177270 218068
rect 177362 217920 177390 218300
rect 185578 218288 185584 218300
rect 185636 218288 185642 218340
rect 185762 218288 185768 218340
rect 185820 218328 185826 218340
rect 192294 218328 192300 218340
rect 185820 218300 192300 218328
rect 185820 218288 185826 218300
rect 192294 218288 192300 218300
rect 192352 218288 192358 218340
rect 193766 218288 193772 218340
rect 193824 218328 193830 218340
rect 229370 218328 229376 218340
rect 193824 218300 229376 218328
rect 193824 218288 193830 218300
rect 229370 218288 229376 218300
rect 229428 218288 229434 218340
rect 229554 218288 229560 218340
rect 229612 218328 229618 218340
rect 231118 218328 231124 218340
rect 229612 218300 231124 218328
rect 229612 218288 229618 218300
rect 231118 218288 231124 218300
rect 231176 218288 231182 218340
rect 232866 218288 232872 218340
rect 232924 218328 232930 218340
rect 234798 218328 234804 218340
rect 232924 218300 234804 218328
rect 232924 218288 232930 218300
rect 234798 218288 234804 218300
rect 234856 218288 234862 218340
rect 365346 218288 365352 218340
rect 365404 218328 365410 218340
rect 373258 218328 373264 218340
rect 365404 218300 373264 218328
rect 365404 218288 365410 218300
rect 373258 218288 373264 218300
rect 373316 218288 373322 218340
rect 426618 218288 426624 218340
rect 426676 218328 426682 218340
rect 429562 218328 429568 218340
rect 426676 218300 429568 218328
rect 426676 218288 426682 218300
rect 429562 218288 429568 218300
rect 429620 218288 429626 218340
rect 434898 218288 434904 218340
rect 434956 218328 434962 218340
rect 436646 218328 436652 218340
rect 434956 218300 436652 218328
rect 434956 218288 434962 218300
rect 436646 218288 436652 218300
rect 436704 218288 436710 218340
rect 500034 218288 500040 218340
rect 500092 218328 500098 218340
rect 507118 218328 507124 218340
rect 500092 218300 507124 218328
rect 500092 218288 500098 218300
rect 507118 218288 507124 218300
rect 507176 218288 507182 218340
rect 507670 218288 507676 218340
rect 507728 218328 507734 218340
rect 529198 218328 529204 218340
rect 507728 218300 529204 218328
rect 507728 218288 507734 218300
rect 529198 218288 529204 218300
rect 529256 218288 529262 218340
rect 529566 218288 529572 218340
rect 529624 218328 529630 218340
rect 571150 218328 571156 218340
rect 529624 218300 571156 218328
rect 529624 218288 529630 218300
rect 571150 218288 571156 218300
rect 571208 218288 571214 218340
rect 572530 218328 572536 218340
rect 571444 218300 572536 218328
rect 179874 218152 179880 218204
rect 179932 218192 179938 218204
rect 221090 218192 221096 218204
rect 179932 218164 221096 218192
rect 179932 218152 179938 218164
rect 221090 218152 221096 218164
rect 221148 218152 221154 218204
rect 221274 218152 221280 218204
rect 221332 218192 221338 218204
rect 221826 218192 221832 218204
rect 221332 218164 221832 218192
rect 221332 218152 221338 218164
rect 221826 218152 221832 218164
rect 221884 218152 221890 218204
rect 222930 218152 222936 218204
rect 222988 218192 222994 218204
rect 223390 218192 223396 218204
rect 222988 218164 223396 218192
rect 222988 218152 222994 218164
rect 223390 218152 223396 218164
rect 223448 218152 223454 218204
rect 223758 218152 223764 218204
rect 223816 218192 223822 218204
rect 224862 218192 224868 218204
rect 223816 218164 224868 218192
rect 223816 218152 223822 218164
rect 224862 218152 224868 218164
rect 224920 218152 224926 218204
rect 227898 218152 227904 218204
rect 227956 218192 227962 218204
rect 229738 218192 229744 218204
rect 227956 218164 229744 218192
rect 227956 218152 227962 218164
rect 229738 218152 229744 218164
rect 229796 218152 229802 218204
rect 235350 218152 235356 218204
rect 235408 218192 235414 218204
rect 235902 218192 235908 218204
rect 235408 218164 235908 218192
rect 235408 218152 235414 218164
rect 235902 218152 235908 218164
rect 235960 218152 235966 218204
rect 236178 218152 236184 218204
rect 236236 218192 236242 218204
rect 236914 218192 236920 218204
rect 236236 218164 236920 218192
rect 236236 218152 236242 218164
rect 236914 218152 236920 218164
rect 236972 218152 236978 218204
rect 249058 218192 249064 218204
rect 238726 218164 249064 218192
rect 177574 218016 177580 218068
rect 177632 218056 177638 218068
rect 181346 218056 181352 218068
rect 177632 218028 181352 218056
rect 177632 218016 177638 218028
rect 181346 218016 181352 218028
rect 181404 218016 181410 218068
rect 182358 218016 182364 218068
rect 182416 218056 182422 218068
rect 183278 218056 183284 218068
rect 182416 218028 183284 218056
rect 182416 218016 182422 218028
rect 183278 218016 183284 218028
rect 183336 218016 183342 218068
rect 184014 218016 184020 218068
rect 184072 218056 184078 218068
rect 184658 218056 184664 218068
rect 184072 218028 184664 218056
rect 184072 218016 184078 218028
rect 184658 218016 184664 218028
rect 184716 218016 184722 218068
rect 185670 218016 185676 218068
rect 185728 218056 185734 218068
rect 186130 218056 186136 218068
rect 185728 218028 186136 218056
rect 185728 218016 185734 218028
rect 186130 218016 186136 218028
rect 186188 218016 186194 218068
rect 186498 218016 186504 218068
rect 186556 218056 186562 218068
rect 186556 218028 189672 218056
rect 186556 218016 186562 218028
rect 173912 217892 177390 217920
rect 189644 217920 189672 218028
rect 189810 218016 189816 218068
rect 189868 218056 189874 218068
rect 190270 218056 190276 218068
rect 189868 218028 190276 218056
rect 189868 218016 189874 218028
rect 190270 218016 190276 218028
rect 190328 218016 190334 218068
rect 193766 218056 193772 218068
rect 190426 218028 193772 218056
rect 190426 217920 190454 218028
rect 193766 218016 193772 218028
rect 193824 218016 193830 218068
rect 193950 218016 193956 218068
rect 194008 218056 194014 218068
rect 194502 218056 194508 218068
rect 194008 218028 194508 218056
rect 194008 218016 194014 218028
rect 194502 218016 194508 218028
rect 194560 218016 194566 218068
rect 194778 218016 194784 218068
rect 194836 218056 194842 218068
rect 195882 218056 195888 218068
rect 194836 218028 195888 218056
rect 194836 218016 194842 218028
rect 195882 218016 195888 218028
rect 195940 218016 195946 218068
rect 196434 218016 196440 218068
rect 196492 218056 196498 218068
rect 197078 218056 197084 218068
rect 196492 218028 197084 218056
rect 196492 218016 196498 218028
rect 197078 218016 197084 218028
rect 197136 218016 197142 218068
rect 198918 218016 198924 218068
rect 198976 218056 198982 218068
rect 200022 218056 200028 218068
rect 198976 218028 200028 218056
rect 198976 218016 198982 218028
rect 200022 218016 200028 218028
rect 200080 218016 200086 218068
rect 202230 218016 202236 218068
rect 202288 218056 202294 218068
rect 202690 218056 202696 218068
rect 202288 218028 202696 218056
rect 202288 218016 202294 218028
rect 202690 218016 202696 218028
rect 202748 218016 202754 218068
rect 203058 218016 203064 218068
rect 203116 218056 203122 218068
rect 203702 218056 203708 218068
rect 203116 218028 203708 218056
rect 203116 218016 203122 218028
rect 203702 218016 203708 218028
rect 203760 218016 203766 218068
rect 204714 218016 204720 218068
rect 204772 218056 204778 218068
rect 206002 218056 206008 218068
rect 204772 218028 206008 218056
rect 204772 218016 204778 218028
rect 206002 218016 206008 218028
rect 206060 218016 206066 218068
rect 210510 218016 210516 218068
rect 210568 218056 210574 218068
rect 210970 218056 210976 218068
rect 210568 218028 210976 218056
rect 210568 218016 210574 218028
rect 210970 218016 210976 218028
rect 211028 218016 211034 218068
rect 212994 218016 213000 218068
rect 213052 218056 213058 218068
rect 213052 218028 215340 218056
rect 213052 218016 213058 218028
rect 189644 217892 190454 217920
rect 215312 217920 215340 218028
rect 215478 218016 215484 218068
rect 215536 218056 215542 218068
rect 216490 218056 216496 218068
rect 215536 218028 216496 218056
rect 215536 218016 215542 218028
rect 216490 218016 216496 218028
rect 216548 218016 216554 218068
rect 238726 218056 238754 218164
rect 249058 218152 249064 218164
rect 249116 218152 249122 218204
rect 249426 218152 249432 218204
rect 249484 218192 249490 218204
rect 251726 218192 251732 218204
rect 249484 218164 251732 218192
rect 249484 218152 249490 218164
rect 251726 218152 251732 218164
rect 251784 218152 251790 218204
rect 269298 218152 269304 218204
rect 269356 218192 269362 218204
rect 273898 218192 273904 218204
rect 269356 218164 273904 218192
rect 269356 218152 269362 218164
rect 273898 218152 273904 218164
rect 273956 218152 273962 218204
rect 299106 218152 299112 218204
rect 299164 218192 299170 218204
rect 300302 218192 300308 218204
rect 299164 218164 300308 218192
rect 299164 218152 299170 218164
rect 300302 218152 300308 218164
rect 300360 218152 300366 218204
rect 304074 218152 304080 218204
rect 304132 218192 304138 218204
rect 305638 218192 305644 218204
rect 304132 218164 305644 218192
rect 304132 218152 304138 218164
rect 305638 218152 305644 218164
rect 305696 218152 305702 218204
rect 310698 218152 310704 218204
rect 310756 218192 310762 218204
rect 315298 218192 315304 218204
rect 310756 218164 315304 218192
rect 310756 218152 310762 218164
rect 315298 218152 315304 218164
rect 315356 218152 315362 218204
rect 330662 218152 330668 218204
rect 330720 218192 330726 218204
rect 333238 218192 333244 218204
rect 330720 218164 333244 218192
rect 330720 218152 330726 218164
rect 333238 218152 333244 218164
rect 333296 218152 333302 218204
rect 348786 218152 348792 218204
rect 348844 218192 348850 218204
rect 351178 218192 351184 218204
rect 348844 218164 351184 218192
rect 348844 218152 348850 218164
rect 351178 218152 351184 218164
rect 351236 218152 351242 218204
rect 364518 218152 364524 218204
rect 364576 218192 364582 218204
rect 367646 218192 367652 218204
rect 364576 218164 367652 218192
rect 364576 218152 364582 218164
rect 367646 218152 367652 218164
rect 367704 218152 367710 218204
rect 369486 218152 369492 218204
rect 369544 218192 369550 218204
rect 370498 218192 370504 218204
rect 369544 218164 370504 218192
rect 369544 218152 369550 218164
rect 370498 218152 370504 218164
rect 370556 218152 370562 218204
rect 376938 218152 376944 218204
rect 376996 218192 377002 218204
rect 382918 218192 382924 218204
rect 376996 218164 382924 218192
rect 376996 218152 377002 218164
rect 382918 218152 382924 218164
rect 382976 218152 382982 218204
rect 386874 218152 386880 218204
rect 386932 218192 386938 218204
rect 388438 218192 388444 218204
rect 386932 218164 388444 218192
rect 386932 218152 386938 218164
rect 388438 218152 388444 218164
rect 388496 218152 388502 218204
rect 394326 218152 394332 218204
rect 394384 218192 394390 218204
rect 402238 218192 402244 218204
rect 394384 218164 402244 218192
rect 394384 218152 394390 218164
rect 402238 218152 402244 218164
rect 402296 218152 402302 218204
rect 407574 218152 407580 218204
rect 407632 218192 407638 218204
rect 411898 218192 411904 218204
rect 407632 218164 411904 218192
rect 407632 218152 407638 218164
rect 411898 218152 411904 218164
rect 411956 218152 411962 218204
rect 422478 218152 422484 218204
rect 422536 218192 422542 218204
rect 425422 218192 425428 218204
rect 422536 218164 425428 218192
rect 422536 218152 422542 218164
rect 425422 218152 425428 218164
rect 425480 218152 425486 218204
rect 425790 218152 425796 218204
rect 425848 218192 425854 218204
rect 428458 218192 428464 218204
rect 425848 218164 428464 218192
rect 425848 218152 425854 218164
rect 428458 218152 428464 218164
rect 428516 218152 428522 218204
rect 433242 218152 433248 218204
rect 433300 218192 433306 218204
rect 435266 218192 435272 218204
rect 433300 218164 435272 218192
rect 433300 218152 433306 218164
rect 435266 218152 435272 218164
rect 435324 218152 435330 218204
rect 455046 218152 455052 218204
rect 455104 218192 455110 218204
rect 460474 218192 460480 218204
rect 455104 218164 460480 218192
rect 455104 218152 455110 218164
rect 460474 218152 460480 218164
rect 460532 218152 460538 218204
rect 461946 218152 461952 218204
rect 462004 218192 462010 218204
rect 466270 218192 466276 218204
rect 462004 218164 466276 218192
rect 462004 218152 462010 218164
rect 466270 218152 466276 218164
rect 466328 218152 466334 218204
rect 494606 218152 494612 218204
rect 494664 218192 494670 218204
rect 495250 218192 495256 218204
rect 494664 218164 495256 218192
rect 494664 218152 494670 218164
rect 495250 218152 495256 218164
rect 495308 218192 495314 218204
rect 519722 218192 519728 218204
rect 495308 218164 519728 218192
rect 495308 218152 495314 218164
rect 519722 218152 519728 218164
rect 519780 218152 519786 218204
rect 519906 218152 519912 218204
rect 519964 218192 519970 218204
rect 524598 218192 524604 218204
rect 519964 218164 524604 218192
rect 519964 218152 519970 218164
rect 524598 218152 524604 218164
rect 524656 218152 524662 218204
rect 527542 218152 527548 218204
rect 527600 218192 527606 218204
rect 571444 218192 571472 218300
rect 572530 218288 572536 218300
rect 572588 218288 572594 218340
rect 572714 218288 572720 218340
rect 572772 218328 572778 218340
rect 574830 218328 574836 218340
rect 572772 218300 574836 218328
rect 572772 218288 572778 218300
rect 574830 218288 574836 218300
rect 574888 218288 574894 218340
rect 575032 218328 575060 218436
rect 575750 218424 575756 218436
rect 575808 218424 575814 218476
rect 576578 218424 576584 218476
rect 576636 218464 576642 218476
rect 607122 218464 607128 218476
rect 576636 218436 607128 218464
rect 576636 218424 576642 218436
rect 607122 218424 607128 218436
rect 607180 218424 607186 218476
rect 604454 218328 604460 218340
rect 575032 218300 604460 218328
rect 604454 218288 604460 218300
rect 604512 218288 604518 218340
rect 527600 218164 571472 218192
rect 527600 218152 527606 218164
rect 571610 218152 571616 218204
rect 571668 218192 571674 218204
rect 581914 218192 581920 218204
rect 571668 218164 581920 218192
rect 571668 218152 571674 218164
rect 581914 218152 581920 218164
rect 581972 218152 581978 218204
rect 582098 218152 582104 218204
rect 582156 218192 582162 218204
rect 582558 218192 582564 218204
rect 582156 218164 582564 218192
rect 582156 218152 582162 218164
rect 582558 218152 582564 218164
rect 582616 218152 582622 218204
rect 582742 218152 582748 218204
rect 582800 218192 582806 218204
rect 592310 218192 592316 218204
rect 582800 218164 592316 218192
rect 582800 218152 582806 218164
rect 592310 218152 592316 218164
rect 592368 218152 592374 218204
rect 676398 218084 676404 218136
rect 676456 218124 676462 218136
rect 677594 218124 677600 218136
rect 676456 218096 677600 218124
rect 676456 218084 676462 218096
rect 677594 218084 677600 218096
rect 677652 218084 677658 218136
rect 216692 218028 238754 218056
rect 216692 217920 216720 218028
rect 244458 218016 244464 218068
rect 244516 218056 244522 218068
rect 247586 218056 247592 218068
rect 244516 218028 247592 218056
rect 244516 218016 244522 218028
rect 247586 218016 247592 218028
rect 247644 218016 247650 218068
rect 247770 218016 247776 218068
rect 247828 218056 247834 218068
rect 248230 218056 248236 218068
rect 247828 218028 248236 218056
rect 247828 218016 247834 218028
rect 248230 218016 248236 218028
rect 248288 218016 248294 218068
rect 248598 218016 248604 218068
rect 248656 218056 248662 218068
rect 249702 218056 249708 218068
rect 248656 218028 249708 218056
rect 248656 218016 248662 218028
rect 249702 218016 249708 218028
rect 249760 218016 249766 218068
rect 250254 218016 250260 218068
rect 250312 218056 250318 218068
rect 251174 218056 251180 218068
rect 250312 218028 251180 218056
rect 250312 218016 250318 218028
rect 251174 218016 251180 218028
rect 251232 218016 251238 218068
rect 251910 218016 251916 218068
rect 251968 218056 251974 218068
rect 252462 218056 252468 218068
rect 251968 218028 252468 218056
rect 251968 218016 251974 218028
rect 252462 218016 252468 218028
rect 252520 218016 252526 218068
rect 262674 218016 262680 218068
rect 262732 218056 262738 218068
rect 263594 218056 263600 218068
rect 262732 218028 263600 218056
rect 262732 218016 262738 218028
rect 263594 218016 263600 218028
rect 263652 218016 263658 218068
rect 264330 218016 264336 218068
rect 264388 218056 264394 218068
rect 264790 218056 264796 218068
rect 264388 218028 264796 218056
rect 264388 218016 264394 218028
rect 264790 218016 264796 218028
rect 264848 218016 264854 218068
rect 265158 218016 265164 218068
rect 265216 218056 265222 218068
rect 266262 218056 266268 218068
rect 265216 218028 266268 218056
rect 265216 218016 265222 218028
rect 266262 218016 266268 218028
rect 266320 218016 266326 218068
rect 266814 218016 266820 218068
rect 266872 218056 266878 218068
rect 267688 218056 267694 218068
rect 266872 218028 267694 218056
rect 266872 218016 266878 218028
rect 267688 218016 267694 218028
rect 267746 218016 267752 218068
rect 268470 218016 268476 218068
rect 268528 218056 268534 218068
rect 269022 218056 269028 218068
rect 268528 218028 269028 218056
rect 268528 218016 268534 218028
rect 269022 218016 269028 218028
rect 269080 218016 269086 218068
rect 270954 218016 270960 218068
rect 271012 218056 271018 218068
rect 271598 218056 271604 218068
rect 271012 218028 271604 218056
rect 271012 218016 271018 218028
rect 271598 218016 271604 218028
rect 271656 218016 271662 218068
rect 276750 218016 276756 218068
rect 276808 218056 276814 218068
rect 277210 218056 277216 218068
rect 276808 218028 277216 218056
rect 276808 218016 276814 218028
rect 277210 218016 277216 218028
rect 277268 218016 277274 218068
rect 277578 218016 277584 218068
rect 277636 218056 277642 218068
rect 278498 218056 278504 218068
rect 277636 218028 278504 218056
rect 277636 218016 277642 218028
rect 278498 218016 278504 218028
rect 278556 218016 278562 218068
rect 281718 218016 281724 218068
rect 281776 218056 281782 218068
rect 282546 218056 282552 218068
rect 281776 218028 282552 218056
rect 281776 218016 281782 218028
rect 282546 218016 282552 218028
rect 282604 218016 282610 218068
rect 285030 218016 285036 218068
rect 285088 218056 285094 218068
rect 285490 218056 285496 218068
rect 285088 218028 285496 218056
rect 285088 218016 285094 218028
rect 285490 218016 285496 218028
rect 285548 218016 285554 218068
rect 287514 218016 287520 218068
rect 287572 218056 287578 218068
rect 288434 218056 288440 218068
rect 287572 218028 288440 218056
rect 287572 218016 287578 218028
rect 288434 218016 288440 218028
rect 288492 218016 288498 218068
rect 289170 218016 289176 218068
rect 289228 218056 289234 218068
rect 289630 218056 289636 218068
rect 289228 218028 289636 218056
rect 289228 218016 289234 218028
rect 289630 218016 289636 218028
rect 289688 218016 289694 218068
rect 293310 218016 293316 218068
rect 293368 218056 293374 218068
rect 293770 218056 293776 218068
rect 293368 218028 293776 218056
rect 293368 218016 293374 218028
rect 293770 218016 293776 218028
rect 293828 218016 293834 218068
rect 295794 218016 295800 218068
rect 295852 218056 295858 218068
rect 296438 218056 296444 218068
rect 295852 218028 296444 218056
rect 295852 218016 295858 218028
rect 296438 218016 296444 218028
rect 296496 218016 296502 218068
rect 297450 218016 297456 218068
rect 297508 218056 297514 218068
rect 298002 218056 298008 218068
rect 297508 218028 298008 218056
rect 297508 218016 297514 218028
rect 298002 218016 298008 218028
rect 298060 218016 298066 218068
rect 298278 218016 298284 218068
rect 298336 218056 298342 218068
rect 299290 218056 299296 218068
rect 298336 218028 299296 218056
rect 298336 218016 298342 218028
rect 299290 218016 299296 218028
rect 299348 218016 299354 218068
rect 301590 218016 301596 218068
rect 301648 218056 301654 218068
rect 302142 218056 302148 218068
rect 301648 218028 302148 218056
rect 301648 218016 301654 218028
rect 302142 218016 302148 218028
rect 302200 218016 302206 218068
rect 302418 218016 302424 218068
rect 302476 218056 302482 218068
rect 303706 218056 303712 218068
rect 302476 218028 303712 218056
rect 302476 218016 302482 218028
rect 303706 218016 303712 218028
rect 303764 218016 303770 218068
rect 305730 218016 305736 218068
rect 305788 218056 305794 218068
rect 306282 218056 306288 218068
rect 305788 218028 306288 218056
rect 305788 218016 305794 218028
rect 306282 218016 306288 218028
rect 306340 218016 306346 218068
rect 306558 218016 306564 218068
rect 306616 218056 306622 218068
rect 307662 218056 307668 218068
rect 306616 218028 307668 218056
rect 306616 218016 306622 218028
rect 307662 218016 307668 218028
rect 307720 218016 307726 218068
rect 308214 218016 308220 218068
rect 308272 218056 308278 218068
rect 308766 218056 308772 218068
rect 308272 218028 308772 218056
rect 308272 218016 308278 218028
rect 308766 218016 308772 218028
rect 308824 218016 308830 218068
rect 312354 218016 312360 218068
rect 312412 218056 312418 218068
rect 314470 218056 314476 218068
rect 312412 218028 314476 218056
rect 312412 218016 312418 218028
rect 314470 218016 314476 218028
rect 314528 218016 314534 218068
rect 314838 218016 314844 218068
rect 314896 218056 314902 218068
rect 315850 218056 315856 218068
rect 314896 218028 315856 218056
rect 314896 218016 314902 218028
rect 315850 218016 315856 218028
rect 315908 218016 315914 218068
rect 316494 218016 316500 218068
rect 316552 218056 316558 218068
rect 317138 218056 317144 218068
rect 316552 218028 317144 218056
rect 316552 218016 316558 218028
rect 317138 218016 317144 218028
rect 317196 218016 317202 218068
rect 318978 218016 318984 218068
rect 319036 218056 319042 218068
rect 319990 218056 319996 218068
rect 319036 218028 319996 218056
rect 319036 218016 319042 218028
rect 319990 218016 319996 218028
rect 320048 218016 320054 218068
rect 322290 218016 322296 218068
rect 322348 218056 322354 218068
rect 322842 218056 322848 218068
rect 322348 218028 322848 218056
rect 322348 218016 322354 218028
rect 322842 218016 322848 218028
rect 322900 218016 322906 218068
rect 324774 218016 324780 218068
rect 324832 218056 324838 218068
rect 325418 218056 325424 218068
rect 324832 218028 325424 218056
rect 324832 218016 324838 218028
rect 325418 218016 325424 218028
rect 325476 218016 325482 218068
rect 326430 218016 326436 218068
rect 326488 218056 326494 218068
rect 326890 218056 326896 218068
rect 326488 218028 326896 218056
rect 326488 218016 326494 218028
rect 326890 218016 326896 218028
rect 326948 218016 326954 218068
rect 328914 218016 328920 218068
rect 328972 218056 328978 218068
rect 330478 218056 330484 218068
rect 328972 218028 330484 218056
rect 328972 218016 328978 218028
rect 330478 218016 330484 218028
rect 330536 218016 330542 218068
rect 333054 218016 333060 218068
rect 333112 218056 333118 218068
rect 333882 218056 333888 218068
rect 333112 218028 333888 218056
rect 333112 218016 333118 218028
rect 333882 218016 333888 218028
rect 333940 218016 333946 218068
rect 334710 218016 334716 218068
rect 334768 218056 334774 218068
rect 335262 218056 335268 218068
rect 334768 218028 335268 218056
rect 334768 218016 334774 218028
rect 335262 218016 335268 218028
rect 335320 218016 335326 218068
rect 335538 218016 335544 218068
rect 335596 218056 335602 218068
rect 336366 218056 336372 218068
rect 335596 218028 336372 218056
rect 335596 218016 335602 218028
rect 336366 218016 336372 218028
rect 336424 218016 336430 218068
rect 339678 218016 339684 218068
rect 339736 218056 339742 218068
rect 340690 218056 340696 218068
rect 339736 218028 340696 218056
rect 339736 218016 339742 218028
rect 340690 218016 340696 218028
rect 340748 218016 340754 218068
rect 342990 218016 342996 218068
rect 343048 218056 343054 218068
rect 343542 218056 343548 218068
rect 343048 218028 343548 218056
rect 343048 218016 343054 218028
rect 343542 218016 343548 218028
rect 343600 218016 343606 218068
rect 347130 218016 347136 218068
rect 347188 218056 347194 218068
rect 347590 218056 347596 218068
rect 347188 218028 347596 218056
rect 347188 218016 347194 218028
rect 347590 218016 347596 218028
rect 347648 218016 347654 218068
rect 347958 218016 347964 218068
rect 348016 218056 348022 218068
rect 349062 218056 349068 218068
rect 348016 218028 349068 218056
rect 348016 218016 348022 218028
rect 349062 218016 349068 218028
rect 349120 218016 349126 218068
rect 349614 218016 349620 218068
rect 349672 218056 349678 218068
rect 350166 218056 350172 218068
rect 349672 218028 350172 218056
rect 349672 218016 349678 218028
rect 350166 218016 350172 218028
rect 350224 218016 350230 218068
rect 353754 218016 353760 218068
rect 353812 218056 353818 218068
rect 354582 218056 354588 218068
rect 353812 218028 354588 218056
rect 353812 218016 353818 218028
rect 354582 218016 354588 218028
rect 354640 218016 354646 218068
rect 356238 218016 356244 218068
rect 356296 218056 356302 218068
rect 357342 218056 357348 218068
rect 356296 218028 357348 218056
rect 356296 218016 356302 218028
rect 357342 218016 357348 218028
rect 357400 218016 357406 218068
rect 357894 218016 357900 218068
rect 357952 218056 357958 218068
rect 359366 218056 359372 218068
rect 357952 218028 359372 218056
rect 357952 218016 357958 218028
rect 359366 218016 359372 218028
rect 359424 218016 359430 218068
rect 363690 218016 363696 218068
rect 363748 218056 363754 218068
rect 364150 218056 364156 218068
rect 363748 218028 364156 218056
rect 363748 218016 363754 218028
rect 364150 218016 364156 218028
rect 364208 218016 364214 218068
rect 366174 218016 366180 218068
rect 366232 218056 366238 218068
rect 366910 218056 366916 218068
rect 366232 218028 366916 218056
rect 366232 218016 366238 218028
rect 366910 218016 366916 218028
rect 366968 218016 366974 218068
rect 368658 218016 368664 218068
rect 368716 218056 368722 218068
rect 369762 218056 369768 218068
rect 368716 218028 369768 218056
rect 368716 218016 368722 218028
rect 369762 218016 369768 218028
rect 369820 218016 369826 218068
rect 370314 218016 370320 218068
rect 370372 218056 370378 218068
rect 370958 218056 370964 218068
rect 370372 218028 370964 218056
rect 370372 218016 370378 218028
rect 370958 218016 370964 218028
rect 371016 218016 371022 218068
rect 371970 218016 371976 218068
rect 372028 218056 372034 218068
rect 372522 218056 372528 218068
rect 372028 218028 372528 218056
rect 372028 218016 372034 218028
rect 372522 218016 372528 218028
rect 372580 218016 372586 218068
rect 372798 218016 372804 218068
rect 372856 218056 372862 218068
rect 373810 218056 373816 218068
rect 372856 218028 373816 218056
rect 372856 218016 372862 218028
rect 373810 218016 373816 218028
rect 373868 218016 373874 218068
rect 376110 218016 376116 218068
rect 376168 218056 376174 218068
rect 376570 218056 376576 218068
rect 376168 218028 376576 218056
rect 376168 218016 376174 218028
rect 376570 218016 376576 218028
rect 376628 218016 376634 218068
rect 378594 218016 378600 218068
rect 378652 218056 378658 218068
rect 379330 218056 379336 218068
rect 378652 218028 379336 218056
rect 378652 218016 378658 218028
rect 379330 218016 379336 218028
rect 379388 218016 379394 218068
rect 381078 218016 381084 218068
rect 381136 218056 381142 218068
rect 381722 218056 381728 218068
rect 381136 218028 381728 218056
rect 381136 218016 381142 218028
rect 381722 218016 381728 218028
rect 381780 218016 381786 218068
rect 385218 218016 385224 218068
rect 385276 218056 385282 218068
rect 386322 218056 386328 218068
rect 385276 218028 386328 218056
rect 385276 218016 385282 218028
rect 386322 218016 386328 218028
rect 386380 218016 386386 218068
rect 388530 218016 388536 218068
rect 388588 218056 388594 218068
rect 389082 218056 389088 218068
rect 388588 218028 389088 218056
rect 388588 218016 388594 218028
rect 389082 218016 389088 218028
rect 389140 218016 389146 218068
rect 389358 218016 389364 218068
rect 389416 218056 389422 218068
rect 390278 218056 390284 218068
rect 389416 218028 390284 218056
rect 389416 218016 389422 218028
rect 390278 218016 390284 218028
rect 390336 218016 390342 218068
rect 392670 218016 392676 218068
rect 392728 218056 392734 218068
rect 393222 218056 393228 218068
rect 392728 218028 393228 218056
rect 392728 218016 392734 218028
rect 393222 218016 393228 218028
rect 393280 218016 393286 218068
rect 393498 218016 393504 218068
rect 393556 218056 393562 218068
rect 394602 218056 394608 218068
rect 393556 218028 394608 218056
rect 393556 218016 393562 218028
rect 394602 218016 394608 218028
rect 394660 218016 394666 218068
rect 395154 218016 395160 218068
rect 395212 218056 395218 218068
rect 395982 218056 395988 218068
rect 395212 218028 395988 218056
rect 395212 218016 395218 218028
rect 395982 218016 395988 218028
rect 396040 218016 396046 218068
rect 396810 218016 396816 218068
rect 396868 218056 396874 218068
rect 397362 218056 397368 218068
rect 396868 218028 397368 218056
rect 396868 218016 396874 218028
rect 397362 218016 397368 218028
rect 397420 218016 397426 218068
rect 400950 218016 400956 218068
rect 401008 218056 401014 218068
rect 401410 218056 401416 218068
rect 401008 218028 401416 218056
rect 401008 218016 401014 218028
rect 401410 218016 401416 218028
rect 401468 218016 401474 218068
rect 409230 218016 409236 218068
rect 409288 218056 409294 218068
rect 409782 218056 409788 218068
rect 409288 218028 409788 218056
rect 409288 218016 409294 218028
rect 409782 218016 409788 218028
rect 409840 218016 409846 218068
rect 410058 218016 410064 218068
rect 410116 218056 410122 218068
rect 411162 218056 411168 218068
rect 410116 218028 411168 218056
rect 410116 218016 410122 218028
rect 411162 218016 411168 218028
rect 411220 218016 411226 218068
rect 413370 218016 413376 218068
rect 413428 218056 413434 218068
rect 413830 218056 413836 218068
rect 413428 218028 413836 218056
rect 413428 218016 413434 218028
rect 413830 218016 413836 218028
rect 413888 218016 413894 218068
rect 418338 218016 418344 218068
rect 418396 218056 418402 218068
rect 419442 218056 419448 218068
rect 418396 218028 419448 218056
rect 418396 218016 418402 218028
rect 419442 218016 419448 218028
rect 419500 218016 419506 218068
rect 419994 218016 420000 218068
rect 420052 218056 420058 218068
rect 420914 218056 420920 218068
rect 420052 218028 420920 218056
rect 420052 218016 420058 218028
rect 420914 218016 420920 218028
rect 420972 218016 420978 218068
rect 424134 218016 424140 218068
rect 424192 218056 424198 218068
rect 426986 218056 426992 218068
rect 424192 218028 426992 218056
rect 424192 218016 424198 218028
rect 426986 218016 426992 218028
rect 427044 218016 427050 218068
rect 427446 218016 427452 218068
rect 427504 218056 427510 218068
rect 427906 218056 427912 218068
rect 427504 218028 427912 218056
rect 427504 218016 427510 218028
rect 427906 218016 427912 218028
rect 427964 218016 427970 218068
rect 429102 218016 429108 218068
rect 429160 218056 429166 218068
rect 430574 218056 430580 218068
rect 429160 218028 430580 218056
rect 429160 218016 429166 218028
rect 430574 218016 430580 218028
rect 430632 218016 430638 218068
rect 432414 218016 432420 218068
rect 432472 218056 432478 218068
rect 433794 218056 433800 218068
rect 432472 218028 433800 218056
rect 432472 218016 432478 218028
rect 433794 218016 433800 218028
rect 433852 218016 433858 218068
rect 435726 218016 435732 218068
rect 435784 218056 435790 218068
rect 436278 218056 436284 218068
rect 435784 218028 436284 218056
rect 435784 218016 435790 218028
rect 436278 218016 436284 218028
rect 436336 218016 436342 218068
rect 436554 218016 436560 218068
rect 436612 218056 436618 218068
rect 437474 218056 437480 218068
rect 436612 218028 437480 218056
rect 436612 218016 436618 218028
rect 437474 218016 437480 218028
rect 437532 218016 437538 218068
rect 438210 218016 438216 218068
rect 438268 218056 438274 218068
rect 438854 218056 438860 218068
rect 438268 218028 438860 218056
rect 438268 218016 438274 218028
rect 438854 218016 438860 218028
rect 438912 218016 438918 218068
rect 439866 218016 439872 218068
rect 439924 218056 439930 218068
rect 440326 218056 440332 218068
rect 439924 218028 440332 218056
rect 439924 218016 439930 218028
rect 440326 218016 440332 218028
rect 440384 218016 440390 218068
rect 453298 218016 453304 218068
rect 453356 218056 453362 218068
rect 455506 218056 455512 218068
rect 453356 218028 455512 218056
rect 453356 218016 453362 218028
rect 455506 218016 455512 218028
rect 455564 218016 455570 218068
rect 456702 218016 456708 218068
rect 456760 218056 456766 218068
rect 457162 218056 457168 218068
rect 456760 218028 457168 218056
rect 456760 218016 456766 218028
rect 457162 218016 457168 218028
rect 457220 218016 457226 218068
rect 463142 218016 463148 218068
rect 463200 218056 463206 218068
rect 464614 218056 464620 218068
rect 463200 218028 464620 218056
rect 463200 218016 463206 218028
rect 464614 218016 464620 218028
rect 464672 218016 464678 218068
rect 467282 218016 467288 218068
rect 467340 218056 467346 218068
rect 467926 218056 467932 218068
rect 467340 218028 467932 218056
rect 467340 218016 467346 218028
rect 467926 218016 467932 218028
rect 467984 218016 467990 218068
rect 470594 218016 470600 218068
rect 470652 218056 470658 218068
rect 472894 218056 472900 218068
rect 470652 218028 472900 218056
rect 470652 218016 470658 218028
rect 472894 218016 472900 218028
rect 472952 218016 472958 218068
rect 488718 218016 488724 218068
rect 488776 218056 488782 218068
rect 497550 218056 497556 218068
rect 488776 218028 497556 218056
rect 488776 218016 488782 218028
rect 497550 218016 497556 218028
rect 497608 218016 497614 218068
rect 505278 218016 505284 218068
rect 505336 218056 505342 218068
rect 505646 218056 505652 218068
rect 505336 218028 505652 218056
rect 505336 218016 505342 218028
rect 505646 218016 505652 218028
rect 505704 218056 505710 218068
rect 613838 218056 613844 218068
rect 505704 218028 567194 218056
rect 505704 218016 505710 218028
rect 567166 217988 567194 218028
rect 576826 218028 613844 218056
rect 576826 217988 576854 218028
rect 613838 218016 613844 218028
rect 613896 218016 613902 218068
rect 567166 217960 576854 217988
rect 215312 217892 216720 217920
rect 550606 217892 560294 217920
rect 505462 217812 505468 217864
rect 505520 217852 505526 217864
rect 514662 217852 514668 217864
rect 505520 217824 514668 217852
rect 505520 217812 505526 217824
rect 514662 217812 514668 217824
rect 514720 217812 514726 217864
rect 528370 217812 528376 217864
rect 528428 217852 528434 217864
rect 550606 217852 550634 217892
rect 528428 217824 550634 217852
rect 560266 217852 560294 217892
rect 602890 217852 602896 217864
rect 560266 217824 602896 217852
rect 528428 217812 528434 217824
rect 602890 217812 602896 217824
rect 602948 217812 602954 217864
rect 603074 217812 603080 217864
rect 603132 217852 603138 217864
rect 612274 217852 612280 217864
rect 603132 217824 612280 217852
rect 603132 217812 603138 217824
rect 612274 217812 612280 217824
rect 612332 217812 612338 217864
rect 551002 217784 551008 217796
rect 550744 217756 551008 217784
rect 514478 217676 514484 217728
rect 514536 217716 514542 217728
rect 519906 217716 519912 217728
rect 514536 217688 519912 217716
rect 514536 217676 514542 217688
rect 519906 217676 519912 217688
rect 519964 217676 519970 217728
rect 533430 217676 533436 217728
rect 533488 217716 533494 217728
rect 542170 217716 542176 217728
rect 533488 217688 542176 217716
rect 533488 217676 533494 217688
rect 542170 217676 542176 217688
rect 542228 217676 542234 217728
rect 542354 217676 542360 217728
rect 542412 217716 542418 217728
rect 550744 217716 550772 217756
rect 551002 217744 551008 217756
rect 551060 217744 551066 217796
rect 542412 217688 550772 217716
rect 542412 217676 542418 217688
rect 551186 217676 551192 217728
rect 551244 217716 551250 217728
rect 603442 217716 603448 217728
rect 551244 217688 603448 217716
rect 551244 217676 551250 217688
rect 603442 217676 603448 217688
rect 603500 217676 603506 217728
rect 604454 217676 604460 217728
rect 604512 217716 604518 217728
rect 615678 217716 615684 217728
rect 604512 217688 615684 217716
rect 604512 217676 604518 217688
rect 615678 217676 615684 217688
rect 615736 217676 615742 217728
rect 523770 217540 523776 217592
rect 523828 217580 523834 217592
rect 524598 217580 524604 217592
rect 523828 217552 524604 217580
rect 523828 217540 523834 217552
rect 524598 217540 524604 217552
rect 524656 217540 524662 217592
rect 533706 217540 533712 217592
rect 533764 217580 533770 217592
rect 534258 217580 534264 217592
rect 533764 217552 534264 217580
rect 533764 217540 533770 217552
rect 534258 217540 534264 217552
rect 534316 217540 534322 217592
rect 538398 217540 538404 217592
rect 538456 217580 538462 217592
rect 542906 217580 542912 217592
rect 538456 217552 542912 217580
rect 538456 217540 538462 217552
rect 542906 217540 542912 217552
rect 542964 217540 542970 217592
rect 543458 217540 543464 217592
rect 543516 217580 543522 217592
rect 543688 217580 543694 217592
rect 543516 217552 543694 217580
rect 543516 217540 543522 217552
rect 543688 217540 543694 217552
rect 543746 217540 543752 217592
rect 543826 217540 543832 217592
rect 543884 217580 543890 217592
rect 557258 217580 557264 217592
rect 543884 217552 557264 217580
rect 543884 217540 543890 217552
rect 557258 217540 557264 217552
rect 557316 217540 557322 217592
rect 557534 217540 557540 217592
rect 557592 217580 557598 217592
rect 572714 217580 572720 217592
rect 557592 217552 572720 217580
rect 557592 217540 557598 217552
rect 572714 217540 572720 217552
rect 572772 217540 572778 217592
rect 575198 217580 575204 217592
rect 573100 217552 575204 217580
rect 573100 217512 573128 217552
rect 575198 217540 575204 217552
rect 575256 217540 575262 217592
rect 576026 217540 576032 217592
rect 576084 217580 576090 217592
rect 593506 217580 593512 217592
rect 576084 217552 593512 217580
rect 576084 217540 576090 217552
rect 593506 217540 593512 217552
rect 593564 217540 593570 217592
rect 596818 217540 596824 217592
rect 596876 217580 596882 217592
rect 623314 217580 623320 217592
rect 596876 217552 623320 217580
rect 596876 217540 596882 217552
rect 623314 217540 623320 217552
rect 623372 217540 623378 217592
rect 572916 217484 573128 217512
rect 524414 217404 524420 217456
rect 524472 217444 524478 217456
rect 541986 217444 541992 217456
rect 524472 217416 541992 217444
rect 524472 217404 524478 217416
rect 541986 217404 541992 217416
rect 542044 217404 542050 217456
rect 542170 217404 542176 217456
rect 542228 217444 542234 217456
rect 549070 217444 549076 217456
rect 542228 217416 549076 217444
rect 542228 217404 542234 217416
rect 549070 217404 549076 217416
rect 549128 217404 549134 217456
rect 549254 217404 549260 217456
rect 549312 217444 549318 217456
rect 551738 217444 551744 217456
rect 549312 217416 551744 217444
rect 549312 217404 549318 217416
rect 551738 217404 551744 217416
rect 551796 217404 551802 217456
rect 553486 217404 553492 217456
rect 553544 217444 553550 217456
rect 564158 217444 564164 217456
rect 553544 217416 564164 217444
rect 553544 217404 553550 217416
rect 564158 217404 564164 217416
rect 564216 217404 564222 217456
rect 564342 217404 564348 217456
rect 564400 217444 564406 217456
rect 571794 217444 571800 217456
rect 564400 217416 571800 217444
rect 564400 217404 564406 217416
rect 571794 217404 571800 217416
rect 571852 217404 571858 217456
rect 571978 217404 571984 217456
rect 572036 217444 572042 217456
rect 572530 217444 572536 217456
rect 572036 217416 572536 217444
rect 572036 217404 572042 217416
rect 572530 217404 572536 217416
rect 572588 217404 572594 217456
rect 572714 217404 572720 217456
rect 572772 217444 572778 217456
rect 572916 217444 572944 217484
rect 572772 217416 572944 217444
rect 572772 217404 572778 217416
rect 573266 217404 573272 217456
rect 573324 217444 573330 217456
rect 609054 217444 609060 217456
rect 573324 217416 609060 217444
rect 573324 217404 573330 217416
rect 609054 217404 609060 217416
rect 609112 217404 609118 217456
rect 542354 217308 542360 217320
rect 534046 217280 542360 217308
rect 436094 217200 436100 217252
rect 436152 217240 436158 217252
rect 437336 217240 437342 217252
rect 436152 217212 437342 217240
rect 436152 217200 436158 217212
rect 437336 217200 437342 217212
rect 437394 217200 437400 217252
rect 447134 217200 447140 217252
rect 447192 217240 447198 217252
rect 448100 217240 448106 217252
rect 447192 217212 448106 217240
rect 447192 217200 447198 217212
rect 448100 217200 448106 217212
rect 448158 217200 448164 217252
rect 448606 217200 448612 217252
rect 448664 217240 448670 217252
rect 449756 217240 449762 217252
rect 448664 217212 449762 217240
rect 448664 217200 448670 217212
rect 449756 217200 449762 217212
rect 449814 217200 449820 217252
rect 469306 217200 469312 217252
rect 469364 217240 469370 217252
rect 470456 217240 470462 217252
rect 469364 217212 470462 217240
rect 469364 217200 469370 217212
rect 470456 217200 470462 217212
rect 470514 217200 470520 217252
rect 530486 217200 530492 217252
rect 530544 217240 530550 217252
rect 530900 217240 530906 217252
rect 530544 217212 530906 217240
rect 530544 217200 530550 217212
rect 530900 217200 530906 217212
rect 530958 217240 530964 217252
rect 534046 217240 534074 217280
rect 542354 217268 542360 217280
rect 542412 217268 542418 217320
rect 548426 217308 548432 217320
rect 545776 217280 548432 217308
rect 530958 217212 534074 217240
rect 530958 217200 530964 217212
rect 535868 217132 535874 217184
rect 535926 217172 535932 217184
rect 545776 217172 545804 217280
rect 548426 217268 548432 217280
rect 548484 217268 548490 217320
rect 550266 217268 550272 217320
rect 550324 217308 550330 217320
rect 550324 217280 550496 217308
rect 550324 217268 550330 217280
rect 550468 217240 550496 217280
rect 551002 217268 551008 217320
rect 551060 217308 551066 217320
rect 557534 217308 557540 217320
rect 551060 217280 557540 217308
rect 551060 217268 551066 217280
rect 557534 217268 557540 217280
rect 557592 217268 557598 217320
rect 558362 217268 558368 217320
rect 558420 217308 558426 217320
rect 562870 217308 562876 217320
rect 558420 217280 562876 217308
rect 558420 217268 558426 217280
rect 562870 217268 562876 217280
rect 562928 217268 562934 217320
rect 563422 217268 563428 217320
rect 563480 217308 563486 217320
rect 570782 217308 570788 217320
rect 563480 217280 570788 217308
rect 563480 217268 563486 217280
rect 570782 217268 570788 217280
rect 570840 217268 570846 217320
rect 571150 217268 571156 217320
rect 571208 217308 571214 217320
rect 571208 217280 572714 217308
rect 571208 217268 571214 217280
rect 550468 217212 550772 217240
rect 535926 217144 545804 217172
rect 535926 217132 535932 217144
rect 547874 217132 547880 217184
rect 547932 217172 547938 217184
rect 547932 217144 548840 217172
rect 547932 217132 547938 217144
rect 520964 217064 520970 217116
rect 521022 217104 521028 217116
rect 546126 217104 546132 217116
rect 521022 217076 524414 217104
rect 521022 217064 521028 217076
rect 524386 217036 524414 217076
rect 545868 217076 546132 217104
rect 545868 217036 545896 217076
rect 546126 217064 546132 217076
rect 546184 217064 546190 217116
rect 548812 217104 548840 217144
rect 549116 217104 549122 217116
rect 548812 217076 549122 217104
rect 549116 217064 549122 217076
rect 549174 217064 549180 217116
rect 549438 217064 549444 217116
rect 549496 217104 549502 217116
rect 550358 217104 550364 217116
rect 549496 217076 550364 217104
rect 549496 217064 549502 217076
rect 550358 217064 550364 217076
rect 550416 217064 550422 217116
rect 524386 217008 545896 217036
rect 550744 217036 550772 217212
rect 550910 217132 550916 217184
rect 550968 217172 550974 217184
rect 551370 217172 551376 217184
rect 550968 217144 551376 217172
rect 550968 217132 550974 217144
rect 551370 217132 551376 217144
rect 551428 217132 551434 217184
rect 551738 217132 551744 217184
rect 551796 217172 551802 217184
rect 571978 217172 571984 217184
rect 551796 217144 571984 217172
rect 551796 217132 551802 217144
rect 571978 217132 571984 217144
rect 572036 217132 572042 217184
rect 572438 217104 572444 217116
rect 572180 217076 572444 217104
rect 572180 217036 572208 217076
rect 572438 217064 572444 217076
rect 572496 217064 572502 217116
rect 550744 217008 572208 217036
rect 572686 217036 572714 217280
rect 573266 217268 573272 217320
rect 573324 217308 573330 217320
rect 604546 217308 604552 217320
rect 573324 217280 604552 217308
rect 573324 217268 573330 217280
rect 604546 217268 604552 217280
rect 604604 217268 604610 217320
rect 607122 217268 607128 217320
rect 607180 217308 607186 217320
rect 616138 217308 616144 217320
rect 607180 217280 616144 217308
rect 607180 217268 607186 217280
rect 616138 217268 616144 217280
rect 616196 217268 616202 217320
rect 573082 217132 573088 217184
rect 573140 217172 573146 217184
rect 574186 217172 574192 217184
rect 573140 217144 574192 217172
rect 573140 217132 573146 217144
rect 574186 217132 574192 217144
rect 574244 217132 574250 217184
rect 575198 217132 575204 217184
rect 575256 217172 575262 217184
rect 603994 217172 604000 217184
rect 575256 217144 578234 217172
rect 575256 217132 575262 217144
rect 578206 217104 578234 217144
rect 579586 217144 604000 217172
rect 579586 217104 579614 217144
rect 603994 217132 604000 217144
rect 604052 217132 604058 217184
rect 578206 217076 579614 217104
rect 572686 217008 576854 217036
rect 576826 216900 576854 217008
rect 582650 216996 582656 217048
rect 582708 217036 582714 217048
rect 590286 217036 590292 217048
rect 582708 217008 590292 217036
rect 582708 216996 582714 217008
rect 590286 216996 590292 217008
rect 590344 216996 590350 217048
rect 591758 216996 591764 217048
rect 591816 217036 591822 217048
rect 592218 217036 592224 217048
rect 591816 217008 592224 217036
rect 591816 216996 591822 217008
rect 592218 216996 592224 217008
rect 592276 216996 592282 217048
rect 592586 216996 592592 217048
rect 592644 217036 592650 217048
rect 614114 217036 614120 217048
rect 592644 217008 614120 217036
rect 592644 216996 592650 217008
rect 614114 216996 614120 217008
rect 614172 216996 614178 217048
rect 576826 216872 582374 216900
rect 582346 216764 582374 216872
rect 582466 216860 582472 216912
rect 582524 216900 582530 216912
rect 590746 216900 590752 216912
rect 582524 216872 590752 216900
rect 582524 216860 582530 216872
rect 590746 216860 590752 216872
rect 590804 216860 590810 216912
rect 593506 216860 593512 216912
rect 593564 216900 593570 216912
rect 605098 216900 605104 216912
rect 593564 216872 605104 216900
rect 593564 216860 593570 216872
rect 605098 216860 605104 216872
rect 605156 216860 605162 216912
rect 605834 216764 605840 216776
rect 582346 216736 605840 216764
rect 605834 216724 605840 216736
rect 605892 216724 605898 216776
rect 574646 216588 574652 216640
rect 574704 216628 574710 216640
rect 582558 216628 582564 216640
rect 574704 216600 582564 216628
rect 574704 216588 574710 216600
rect 582558 216588 582564 216600
rect 582616 216588 582622 216640
rect 591758 216588 591764 216640
rect 591816 216628 591822 216640
rect 595898 216628 595904 216640
rect 591816 216600 595904 216628
rect 591816 216588 591822 216600
rect 595898 216588 595904 216600
rect 595956 216588 595962 216640
rect 576854 216452 576860 216504
rect 576912 216492 576918 216504
rect 582742 216492 582748 216504
rect 576912 216464 582748 216492
rect 576912 216452 576918 216464
rect 582742 216452 582748 216464
rect 582800 216452 582806 216504
rect 592034 216452 592040 216504
rect 592092 216492 592098 216504
rect 596818 216492 596824 216504
rect 592092 216464 596824 216492
rect 592092 216452 592098 216464
rect 596818 216452 596824 216464
rect 596876 216452 596882 216504
rect 582374 216248 582380 216300
rect 582432 216288 582438 216300
rect 592218 216288 592224 216300
rect 582432 216260 592224 216288
rect 582432 216248 582438 216260
rect 592218 216248 592224 216260
rect 592276 216248 592282 216300
rect 590102 216112 590108 216164
rect 590160 216152 590166 216164
rect 597922 216152 597928 216164
rect 590160 216124 597928 216152
rect 590160 216112 590166 216124
rect 597922 216112 597928 216124
rect 597980 216112 597986 216164
rect 590746 215976 590752 216028
rect 590804 216016 590810 216028
rect 596358 216016 596364 216028
rect 590804 215988 596364 216016
rect 590804 215976 590810 215988
rect 596358 215976 596364 215988
rect 596416 215976 596422 216028
rect 599210 215908 599216 215960
rect 599268 215948 599274 215960
rect 613378 215948 613384 215960
rect 599268 215920 613384 215948
rect 599268 215908 599274 215920
rect 613378 215908 613384 215920
rect 613436 215908 613442 215960
rect 652846 215908 652852 215960
rect 652904 215948 652910 215960
rect 654778 215948 654784 215960
rect 652904 215920 654784 215948
rect 652904 215908 652910 215920
rect 654778 215908 654784 215920
rect 654836 215908 654842 215960
rect 590286 215568 590292 215620
rect 590344 215608 590350 215620
rect 598474 215608 598480 215620
rect 590344 215580 598480 215608
rect 590344 215568 590350 215580
rect 598474 215568 598480 215580
rect 598532 215568 598538 215620
rect 613838 215364 613844 215416
rect 613896 215404 613902 215416
rect 615034 215404 615040 215416
rect 613896 215376 615040 215404
rect 613896 215364 613902 215376
rect 615034 215364 615040 215376
rect 615092 215364 615098 215416
rect 636654 215296 636660 215348
rect 636712 215336 636718 215348
rect 639598 215336 639604 215348
rect 636712 215308 639604 215336
rect 636712 215296 636718 215308
rect 639598 215296 639604 215308
rect 639656 215296 639662 215348
rect 575566 215228 575572 215280
rect 575624 215268 575630 215280
rect 621658 215268 621664 215280
rect 575624 215240 621664 215268
rect 575624 215228 575630 215240
rect 621658 215228 621664 215240
rect 621716 215228 621722 215280
rect 574370 215092 574376 215144
rect 574428 215132 574434 215144
rect 619634 215132 619640 215144
rect 574428 215104 619640 215132
rect 574428 215092 574434 215104
rect 619634 215092 619640 215104
rect 619692 215092 619698 215144
rect 675938 215092 675944 215144
rect 675996 215132 676002 215144
rect 677226 215132 677232 215144
rect 675996 215104 677232 215132
rect 675996 215092 676002 215104
rect 677226 215092 677232 215104
rect 677284 215092 677290 215144
rect 577682 214956 577688 215008
rect 577740 214996 577746 215008
rect 626074 214996 626080 215008
rect 577740 214968 626080 214996
rect 577740 214956 577746 214968
rect 626074 214956 626080 214968
rect 626132 214956 626138 215008
rect 576394 214820 576400 214872
rect 576452 214860 576458 214872
rect 622394 214860 622400 214872
rect 576452 214832 622400 214860
rect 576452 214820 576458 214832
rect 622394 214820 622400 214832
rect 622452 214820 622458 214872
rect 574830 214684 574836 214736
rect 574888 214724 574894 214736
rect 616690 214724 616696 214736
rect 574888 214696 616696 214724
rect 574888 214684 574894 214696
rect 616690 214684 616696 214696
rect 616748 214684 616754 214736
rect 616874 214684 616880 214736
rect 616932 214724 616938 214736
rect 617794 214724 617800 214736
rect 616932 214696 617800 214724
rect 616932 214684 616938 214696
rect 617794 214684 617800 214696
rect 617852 214684 617858 214736
rect 624418 214684 624424 214736
rect 624476 214724 624482 214736
rect 633802 214724 633808 214736
rect 624476 214696 633808 214724
rect 624476 214684 624482 214696
rect 633802 214684 633808 214696
rect 633860 214684 633866 214736
rect 577866 214548 577872 214600
rect 577924 214588 577930 214600
rect 577924 214560 625154 214588
rect 577924 214548 577930 214560
rect 575750 214412 575756 214464
rect 575808 214452 575814 214464
rect 620002 214452 620008 214464
rect 575808 214424 620008 214452
rect 575808 214412 575814 214424
rect 620002 214412 620008 214424
rect 620060 214412 620066 214464
rect 625126 214452 625154 214560
rect 626626 214548 626632 214600
rect 626684 214588 626690 214600
rect 627178 214588 627184 214600
rect 626684 214560 627184 214588
rect 626684 214548 626690 214560
rect 627178 214548 627184 214560
rect 627236 214548 627242 214600
rect 628006 214548 628012 214600
rect 628064 214588 628070 214600
rect 628834 214588 628840 214600
rect 628064 214560 628840 214588
rect 628064 214548 628070 214560
rect 628834 214548 628840 214560
rect 628892 214548 628898 214600
rect 630766 214548 630772 214600
rect 630824 214588 630830 214600
rect 631594 214588 631600 214600
rect 630824 214560 631600 214588
rect 630824 214548 630830 214560
rect 631594 214548 631600 214560
rect 631652 214548 631658 214600
rect 628374 214452 628380 214464
rect 625126 214424 628380 214452
rect 628374 214412 628380 214424
rect 628432 214412 628438 214464
rect 600406 214276 600412 214328
rect 600464 214316 600470 214328
rect 600774 214316 600780 214328
rect 600464 214288 600780 214316
rect 600464 214276 600470 214288
rect 600774 214276 600780 214288
rect 600832 214276 600838 214328
rect 607306 214276 607312 214328
rect 607364 214316 607370 214328
rect 607858 214316 607864 214328
rect 607364 214288 607864 214316
rect 607364 214276 607370 214288
rect 607858 214276 607864 214288
rect 607916 214276 607922 214328
rect 608686 214276 608692 214328
rect 608744 214316 608750 214328
rect 609514 214316 609520 214328
rect 608744 214288 609520 214316
rect 608744 214276 608750 214288
rect 609514 214276 609520 214288
rect 609572 214276 609578 214328
rect 616690 214276 616696 214328
rect 616748 214316 616754 214328
rect 624418 214316 624424 214328
rect 616748 214288 624424 214316
rect 616748 214276 616754 214288
rect 624418 214276 624424 214288
rect 624476 214276 624482 214328
rect 658734 214140 658740 214192
rect 658792 214180 658798 214192
rect 661678 214180 661684 214192
rect 658792 214152 661684 214180
rect 658792 214140 658798 214152
rect 661678 214140 661684 214152
rect 661736 214140 661742 214192
rect 662046 214004 662052 214056
rect 662104 214044 662110 214056
rect 665818 214044 665824 214056
rect 662104 214016 665824 214044
rect 662104 214004 662110 214016
rect 665818 214004 665824 214016
rect 665876 214004 665882 214056
rect 35802 213936 35808 213988
rect 35860 213976 35866 213988
rect 40678 213976 40684 213988
rect 35860 213948 40684 213976
rect 35860 213936 35866 213948
rect 40678 213936 40684 213948
rect 40736 213936 40742 213988
rect 675846 213936 675852 213988
rect 675904 213976 675910 213988
rect 676490 213976 676496 213988
rect 675904 213948 676496 213976
rect 675904 213936 675910 213948
rect 676490 213936 676496 213948
rect 676548 213936 676554 213988
rect 626442 213868 626448 213920
rect 626500 213908 626506 213920
rect 629386 213908 629392 213920
rect 626500 213880 629392 213908
rect 626500 213868 626506 213880
rect 629386 213868 629392 213880
rect 629444 213868 629450 213920
rect 638310 213868 638316 213920
rect 638368 213908 638374 213920
rect 640058 213908 640064 213920
rect 638368 213880 640064 213908
rect 638368 213868 638374 213880
rect 640058 213868 640064 213880
rect 640116 213868 640122 213920
rect 648522 213868 648528 213920
rect 648580 213908 648586 213920
rect 650638 213908 650644 213920
rect 648580 213880 650644 213908
rect 648580 213868 648586 213880
rect 650638 213868 650644 213880
rect 650696 213868 650702 213920
rect 655698 213868 655704 213920
rect 655756 213908 655762 213920
rect 656802 213908 656808 213920
rect 655756 213880 656808 213908
rect 655756 213868 655762 213880
rect 656802 213868 656808 213880
rect 656860 213868 656866 213920
rect 660390 213868 660396 213920
rect 660448 213908 660454 213920
rect 660942 213908 660948 213920
rect 660448 213880 660948 213908
rect 660448 213868 660454 213880
rect 660942 213868 660948 213880
rect 661000 213868 661006 213920
rect 651834 213732 651840 213784
rect 651892 213772 651898 213784
rect 657998 213772 658004 213784
rect 651892 213744 658004 213772
rect 651892 213732 651898 213744
rect 657998 213732 658004 213744
rect 658056 213732 658062 213784
rect 660942 213732 660948 213784
rect 661000 213772 661006 213784
rect 662966 213772 662972 213784
rect 661000 213744 662972 213772
rect 661000 213732 661006 213744
rect 662966 213732 662972 213744
rect 663024 213732 663030 213784
rect 663150 213732 663156 213784
rect 663208 213772 663214 213784
rect 664438 213772 664444 213784
rect 663208 213744 664444 213772
rect 663208 213732 663214 213744
rect 664438 213732 664444 213744
rect 664496 213732 664502 213784
rect 576210 213596 576216 213648
rect 576268 213636 576274 213648
rect 601786 213636 601792 213648
rect 576268 213608 601792 213636
rect 576268 213596 576274 213608
rect 601786 213596 601792 213608
rect 601844 213596 601850 213648
rect 645486 213596 645492 213648
rect 645544 213636 645550 213648
rect 659470 213636 659476 213648
rect 645544 213608 659476 213636
rect 645544 213596 645550 213608
rect 659470 213596 659476 213608
rect 659528 213596 659534 213648
rect 574186 213460 574192 213512
rect 574244 213500 574250 213512
rect 601234 213500 601240 213512
rect 574244 213472 601240 213500
rect 574244 213460 574250 213472
rect 601234 213460 601240 213472
rect 601292 213460 601298 213512
rect 639966 213460 639972 213512
rect 640024 213500 640030 213512
rect 642082 213500 642088 213512
rect 640024 213472 642088 213500
rect 640024 213460 640030 213472
rect 642082 213460 642088 213472
rect 642140 213460 642146 213512
rect 650454 213460 650460 213512
rect 650512 213500 650518 213512
rect 650512 213472 654134 213500
rect 650512 213460 650518 213472
rect 575658 213324 575664 213376
rect 575716 213364 575722 213376
rect 612826 213364 612832 213376
rect 575716 213336 612832 213364
rect 575716 213324 575722 213336
rect 612826 213324 612832 213336
rect 612884 213324 612890 213376
rect 635550 213324 635556 213376
rect 635608 213364 635614 213376
rect 652018 213364 652024 213376
rect 635608 213336 652024 213364
rect 635608 213324 635614 213336
rect 652018 213324 652024 213336
rect 652076 213324 652082 213376
rect 654106 213364 654134 213472
rect 666002 213364 666008 213376
rect 654106 213336 666008 213364
rect 666002 213324 666008 213336
rect 666060 213324 666066 213376
rect 575382 213188 575388 213240
rect 575440 213228 575446 213240
rect 623866 213228 623872 213240
rect 575440 213200 623872 213228
rect 575440 213188 575446 213200
rect 623866 213188 623872 213200
rect 623924 213188 623930 213240
rect 641622 213188 641628 213240
rect 641680 213228 641686 213240
rect 658918 213228 658924 213240
rect 641680 213200 658924 213228
rect 641680 213188 641686 213200
rect 658918 213188 658924 213200
rect 658976 213188 658982 213240
rect 654042 212984 654048 213036
rect 654100 213024 654106 213036
rect 654778 213024 654784 213036
rect 654100 212996 654784 213024
rect 654100 212984 654106 212996
rect 654778 212984 654784 212996
rect 654836 212984 654842 213036
rect 664254 212984 664260 213036
rect 664312 213024 664318 213036
rect 665082 213024 665088 213036
rect 664312 212996 665088 213024
rect 664312 212984 664318 212996
rect 665082 212984 665088 212996
rect 665140 212984 665146 213036
rect 632698 212848 632704 212900
rect 632756 212888 632762 212900
rect 634354 212888 634360 212900
rect 632756 212860 634360 212888
rect 632756 212848 632762 212860
rect 634354 212848 634360 212860
rect 634412 212848 634418 212900
rect 628558 212712 628564 212764
rect 628616 212752 628622 212764
rect 632698 212752 632704 212764
rect 628616 212724 632704 212752
rect 628616 212712 628622 212724
rect 632698 212712 632704 212724
rect 632756 212712 632762 212764
rect 637206 212712 637212 212764
rect 637264 212752 637270 212764
rect 641438 212752 641444 212764
rect 637264 212724 641444 212752
rect 637264 212712 637270 212724
rect 641438 212712 641444 212724
rect 641496 212712 641502 212764
rect 578510 211624 578516 211676
rect 578568 211664 578574 211676
rect 580442 211664 580448 211676
rect 578568 211636 580448 211664
rect 578568 211624 578574 211636
rect 580442 211624 580448 211636
rect 580500 211624 580506 211676
rect 35802 211148 35808 211200
rect 35860 211188 35866 211200
rect 41690 211188 41696 211200
rect 35860 211160 41696 211188
rect 35860 211148 35866 211160
rect 41690 211148 41696 211160
rect 41748 211148 41754 211200
rect 579246 209788 579252 209840
rect 579304 209828 579310 209840
rect 581730 209828 581736 209840
rect 579304 209800 581736 209828
rect 579304 209788 579310 209800
rect 581730 209788 581736 209800
rect 581788 209788 581794 209840
rect 632146 209556 632152 209568
rect 625126 209528 632152 209556
rect 581546 208564 581552 208616
rect 581604 208604 581610 208616
rect 625126 208604 625154 209528
rect 632146 209516 632152 209528
rect 632204 209516 632210 209568
rect 652202 209516 652208 209568
rect 652260 209556 652266 209568
rect 652260 209528 654134 209556
rect 652260 209516 652266 209528
rect 654106 209080 654134 209528
rect 666830 209080 666836 209092
rect 654106 209052 666836 209080
rect 666830 209040 666836 209052
rect 666888 209040 666894 209092
rect 581604 208576 625154 208604
rect 581604 208564 581610 208576
rect 35802 208360 35808 208412
rect 35860 208400 35866 208412
rect 40034 208400 40040 208412
rect 35860 208372 40040 208400
rect 35860 208360 35866 208372
rect 40034 208360 40040 208372
rect 40092 208360 40098 208412
rect 578878 208292 578884 208344
rect 578936 208332 578942 208344
rect 589458 208332 589464 208344
rect 578936 208304 589464 208332
rect 578936 208292 578942 208304
rect 589458 208292 589464 208304
rect 589516 208292 589522 208344
rect 580442 207612 580448 207664
rect 580500 207652 580506 207664
rect 589458 207652 589464 207664
rect 580500 207624 589464 207652
rect 580500 207612 580506 207624
rect 589458 207612 589464 207624
rect 589516 207612 589522 207664
rect 581730 206252 581736 206304
rect 581788 206292 581794 206304
rect 589642 206292 589648 206304
rect 581788 206264 589648 206292
rect 581788 206252 581794 206264
rect 589642 206252 589648 206264
rect 589700 206252 589706 206304
rect 579522 205776 579528 205828
rect 579580 205816 579586 205828
rect 580994 205816 581000 205828
rect 579580 205788 581000 205816
rect 579580 205776 579586 205788
rect 580994 205776 581000 205788
rect 581052 205776 581058 205828
rect 579706 204212 579712 204264
rect 579764 204252 579770 204264
rect 589458 204252 589464 204264
rect 579764 204224 589464 204252
rect 579764 204212 579770 204224
rect 589458 204212 589464 204224
rect 589516 204212 589522 204264
rect 35802 202852 35808 202904
rect 35860 202892 35866 202904
rect 37918 202892 37924 202904
rect 35860 202864 37924 202892
rect 35860 202852 35866 202864
rect 37918 202852 37924 202864
rect 37976 202852 37982 202904
rect 578326 202852 578332 202904
rect 578384 202892 578390 202904
rect 580258 202892 580264 202904
rect 578384 202864 580264 202892
rect 578384 202852 578390 202864
rect 580258 202852 580264 202864
rect 580316 202852 580322 202904
rect 580994 202784 581000 202836
rect 581052 202824 581058 202836
rect 589458 202824 589464 202836
rect 581052 202796 589464 202824
rect 581052 202784 581058 202796
rect 589458 202784 589464 202796
rect 589516 202784 589522 202836
rect 578786 200132 578792 200184
rect 578844 200172 578850 200184
rect 590378 200172 590384 200184
rect 578844 200144 590384 200172
rect 578844 200132 578850 200144
rect 590378 200132 590384 200144
rect 590436 200132 590442 200184
rect 580258 199996 580264 200048
rect 580316 200036 580322 200048
rect 589458 200036 589464 200048
rect 580316 200008 589464 200036
rect 580316 199996 580322 200008
rect 589458 199996 589464 200008
rect 589516 199996 589522 200048
rect 669130 199316 669136 199368
rect 669188 199356 669194 199368
rect 670786 199356 670792 199368
rect 669188 199328 670792 199356
rect 669188 199316 669194 199328
rect 670786 199316 670792 199328
rect 670844 199316 670850 199368
rect 579522 198704 579528 198756
rect 579580 198744 579586 198756
rect 589458 198744 589464 198756
rect 579580 198716 589464 198744
rect 579580 198704 579586 198716
rect 589458 198704 589464 198716
rect 589516 198704 589522 198756
rect 578510 195984 578516 196036
rect 578568 196024 578574 196036
rect 589274 196024 589280 196036
rect 578568 195996 589280 196024
rect 578568 195984 578574 195996
rect 589274 195984 589280 195996
rect 589332 195984 589338 196036
rect 579522 194556 579528 194608
rect 579580 194596 579586 194608
rect 589458 194596 589464 194608
rect 579580 194568 589464 194596
rect 579580 194556 579586 194568
rect 589458 194556 589464 194568
rect 589516 194556 589522 194608
rect 669130 194284 669136 194336
rect 669188 194324 669194 194336
rect 670786 194324 670792 194336
rect 669188 194296 670792 194324
rect 669188 194284 669194 194296
rect 670786 194284 670792 194296
rect 670844 194284 670850 194336
rect 579522 191836 579528 191888
rect 579580 191876 579586 191888
rect 589458 191876 589464 191888
rect 579580 191848 589464 191876
rect 579580 191836 579586 191848
rect 589458 191836 589464 191848
rect 589516 191836 589522 191888
rect 579522 190476 579528 190528
rect 579580 190516 579586 190528
rect 590562 190516 590568 190528
rect 579580 190488 590568 190516
rect 579580 190476 579586 190488
rect 590562 190476 590568 190488
rect 590620 190476 590626 190528
rect 667934 189388 667940 189440
rect 667992 189428 667998 189440
rect 670786 189428 670792 189440
rect 667992 189400 670792 189428
rect 667992 189388 667998 189400
rect 670786 189388 670792 189400
rect 670844 189388 670850 189440
rect 579522 187688 579528 187740
rect 579580 187728 579586 187740
rect 589458 187728 589464 187740
rect 579580 187700 589464 187728
rect 579580 187688 579586 187700
rect 589458 187688 589464 187700
rect 589516 187688 589522 187740
rect 579522 186260 579528 186312
rect 579580 186300 579586 186312
rect 589642 186300 589648 186312
rect 579580 186272 589648 186300
rect 579580 186260 579586 186272
rect 589642 186260 589648 186272
rect 589700 186260 589706 186312
rect 579522 184832 579528 184884
rect 579580 184872 579586 184884
rect 589458 184872 589464 184884
rect 579580 184844 589464 184872
rect 579580 184832 579586 184844
rect 589458 184832 589464 184844
rect 589516 184832 589522 184884
rect 579522 182112 579528 182164
rect 579580 182152 579586 182164
rect 589458 182152 589464 182164
rect 579580 182124 589464 182152
rect 579580 182112 579586 182124
rect 589458 182112 589464 182124
rect 589516 182112 589522 182164
rect 578786 180752 578792 180804
rect 578844 180792 578850 180804
rect 590562 180792 590568 180804
rect 578844 180764 590568 180792
rect 578844 180752 578850 180764
rect 590562 180752 590568 180764
rect 590620 180752 590626 180804
rect 578786 178032 578792 178084
rect 578844 178072 578850 178084
rect 589458 178072 589464 178084
rect 578844 178044 589464 178072
rect 578844 178032 578850 178044
rect 589458 178032 589464 178044
rect 589516 178032 589522 178084
rect 579522 177896 579528 177948
rect 579580 177936 579586 177948
rect 589642 177936 589648 177948
rect 579580 177908 589648 177936
rect 579580 177896 579586 177908
rect 589642 177896 589648 177908
rect 589700 177896 589706 177948
rect 589458 175352 589464 175364
rect 586486 175324 589464 175352
rect 579982 175244 579988 175296
rect 580040 175284 580046 175296
rect 586486 175284 586514 175324
rect 589458 175312 589464 175324
rect 589516 175312 589522 175364
rect 580040 175256 586514 175284
rect 580040 175244 580046 175256
rect 667934 174700 667940 174752
rect 667992 174740 667998 174752
rect 669774 174740 669780 174752
rect 667992 174712 669780 174740
rect 667992 174700 667998 174712
rect 669774 174700 669780 174712
rect 669832 174700 669838 174752
rect 578418 174496 578424 174548
rect 578476 174536 578482 174548
rect 589642 174536 589648 174548
rect 578476 174508 589648 174536
rect 578476 174496 578482 174508
rect 589642 174496 589648 174508
rect 589700 174496 589706 174548
rect 578234 172864 578240 172916
rect 578292 172904 578298 172916
rect 579982 172904 579988 172916
rect 578292 172876 579988 172904
rect 578292 172864 578298 172876
rect 579982 172864 579988 172876
rect 580040 172864 580046 172916
rect 580902 172524 580908 172576
rect 580960 172564 580966 172576
rect 589458 172564 589464 172576
rect 580960 172536 589464 172564
rect 580960 172524 580966 172536
rect 589458 172524 589464 172536
rect 589516 172524 589522 172576
rect 579890 171096 579896 171148
rect 579948 171136 579954 171148
rect 589458 171136 589464 171148
rect 579948 171108 589464 171136
rect 579948 171096 579954 171108
rect 589458 171096 589464 171108
rect 589516 171096 589522 171148
rect 578694 169736 578700 169788
rect 578752 169776 578758 169788
rect 580902 169776 580908 169788
rect 578752 169748 580908 169776
rect 578752 169736 578758 169748
rect 580902 169736 580908 169748
rect 580960 169736 580966 169788
rect 582374 169736 582380 169788
rect 582432 169776 582438 169788
rect 589458 169776 589464 169788
rect 582432 169748 589464 169776
rect 582432 169736 582438 169748
rect 589458 169736 589464 169748
rect 589516 169736 589522 169788
rect 668026 169668 668032 169720
rect 668084 169708 668090 169720
rect 670326 169708 670332 169720
rect 668084 169680 670332 169708
rect 668084 169668 668090 169680
rect 670326 169668 670332 169680
rect 670384 169668 670390 169720
rect 579706 168376 579712 168428
rect 579764 168416 579770 168428
rect 589458 168416 589464 168428
rect 579764 168388 589464 168416
rect 579764 168376 579770 168388
rect 589458 168376 589464 168388
rect 589516 168376 589522 168428
rect 583754 167016 583760 167068
rect 583812 167056 583818 167068
rect 589458 167056 589464 167068
rect 583812 167028 589464 167056
rect 583812 167016 583818 167028
rect 589458 167016 589464 167028
rect 589516 167016 589522 167068
rect 578878 165520 578884 165572
rect 578936 165560 578942 165572
rect 582374 165560 582380 165572
rect 578936 165532 582380 165560
rect 578936 165520 578942 165532
rect 582374 165520 582380 165532
rect 582432 165520 582438 165572
rect 667934 164908 667940 164960
rect 667992 164948 667998 164960
rect 670142 164948 670148 164960
rect 667992 164920 670148 164948
rect 667992 164908 667998 164920
rect 670142 164908 670148 164920
rect 670200 164908 670206 164960
rect 582466 164228 582472 164280
rect 582524 164268 582530 164280
rect 589458 164268 589464 164280
rect 582524 164240 589464 164268
rect 582524 164228 582530 164240
rect 589458 164228 589464 164240
rect 589516 164228 589522 164280
rect 580902 162868 580908 162920
rect 580960 162908 580966 162920
rect 589458 162908 589464 162920
rect 580960 162880 589464 162908
rect 580960 162868 580966 162880
rect 589458 162868 589464 162880
rect 589516 162868 589522 162920
rect 676122 162800 676128 162852
rect 676180 162840 676186 162852
rect 678238 162840 678244 162852
rect 676180 162812 678244 162840
rect 676180 162800 676186 162812
rect 678238 162800 678244 162812
rect 678296 162800 678302 162852
rect 578418 162664 578424 162716
rect 578476 162704 578482 162716
rect 582466 162704 582472 162716
rect 578476 162676 582472 162704
rect 578476 162664 578482 162676
rect 582466 162664 582472 162676
rect 582524 162664 582530 162716
rect 675938 162596 675944 162648
rect 675996 162636 676002 162648
rect 679618 162636 679624 162648
rect 675996 162608 679624 162636
rect 675996 162596 676002 162608
rect 679618 162596 679624 162608
rect 679676 162596 679682 162648
rect 578234 162528 578240 162580
rect 578292 162568 578298 162580
rect 583754 162568 583760 162580
rect 578292 162540 583760 162568
rect 578292 162528 578298 162540
rect 583754 162528 583760 162540
rect 583812 162528 583818 162580
rect 675846 161712 675852 161764
rect 675904 161752 675910 161764
rect 680998 161752 681004 161764
rect 675904 161724 681004 161752
rect 675904 161712 675910 161724
rect 680998 161712 681004 161724
rect 681056 161712 681062 161764
rect 580534 161440 580540 161492
rect 580592 161480 580598 161492
rect 589458 161480 589464 161492
rect 580592 161452 589464 161480
rect 580592 161440 580598 161452
rect 589458 161440 589464 161452
rect 589516 161440 589522 161492
rect 580718 160080 580724 160132
rect 580776 160120 580782 160132
rect 589458 160120 589464 160132
rect 580776 160092 589464 160120
rect 580776 160080 580782 160092
rect 589458 160080 589464 160092
rect 589516 160080 589522 160132
rect 578878 158720 578884 158772
rect 578936 158760 578942 158772
rect 580902 158760 580908 158772
rect 578936 158732 580908 158760
rect 578936 158720 578942 158732
rect 580902 158720 580908 158732
rect 580960 158720 580966 158772
rect 587158 158720 587164 158772
rect 587216 158760 587222 158772
rect 589826 158760 589832 158772
rect 587216 158732 589832 158760
rect 587216 158720 587222 158732
rect 589826 158720 589832 158732
rect 589884 158720 589890 158772
rect 585778 157360 585784 157412
rect 585836 157400 585842 157412
rect 589458 157400 589464 157412
rect 585836 157372 589464 157400
rect 585836 157360 585842 157372
rect 589458 157360 589464 157372
rect 589516 157360 589522 157412
rect 578326 154640 578332 154692
rect 578384 154680 578390 154692
rect 580534 154680 580540 154692
rect 578384 154652 580540 154680
rect 578384 154640 578390 154652
rect 580534 154640 580540 154652
rect 580592 154640 580598 154692
rect 584398 154572 584404 154624
rect 584456 154612 584462 154624
rect 589458 154612 589464 154624
rect 584456 154584 589464 154612
rect 584456 154572 584462 154584
rect 589458 154572 589464 154584
rect 589516 154572 589522 154624
rect 583018 153212 583024 153264
rect 583076 153252 583082 153264
rect 589458 153252 589464 153264
rect 583076 153224 589464 153252
rect 583076 153212 583082 153224
rect 589458 153212 589464 153224
rect 589516 153212 589522 153264
rect 578234 152736 578240 152788
rect 578292 152776 578298 152788
rect 580718 152776 580724 152788
rect 578292 152748 580724 152776
rect 578292 152736 578298 152748
rect 580718 152736 580724 152748
rect 580776 152736 580782 152788
rect 580442 151784 580448 151836
rect 580500 151824 580506 151836
rect 589458 151824 589464 151836
rect 580500 151796 589464 151824
rect 580500 151784 580506 151796
rect 589458 151784 589464 151796
rect 589516 151784 589522 151836
rect 578326 151036 578332 151088
rect 578384 151076 578390 151088
rect 587158 151076 587164 151088
rect 578384 151048 587164 151076
rect 578384 151036 578390 151048
rect 587158 151036 587164 151048
rect 587216 151036 587222 151088
rect 578878 149064 578884 149116
rect 578936 149104 578942 149116
rect 589458 149104 589464 149116
rect 578936 149076 589464 149104
rect 578936 149064 578942 149076
rect 589458 149064 589464 149076
rect 589516 149064 589522 149116
rect 578694 147228 578700 147280
rect 578752 147268 578758 147280
rect 585778 147268 585784 147280
rect 578752 147240 585784 147268
rect 578752 147228 578758 147240
rect 585778 147228 585784 147240
rect 585836 147228 585842 147280
rect 668578 145528 668584 145580
rect 668636 145568 668642 145580
rect 670786 145568 670792 145580
rect 668636 145540 670792 145568
rect 668636 145528 668642 145540
rect 670786 145528 670792 145540
rect 670844 145528 670850 145580
rect 585962 144916 585968 144968
rect 586020 144956 586026 144968
rect 589458 144956 589464 144968
rect 586020 144928 589464 144956
rect 586020 144916 586026 144928
rect 589458 144916 589464 144928
rect 589516 144916 589522 144968
rect 579246 144644 579252 144696
rect 579304 144684 579310 144696
rect 584398 144684 584404 144696
rect 579304 144656 584404 144684
rect 579304 144644 579310 144656
rect 584398 144644 584404 144656
rect 584456 144644 584462 144696
rect 584582 143556 584588 143608
rect 584640 143596 584646 143608
rect 589458 143596 589464 143608
rect 584640 143568 589464 143596
rect 584640 143556 584646 143568
rect 589458 143556 589464 143568
rect 589516 143556 589522 143608
rect 579522 143420 579528 143472
rect 579580 143460 579586 143472
rect 583018 143460 583024 143472
rect 579580 143432 583024 143460
rect 579580 143420 579586 143432
rect 583018 143420 583024 143432
rect 583076 143420 583082 143472
rect 587158 142400 587164 142452
rect 587216 142440 587222 142452
rect 589826 142440 589832 142452
rect 587216 142412 589832 142440
rect 587216 142400 587222 142412
rect 589826 142400 589832 142412
rect 589884 142400 589890 142452
rect 583018 140768 583024 140820
rect 583076 140808 583082 140820
rect 589458 140808 589464 140820
rect 583076 140780 589464 140808
rect 583076 140768 583082 140780
rect 589458 140768 589464 140780
rect 589516 140768 589522 140820
rect 578602 140700 578608 140752
rect 578660 140740 578666 140752
rect 580442 140740 580448 140752
rect 578660 140712 580448 140740
rect 578660 140700 578666 140712
rect 580442 140700 580448 140712
rect 580500 140700 580506 140752
rect 580258 139408 580264 139460
rect 580316 139448 580322 139460
rect 589458 139448 589464 139460
rect 580316 139420 589464 139448
rect 580316 139408 580322 139420
rect 589458 139408 589464 139420
rect 589516 139408 589522 139460
rect 578602 139272 578608 139324
rect 578660 139312 578666 139324
rect 589918 139312 589924 139324
rect 578660 139284 589924 139312
rect 578660 139272 578666 139284
rect 589918 139272 589924 139284
rect 589976 139272 589982 139324
rect 578694 137232 578700 137284
rect 578752 137272 578758 137284
rect 588538 137272 588544 137284
rect 578752 137244 588544 137272
rect 578752 137232 578758 137244
rect 588538 137232 588544 137244
rect 588596 137232 588602 137284
rect 579062 137096 579068 137148
rect 579120 137136 579126 137148
rect 585962 137136 585968 137148
rect 579120 137108 585968 137136
rect 579120 137096 579126 137108
rect 585962 137096 585968 137108
rect 586020 137096 586026 137148
rect 585778 136620 585784 136672
rect 585836 136660 585842 136672
rect 589458 136660 589464 136672
rect 585836 136632 589464 136660
rect 585836 136620 585842 136632
rect 589458 136620 589464 136632
rect 589516 136620 589522 136672
rect 667934 136348 667940 136400
rect 667992 136388 667998 136400
rect 669958 136388 669964 136400
rect 667992 136360 669964 136388
rect 667992 136348 667998 136360
rect 669958 136348 669964 136360
rect 670016 136348 670022 136400
rect 584398 135260 584404 135312
rect 584456 135300 584462 135312
rect 589458 135300 589464 135312
rect 584456 135272 589464 135300
rect 584456 135260 584462 135272
rect 589458 135260 589464 135272
rect 589516 135260 589522 135312
rect 675846 133900 675852 133952
rect 675904 133940 675910 133952
rect 676490 133940 676496 133952
rect 675904 133912 676496 133940
rect 675904 133900 675910 133912
rect 676490 133900 676496 133912
rect 676548 133900 676554 133952
rect 580626 131724 580632 131776
rect 580684 131764 580690 131776
rect 590286 131764 590292 131776
rect 580684 131736 590292 131764
rect 580684 131724 580690 131736
rect 590286 131724 590292 131736
rect 590344 131724 590350 131776
rect 578878 131248 578884 131300
rect 578936 131288 578942 131300
rect 589458 131288 589464 131300
rect 578936 131260 589464 131288
rect 578936 131248 578942 131260
rect 589458 131248 589464 131260
rect 589516 131248 589522 131300
rect 579062 131112 579068 131164
rect 579120 131152 579126 131164
rect 584582 131152 584588 131164
rect 579120 131124 584588 131152
rect 579120 131112 579126 131124
rect 584582 131112 584588 131124
rect 584640 131112 584646 131164
rect 579154 128256 579160 128308
rect 579212 128296 579218 128308
rect 587158 128296 587164 128308
rect 579212 128268 587164 128296
rect 579212 128256 579218 128268
rect 587158 128256 587164 128268
rect 587216 128256 587222 128308
rect 587618 127168 587624 127220
rect 587676 127208 587682 127220
rect 589458 127208 589464 127220
rect 587676 127180 589464 127208
rect 587676 127168 587682 127180
rect 589458 127168 589464 127180
rect 589516 127168 589522 127220
rect 579062 126216 579068 126268
rect 579120 126256 579126 126268
rect 587618 126256 587624 126268
rect 579120 126228 587624 126256
rect 579120 126216 579126 126228
rect 587618 126216 587624 126228
rect 587676 126216 587682 126268
rect 667934 125536 667940 125588
rect 667992 125576 667998 125588
rect 669774 125576 669780 125588
rect 667992 125548 669780 125576
rect 667992 125536 667998 125548
rect 669774 125536 669780 125548
rect 669832 125536 669838 125588
rect 579522 125332 579528 125384
rect 579580 125372 579586 125384
rect 583018 125372 583024 125384
rect 579580 125344 583024 125372
rect 579580 125332 579586 125344
rect 583018 125332 583024 125344
rect 583076 125332 583082 125384
rect 583202 124856 583208 124908
rect 583260 124896 583266 124908
rect 589642 124896 589648 124908
rect 583260 124868 589648 124896
rect 583260 124856 583266 124868
rect 589642 124856 589648 124868
rect 589700 124856 589706 124908
rect 578326 124108 578332 124160
rect 578384 124148 578390 124160
rect 580258 124148 580264 124160
rect 578384 124120 580264 124148
rect 578384 124108 578390 124120
rect 580258 124108 580264 124120
rect 580316 124108 580322 124160
rect 580442 122816 580448 122868
rect 580500 122856 580506 122868
rect 589458 122856 589464 122868
rect 580500 122828 589464 122856
rect 580500 122816 580506 122828
rect 589458 122816 589464 122828
rect 589516 122816 589522 122868
rect 581822 122068 581828 122120
rect 581880 122108 581886 122120
rect 590102 122108 590108 122120
rect 581880 122080 590108 122108
rect 581880 122068 581886 122080
rect 590102 122068 590108 122080
rect 590160 122068 590166 122120
rect 587342 121456 587348 121508
rect 587400 121496 587406 121508
rect 589274 121496 589280 121508
rect 587400 121468 589280 121496
rect 587400 121456 587406 121468
rect 589274 121456 589280 121468
rect 589332 121456 589338 121508
rect 579522 121388 579528 121440
rect 579580 121428 579586 121440
rect 585778 121428 585784 121440
rect 579580 121400 585784 121428
rect 579580 121388 579586 121400
rect 585778 121388 585784 121400
rect 585836 121388 585842 121440
rect 584582 118668 584588 118720
rect 584640 118708 584646 118720
rect 589458 118708 589464 118720
rect 584640 118680 589464 118708
rect 584640 118668 584646 118680
rect 589458 118668 589464 118680
rect 589516 118668 589522 118720
rect 578694 118532 578700 118584
rect 578752 118572 578758 118584
rect 584398 118572 584404 118584
rect 578752 118544 584404 118572
rect 578752 118532 578758 118544
rect 584398 118532 584404 118544
rect 584456 118532 584462 118584
rect 668026 118464 668032 118516
rect 668084 118504 668090 118516
rect 670326 118504 670332 118516
rect 668084 118476 670332 118504
rect 668084 118464 668090 118476
rect 670326 118464 670332 118476
rect 670384 118464 670390 118516
rect 585962 117308 585968 117360
rect 586020 117348 586026 117360
rect 589458 117348 589464 117360
rect 586020 117320 589464 117348
rect 586020 117308 586026 117320
rect 589458 117308 589464 117320
rect 589516 117308 589522 117360
rect 675846 117240 675852 117292
rect 675904 117280 675910 117292
rect 682378 117280 682384 117292
rect 675904 117252 682384 117280
rect 675904 117240 675910 117252
rect 682378 117240 682384 117252
rect 682436 117240 682442 117292
rect 578694 117172 578700 117224
rect 578752 117212 578758 117224
rect 580626 117212 580632 117224
rect 578752 117184 580632 117212
rect 578752 117172 578758 117184
rect 580626 117172 580632 117184
rect 580684 117172 580690 117224
rect 585778 115948 585784 116000
rect 585836 115988 585842 116000
rect 589458 115988 589464 116000
rect 585836 115960 589464 115988
rect 585836 115948 585842 115960
rect 589458 115948 589464 115960
rect 589516 115948 589522 116000
rect 579246 114452 579252 114504
rect 579304 114492 579310 114504
rect 581638 114492 581644 114504
rect 579304 114464 581644 114492
rect 579304 114452 579310 114464
rect 581638 114452 581644 114464
rect 581696 114452 581702 114504
rect 668118 114112 668124 114164
rect 668176 114152 668182 114164
rect 669958 114152 669964 114164
rect 668176 114124 669964 114152
rect 668176 114112 668182 114124
rect 669958 114112 669964 114124
rect 670016 114112 670022 114164
rect 584398 113160 584404 113212
rect 584456 113200 584462 113212
rect 589458 113200 589464 113212
rect 584456 113172 589464 113200
rect 584456 113160 584462 113172
rect 589458 113160 589464 113172
rect 589516 113160 589522 113212
rect 579154 113024 579160 113076
rect 579212 113064 579218 113076
rect 588722 113064 588728 113076
rect 579212 113036 588728 113064
rect 579212 113024 579218 113036
rect 588722 113024 588728 113036
rect 588780 113024 588786 113076
rect 581638 111052 581644 111104
rect 581696 111092 581702 111104
rect 589918 111092 589924 111104
rect 581696 111064 589924 111092
rect 581696 111052 581702 111064
rect 589918 111052 589924 111064
rect 589976 111052 589982 111104
rect 583018 109692 583024 109744
rect 583076 109732 583082 109744
rect 589366 109732 589372 109744
rect 583076 109704 589372 109732
rect 583076 109692 583082 109704
rect 589366 109692 589372 109704
rect 589424 109692 589430 109744
rect 578878 108944 578884 108996
rect 578936 108984 578942 108996
rect 581822 108984 581828 108996
rect 578936 108956 581828 108984
rect 578936 108944 578942 108956
rect 581822 108944 581828 108956
rect 581880 108944 581886 108996
rect 589458 107692 589464 107704
rect 581012 107664 589464 107692
rect 578878 107584 578884 107636
rect 578936 107624 578942 107636
rect 581012 107624 581040 107664
rect 589458 107652 589464 107664
rect 589516 107652 589522 107704
rect 578936 107596 581040 107624
rect 578936 107584 578942 107596
rect 581822 106292 581828 106344
rect 581880 106332 581886 106344
rect 589458 106332 589464 106344
rect 581880 106304 589464 106332
rect 581880 106292 581886 106304
rect 589458 106292 589464 106304
rect 589516 106292 589522 106344
rect 668394 106156 668400 106208
rect 668452 106196 668458 106208
rect 670786 106196 670792 106208
rect 668452 106168 670792 106196
rect 668452 106156 668458 106168
rect 670786 106156 670792 106168
rect 670844 106156 670850 106208
rect 580258 104864 580264 104916
rect 580316 104904 580322 104916
rect 589458 104904 589464 104916
rect 580316 104876 589464 104904
rect 580316 104864 580322 104876
rect 589458 104864 589464 104876
rect 589516 104864 589522 104916
rect 578326 103300 578332 103352
rect 578384 103340 578390 103352
rect 583202 103340 583208 103352
rect 578384 103312 583208 103340
rect 578384 103300 578390 103312
rect 583202 103300 583208 103312
rect 583260 103300 583266 103352
rect 578510 102076 578516 102128
rect 578568 102116 578574 102128
rect 580442 102116 580448 102128
rect 578568 102088 580448 102116
rect 578568 102076 578574 102088
rect 580442 102076 580448 102088
rect 580500 102076 580506 102128
rect 587158 100716 587164 100768
rect 587216 100756 587222 100768
rect 589550 100756 589556 100768
rect 587216 100728 589556 100756
rect 587216 100716 587222 100728
rect 589550 100716 589556 100728
rect 589608 100716 589614 100768
rect 624786 100104 624792 100156
rect 624844 100144 624850 100156
rect 668118 100144 668124 100156
rect 624844 100116 668124 100144
rect 624844 100104 624850 100116
rect 668118 100104 668124 100116
rect 668176 100104 668182 100156
rect 580442 99968 580448 100020
rect 580500 100008 580506 100020
rect 590102 100008 590108 100020
rect 580500 99980 590108 100008
rect 580500 99968 580506 99980
rect 590102 99968 590108 99980
rect 590160 99968 590166 100020
rect 667934 100008 667940 100020
rect 615466 99980 667940 100008
rect 614850 99900 614856 99952
rect 614908 99940 614914 99952
rect 615466 99940 615494 99980
rect 667934 99968 667940 99980
rect 667992 99968 667998 100020
rect 614908 99912 615494 99940
rect 614908 99900 614914 99912
rect 622302 99288 622308 99340
rect 622360 99328 622366 99340
rect 630766 99328 630772 99340
rect 622360 99300 630772 99328
rect 622360 99288 622366 99300
rect 630766 99288 630772 99300
rect 630824 99288 630830 99340
rect 579246 99220 579252 99272
rect 579304 99260 579310 99272
rect 581638 99260 581644 99272
rect 579304 99232 581644 99260
rect 579304 99220 579310 99232
rect 581638 99220 581644 99232
rect 581696 99220 581702 99272
rect 623682 99152 623688 99204
rect 623740 99192 623746 99204
rect 633434 99192 633440 99204
rect 623740 99164 633440 99192
rect 623740 99152 623746 99164
rect 633434 99152 633440 99164
rect 633492 99152 633498 99204
rect 577498 99084 577504 99136
rect 577556 99124 577562 99136
rect 595254 99124 595260 99136
rect 577556 99096 595260 99124
rect 577556 99084 577562 99096
rect 595254 99084 595260 99096
rect 595312 99084 595318 99136
rect 625062 99016 625068 99068
rect 625120 99056 625126 99068
rect 636286 99056 636292 99068
rect 625120 99028 636292 99056
rect 625120 99016 625126 99028
rect 636286 99016 636292 99028
rect 636344 99016 636350 99068
rect 629018 98880 629024 98932
rect 629076 98920 629082 98932
rect 643646 98920 643652 98932
rect 629076 98892 643652 98920
rect 629076 98880 629082 98892
rect 643646 98880 643652 98892
rect 643704 98880 643710 98932
rect 629754 98744 629760 98796
rect 629812 98784 629818 98796
rect 645118 98784 645124 98796
rect 629812 98756 645124 98784
rect 629812 98744 629818 98756
rect 645118 98744 645124 98756
rect 645176 98744 645182 98796
rect 630490 98608 630496 98660
rect 630548 98648 630554 98660
rect 646590 98648 646596 98660
rect 630548 98620 646596 98648
rect 630548 98608 630554 98620
rect 646590 98608 646596 98620
rect 646648 98608 646654 98660
rect 642174 98172 642180 98184
rect 631428 98144 642180 98172
rect 578326 97928 578332 97980
rect 578384 97968 578390 97980
rect 587342 97968 587348 97980
rect 578384 97940 587348 97968
rect 578384 97928 578390 97940
rect 587342 97928 587348 97940
rect 587400 97928 587406 97980
rect 605466 97928 605472 97980
rect 605524 97968 605530 97980
rect 606478 97968 606484 97980
rect 605524 97940 606484 97968
rect 605524 97928 605530 97940
rect 606478 97928 606484 97940
rect 606536 97928 606542 97980
rect 618714 97928 618720 97980
rect 618772 97968 618778 97980
rect 625798 97968 625804 97980
rect 618772 97940 625804 97968
rect 618772 97928 618778 97940
rect 625798 97928 625804 97940
rect 625856 97928 625862 97980
rect 628282 97928 628288 97980
rect 628340 97968 628346 97980
rect 631428 97968 631456 98144
rect 642174 98132 642180 98144
rect 642232 98132 642238 98184
rect 640702 98036 640708 98048
rect 628340 97940 631456 97968
rect 631520 98008 640708 98036
rect 628340 97928 628346 97940
rect 627546 97792 627552 97844
rect 627604 97832 627610 97844
rect 631520 97832 631548 98008
rect 640702 97996 640708 98008
rect 640760 97996 640766 98048
rect 650730 97968 650736 97980
rect 645136 97940 650736 97968
rect 627604 97804 631548 97832
rect 627604 97792 627610 97804
rect 634170 97792 634176 97844
rect 634228 97832 634234 97844
rect 645136 97832 645164 97940
rect 650730 97928 650736 97940
rect 650788 97928 650794 97980
rect 655422 97928 655428 97980
rect 655480 97968 655486 97980
rect 662506 97968 662512 97980
rect 655480 97940 662512 97968
rect 655480 97928 655486 97940
rect 662506 97928 662512 97940
rect 662564 97928 662570 97980
rect 634228 97804 645164 97832
rect 634228 97792 634234 97804
rect 647142 97792 647148 97844
rect 647200 97832 647206 97844
rect 659010 97832 659016 97844
rect 647200 97804 659016 97832
rect 647200 97792 647206 97804
rect 659010 97792 659016 97804
rect 659068 97792 659074 97844
rect 659194 97792 659200 97844
rect 659252 97832 659258 97844
rect 663886 97832 663892 97844
rect 659252 97804 663892 97832
rect 659252 97792 659258 97804
rect 663886 97792 663892 97804
rect 663944 97792 663950 97844
rect 621658 97656 621664 97708
rect 621716 97696 621722 97708
rect 629294 97696 629300 97708
rect 621716 97668 629300 97696
rect 621716 97656 621722 97668
rect 629294 97656 629300 97668
rect 629352 97656 629358 97708
rect 631962 97656 631968 97708
rect 632020 97696 632026 97708
rect 648614 97696 648620 97708
rect 632020 97668 648620 97696
rect 632020 97656 632026 97668
rect 648614 97656 648620 97668
rect 648672 97656 648678 97708
rect 653950 97656 653956 97708
rect 654008 97696 654014 97708
rect 655054 97696 655060 97708
rect 654008 97668 655060 97696
rect 654008 97656 654014 97668
rect 655054 97656 655060 97668
rect 655112 97656 655118 97708
rect 659930 97656 659936 97708
rect 659988 97696 659994 97708
rect 665358 97696 665364 97708
rect 659988 97668 665364 97696
rect 659988 97656 659994 97668
rect 665358 97656 665364 97668
rect 665416 97656 665422 97708
rect 659746 97628 659752 97640
rect 657418 97600 659752 97628
rect 626074 97520 626080 97572
rect 626132 97560 626138 97572
rect 637758 97560 637764 97572
rect 626132 97532 637764 97560
rect 626132 97520 626138 97532
rect 637758 97520 637764 97532
rect 637816 97520 637822 97572
rect 639046 97520 639052 97572
rect 639104 97560 639110 97572
rect 639104 97532 640012 97560
rect 639104 97520 639110 97532
rect 613562 97384 613568 97436
rect 613620 97424 613626 97436
rect 618898 97424 618904 97436
rect 613620 97396 618904 97424
rect 613620 97384 613626 97396
rect 618898 97384 618904 97396
rect 618956 97384 618962 97436
rect 620186 97384 620192 97436
rect 620244 97424 620250 97436
rect 625982 97424 625988 97436
rect 620244 97396 625988 97424
rect 620244 97384 620250 97396
rect 625982 97384 625988 97396
rect 626040 97384 626046 97436
rect 631226 97384 631232 97436
rect 631284 97424 631290 97436
rect 639782 97424 639788 97436
rect 631284 97396 639788 97424
rect 631284 97384 631290 97396
rect 639782 97384 639788 97396
rect 639840 97384 639846 97436
rect 639984 97424 640012 97532
rect 643002 97520 643008 97572
rect 643060 97560 643066 97572
rect 657418 97560 657446 97600
rect 659746 97588 659752 97600
rect 659804 97588 659810 97640
rect 643060 97532 657446 97560
rect 643060 97520 643066 97532
rect 658182 97452 658188 97504
rect 658240 97492 658246 97504
rect 663058 97492 663064 97504
rect 658240 97464 663064 97492
rect 658240 97452 658246 97464
rect 663058 97452 663064 97464
rect 663116 97452 663122 97504
rect 647050 97424 647056 97436
rect 639984 97396 647056 97424
rect 647050 97384 647056 97396
rect 647108 97384 647114 97436
rect 651098 97384 651104 97436
rect 651156 97424 651162 97436
rect 654594 97424 654600 97436
rect 651156 97396 654600 97424
rect 651156 97384 651162 97396
rect 654594 97384 654600 97396
rect 654652 97384 654658 97436
rect 656802 97316 656808 97368
rect 656860 97356 656866 97368
rect 661402 97356 661408 97368
rect 656860 97328 661408 97356
rect 656860 97316 656866 97328
rect 661402 97316 661408 97328
rect 661460 97316 661466 97368
rect 623130 97248 623136 97300
rect 623188 97288 623194 97300
rect 632054 97288 632060 97300
rect 623188 97260 632060 97288
rect 623188 97248 623194 97260
rect 632054 97248 632060 97260
rect 632112 97248 632118 97300
rect 632698 97248 632704 97300
rect 632756 97288 632762 97300
rect 650546 97288 650552 97300
rect 632756 97260 650552 97288
rect 632756 97248 632762 97260
rect 650546 97248 650552 97260
rect 650604 97248 650610 97300
rect 651834 97248 651840 97300
rect 651892 97288 651898 97300
rect 654318 97288 654324 97300
rect 651892 97260 654324 97288
rect 651892 97248 651898 97260
rect 654318 97248 654324 97260
rect 654376 97248 654382 97300
rect 658826 97220 658832 97232
rect 654520 97192 658832 97220
rect 626810 97112 626816 97164
rect 626868 97152 626874 97164
rect 639230 97152 639236 97164
rect 626868 97124 639236 97152
rect 626868 97112 626874 97124
rect 639230 97112 639236 97124
rect 639288 97112 639294 97164
rect 644290 97112 644296 97164
rect 644348 97152 644354 97164
rect 654520 97152 654548 97192
rect 658826 97180 658832 97192
rect 658884 97180 658890 97232
rect 659010 97180 659016 97232
rect 659068 97220 659074 97232
rect 661954 97220 661960 97232
rect 659068 97192 661960 97220
rect 659068 97180 659074 97192
rect 661954 97180 661960 97192
rect 662012 97180 662018 97232
rect 644348 97124 654548 97152
rect 644348 97112 644354 97124
rect 612642 97044 612648 97096
rect 612700 97084 612706 97096
rect 621658 97084 621664 97096
rect 612700 97056 621664 97084
rect 612700 97044 612706 97056
rect 621658 97044 621664 97056
rect 621716 97044 621722 97096
rect 658274 97084 658280 97096
rect 654612 97056 658280 97084
rect 624602 96976 624608 97028
rect 624660 97016 624666 97028
rect 634998 97016 635004 97028
rect 624660 96988 635004 97016
rect 624660 96976 624666 96988
rect 634998 96976 635004 96988
rect 635056 96976 635062 97028
rect 635550 96976 635556 97028
rect 635608 97016 635614 97028
rect 639046 97016 639052 97028
rect 635608 96988 639052 97016
rect 635608 96976 635614 96988
rect 639046 96976 639052 96988
rect 639104 96976 639110 97028
rect 639414 96976 639420 97028
rect 639472 97016 639478 97028
rect 647510 97016 647516 97028
rect 639472 96988 647516 97016
rect 639472 96976 639478 96988
rect 647510 96976 647516 96988
rect 647568 96976 647574 97028
rect 650362 96976 650368 97028
rect 650420 97016 650426 97028
rect 654612 97016 654640 97056
rect 658274 97044 658280 97056
rect 658332 97044 658338 97096
rect 650420 96988 654640 97016
rect 650420 96976 650426 96988
rect 596174 96908 596180 96960
rect 596232 96948 596238 96960
rect 596726 96948 596732 96960
rect 596232 96920 596732 96948
rect 596232 96908 596238 96920
rect 596726 96908 596732 96920
rect 596784 96908 596790 96960
rect 615770 96908 615776 96960
rect 615828 96948 615834 96960
rect 616782 96948 616788 96960
rect 615828 96920 616788 96948
rect 615828 96908 615834 96920
rect 616782 96908 616788 96920
rect 616840 96908 616846 96960
rect 654778 96908 654784 96960
rect 654836 96948 654842 96960
rect 655422 96948 655428 96960
rect 654836 96920 655428 96948
rect 654836 96908 654842 96920
rect 655422 96908 655428 96920
rect 655480 96908 655486 96960
rect 660666 96908 660672 96960
rect 660724 96948 660730 96960
rect 663242 96948 663248 96960
rect 660724 96920 663248 96948
rect 660724 96908 660730 96920
rect 663242 96908 663248 96920
rect 663300 96908 663306 96960
rect 612090 96840 612096 96892
rect 612148 96880 612154 96892
rect 612642 96880 612648 96892
rect 612148 96852 612648 96880
rect 612148 96840 612154 96852
rect 612642 96840 612648 96852
rect 612700 96840 612706 96892
rect 617242 96840 617248 96892
rect 617300 96880 617306 96892
rect 618162 96880 618168 96892
rect 617300 96852 618168 96880
rect 617300 96840 617306 96852
rect 618162 96840 618168 96852
rect 618220 96840 618226 96892
rect 633250 96840 633256 96892
rect 633308 96880 633314 96892
rect 633308 96852 639644 96880
rect 633308 96840 633314 96852
rect 606202 96704 606208 96756
rect 606260 96744 606266 96756
rect 611998 96744 612004 96756
rect 606260 96716 612004 96744
rect 606260 96704 606266 96716
rect 611998 96704 612004 96716
rect 612056 96704 612062 96756
rect 634722 96704 634728 96756
rect 634780 96744 634786 96756
rect 639414 96744 639420 96756
rect 634780 96716 639420 96744
rect 634780 96704 634786 96716
rect 639414 96704 639420 96716
rect 639472 96704 639478 96756
rect 639616 96744 639644 96852
rect 639782 96840 639788 96892
rect 639840 96880 639846 96892
rect 647326 96880 647332 96892
rect 639840 96852 647332 96880
rect 639840 96840 639846 96852
rect 647326 96840 647332 96852
rect 647384 96840 647390 96892
rect 654318 96772 654324 96824
rect 654376 96812 654382 96824
rect 659562 96812 659568 96824
rect 654376 96784 659568 96812
rect 654376 96772 654382 96784
rect 659562 96772 659568 96784
rect 659620 96772 659626 96824
rect 650178 96744 650184 96756
rect 639616 96716 650184 96744
rect 650178 96704 650184 96716
rect 650236 96704 650242 96756
rect 638586 96568 638592 96620
rect 638644 96608 638650 96620
rect 638644 96580 642864 96608
rect 638644 96568 638650 96580
rect 639598 96432 639604 96484
rect 639656 96472 639662 96484
rect 642634 96472 642640 96484
rect 639656 96444 642640 96472
rect 639656 96432 639662 96444
rect 642634 96432 642640 96444
rect 642692 96432 642698 96484
rect 642836 96472 642864 96580
rect 645762 96568 645768 96620
rect 645820 96608 645826 96620
rect 652018 96608 652024 96620
rect 645820 96580 652024 96608
rect 645820 96568 645826 96580
rect 652018 96568 652024 96580
rect 652076 96568 652082 96620
rect 652570 96568 652576 96620
rect 652628 96608 652634 96620
rect 664346 96608 664352 96620
rect 652628 96580 664352 96608
rect 652628 96568 652634 96580
rect 664346 96568 664352 96580
rect 664404 96568 664410 96620
rect 652202 96472 652208 96484
rect 642836 96444 652208 96472
rect 652202 96432 652208 96444
rect 652260 96432 652266 96484
rect 653306 96432 653312 96484
rect 653364 96472 653370 96484
rect 665174 96472 665180 96484
rect 653364 96444 665180 96472
rect 653364 96432 653370 96444
rect 665174 96432 665180 96444
rect 665232 96432 665238 96484
rect 640058 96296 640064 96348
rect 640116 96336 640122 96348
rect 647878 96336 647884 96348
rect 640116 96308 647884 96336
rect 640116 96296 640122 96308
rect 647878 96296 647884 96308
rect 647936 96296 647942 96348
rect 648890 96296 648896 96348
rect 648948 96336 648954 96348
rect 664162 96336 664168 96348
rect 648948 96308 664168 96336
rect 648948 96296 648954 96308
rect 664162 96296 664168 96308
rect 664220 96296 664226 96348
rect 637574 96160 637580 96212
rect 637632 96200 637638 96212
rect 660666 96200 660672 96212
rect 637632 96172 660672 96200
rect 637632 96160 637638 96172
rect 660666 96160 660672 96172
rect 660724 96160 660730 96212
rect 610618 96024 610624 96076
rect 610676 96064 610682 96076
rect 623038 96064 623044 96076
rect 610676 96036 623044 96064
rect 610676 96024 610682 96036
rect 623038 96024 623044 96036
rect 623096 96024 623102 96076
rect 641530 96024 641536 96076
rect 641588 96064 641594 96076
rect 663702 96064 663708 96076
rect 641588 96036 663708 96064
rect 641588 96024 641594 96036
rect 663702 96024 663708 96036
rect 663760 96024 663766 96076
rect 577498 95888 577504 95940
rect 577556 95928 577562 95940
rect 601878 95928 601884 95940
rect 577556 95900 601884 95928
rect 577556 95888 577562 95900
rect 601878 95888 601884 95900
rect 601936 95888 601942 95940
rect 607674 95888 607680 95940
rect 607732 95928 607738 95940
rect 622302 95928 622308 95940
rect 607732 95900 622308 95928
rect 607732 95888 607738 95900
rect 622302 95888 622308 95900
rect 622360 95888 622366 95940
rect 645302 95888 645308 95940
rect 645360 95928 645366 95940
rect 649442 95928 649448 95940
rect 645360 95900 649448 95928
rect 645360 95888 645366 95900
rect 649442 95888 649448 95900
rect 649500 95888 649506 95940
rect 649948 95888 649954 95940
rect 650006 95928 650012 95940
rect 664530 95928 664536 95940
rect 650006 95900 664536 95928
rect 650006 95888 650012 95900
rect 664530 95888 664536 95900
rect 664588 95888 664594 95940
rect 642634 95684 642640 95736
rect 642692 95724 642698 95736
rect 651834 95724 651840 95736
rect 642692 95696 651840 95724
rect 642692 95684 642698 95696
rect 651834 95684 651840 95696
rect 651892 95684 651898 95736
rect 641990 95548 641996 95600
rect 642048 95588 642054 95600
rect 646222 95588 646228 95600
rect 642048 95560 646228 95588
rect 642048 95548 642054 95560
rect 646222 95548 646228 95560
rect 646280 95548 646286 95600
rect 646406 95548 646412 95600
rect 646464 95588 646470 95600
rect 646464 95560 649488 95588
rect 646464 95548 646470 95560
rect 649460 95520 649488 95560
rect 649460 95492 649994 95520
rect 640518 95412 640524 95464
rect 640576 95412 640582 95464
rect 643462 95412 643468 95464
rect 643520 95452 643526 95464
rect 649258 95452 649264 95464
rect 643520 95424 649264 95452
rect 643520 95412 643526 95424
rect 649258 95412 649264 95424
rect 649316 95412 649322 95464
rect 640536 95316 640564 95412
rect 649966 95316 649994 95492
rect 653398 95316 653404 95328
rect 640536 95288 649764 95316
rect 649966 95288 653404 95316
rect 620922 95140 620928 95192
rect 620980 95180 620986 95192
rect 626442 95180 626448 95192
rect 620980 95152 626448 95180
rect 620980 95140 620986 95152
rect 626442 95140 626448 95152
rect 626500 95140 626506 95192
rect 647050 95140 647056 95192
rect 647108 95180 647114 95192
rect 648890 95180 648896 95192
rect 647108 95152 648896 95180
rect 647108 95140 647114 95152
rect 648890 95140 648896 95152
rect 648948 95140 648954 95192
rect 649736 95180 649764 95288
rect 653398 95276 653404 95288
rect 653456 95276 653462 95328
rect 649902 95180 649908 95192
rect 649736 95152 649908 95180
rect 649902 95140 649908 95152
rect 649960 95140 649966 95192
rect 579430 95004 579436 95056
rect 579488 95044 579494 95056
rect 584582 95044 584588 95056
rect 579488 95016 584588 95044
rect 579488 95004 579494 95016
rect 584582 95004 584588 95016
rect 584640 95004 584646 95056
rect 649442 94800 649448 94852
rect 649500 94840 649506 94852
rect 656158 94840 656164 94852
rect 649500 94812 656164 94840
rect 649500 94800 649506 94812
rect 656158 94800 656164 94812
rect 656216 94800 656222 94852
rect 609146 94460 609152 94512
rect 609204 94500 609210 94512
rect 620278 94500 620284 94512
rect 609204 94472 620284 94500
rect 609204 94460 609210 94472
rect 620278 94460 620284 94472
rect 620336 94460 620342 94512
rect 648154 93848 648160 93900
rect 648212 93888 648218 93900
rect 654410 93888 654416 93900
rect 648212 93860 654416 93888
rect 648212 93848 648218 93860
rect 654410 93848 654416 93860
rect 654468 93848 654474 93900
rect 619542 93780 619548 93832
rect 619600 93820 619606 93832
rect 626442 93820 626448 93832
rect 619600 93792 626448 93820
rect 619600 93780 619606 93792
rect 626442 93780 626448 93792
rect 626500 93780 626506 93832
rect 579522 93372 579528 93424
rect 579580 93412 579586 93424
rect 585962 93412 585968 93424
rect 579580 93384 585968 93412
rect 579580 93372 579586 93384
rect 585962 93372 585968 93384
rect 586020 93372 586026 93424
rect 611262 93100 611268 93152
rect 611320 93140 611326 93152
rect 619542 93140 619548 93152
rect 611320 93112 619548 93140
rect 611320 93100 611326 93112
rect 619542 93100 619548 93112
rect 619600 93100 619606 93152
rect 647694 92760 647700 92812
rect 647752 92800 647758 92812
rect 655422 92800 655428 92812
rect 647752 92772 655428 92800
rect 647752 92760 647758 92772
rect 655422 92760 655428 92772
rect 655480 92760 655486 92812
rect 607122 92556 607128 92608
rect 607180 92596 607186 92608
rect 610066 92596 610072 92608
rect 607180 92568 610072 92596
rect 607180 92556 607186 92568
rect 610066 92556 610072 92568
rect 610124 92556 610130 92608
rect 617978 92420 617984 92472
rect 618036 92460 618042 92472
rect 626442 92460 626448 92472
rect 618036 92432 626448 92460
rect 618036 92420 618042 92432
rect 626442 92420 626448 92432
rect 626500 92420 626506 92472
rect 652202 92420 652208 92472
rect 652260 92460 652266 92472
rect 655238 92460 655244 92472
rect 652260 92432 655244 92460
rect 652260 92420 652266 92432
rect 655238 92420 655244 92432
rect 655296 92420 655302 92472
rect 579338 91944 579344 91996
rect 579396 91984 579402 91996
rect 585778 91984 585784 91996
rect 579396 91956 585784 91984
rect 579396 91944 579402 91956
rect 585778 91944 585784 91956
rect 585836 91944 585842 91996
rect 579522 91740 579528 91792
rect 579580 91780 579586 91792
rect 588538 91780 588544 91792
rect 579580 91752 588544 91780
rect 579580 91740 579586 91752
rect 588538 91740 588544 91752
rect 588596 91740 588602 91792
rect 616598 91740 616604 91792
rect 616656 91780 616662 91792
rect 626258 91780 626264 91792
rect 616656 91752 626264 91780
rect 616656 91740 616662 91752
rect 626258 91740 626264 91752
rect 626316 91740 626322 91792
rect 618162 90992 618168 91044
rect 618220 91032 618226 91044
rect 626442 91032 626448 91044
rect 618220 91004 626448 91032
rect 618220 90992 618226 91004
rect 626442 90992 626448 91004
rect 626500 90992 626506 91044
rect 622302 89632 622308 89684
rect 622360 89672 622366 89684
rect 626442 89672 626448 89684
rect 622360 89644 626448 89672
rect 622360 89632 622366 89644
rect 626442 89632 626448 89644
rect 626500 89632 626506 89684
rect 581638 88952 581644 89004
rect 581696 88992 581702 89004
rect 600314 88992 600320 89004
rect 581696 88964 600320 88992
rect 581696 88952 581702 88964
rect 600314 88952 600320 88964
rect 600372 88952 600378 89004
rect 649718 88748 649724 88800
rect 649776 88788 649782 88800
rect 658550 88788 658556 88800
rect 649776 88760 658556 88788
rect 649776 88748 649782 88760
rect 658550 88748 658556 88760
rect 658608 88748 658614 88800
rect 662322 88748 662328 88800
rect 662380 88788 662386 88800
rect 663886 88788 663892 88800
rect 662380 88760 663892 88788
rect 662380 88748 662386 88760
rect 663886 88748 663892 88760
rect 663944 88748 663950 88800
rect 610066 88272 610072 88324
rect 610124 88312 610130 88324
rect 626442 88312 626448 88324
rect 610124 88284 626448 88312
rect 610124 88272 610130 88284
rect 626442 88272 626448 88284
rect 626500 88272 626506 88324
rect 655054 88272 655060 88324
rect 655112 88312 655118 88324
rect 658458 88312 658464 88324
rect 655112 88284 658464 88312
rect 655112 88272 655118 88284
rect 658458 88272 658464 88284
rect 658516 88272 658522 88324
rect 619542 88136 619548 88188
rect 619600 88176 619606 88188
rect 626258 88176 626264 88188
rect 619600 88148 626264 88176
rect 619600 88136 619606 88148
rect 626258 88136 626264 88148
rect 626316 88136 626322 88188
rect 578326 86912 578332 86964
rect 578384 86952 578390 86964
rect 580442 86952 580448 86964
rect 578384 86924 580448 86952
rect 578384 86912 578390 86924
rect 580442 86912 580448 86924
rect 580500 86912 580506 86964
rect 659562 86912 659568 86964
rect 659620 86952 659626 86964
rect 663242 86952 663248 86964
rect 659620 86924 663248 86952
rect 659620 86912 659626 86924
rect 663242 86912 663248 86924
rect 663300 86912 663306 86964
rect 652018 86844 652024 86896
rect 652076 86884 652082 86896
rect 657722 86884 657728 86896
rect 652076 86856 657728 86884
rect 652076 86844 652082 86856
rect 657722 86844 657728 86856
rect 657780 86844 657786 86896
rect 649258 86708 649264 86760
rect 649316 86748 649322 86760
rect 661402 86748 661408 86760
rect 649316 86720 661408 86748
rect 649316 86708 649322 86720
rect 661402 86708 661408 86720
rect 661460 86708 661466 86760
rect 647878 86572 647884 86624
rect 647936 86612 647942 86624
rect 660114 86612 660120 86624
rect 647936 86584 660120 86612
rect 647936 86572 647942 86584
rect 660114 86572 660120 86584
rect 660172 86572 660178 86624
rect 656158 86436 656164 86488
rect 656216 86476 656222 86488
rect 660666 86476 660672 86488
rect 656216 86448 660672 86476
rect 656216 86436 656222 86448
rect 660666 86436 660672 86448
rect 660724 86436 660730 86488
rect 623038 86300 623044 86352
rect 623096 86340 623102 86352
rect 626442 86340 626448 86352
rect 623096 86312 626448 86340
rect 623096 86300 623102 86312
rect 626442 86300 626448 86312
rect 626500 86300 626506 86352
rect 654410 86300 654416 86352
rect 654468 86340 654474 86352
rect 662506 86340 662512 86352
rect 654468 86312 662512 86340
rect 654468 86300 654474 86312
rect 662506 86300 662512 86312
rect 662564 86300 662570 86352
rect 653398 86164 653404 86216
rect 653456 86204 653462 86216
rect 657170 86204 657176 86216
rect 653456 86176 657176 86204
rect 653456 86164 653462 86176
rect 657170 86164 657176 86176
rect 657228 86164 657234 86216
rect 609882 85484 609888 85536
rect 609940 85524 609946 85536
rect 626442 85524 626448 85536
rect 609940 85496 626448 85524
rect 609940 85484 609946 85496
rect 626442 85484 626448 85496
rect 626500 85484 626506 85536
rect 578418 85416 578424 85468
rect 578476 85456 578482 85468
rect 581822 85456 581828 85468
rect 578476 85428 581828 85456
rect 578476 85416 578482 85428
rect 581822 85416 581828 85428
rect 581880 85416 581886 85468
rect 620278 85348 620284 85400
rect 620336 85388 620342 85400
rect 625246 85388 625252 85400
rect 620336 85360 625252 85388
rect 620336 85348 620342 85360
rect 625246 85348 625252 85360
rect 625304 85348 625310 85400
rect 608502 84124 608508 84176
rect 608560 84164 608566 84176
rect 625798 84164 625804 84176
rect 608560 84136 625804 84164
rect 608560 84124 608566 84136
rect 625798 84124 625804 84136
rect 625856 84124 625862 84176
rect 579522 83988 579528 84040
rect 579580 84028 579586 84040
rect 583018 84028 583024 84040
rect 579580 84000 583024 84028
rect 579580 83988 579586 84000
rect 583018 83988 583024 84000
rect 583076 83988 583082 84040
rect 579430 82424 579436 82476
rect 579488 82464 579494 82476
rect 584398 82464 584404 82476
rect 579488 82436 584404 82464
rect 579488 82424 579494 82436
rect 584398 82424 584404 82436
rect 584456 82424 584462 82476
rect 628742 81064 628748 81116
rect 628800 81104 628806 81116
rect 642450 81104 642456 81116
rect 628800 81076 642456 81104
rect 628800 81064 628806 81076
rect 642450 81064 642456 81076
rect 642508 81064 642514 81116
rect 618898 80928 618904 80980
rect 618956 80968 618962 80980
rect 649074 80968 649080 80980
rect 618956 80940 649080 80968
rect 618956 80928 618962 80940
rect 649074 80928 649080 80940
rect 649132 80928 649138 80980
rect 614022 80792 614028 80844
rect 614080 80832 614086 80844
rect 646038 80832 646044 80844
rect 614080 80804 646044 80832
rect 614080 80792 614086 80804
rect 646038 80792 646044 80804
rect 646096 80792 646102 80844
rect 595438 80656 595444 80708
rect 595496 80696 595502 80708
rect 636102 80696 636108 80708
rect 595496 80668 636108 80696
rect 595496 80656 595502 80668
rect 636102 80656 636108 80668
rect 636160 80656 636166 80708
rect 585778 79432 585784 79484
rect 585836 79472 585842 79484
rect 589918 79472 589924 79484
rect 585836 79444 589924 79472
rect 585836 79432 585842 79444
rect 589918 79432 589924 79444
rect 589976 79432 589982 79484
rect 629202 79432 629208 79484
rect 629260 79472 629266 79484
rect 645302 79472 645308 79484
rect 629260 79444 645308 79472
rect 629260 79432 629266 79444
rect 645302 79432 645308 79444
rect 645360 79432 645366 79484
rect 579062 79296 579068 79348
rect 579120 79336 579126 79348
rect 598934 79336 598940 79348
rect 579120 79308 598940 79336
rect 579120 79296 579126 79308
rect 598934 79296 598940 79308
rect 598992 79296 598998 79348
rect 615402 79296 615408 79348
rect 615460 79336 615466 79348
rect 646222 79336 646228 79348
rect 615460 79308 646228 79336
rect 615460 79296 615466 79308
rect 646222 79296 646228 79308
rect 646280 79296 646286 79348
rect 631042 78072 631048 78124
rect 631100 78112 631106 78124
rect 643094 78112 643100 78124
rect 631100 78084 643100 78112
rect 631100 78072 631106 78084
rect 643094 78072 643100 78084
rect 643152 78072 643158 78124
rect 621658 77936 621664 77988
rect 621716 77976 621722 77988
rect 648706 77976 648712 77988
rect 621716 77948 648712 77976
rect 621716 77936 621722 77948
rect 648706 77936 648712 77948
rect 648764 77936 648770 77988
rect 578326 77664 578332 77716
rect 578384 77704 578390 77716
rect 580258 77704 580264 77716
rect 578384 77676 580264 77704
rect 578384 77664 578390 77676
rect 580258 77664 580264 77676
rect 580316 77664 580322 77716
rect 631042 77432 631048 77444
rect 625126 77404 631048 77432
rect 584398 77256 584404 77308
rect 584456 77296 584462 77308
rect 625126 77296 625154 77404
rect 631042 77392 631048 77404
rect 631100 77392 631106 77444
rect 584456 77268 625154 77296
rect 584456 77256 584462 77268
rect 628466 77256 628472 77308
rect 628524 77296 628530 77308
rect 632790 77296 632796 77308
rect 628524 77268 632796 77296
rect 628524 77256 628530 77268
rect 632790 77256 632796 77268
rect 632848 77256 632854 77308
rect 616782 76644 616788 76696
rect 616840 76684 616846 76696
rect 646774 76684 646780 76696
rect 616840 76656 646780 76684
rect 616840 76644 616846 76656
rect 646774 76644 646780 76656
rect 646832 76644 646838 76696
rect 606478 76508 606484 76560
rect 606536 76548 606542 76560
rect 662414 76548 662420 76560
rect 606536 76520 662420 76548
rect 606536 76508 606542 76520
rect 662414 76508 662420 76520
rect 662472 76508 662478 76560
rect 588538 75896 588544 75948
rect 588596 75936 588602 75948
rect 628466 75936 628472 75948
rect 588596 75908 628472 75936
rect 588596 75896 588602 75908
rect 628466 75896 628472 75908
rect 628524 75896 628530 75948
rect 612642 75420 612648 75472
rect 612700 75460 612706 75472
rect 646590 75460 646596 75472
rect 612700 75432 646596 75460
rect 612700 75420 612706 75432
rect 646590 75420 646596 75432
rect 646648 75420 646654 75472
rect 611998 75284 612004 75336
rect 612056 75324 612062 75336
rect 646406 75324 646412 75336
rect 612056 75296 646412 75324
rect 612056 75284 612062 75296
rect 646406 75284 646412 75296
rect 646464 75284 646470 75336
rect 578878 75148 578884 75200
rect 578936 75188 578942 75200
rect 666554 75188 666560 75200
rect 578936 75160 666560 75188
rect 578936 75148 578942 75160
rect 666554 75148 666560 75160
rect 666612 75148 666618 75200
rect 579522 73108 579528 73160
rect 579580 73148 579586 73160
rect 587158 73148 587164 73160
rect 579580 73120 587164 73148
rect 579580 73108 579586 73120
rect 587158 73108 587164 73120
rect 587216 73108 587222 73160
rect 579522 71204 579528 71256
rect 579580 71244 579586 71256
rect 585778 71244 585784 71256
rect 579580 71216 585784 71244
rect 579580 71204 579586 71216
rect 585778 71204 585784 71216
rect 585836 71204 585842 71256
rect 585778 68280 585784 68332
rect 585836 68320 585842 68332
rect 601878 68320 601884 68332
rect 585836 68292 601884 68320
rect 585836 68280 585842 68292
rect 601878 68280 601884 68292
rect 601936 68280 601942 68332
rect 579522 66240 579528 66292
rect 579580 66280 579586 66292
rect 623038 66280 623044 66292
rect 579580 66252 623044 66280
rect 579580 66240 579586 66252
rect 623038 66240 623044 66252
rect 623096 66240 623102 66292
rect 579522 64812 579528 64864
rect 579580 64852 579586 64864
rect 614850 64852 614856 64864
rect 579580 64824 614856 64852
rect 579580 64812 579586 64824
rect 614850 64812 614856 64824
rect 614908 64812 614914 64864
rect 578510 62024 578516 62076
rect 578568 62064 578574 62076
rect 613378 62064 613384 62076
rect 578568 62036 613384 62064
rect 578568 62024 578574 62036
rect 613378 62024 613384 62036
rect 613436 62024 613442 62076
rect 580258 58624 580264 58676
rect 580316 58664 580322 58676
rect 600498 58664 600504 58676
rect 580316 58636 600504 58664
rect 580316 58624 580322 58636
rect 600498 58624 600504 58636
rect 600556 58624 600562 58676
rect 579522 57876 579528 57928
rect 579580 57916 579586 57928
rect 624418 57916 624424 57928
rect 579580 57888 624424 57916
rect 579580 57876 579586 57888
rect 624418 57876 624424 57888
rect 624476 57876 624482 57928
rect 576854 57196 576860 57248
rect 576912 57236 576918 57248
rect 603074 57236 603080 57248
rect 576912 57208 603080 57236
rect 576912 57196 576918 57208
rect 603074 57196 603080 57208
rect 603132 57196 603138 57248
rect 579522 56516 579528 56568
rect 579580 56556 579586 56568
rect 588538 56556 588544 56568
rect 579580 56528 588544 56556
rect 579580 56516 579586 56528
rect 588538 56516 588544 56528
rect 588596 56516 588602 56568
rect 574554 56108 574560 56160
rect 574612 56148 574618 56160
rect 596450 56148 596456 56160
rect 574612 56120 596456 56148
rect 574612 56108 574618 56120
rect 596450 56108 596456 56120
rect 596508 56108 596514 56160
rect 574922 55972 574928 56024
rect 574980 56012 574986 56024
rect 596174 56012 596180 56024
rect 574980 55984 596180 56012
rect 574980 55972 574986 55984
rect 596174 55972 596180 55984
rect 596232 55972 596238 56024
rect 574738 55836 574744 55888
rect 574796 55876 574802 55888
rect 599118 55876 599124 55888
rect 574796 55848 599124 55876
rect 574796 55836 574802 55848
rect 599118 55836 599124 55848
rect 599176 55836 599182 55888
rect 462286 55576 488534 55604
rect 462286 53644 462314 55576
rect 473924 55372 478874 55400
rect 473924 55264 473952 55372
rect 478846 55332 478874 55372
rect 478846 55304 479012 55332
rect 473326 55236 473952 55264
rect 473326 55060 473354 55236
rect 462222 53592 462228 53644
rect 462280 53604 462314 53644
rect 462378 55032 473354 55060
rect 478984 55060 479012 55304
rect 479260 55236 483796 55264
rect 479260 55060 479288 55236
rect 478984 55032 479288 55060
rect 483768 55060 483796 55236
rect 488506 55196 488534 55576
rect 581638 55196 581644 55208
rect 488506 55168 581644 55196
rect 581638 55156 581644 55168
rect 581696 55156 581702 55208
rect 579062 55060 579068 55072
rect 483768 55032 579068 55060
rect 462280 53592 462286 53604
rect 459462 53456 459468 53508
rect 459520 53496 459526 53508
rect 462378 53496 462406 55032
rect 579062 55020 579068 55032
rect 579120 55020 579126 55072
rect 584398 54924 584404 54936
rect 467116 54896 584404 54924
rect 467116 53904 467144 54896
rect 584398 54884 584404 54896
rect 584456 54884 584462 54936
rect 589918 54788 589924 54800
rect 462792 53876 467144 53904
rect 472728 54760 589924 54788
rect 462792 53644 462820 53876
rect 472728 53644 472756 54760
rect 589918 54748 589924 54760
rect 589976 54748 589982 54800
rect 597646 54652 597652 54664
rect 475672 54624 597652 54652
rect 475672 53904 475700 54624
rect 597646 54612 597652 54624
rect 597704 54612 597710 54664
rect 597922 54516 597928 54528
rect 473188 53876 475700 53904
rect 476776 54488 597928 54516
rect 473188 53644 473216 53876
rect 476776 53644 476804 54488
rect 597922 54476 597928 54488
rect 597980 54476 597986 54528
rect 583018 54380 583024 54392
rect 477880 54352 583024 54380
rect 477880 53644 477908 54352
rect 583018 54340 583024 54352
rect 583076 54340 583082 54392
rect 580258 54244 580264 54256
rect 481744 54216 580264 54244
rect 481744 53644 481772 54216
rect 580258 54204 580264 54216
rect 580316 54204 580322 54256
rect 574738 54108 574744 54120
rect 485148 54080 574744 54108
rect 485148 53768 485176 54080
rect 574738 54068 574744 54080
rect 574796 54068 574802 54120
rect 574554 53972 574560 53984
rect 482296 53740 485176 53768
rect 485240 53944 574560 53972
rect 482296 53644 482324 53740
rect 485240 53644 485268 53944
rect 574554 53932 574560 53944
rect 574612 53932 574618 53984
rect 574922 53836 574928 53848
rect 489886 53808 574928 53836
rect 462774 53592 462780 53644
rect 462832 53592 462838 53644
rect 463602 53592 463608 53644
rect 463660 53632 463666 53644
rect 464338 53632 464344 53644
rect 463660 53604 464344 53632
rect 463660 53592 463666 53604
rect 464338 53592 464344 53604
rect 464396 53592 464402 53644
rect 472710 53592 472716 53644
rect 472768 53592 472774 53644
rect 473170 53592 473176 53644
rect 473228 53592 473234 53644
rect 476758 53592 476764 53644
rect 476816 53592 476822 53644
rect 477862 53592 477868 53644
rect 477920 53592 477926 53644
rect 481726 53592 481732 53644
rect 481784 53592 481790 53644
rect 482278 53592 482284 53644
rect 482336 53592 482342 53644
rect 485222 53592 485228 53644
rect 485280 53592 485286 53644
rect 472526 53564 472532 53576
rect 467806 53536 472532 53564
rect 459520 53468 462406 53496
rect 459520 53456 459526 53468
rect 463142 53456 463148 53508
rect 463200 53496 463206 53508
rect 467806 53496 467834 53536
rect 472526 53524 472532 53536
rect 472584 53524 472590 53576
rect 463200 53468 467834 53496
rect 463200 53456 463206 53468
rect 477126 53456 477132 53508
rect 477184 53496 477190 53508
rect 482094 53496 482100 53508
rect 477184 53468 482100 53496
rect 477184 53456 477190 53468
rect 482094 53456 482100 53468
rect 482152 53456 482158 53508
rect 482462 53456 482468 53508
rect 482520 53496 482526 53508
rect 489886 53496 489914 53808
rect 574922 53796 574928 53808
rect 574980 53796 574986 53848
rect 482520 53468 489914 53496
rect 482520 53456 482526 53468
rect 50338 53320 50344 53372
rect 50396 53360 50402 53372
rect 130378 53360 130384 53372
rect 50396 53332 130384 53360
rect 50396 53320 50402 53332
rect 130378 53320 130384 53332
rect 130436 53320 130442 53372
rect 460382 53320 460388 53372
rect 460440 53360 460446 53372
rect 462774 53360 462780 53372
rect 460440 53332 462780 53360
rect 460440 53320 460446 53332
rect 462774 53320 462780 53332
rect 462832 53320 462838 53372
rect 465442 53320 465448 53372
rect 465500 53360 465506 53372
rect 477862 53360 477868 53372
rect 465500 53332 477868 53360
rect 465500 53320 465506 53332
rect 477862 53320 477868 53332
rect 477920 53320 477926 53372
rect 47762 53184 47768 53236
rect 47820 53224 47826 53236
rect 130562 53224 130568 53236
rect 47820 53196 130568 53224
rect 47820 53184 47826 53196
rect 130562 53184 130568 53196
rect 130620 53184 130626 53236
rect 463418 53184 463424 53236
rect 463476 53224 463482 53236
rect 476758 53224 476764 53236
rect 463476 53196 476764 53224
rect 463476 53184 463482 53196
rect 476758 53184 476764 53196
rect 476816 53184 476822 53236
rect 312354 53116 312360 53168
rect 312412 53156 312418 53168
rect 313734 53156 313740 53168
rect 312412 53128 313740 53156
rect 312412 53116 312418 53128
rect 313734 53116 313740 53128
rect 313792 53116 313798 53168
rect 316310 53116 316316 53168
rect 316368 53156 316374 53168
rect 317690 53156 317696 53168
rect 316368 53128 317696 53156
rect 316368 53116 316374 53128
rect 317690 53116 317696 53128
rect 317748 53116 317754 53168
rect 46198 53048 46204 53100
rect 46256 53088 46262 53100
rect 128998 53088 129004 53100
rect 46256 53060 129004 53088
rect 46256 53048 46262 53060
rect 128998 53048 129004 53060
rect 129056 53048 129062 53100
rect 464522 53048 464528 53100
rect 464580 53088 464586 53100
rect 473170 53088 473176 53100
rect 464580 53060 473176 53088
rect 464580 53048 464586 53060
rect 473170 53048 473176 53060
rect 473228 53048 473234 53100
rect 464062 52912 464068 52964
rect 464120 52952 464126 52964
rect 477126 52952 477132 52964
rect 464120 52924 477132 52952
rect 464120 52912 464126 52924
rect 477126 52912 477132 52924
rect 477184 52912 477190 52964
rect 464660 52776 464666 52828
rect 464718 52816 464724 52828
rect 485222 52816 485228 52828
rect 464718 52788 485228 52816
rect 464718 52776 464724 52788
rect 485222 52776 485228 52788
rect 485280 52776 485286 52828
rect 460980 52708 460986 52760
rect 461038 52748 461044 52760
rect 463602 52748 463608 52760
rect 461038 52720 463608 52748
rect 461038 52708 461044 52720
rect 463602 52708 463608 52720
rect 463660 52708 463666 52760
rect 465902 52640 465908 52692
rect 465960 52680 465966 52692
rect 472710 52680 472716 52692
rect 465960 52652 472716 52680
rect 465960 52640 465966 52652
rect 472710 52640 472716 52652
rect 472768 52640 472774 52692
rect 145374 52436 145380 52488
rect 145432 52476 145438 52488
rect 306006 52476 306012 52488
rect 145432 52448 306012 52476
rect 145432 52436 145438 52448
rect 306006 52436 306012 52448
rect 306064 52436 306070 52488
rect 49142 51960 49148 52012
rect 49200 52000 49206 52012
rect 126422 52000 126428 52012
rect 49200 51972 126428 52000
rect 49200 51960 49206 51972
rect 126422 51960 126428 51972
rect 126480 51960 126486 52012
rect 48958 51824 48964 51876
rect 49016 51864 49022 51876
rect 129458 51864 129464 51876
rect 49016 51836 129464 51864
rect 49016 51824 49022 51836
rect 129458 51824 129464 51836
rect 129516 51824 129522 51876
rect 46382 51688 46388 51740
rect 46440 51728 46446 51740
rect 130746 51728 130752 51740
rect 46440 51700 130752 51728
rect 46440 51688 46446 51700
rect 130746 51688 130752 51700
rect 130804 51688 130810 51740
rect 126422 50736 126428 50788
rect 126480 50776 126486 50788
rect 129274 50776 129280 50788
rect 126480 50748 129280 50776
rect 126480 50736 126486 50748
rect 129274 50736 129280 50748
rect 129332 50736 129338 50788
rect 50522 50464 50528 50516
rect 50580 50504 50586 50516
rect 128630 50504 128636 50516
rect 50580 50476 128636 50504
rect 50580 50464 50586 50476
rect 128630 50464 128636 50476
rect 128688 50464 128694 50516
rect 318334 50464 318340 50516
rect 318392 50504 318398 50516
rect 458358 50504 458364 50516
rect 318392 50476 458364 50504
rect 318392 50464 318398 50476
rect 458358 50464 458364 50476
rect 458416 50464 458422 50516
rect 45462 50328 45468 50380
rect 45520 50368 45526 50380
rect 128998 50368 129004 50380
rect 45520 50340 129004 50368
rect 45520 50328 45526 50340
rect 128998 50328 129004 50340
rect 129056 50328 129062 50380
rect 314010 50328 314016 50380
rect 314068 50368 314074 50380
rect 458174 50368 458180 50380
rect 314068 50340 458180 50368
rect 314068 50328 314074 50340
rect 458174 50328 458180 50340
rect 458232 50328 458238 50380
rect 51718 49104 51724 49156
rect 51776 49144 51782 49156
rect 128446 49144 128452 49156
rect 51776 49116 128452 49144
rect 51776 49104 51782 49116
rect 128446 49104 128452 49116
rect 128504 49104 128510 49156
rect 47578 48968 47584 49020
rect 47636 49008 47642 49020
rect 129642 49008 129648 49020
rect 47636 48980 129648 49008
rect 47636 48968 47642 48980
rect 129642 48968 129648 48980
rect 129700 48968 129706 49020
rect 128630 48084 128636 48136
rect 128688 48124 128694 48136
rect 132126 48124 132132 48136
rect 128688 48096 132132 48124
rect 128688 48084 128694 48096
rect 132126 48084 132132 48096
rect 132184 48084 132190 48136
rect 129182 47676 129188 47728
rect 129240 47716 129246 47728
rect 131850 47716 131856 47728
rect 129240 47688 131856 47716
rect 129240 47676 129246 47688
rect 131850 47676 131856 47688
rect 131908 47676 131914 47728
rect 623038 46452 623044 46504
rect 623096 46492 623102 46504
rect 661586 46492 661592 46504
rect 623096 46464 661592 46492
rect 623096 46452 623102 46464
rect 661586 46452 661592 46464
rect 661644 46452 661650 46504
rect 129550 45024 129556 45076
rect 129608 45064 129614 45076
rect 130856 45064 131146 45076
rect 129608 45048 131146 45064
rect 129608 45036 130884 45048
rect 129608 45024 129614 45036
rect 131316 44964 131376 44992
rect 129734 44888 129740 44940
rect 129792 44928 129798 44940
rect 131316 44928 131344 44964
rect 129792 44900 131344 44928
rect 129792 44888 129798 44900
rect 131592 44792 131620 44894
rect 131546 44764 131620 44792
rect 131730 44796 131790 44824
rect 131546 44740 131574 44764
rect 131500 44724 131574 44740
rect 131408 44712 131574 44724
rect 131408 44696 131528 44712
rect 128446 44616 128452 44668
rect 128504 44656 128510 44668
rect 131408 44656 131436 44696
rect 128504 44628 131436 44656
rect 128504 44616 128510 44628
rect 129366 44480 129372 44532
rect 129424 44520 129430 44532
rect 131730 44520 131758 44796
rect 131960 44724 131988 44726
rect 131868 44696 131988 44724
rect 131868 44600 131896 44696
rect 131850 44548 131856 44600
rect 131908 44548 131914 44600
rect 132236 44520 132264 44642
rect 129424 44492 131758 44520
rect 132144 44500 132264 44520
rect 129424 44480 129430 44492
rect 132126 44448 132132 44500
rect 132184 44492 132264 44500
rect 132184 44448 132190 44492
rect 132420 44464 132448 44558
rect 132402 44412 132408 44464
rect 132460 44412 132466 44464
rect 130746 44276 130752 44328
rect 130804 44316 130810 44328
rect 132604 44316 132632 44474
rect 130804 44288 132632 44316
rect 130804 44276 130810 44288
rect 128998 44140 129004 44192
rect 129056 44180 129062 44192
rect 132218 44180 132224 44192
rect 129056 44152 132224 44180
rect 129056 44140 129062 44152
rect 132218 44140 132224 44152
rect 132276 44140 132282 44192
rect 132788 44180 132816 44362
rect 132420 44152 132816 44180
rect 130378 44004 130384 44056
rect 130436 44044 130442 44056
rect 132420 44044 132448 44152
rect 130436 44016 132448 44044
rect 130436 44004 130442 44016
rect 130562 43868 130568 43920
rect 130620 43908 130626 43920
rect 132972 43908 133000 44250
rect 130620 43880 133000 43908
rect 130620 43868 130626 43880
rect 43438 42780 43444 42832
rect 43496 42820 43502 42832
rect 133156 42820 133184 44138
rect 431218 43636 431224 43648
rect 412606 43608 431224 43636
rect 187326 43528 187332 43580
rect 187384 43568 187390 43580
rect 412606 43568 412634 43608
rect 431218 43596 431224 43608
rect 431276 43596 431282 43648
rect 187384 43540 412634 43568
rect 187384 43528 187390 43540
rect 43496 42792 133184 42820
rect 43496 42780 43502 42792
rect 310422 42712 310428 42764
rect 310480 42752 310486 42764
rect 310480 42724 354674 42752
rect 310480 42712 310486 42724
rect 354646 42616 354674 42724
rect 364886 42712 364892 42764
rect 364944 42752 364950 42764
rect 431218 42752 431224 42764
rect 364944 42724 431224 42752
rect 364944 42712 364950 42724
rect 431218 42712 431224 42724
rect 431276 42712 431282 42764
rect 456058 42712 456064 42764
rect 456116 42752 456122 42764
rect 463878 42752 463884 42764
rect 456116 42724 463884 42752
rect 456116 42712 456122 42724
rect 463878 42712 463884 42724
rect 463936 42712 463942 42764
rect 427078 42616 427084 42628
rect 354646 42588 427084 42616
rect 427078 42576 427084 42588
rect 427136 42576 427142 42628
rect 455414 42440 455420 42492
rect 455472 42480 455478 42492
rect 462958 42480 462964 42492
rect 455472 42452 462964 42480
rect 455472 42440 455478 42452
rect 462958 42440 462964 42452
rect 463016 42440 463022 42492
rect 404446 42304 404452 42356
rect 404504 42344 404510 42356
rect 405182 42344 405188 42356
rect 404504 42316 405188 42344
rect 404504 42304 404510 42316
rect 405182 42304 405188 42316
rect 405240 42304 405246 42356
rect 420730 42304 420736 42356
rect 420788 42344 420794 42356
rect 426894 42344 426900 42356
rect 420788 42316 426900 42344
rect 420788 42304 420794 42316
rect 426894 42304 426900 42316
rect 426952 42304 426958 42356
rect 663794 42173 663800 42225
rect 663852 42173 663858 42225
rect 427078 42032 427084 42084
rect 427136 42072 427142 42084
rect 427136 42044 427814 42072
rect 427136 42032 427142 42044
rect 427786 41936 427814 42044
rect 431218 42032 431224 42084
rect 431276 42072 431282 42084
rect 456058 42072 456064 42084
rect 431276 42044 456064 42072
rect 431276 42032 431282 42044
rect 456058 42032 456064 42044
rect 456116 42032 456122 42084
rect 455414 41936 455420 41948
rect 427786 41908 455420 41936
rect 455414 41896 455420 41908
rect 455472 41896 455478 41948
rect 404446 41420 404452 41472
rect 404504 41460 404510 41472
rect 420730 41460 420736 41472
rect 404504 41432 420736 41460
rect 404504 41420 404510 41432
rect 420730 41420 420736 41432
rect 420788 41420 420794 41472
rect 426894 41420 426900 41472
rect 426952 41460 426958 41472
rect 459186 41460 459192 41472
rect 426952 41432 459192 41460
rect 426952 41420 426958 41432
rect 459186 41420 459192 41432
rect 459244 41420 459250 41472
<< via1 >>
rect 366180 1027828 366232 1027880
rect 366548 1027828 366600 1027880
rect 366180 1024360 366232 1024412
rect 366548 1024360 366600 1024412
rect 426348 1007088 426400 1007140
rect 437480 1007088 437532 1007140
rect 358544 1006952 358596 1007004
rect 373264 1006952 373316 1007004
rect 553952 1006952 554004 1007004
rect 562324 1006952 562376 1007004
rect 505008 1006884 505060 1006936
rect 513380 1006884 513432 1006936
rect 359372 1006816 359424 1006868
rect 380164 1006816 380216 1006868
rect 555976 1006816 556028 1006868
rect 569408 1006816 569460 1006868
rect 429200 1006748 429252 1006800
rect 144184 1006680 144236 1006732
rect 150256 1006680 150308 1006732
rect 161940 1006680 161992 1006732
rect 164884 1006680 164936 1006732
rect 360200 1006680 360252 1006732
rect 94504 1006544 94556 1006596
rect 101956 1006544 102008 1006596
rect 145748 1006544 145800 1006596
rect 153752 1006544 153804 1006596
rect 157432 1006544 157484 1006596
rect 166264 1006544 166316 1006596
rect 93124 1006408 93176 1006460
rect 98276 1006408 98328 1006460
rect 145564 1006408 145616 1006460
rect 152924 1006408 152976 1006460
rect 160284 1006408 160336 1006460
rect 161940 1006408 161992 1006460
rect 162768 1006408 162820 1006460
rect 173164 1006544 173216 1006596
rect 364892 1006544 364944 1006596
rect 371884 1006544 371936 1006596
rect 247684 1006408 247736 1006460
rect 256148 1006408 256200 1006460
rect 354864 1006408 354916 1006460
rect 363604 1006408 363656 1006460
rect 374644 1006408 374696 1006460
rect 101404 1006272 101456 1006324
rect 103980 1006272 104032 1006324
rect 108488 1006272 108540 1006324
rect 126244 1006272 126296 1006324
rect 144368 1006204 144420 1006256
rect 151268 1006204 151320 1006256
rect 92480 1006136 92532 1006188
rect 94688 1006000 94740 1006052
rect 99472 1006000 99524 1006052
rect 101588 1006136 101640 1006188
rect 104808 1006136 104860 1006188
rect 106832 1006136 106884 1006188
rect 113824 1006136 113876 1006188
rect 148876 1006068 148928 1006120
rect 150072 1006068 150124 1006120
rect 150256 1006068 150308 1006120
rect 152096 1006272 152148 1006324
rect 158260 1006272 158312 1006324
rect 171784 1006272 171836 1006324
rect 255964 1006272 256016 1006324
rect 259000 1006272 259052 1006324
rect 301504 1006272 301556 1006324
rect 307760 1006272 307812 1006324
rect 314660 1006272 314712 1006324
rect 320824 1006272 320876 1006324
rect 361396 1006272 361448 1006324
rect 158628 1006136 158680 1006188
rect 162768 1006136 162820 1006188
rect 166264 1006136 166316 1006188
rect 175924 1006136 175976 1006188
rect 210424 1006136 210476 1006188
rect 228364 1006136 228416 1006188
rect 249064 1006136 249116 1006188
rect 257344 1006136 257396 1006188
rect 262680 1006136 262732 1006188
rect 269764 1006136 269816 1006188
rect 298744 1006136 298796 1006188
rect 304908 1006136 304960 1006188
rect 360568 1006136 360620 1006188
rect 103152 1006000 103204 1006052
rect 106004 1006000 106056 1006052
rect 124864 1006000 124916 1006052
rect 153936 1006000 153988 1006052
rect 158260 1006000 158312 1006052
rect 159456 1006000 159508 1006052
rect 177304 1006000 177356 1006052
rect 195152 1006000 195204 1006052
rect 201040 1006000 201092 1006052
rect 208400 1006000 208452 1006052
rect 229744 1006000 229796 1006052
rect 257344 1006000 257396 1006052
rect 258172 1006000 258224 1006052
rect 261852 1006000 261904 1006052
rect 279424 1006000 279476 1006052
rect 298928 1006000 298980 1006052
rect 303252 1006000 303304 1006052
rect 304080 1006000 304132 1006052
rect 311808 1006000 311860 1006052
rect 314660 1006000 314712 1006052
rect 319444 1006000 319496 1006052
rect 358544 1006000 358596 1006052
rect 362224 1006000 362276 1006052
rect 363420 1006136 363472 1006188
rect 402244 1006272 402296 1006324
rect 431684 1006612 431736 1006664
rect 507860 1006680 507912 1006732
rect 520924 1006680 520976 1006732
rect 556804 1006680 556856 1006732
rect 564440 1006680 564492 1006732
rect 469864 1006544 469916 1006596
rect 505376 1006544 505428 1006596
rect 518164 1006544 518216 1006596
rect 428372 1006476 428424 1006528
rect 440884 1006476 440936 1006528
rect 506204 1006408 506256 1006460
rect 427544 1006272 427596 1006324
rect 364892 1006000 364944 1006052
rect 365076 1006000 365128 1006052
rect 367744 1006000 367796 1006052
rect 377404 1006136 377456 1006188
rect 382832 1006000 382884 1006052
rect 400864 1006000 400916 1006052
rect 429200 1006136 429252 1006188
rect 451924 1006136 451976 1006188
rect 425152 1006000 425204 1006052
rect 429752 1006000 429804 1006052
rect 431684 1006000 431736 1006052
rect 471244 1006000 471296 1006052
rect 496728 1006000 496780 1006052
rect 498844 1006000 498896 1006052
rect 555148 1006408 555200 1006460
rect 570328 1006408 570380 1006460
rect 551468 1006272 551520 1006324
rect 556804 1006272 556856 1006324
rect 555424 1006136 555476 1006188
rect 558828 1006136 558880 1006188
rect 562324 1006136 562376 1006188
rect 567844 1006136 567896 1006188
rect 522304 1006000 522356 1006052
rect 549168 1006000 549220 1006052
rect 550272 1006000 550324 1006052
rect 554780 1006000 554832 1006052
rect 573548 1006000 573600 1006052
rect 428372 1005796 428424 1005848
rect 454684 1005796 454736 1005848
rect 423496 1005660 423548 1005712
rect 432420 1005660 432472 1005712
rect 421840 1005524 421892 1005576
rect 425704 1005524 425756 1005576
rect 445024 1005660 445076 1005712
rect 360568 1005388 360620 1005440
rect 378784 1005388 378836 1005440
rect 423496 1005388 423548 1005440
rect 437480 1005524 437532 1005576
rect 467104 1005524 467156 1005576
rect 432420 1005388 432472 1005440
rect 457444 1005388 457496 1005440
rect 499488 1005388 499540 1005440
rect 500500 1005388 500552 1005440
rect 564440 1005388 564492 1005440
rect 570604 1005388 570656 1005440
rect 427176 1005320 427228 1005372
rect 102784 1005252 102836 1005304
rect 108856 1005252 108908 1005304
rect 204904 1005252 204956 1005304
rect 212080 1005252 212132 1005304
rect 355692 1005252 355744 1005304
rect 376024 1005252 376076 1005304
rect 463700 1005252 463752 1005304
rect 498844 1005252 498896 1005304
rect 516784 1005252 516836 1005304
rect 551468 1005252 551520 1005304
rect 569224 1005252 569276 1005304
rect 304264 1005184 304316 1005236
rect 307300 1005184 307352 1005236
rect 151084 1005048 151136 1005100
rect 153752 1005048 153804 1005100
rect 365076 1005048 365128 1005100
rect 370504 1005048 370556 1005100
rect 425520 1005048 425572 1005100
rect 431224 1005048 431276 1005100
rect 149704 1004912 149756 1004964
rect 152924 1004912 152976 1004964
rect 209228 1004912 209280 1004964
rect 211804 1004912 211856 1004964
rect 263048 1004912 263100 1004964
rect 268384 1004912 268436 1004964
rect 303620 1004912 303672 1004964
rect 306932 1004912 306984 1004964
rect 354588 1004912 354640 1004964
rect 356520 1004912 356572 1004964
rect 361396 1004912 361448 1004964
rect 364984 1004912 365036 1004964
rect 428004 1004912 428056 1004964
rect 439504 1005048 439556 1005100
rect 498108 1004912 498160 1004964
rect 500500 1004912 500552 1004964
rect 557172 1004912 557224 1004964
rect 558920 1004912 558972 1004964
rect 151268 1004776 151320 1004828
rect 154120 1004776 154172 1004828
rect 160652 1004776 160704 1004828
rect 163136 1004776 163188 1004828
rect 211252 1004776 211304 1004828
rect 215944 1004776 215996 1004828
rect 258172 1004776 258224 1004828
rect 259460 1004776 259512 1004828
rect 305828 1004776 305880 1004828
rect 308956 1004776 309008 1004828
rect 313832 1004776 313884 1004828
rect 316040 1004776 316092 1004828
rect 353208 1004776 353260 1004828
rect 355692 1004776 355744 1004828
rect 362592 1004776 362644 1004828
rect 365168 1004776 365220 1004828
rect 420460 1004776 420512 1004828
rect 422668 1004776 422720 1004828
rect 497924 1004776 497976 1004828
rect 499672 1004776 499724 1004828
rect 555976 1004776 556028 1004828
rect 558184 1004776 558236 1004828
rect 106188 1004640 106240 1004692
rect 108488 1004640 108540 1004692
rect 149888 1004640 149940 1004692
rect 151728 1004640 151780 1004692
rect 161112 1004640 161164 1004692
rect 162952 1004640 163004 1004692
rect 209228 1004640 209280 1004692
rect 211160 1004640 211212 1004692
rect 305644 1004640 305696 1004692
rect 308128 1004640 308180 1004692
rect 315488 1004640 315540 1004692
rect 318064 1004640 318116 1004692
rect 364248 1004640 364300 1004692
rect 366364 1004640 366416 1004692
rect 432880 1004640 432932 1004692
rect 438124 1004640 438176 1004692
rect 557632 1004640 557684 1004692
rect 559564 1004640 559616 1004692
rect 560852 1004640 560904 1004692
rect 566464 1004640 566516 1004692
rect 570328 1004096 570380 1004148
rect 573364 1004096 573416 1004148
rect 513380 1004028 513432 1004080
rect 518900 1004028 518952 1004080
rect 247132 1003892 247184 1003944
rect 255320 1003892 255372 1003944
rect 424324 1003892 424376 1003944
rect 443644 1003892 443696 1003944
rect 558920 1003892 558972 1003944
rect 570788 1003892 570840 1003944
rect 300308 1003280 300360 1003332
rect 305276 1003280 305328 1003332
rect 553400 1003280 553452 1003332
rect 554596 1003280 554648 1003332
rect 299296 1003144 299348 1003196
rect 308956 1003144 309008 1003196
rect 253112 1002668 253164 1002720
rect 256148 1002668 256200 1002720
rect 424692 1002668 424744 1002720
rect 448980 1002668 449032 1002720
rect 97264 1002600 97316 1002652
rect 100300 1002600 100352 1002652
rect 553124 1002600 553176 1002652
rect 553768 1002600 553820 1002652
rect 558828 1002600 558880 1002652
rect 562508 1002600 562560 1002652
rect 246580 1002532 246632 1002584
rect 254124 1002532 254176 1002584
rect 429752 1002532 429804 1002584
rect 464988 1002532 465040 1002584
rect 98644 1002464 98696 1002516
rect 101956 1002464 102008 1002516
rect 202880 1002464 202932 1002516
rect 206376 1002464 206428 1002516
rect 509884 1002464 509936 1002516
rect 515404 1002464 515456 1002516
rect 560852 1002464 560904 1002516
rect 565084 1002464 565136 1002516
rect 97448 1002328 97500 1002380
rect 100300 1002328 100352 1002380
rect 100484 1002328 100536 1002380
rect 103152 1002328 103204 1002380
rect 107660 1002328 107712 1002380
rect 109500 1002328 109552 1002380
rect 148508 1002328 148560 1002380
rect 150900 1002328 150952 1002380
rect 251824 1002328 251876 1002380
rect 254492 1002328 254544 1002380
rect 261024 1002328 261076 1002380
rect 264244 1002328 264296 1002380
rect 357716 1002328 357768 1002380
rect 360844 1002328 360896 1002380
rect 501696 1002328 501748 1002380
rect 503720 1002328 503772 1002380
rect 560484 1002328 560536 1002380
rect 563060 1002328 563112 1002380
rect 98828 1002192 98880 1002244
rect 101128 1002192 101180 1002244
rect 105636 1002192 105688 1002244
rect 107844 1002192 107896 1002244
rect 108028 1002192 108080 1002244
rect 110420 1002192 110472 1002244
rect 155776 1002192 155828 1002244
rect 157340 1002192 157392 1002244
rect 205088 1002192 205140 1002244
rect 207204 1002192 207256 1002244
rect 254584 1002192 254636 1002244
rect 256516 1002192 256568 1002244
rect 260196 1002192 260248 1002244
rect 262864 1002192 262916 1002244
rect 303068 1002192 303120 1002244
rect 306104 1002192 306156 1002244
rect 308404 1002192 308456 1002244
rect 310612 1002192 310664 1002244
rect 500592 1002192 500644 1002244
rect 503352 1002192 503404 1002244
rect 504180 1002192 504232 1002244
rect 510068 1002192 510120 1002244
rect 558000 1002192 558052 1002244
rect 560944 1002192 560996 1002244
rect 553216 1002124 553268 1002176
rect 553952 1002124 554004 1002176
rect 96068 1002056 96120 1002108
rect 99104 1002056 99156 1002108
rect 100024 1002056 100076 1002108
rect 102324 1002056 102376 1002108
rect 103980 1002056 104032 1002108
rect 106464 1002056 106516 1002108
rect 106832 1002056 106884 1002108
rect 109040 1002056 109092 1002108
rect 109684 1002056 109736 1002108
rect 111800 1002056 111852 1002108
rect 148324 1002056 148376 1002108
rect 150900 1002056 150952 1002108
rect 152464 1002056 152516 1002108
rect 154580 1002056 154632 1002108
rect 157800 1002056 157852 1002108
rect 160100 1002056 160152 1002108
rect 206744 1002056 206796 1002108
rect 208584 1002056 208636 1002108
rect 210884 1002056 210936 1002108
rect 213184 1002056 213236 1002108
rect 253388 1002056 253440 1002108
rect 255320 1002056 255372 1002108
rect 259828 1002056 259880 1002108
rect 262220 1002056 262272 1002108
rect 263876 1002056 263928 1002108
rect 267004 1002056 267056 1002108
rect 300124 1002056 300176 1002108
rect 304080 1002056 304132 1002108
rect 355784 1002056 355836 1002108
rect 357716 1002056 357768 1002108
rect 423588 1002056 423640 1002108
rect 426348 1002056 426400 1002108
rect 502524 1002056 502576 1002108
rect 505744 1002056 505796 1002108
rect 560024 1002056 560076 1002108
rect 562324 1002056 562376 1002108
rect 95884 1001920 95936 1001972
rect 98276 1001920 98328 1001972
rect 99012 1001920 99064 1001972
rect 101128 1001920 101180 1001972
rect 106004 1001920 106056 1001972
rect 107752 1001920 107804 1001972
rect 146944 1001920 146996 1001972
rect 149244 1001920 149296 1001972
rect 156604 1001920 156656 1001972
rect 158720 1001920 158772 1001972
rect 202880 1001920 202932 1001972
rect 204168 1001920 204220 1001972
rect 205548 1001920 205600 1001972
rect 206284 1001920 206336 1001972
rect 207572 1001920 207624 1001972
rect 212540 1001920 212592 1001972
rect 214564 1001920 214616 1001972
rect 254768 1001920 254820 1001972
rect 256976 1001920 257028 1001972
rect 260196 1001920 260248 1001972
rect 260932 1001920 260984 1001972
rect 263508 1001920 263560 1001972
rect 265624 1001920 265676 1001972
rect 302884 1001920 302936 1001972
rect 306104 1001920 306156 1001972
rect 310152 1001920 310204 1001972
rect 311900 1001920 311952 1001972
rect 351828 1001920 351880 1001972
rect 354036 1001920 354088 1001972
rect 365904 1001920 365956 1001972
rect 369124 1001920 369176 1001972
rect 419448 1001920 419500 1001972
rect 421472 1001920 421524 1001972
rect 425520 1001920 425572 1001972
rect 500776 1001920 500828 1001972
rect 501328 1001920 501380 1001972
rect 504548 1001920 504600 1001972
rect 506848 1001920 506900 1001972
rect 558000 1001920 558052 1001972
rect 560300 1001920 560352 1001972
rect 561680 1001920 561732 1001972
rect 563704 1001920 563756 1001972
rect 428188 1001852 428240 1001904
rect 195152 1001716 195204 1001768
rect 439504 1001444 439556 1001496
rect 458180 1001444 458232 1001496
rect 425704 1001308 425756 1001360
rect 446404 1001308 446456 1001360
rect 353208 1001172 353260 1001224
rect 380900 1001172 380952 1001224
rect 423588 1001172 423640 1001224
rect 462228 1001172 462280 1001224
rect 497924 1001172 497976 1001224
rect 521292 1001172 521344 1001224
rect 550272 1001172 550324 1001224
rect 574100 1001172 574152 1001224
rect 298468 1000492 298520 1000544
rect 305828 1000492 305880 1000544
rect 499488 1000492 499540 1000544
rect 500316 1000492 500368 1000544
rect 503720 1000492 503772 1000544
rect 516876 1000492 516928 1000544
rect 617340 1000492 617392 1000544
rect 625436 1000492 625488 1000544
rect 567844 1000084 567896 1000136
rect 571340 1000084 571392 1000136
rect 558184 999948 558236 1000000
rect 565820 999948 565872 1000000
rect 93308 999744 93360 999796
rect 99012 999744 99064 999796
rect 246948 999744 247000 999796
rect 254768 999744 254820 999796
rect 590936 999268 590988 999320
rect 625068 999268 625120 999320
rect 618168 999132 618220 999184
rect 625620 999132 625672 999184
rect 507400 999064 507452 999116
rect 509240 999064 509292 999116
rect 553400 999064 553452 999116
rect 556344 999064 556396 999116
rect 505376 998928 505428 998980
rect 511448 998928 511500 998980
rect 200212 998792 200264 998844
rect 203892 998792 203944 998844
rect 356060 998792 356112 998844
rect 372160 998792 372212 998844
rect 373264 998792 373316 998844
rect 382648 998860 382700 998912
rect 440884 998792 440936 998844
rect 448520 998792 448572 998844
rect 378784 998724 378836 998776
rect 383568 998724 383620 998776
rect 196808 998656 196860 998708
rect 204352 998656 204404 998708
rect 351828 998656 351880 998708
rect 378600 998656 378652 998708
rect 446404 998656 446456 998708
rect 458364 998792 458416 998844
rect 462228 998792 462280 998844
rect 472256 998792 472308 998844
rect 500960 998792 501012 998844
rect 517520 998792 517572 998844
rect 458180 998656 458232 998708
rect 472440 998656 472492 998708
rect 507032 998656 507084 998708
rect 509884 998656 509936 998708
rect 510068 998656 510120 998708
rect 523868 998860 523920 998912
rect 556804 998656 556856 998708
rect 567476 998656 567528 998708
rect 92296 998520 92348 998572
rect 92848 998520 92900 998572
rect 196624 998520 196676 998572
rect 203524 998520 203576 998572
rect 355784 998520 355836 998572
rect 383292 998520 383344 998572
rect 445024 998520 445076 998572
rect 461584 998520 461636 998572
rect 463700 998520 463752 998572
rect 472624 998520 472676 998572
rect 502156 998520 502208 998572
rect 516692 998520 516744 998572
rect 516876 998520 516928 998572
rect 524052 998520 524104 998572
rect 553768 998520 553820 998572
rect 569132 998520 569184 998572
rect 247316 998452 247368 998504
rect 92296 998384 92348 998436
rect 100484 998384 100536 998436
rect 144000 998384 144052 998436
rect 155960 998384 156012 998436
rect 195704 998384 195756 998436
rect 204168 998384 204220 998436
rect 246764 998316 246816 998368
rect 252468 998316 252520 998368
rect 200396 998180 200448 998232
rect 203524 998180 203576 998232
rect 250444 998112 250496 998164
rect 253664 998112 253716 998164
rect 199384 998044 199436 998096
rect 202696 998044 202748 998096
rect 197544 997908 197596 997960
rect 201868 997908 201920 997960
rect 202144 997908 202196 997960
rect 205548 997908 205600 997960
rect 251180 997908 251232 997960
rect 253664 997908 253716 997960
rect 92664 997772 92716 997824
rect 121736 997772 121788 997824
rect 202328 997772 202380 997824
rect 204720 997772 204772 997824
rect 247868 997772 247920 997824
rect 252468 997772 252520 997824
rect 354588 998384 354640 998436
rect 383476 998384 383528 998436
rect 428188 998384 428240 998436
rect 472072 998384 472124 998436
rect 500776 998384 500828 998436
rect 523684 998384 523736 998436
rect 549168 998384 549220 998436
rect 564440 998384 564492 998436
rect 591120 998384 591172 998436
rect 617340 998384 617392 998436
rect 371884 998248 371936 998300
rect 372988 998248 373040 998300
rect 378600 998248 378652 998300
rect 382464 998248 382516 998300
rect 430856 998248 430908 998300
rect 433984 998248 434036 998300
rect 509056 998248 509108 998300
rect 514024 998248 514076 998300
rect 550548 998248 550600 998300
rect 552940 998248 552992 998300
rect 430028 998112 430080 998164
rect 432604 998112 432656 998164
rect 508228 998112 508280 998164
rect 511264 998112 511316 998164
rect 432052 997976 432104 998028
rect 436744 997976 436796 998028
rect 508228 997908 508280 997960
rect 510712 997908 510764 997960
rect 430028 997840 430080 997892
rect 432052 997840 432104 997892
rect 278228 997772 278280 997824
rect 377404 997772 377456 997824
rect 383108 997772 383160 997824
rect 591304 997772 591356 997824
rect 625804 997772 625856 997824
rect 143816 997704 143868 997756
rect 153936 997704 153988 997756
rect 298836 997704 298888 997756
rect 311900 997704 311952 997756
rect 358820 997704 358872 997756
rect 372344 997704 372396 997756
rect 431224 997704 431276 997756
rect 439688 997704 439740 997756
rect 488908 997704 488960 997756
rect 509240 997704 509292 997756
rect 509884 997704 509936 997756
rect 516876 997704 516928 997756
rect 92480 997636 92532 997688
rect 101588 997636 101640 997688
rect 109500 997636 109552 997688
rect 117228 997636 117280 997688
rect 246672 997636 246724 997688
rect 258080 997636 258132 997688
rect 569500 997636 569552 997688
rect 623688 997636 623740 997688
rect 144828 997568 144880 997620
rect 160100 997568 160152 997620
rect 299480 997568 299532 997620
rect 310520 997568 310572 997620
rect 365168 997568 365220 997620
rect 372528 997568 372580 997620
rect 433984 997568 434036 997620
rect 439872 997568 439924 997620
rect 489092 997568 489144 997620
rect 510712 997568 510764 997620
rect 113824 997500 113876 997552
rect 116952 997500 117004 997552
rect 550548 997500 550600 997552
rect 618168 997500 618220 997552
rect 432604 997432 432656 997484
rect 440056 997432 440108 997484
rect 500592 997432 500644 997484
rect 516692 997432 516744 997484
rect 540336 997364 540388 997416
rect 555424 997364 555476 997416
rect 200212 997228 200264 997280
rect 205088 997228 205140 997280
rect 552296 997228 552348 997280
rect 590384 997364 590436 997416
rect 573548 997228 573600 997280
rect 591304 997228 591356 997280
rect 160744 997160 160796 997212
rect 162952 997160 163004 997212
rect 399944 997092 399996 997144
rect 432052 997092 432104 997144
rect 571340 997092 571392 997144
rect 591120 997092 591172 997144
rect 144644 997024 144696 997076
rect 158720 997024 158772 997076
rect 197360 997024 197412 997076
rect 226340 997024 226392 997076
rect 320824 997024 320876 997076
rect 332600 997024 332652 997076
rect 448980 997024 449032 997076
rect 470508 997024 470560 997076
rect 498200 997024 498252 997076
rect 517704 997024 517756 997076
rect 565820 996888 565872 996940
rect 590568 996888 590620 996940
rect 553216 996752 553268 996804
rect 590568 996684 590620 996736
rect 564440 996616 564492 996668
rect 568856 996616 568908 996668
rect 143724 996344 143776 996396
rect 151268 996344 151320 996396
rect 298652 996344 298704 996396
rect 365168 996344 365220 996396
rect 262864 996276 262916 996328
rect 270408 996276 270460 996328
rect 556344 996276 556396 996328
rect 590384 996276 590436 996328
rect 195612 996208 195664 996260
rect 200672 996208 200724 996260
rect 171784 996072 171836 996124
rect 567476 996140 567528 996192
rect 590568 996140 590620 996192
rect 211160 996072 211212 996124
rect 229744 996072 229796 996124
rect 262220 996072 262272 996124
rect 269764 996072 269816 996124
rect 316040 996072 316092 996124
rect 366364 996072 366416 996124
rect 402244 996072 402296 996124
rect 511264 996072 511316 996124
rect 563060 996072 563112 996124
rect 170680 995936 170732 995988
rect 171232 995936 171284 995988
rect 195888 995936 195940 995988
rect 202512 995936 202564 995988
rect 213184 995936 213236 995988
rect 261116 995936 261168 995988
rect 264244 995936 264296 995988
rect 299204 995936 299256 995988
rect 364984 995936 365036 995988
rect 400864 995936 400916 995988
rect 522304 995936 522356 995988
rect 560300 995936 560352 995988
rect 92664 995800 92716 995852
rect 97448 995800 97500 995852
rect 140780 995800 140832 995852
rect 144000 995800 144052 995852
rect 169392 995800 169444 995852
rect 171508 995800 171560 995852
rect 211804 995800 211856 995852
rect 260932 995800 260984 995852
rect 360844 995800 360896 995852
rect 399852 995800 399904 995852
rect 517520 995800 517572 995852
rect 523316 995800 523368 995852
rect 92480 995528 92532 995580
rect 98828 995528 98880 995580
rect 143724 995528 143776 995580
rect 145748 995528 145800 995580
rect 171048 995528 171100 995580
rect 297824 995528 297876 995580
rect 298468 995528 298520 995580
rect 383108 995528 383160 995580
rect 385684 995528 385736 995580
rect 472440 995528 472492 995580
rect 473360 995528 473412 995580
rect 623688 995528 623740 995580
rect 626540 995528 626592 995580
rect 194876 995460 194928 995512
rect 195704 995460 195756 995512
rect 246212 995460 246264 995512
rect 247132 995460 247184 995512
rect 507032 995460 507084 995512
rect 527916 995460 527968 995512
rect 629208 995460 629260 995512
rect 631508 995460 631560 995512
rect 380164 995392 380216 995444
rect 383108 995392 383160 995444
rect 383292 995392 383344 995444
rect 388628 995392 388680 995444
rect 389088 995392 389140 995444
rect 389732 995392 389784 995444
rect 415400 995392 415452 995444
rect 171692 995277 171744 995329
rect 180708 995324 180760 995376
rect 202144 995324 202196 995376
rect 236552 995324 236604 995376
rect 251824 995324 251876 995376
rect 293592 995324 293644 995376
rect 295984 995324 296036 995376
rect 296168 995324 296220 995376
rect 298100 995324 298152 995376
rect 395252 995324 395304 995376
rect 399852 995324 399904 995376
rect 382188 995256 382240 995308
rect 386328 995256 386380 995308
rect 386512 995256 386564 995308
rect 171508 995165 171560 995217
rect 182962 995188 183014 995240
rect 208584 995188 208636 995240
rect 234390 995188 234442 995240
rect 259460 995188 259512 995240
rect 285956 995188 286008 995240
rect 309140 995188 309192 995240
rect 398840 995188 398892 995240
rect 416136 995235 416188 995287
rect 362224 995120 362276 995172
rect 388352 995120 388404 995172
rect 528928 995120 528980 995172
rect 532884 995120 532936 995172
rect 533344 995120 533396 995172
rect 534080 995120 534132 995172
rect 625252 995120 625304 995172
rect 633992 995120 634044 995172
rect 171232 995053 171284 995105
rect 180156 995052 180208 995104
rect 207020 995052 207072 995104
rect 231584 995052 231636 995104
rect 257344 995052 257396 995104
rect 284116 995052 284168 995104
rect 308404 995052 308456 995104
rect 454684 995052 454736 995104
rect 485964 995052 486016 995104
rect 505744 995052 505796 995104
rect 528744 995052 528796 995104
rect 569132 995052 569184 995104
rect 625114 995052 625166 995104
rect 638868 995052 638920 995104
rect 640800 995052 640852 995104
rect 660304 995095 660356 995147
rect 358084 994984 358136 995036
rect 393320 994984 393372 995036
rect 181444 994916 181496 994968
rect 206284 994916 206336 994968
rect 232872 994916 232924 994968
rect 255964 994916 256016 994968
rect 287152 994916 287204 994968
rect 304264 994916 304316 994968
rect 420460 994916 420512 994968
rect 80152 994780 80204 994832
rect 106464 994780 106516 994832
rect 129740 994780 129792 994832
rect 137100 994780 137152 994832
rect 137284 994780 137336 994832
rect 77668 994644 77720 994696
rect 100024 994644 100076 994696
rect 129096 994644 129148 994696
rect 151084 994644 151136 994696
rect 170496 994712 170548 994764
rect 171232 994829 171284 994881
rect 363604 994848 363656 994900
rect 397644 994848 397696 994900
rect 461584 994780 461636 994832
rect 490012 994780 490064 994832
rect 496728 994780 496780 994832
rect 513656 994780 513708 994832
rect 513840 994780 513892 994832
rect 539232 994780 539284 994832
rect 551928 994780 551980 994832
rect 634820 994780 634872 994832
rect 171048 994712 171100 994764
rect 295064 994712 295116 994764
rect 376024 994712 376076 994764
rect 393964 994712 394016 994764
rect 157340 994644 157392 994696
rect 419448 994644 419500 994696
rect 660304 994644 660356 994696
rect 170680 994576 170732 994628
rect 250444 994576 250496 994628
rect 283472 994576 283524 994628
rect 305644 994576 305696 994628
rect 372988 994576 373040 994628
rect 397000 994576 397052 994628
rect 660764 994576 660816 994628
rect 81348 994508 81400 994560
rect 98644 994508 98696 994560
rect 132408 994508 132460 994560
rect 149888 994508 149940 994560
rect 470508 994508 470560 994560
rect 482284 994508 482336 994560
rect 482928 994508 482980 994560
rect 489828 994508 489880 994560
rect 502340 994508 502392 994560
rect 513840 994508 513892 994560
rect 514208 994508 514260 994560
rect 523500 994508 523552 994560
rect 523684 994508 523736 994560
rect 534356 994508 534408 994560
rect 573364 994508 573416 994560
rect 590936 994508 590988 994560
rect 591304 994508 591356 994560
rect 639052 994508 639104 994560
rect 660948 994508 661000 994560
rect 170864 994440 170916 994492
rect 298836 994440 298888 994492
rect 80704 994372 80756 994424
rect 94504 994372 94556 994424
rect 128452 994372 128504 994424
rect 137284 994372 137336 994424
rect 471428 994372 471480 994424
rect 484584 994372 484636 994424
rect 500316 994372 500368 994424
rect 534080 994372 534132 994424
rect 568856 994372 568908 994424
rect 639512 994372 639564 994424
rect 184480 994304 184532 994356
rect 191104 994304 191156 994356
rect 191748 994304 191800 994356
rect 197360 994304 197412 994356
rect 137100 994236 137152 994288
rect 144644 994236 144696 994288
rect 226340 994236 226392 994288
rect 251456 994236 251508 994288
rect 278228 994236 278280 994288
rect 316408 994236 316460 994288
rect 365168 994236 365220 994288
rect 381176 994236 381228 994288
rect 414480 994236 414532 994288
rect 446128 994236 446180 994288
rect 472072 994236 472124 994288
rect 477960 994236 478012 994288
rect 513656 994236 513708 994288
rect 514208 994236 514260 994288
rect 517704 994236 517756 994288
rect 523684 994236 523736 994288
rect 139216 994100 139268 994152
rect 142068 994100 142120 994152
rect 169392 994100 169444 994152
rect 247868 994100 247920 994152
rect 295064 994100 295116 994152
rect 300124 994100 300176 994152
rect 523500 994100 523552 994152
rect 538036 994236 538088 994288
rect 570604 994236 570656 994288
rect 591304 994236 591356 994288
rect 625436 994236 625488 994288
rect 630864 994236 630916 994288
rect 574100 994032 574152 994084
rect 141884 993964 141936 994016
rect 142344 993964 142396 994016
rect 191104 993964 191156 994016
rect 196808 993964 196860 994016
rect 232228 993964 232280 994016
rect 254584 993964 254636 994016
rect 569316 993896 569368 993948
rect 171232 993760 171284 993812
rect 195520 993760 195572 993812
rect 521292 993760 521344 993812
rect 660948 993760 661000 993812
rect 142160 993692 142212 993744
rect 143908 993692 143960 993744
rect 170496 993624 170548 993676
rect 197544 993624 197596 993676
rect 517060 993624 517112 993676
rect 660764 993624 660816 993676
rect 188160 993488 188212 993540
rect 195888 993488 195940 993540
rect 50344 993148 50396 993200
rect 107752 993148 107804 993200
rect 44824 993012 44876 993064
rect 109040 993012 109092 993064
rect 318064 993012 318116 993064
rect 349160 993012 349212 993064
rect 562508 993012 562560 993064
rect 660304 993012 660356 993064
rect 54484 992876 54536 992928
rect 148324 992876 148376 992928
rect 319444 992876 319496 992928
rect 364984 992876 365036 992928
rect 560944 992876 560996 992928
rect 667204 992876 667256 992928
rect 47584 991720 47636 991772
rect 96068 991720 96120 991772
rect 51724 991584 51776 991636
rect 110420 991584 110472 991636
rect 138296 991584 138348 991636
rect 163136 991584 163188 991636
rect 369124 991584 369176 991636
rect 414112 991584 414164 991636
rect 55864 991448 55916 991500
rect 146944 991448 146996 991500
rect 267004 991448 267056 991500
rect 284300 991448 284352 991500
rect 367744 991448 367796 991500
rect 430304 991448 430356 991500
rect 435364 991448 435416 991500
rect 478972 991448 479024 991500
rect 559564 991448 559616 991500
rect 658924 991448 658976 991500
rect 214564 991176 214616 991228
rect 219440 991176 219492 991228
rect 164884 990836 164936 990888
rect 170772 990836 170824 990888
rect 265624 990836 265676 990888
rect 267648 990836 267700 990888
rect 572812 990836 572864 990888
rect 576308 990836 576360 990888
rect 53288 990224 53340 990276
rect 95884 990224 95936 990276
rect 48964 990088 49016 990140
rect 108120 990088 108172 990140
rect 512644 990088 512696 990140
rect 543832 990088 543884 990140
rect 562324 990088 562376 990140
rect 668584 990088 668636 990140
rect 563704 987368 563756 987420
rect 608784 987368 608836 987420
rect 203156 986620 203208 986672
rect 204904 986620 204956 986672
rect 89628 986076 89680 986128
rect 111800 986076 111852 986128
rect 438124 986076 438176 986128
rect 462780 986076 462832 986128
rect 515404 986076 515456 986128
rect 527640 986076 527692 986128
rect 566464 986076 566516 986128
rect 592500 986076 592552 986128
rect 73436 985940 73488 985992
rect 102784 985940 102836 985992
rect 215944 985940 215996 985992
rect 235632 985940 235684 985992
rect 268384 985940 268436 985992
rect 300492 985940 300544 985992
rect 370504 985940 370556 985992
rect 397828 985940 397880 985992
rect 436744 985940 436796 985992
rect 495164 985940 495216 985992
rect 514024 985940 514076 985992
rect 560116 985940 560168 985992
rect 565084 985940 565136 985992
rect 624976 985940 625028 985992
rect 154488 985668 154540 985720
rect 160744 985668 160796 985720
rect 43444 975672 43496 975724
rect 62120 975672 62172 975724
rect 651656 975672 651708 975724
rect 664444 975672 664496 975724
rect 46204 961868 46256 961920
rect 62120 961868 62172 961920
rect 651472 961868 651524 961920
rect 665824 961868 665876 961920
rect 36544 952348 36596 952400
rect 41696 952348 41748 952400
rect 33784 951464 33836 951516
rect 41512 951464 41564 951516
rect 675852 949424 675904 949476
rect 682384 949424 682436 949476
rect 652208 948064 652260 948116
rect 663064 948064 663116 948116
rect 676036 947996 676088 948048
rect 681004 947996 681056 948048
rect 45560 945956 45612 946008
rect 62120 945956 62172 946008
rect 28724 945276 28776 945328
rect 31760 945276 31812 945328
rect 35808 942556 35860 942608
rect 41696 942556 41748 942608
rect 35808 941196 35860 941248
rect 41420 941196 41472 941248
rect 35808 939768 35860 939820
rect 41604 939768 41656 939820
rect 651472 936980 651524 937032
rect 661684 936980 661736 937032
rect 675852 928752 675904 928804
rect 683120 928752 683172 928804
rect 53104 923244 53156 923296
rect 62120 923244 62172 923296
rect 651472 921816 651524 921868
rect 661684 921816 661736 921868
rect 50344 909440 50396 909492
rect 62120 909440 62172 909492
rect 652392 909440 652444 909492
rect 663064 909440 663116 909492
rect 47768 896996 47820 897048
rect 62120 896996 62172 897048
rect 651472 895636 651524 895688
rect 671344 895636 671396 895688
rect 42846 892440 42898 892492
rect 43076 892304 43128 892356
rect 42938 892202 42990 892254
rect 44088 891896 44140 891948
rect 651656 881832 651708 881884
rect 664444 881832 664496 881884
rect 46204 870816 46256 870868
rect 62120 870816 62172 870868
rect 651472 869388 651524 869440
rect 658924 869388 658976 869440
rect 652392 855584 652444 855636
rect 664444 855584 664496 855636
rect 54484 844568 54536 844620
rect 62120 844568 62172 844620
rect 55864 832124 55916 832176
rect 62120 832124 62172 832176
rect 651472 829404 651524 829456
rect 660304 829404 660356 829456
rect 47584 818320 47636 818372
rect 62120 818320 62172 818372
rect 35808 817028 35860 817080
rect 41696 817028 41748 817080
rect 35808 815600 35860 815652
rect 41420 815600 41472 815652
rect 651472 815600 651524 815652
rect 669964 815600 670016 815652
rect 35808 814240 35860 814292
rect 41604 814240 41656 814292
rect 41328 811452 41380 811504
rect 41696 811452 41748 811504
rect 40592 808256 40644 808308
rect 41604 808256 41656 808308
rect 50344 805944 50396 805996
rect 62120 805944 62172 805996
rect 651472 803224 651524 803276
rect 667204 803156 667256 803208
rect 35164 802408 35216 802460
rect 41696 802408 41748 802460
rect 35900 802272 35952 802324
rect 41696 802272 41748 802324
rect 651472 789352 651524 789404
rect 668584 789352 668636 789404
rect 651472 775548 651524 775600
rect 668768 775548 668820 775600
rect 35808 772828 35860 772880
rect 41696 772828 41748 772880
rect 35808 768952 35860 769004
rect 41328 768952 41380 769004
rect 35624 768816 35676 768868
rect 41696 768816 41748 768868
rect 35440 768680 35492 768732
rect 40040 768680 40092 768732
rect 35808 767524 35860 767576
rect 37924 767456 37976 767508
rect 35808 767320 35860 767372
rect 36544 767320 36596 767372
rect 48964 767320 49016 767372
rect 62120 767320 62172 767372
rect 37096 763240 37148 763292
rect 39304 763240 39356 763292
rect 651472 763240 651524 763292
rect 660304 763172 660356 763224
rect 37924 759092 37976 759144
rect 40868 759092 40920 759144
rect 35164 758956 35216 759008
rect 40316 758956 40368 759008
rect 31024 758276 31076 758328
rect 40592 758276 40644 758328
rect 676036 757120 676088 757172
rect 683120 757120 683172 757172
rect 51724 753516 51776 753568
rect 62120 753516 62172 753568
rect 651472 749368 651524 749420
rect 665824 749368 665876 749420
rect 54484 741072 54536 741124
rect 62120 741072 62172 741124
rect 652576 735564 652628 735616
rect 671344 735564 671396 735616
rect 673552 732096 673604 732148
rect 674012 732096 674064 732148
rect 35624 730192 35676 730244
rect 41696 730192 41748 730244
rect 35808 730056 35860 730108
rect 41512 730056 41564 730108
rect 673828 728560 673880 728612
rect 673368 728424 673420 728476
rect 673000 728084 673052 728136
rect 674150 728084 674202 728136
rect 41328 726044 41380 726096
rect 41696 726044 41748 726096
rect 41328 724480 41380 724532
rect 41696 724480 41748 724532
rect 677324 724208 677376 724260
rect 683304 724208 683356 724260
rect 651472 723120 651524 723172
rect 663064 723120 663116 723172
rect 31024 716864 31076 716916
rect 41512 716864 41564 716916
rect 33784 715640 33836 715692
rect 39856 715640 39908 715692
rect 33048 715504 33100 715556
rect 40224 715504 40276 715556
rect 36544 715300 36596 715352
rect 41696 715300 41748 715352
rect 50344 714824 50396 714876
rect 62120 714824 62172 714876
rect 652576 709316 652628 709368
rect 664444 709316 664496 709368
rect 672448 707208 672500 707260
rect 673000 707208 673052 707260
rect 55864 701020 55916 701072
rect 62120 701020 62172 701072
rect 652392 696940 652444 696992
rect 661684 696940 661736 696992
rect 53104 688644 53156 688696
rect 62120 688644 62172 688696
rect 35808 687216 35860 687268
rect 41696 687216 41748 687268
rect 44548 685040 44600 685092
rect 45376 685040 45428 685092
rect 35808 683136 35860 683188
rect 41696 683136 41748 683188
rect 35624 681844 35676 681896
rect 41696 681844 41748 681896
rect 35808 681708 35860 681760
rect 41328 681708 41380 681760
rect 35440 681028 35492 681080
rect 41604 681028 41656 681080
rect 35624 680620 35676 680672
rect 36544 680620 36596 680672
rect 35808 680348 35860 680400
rect 37924 680348 37976 680400
rect 51724 674840 51776 674892
rect 62120 674840 62172 674892
rect 35164 672732 35216 672784
rect 38936 672732 38988 672784
rect 36544 672052 36596 672104
rect 39580 672052 39632 672104
rect 651472 669332 651524 669384
rect 661868 669332 661920 669384
rect 671068 666204 671120 666256
rect 673368 666204 673420 666256
rect 47584 662396 47636 662448
rect 62120 662396 62172 662448
rect 651472 656888 651524 656940
rect 670148 656888 670200 656940
rect 54484 647844 54536 647896
rect 62120 647844 62172 647896
rect 651472 643084 651524 643136
rect 668584 643084 668636 643136
rect 35808 639140 35860 639192
rect 41696 639072 41748 639124
rect 35808 638936 35860 638988
rect 40040 638936 40092 638988
rect 35808 637576 35860 637628
rect 41328 637576 41380 637628
rect 51724 636216 51776 636268
rect 62120 636216 62172 636268
rect 44916 635944 44968 635996
rect 45100 635672 45152 635724
rect 32404 629892 32456 629944
rect 41696 629892 41748 629944
rect 651472 629280 651524 629332
rect 667204 629280 667256 629332
rect 670976 627104 671028 627156
rect 672172 627104 672224 627156
rect 672908 626696 672960 626748
rect 673552 626696 673604 626748
rect 673092 626560 673144 626612
rect 675852 626560 675904 626612
rect 676496 626560 676548 626612
rect 672908 626356 672960 626408
rect 44088 626084 44140 626136
rect 44916 626084 44968 626136
rect 48964 623772 49016 623824
rect 62120 623772 62172 623824
rect 651472 616836 651524 616888
rect 660304 616836 660356 616888
rect 671436 616156 671488 616208
rect 671896 616156 671948 616208
rect 43536 612892 43588 612944
rect 43371 612688 43423 612740
rect 43720 612484 43772 612536
rect 43582 612280 43634 612332
rect 46388 612348 46440 612400
rect 45560 612144 45612 612196
rect 46940 611668 46992 611720
rect 44180 611532 44232 611584
rect 45744 611260 45796 611312
rect 47216 611056 47268 611108
rect 45376 610852 45428 610904
rect 44502 610580 44554 610632
rect 56048 608608 56100 608660
rect 62120 608608 62172 608660
rect 651472 603100 651524 603152
rect 664628 603100 664680 603152
rect 48964 597524 49016 597576
rect 62120 597524 62172 597576
rect 40316 596164 40368 596216
rect 41696 596164 41748 596216
rect 40868 596028 40920 596080
rect 41328 596028 41380 596080
rect 40684 593240 40736 593292
rect 41604 593240 41656 593292
rect 40960 593036 41012 593088
rect 41604 593036 41656 593088
rect 675944 591336 675996 591388
rect 679624 591336 679676 591388
rect 676128 591200 676180 591252
rect 682384 591200 682436 591252
rect 651472 590656 651524 590708
rect 662052 590656 662104 590708
rect 35164 585896 35216 585948
rect 40500 585896 40552 585948
rect 32404 585760 32456 585812
rect 39488 585760 39540 585812
rect 36544 585148 36596 585200
rect 41420 585148 41472 585200
rect 51724 583720 51776 583772
rect 62120 583720 62172 583772
rect 672356 579504 672408 579556
rect 673000 579504 673052 579556
rect 651472 576852 651524 576904
rect 665824 576852 665876 576904
rect 672448 572704 672500 572756
rect 672908 572704 672960 572756
rect 679624 571276 679676 571328
rect 683120 571276 683172 571328
rect 672264 567264 672316 567316
rect 672908 567264 672960 567316
rect 651656 563048 651708 563100
rect 658924 563048 658976 563100
rect 55864 558084 55916 558136
rect 62120 558084 62172 558136
rect 35808 557540 35860 557592
rect 41512 557540 41564 557592
rect 35808 554752 35860 554804
rect 41696 554752 41748 554804
rect 35808 553528 35860 553580
rect 41420 553528 41472 553580
rect 35624 553392 35676 553444
rect 41696 553392 41748 553444
rect 41052 552100 41104 552152
rect 41696 552032 41748 552084
rect 41236 550604 41288 550656
rect 41696 550604 41748 550656
rect 651472 550604 651524 550656
rect 660304 550604 660356 550656
rect 41328 547884 41380 547936
rect 41696 547884 41748 547936
rect 675852 547612 675904 547664
rect 678244 547612 678296 547664
rect 31760 547408 31812 547460
rect 37096 547408 37148 547460
rect 47584 545096 47636 545148
rect 62120 545096 62172 545148
rect 33784 542988 33836 543040
rect 41512 542988 41564 543040
rect 37096 542308 37148 542360
rect 41696 542308 41748 542360
rect 651472 536800 651524 536852
rect 669964 536800 670016 536852
rect 671252 533128 671304 533180
rect 670884 532856 670936 532908
rect 50344 532720 50396 532772
rect 62120 532720 62172 532772
rect 675852 532244 675904 532296
rect 676588 532244 676640 532296
rect 651840 522996 651892 523048
rect 661868 522996 661920 523048
rect 54484 518916 54536 518968
rect 62120 518916 62172 518968
rect 675852 518780 675904 518832
rect 677876 518780 677928 518832
rect 651472 510620 651524 510672
rect 659108 510620 659160 510672
rect 46204 506472 46256 506524
rect 62120 506472 62172 506524
rect 675852 503616 675904 503668
rect 679624 503616 679676 503668
rect 676036 503480 676088 503532
rect 682384 503480 682436 503532
rect 675852 502324 675904 502376
rect 676864 502324 676916 502376
rect 676036 500896 676088 500948
rect 681004 500896 681056 500948
rect 651472 496816 651524 496868
rect 663248 496816 663300 496868
rect 676036 492668 676088 492720
rect 683396 492668 683448 492720
rect 48964 491920 49016 491972
rect 62120 491920 62172 491972
rect 651472 484440 651524 484492
rect 667204 484372 667256 484424
rect 51724 480224 51776 480276
rect 62120 480224 62172 480276
rect 651472 470568 651524 470620
rect 665824 470568 665876 470620
rect 51908 466420 51960 466472
rect 62120 466420 62172 466472
rect 652392 456764 652444 456816
rect 661684 456764 661736 456816
rect 673948 456424 674000 456476
rect 673828 456016 673880 456068
rect 673460 455812 673512 455864
rect 673598 455608 673650 455660
rect 673506 455336 673558 455388
rect 673388 455132 673440 455184
rect 671068 454996 671120 455048
rect 673164 454792 673216 454844
rect 673046 454588 673098 454640
rect 672954 454316 673006 454368
rect 53104 454044 53156 454096
rect 62120 454044 62172 454096
rect 672816 454044 672868 454096
rect 672264 453908 672316 453960
rect 651472 444456 651524 444508
rect 668584 444388 668636 444440
rect 50528 440240 50580 440292
rect 62120 440240 62172 440292
rect 651472 430584 651524 430636
rect 671344 430584 671396 430636
rect 54484 427796 54536 427848
rect 62120 427796 62172 427848
rect 41328 423648 41380 423700
rect 41696 423648 41748 423700
rect 651840 416780 651892 416832
rect 663064 416780 663116 416832
rect 47584 415420 47636 415472
rect 62120 415420 62172 415472
rect 36544 415352 36596 415404
rect 41696 415352 41748 415404
rect 651472 404336 651524 404388
rect 664444 404336 664496 404388
rect 55864 401616 55916 401668
rect 62120 401616 62172 401668
rect 675852 395700 675904 395752
rect 676404 395700 676456 395752
rect 652576 390532 652628 390584
rect 658924 390532 658976 390584
rect 47768 389240 47820 389292
rect 62120 389240 62172 389292
rect 41144 387064 41196 387116
rect 41696 387064 41748 387116
rect 41328 382372 41380 382424
rect 41512 382372 41564 382424
rect 35808 379516 35860 379568
rect 41696 379516 41748 379568
rect 40224 378496 40276 378548
rect 41696 378496 41748 378548
rect 35808 375368 35860 375420
rect 41696 375368 41748 375420
rect 51724 375368 51776 375420
rect 62120 375368 62172 375420
rect 37924 372580 37976 372632
rect 41696 372580 41748 372632
rect 651656 364352 651708 364404
rect 661868 364352 661920 364404
rect 46388 362924 46440 362976
rect 62120 362924 62172 362976
rect 45008 355784 45060 355836
rect 45652 355784 45704 355836
rect 44640 355648 44692 355700
rect 44575 354832 44627 354884
rect 44575 354628 44627 354680
rect 44799 354424 44851 354476
rect 44686 354288 44738 354340
rect 45652 354016 45704 354068
rect 45928 353744 45980 353796
rect 45560 353200 45612 353252
rect 651472 350548 651524 350600
rect 667388 350548 667440 350600
rect 28908 345040 28960 345092
rect 40224 345040 40276 345092
rect 35808 339464 35860 339516
rect 37924 339464 37976 339516
rect 35808 338104 35860 338156
rect 36544 338104 36596 338156
rect 651472 338104 651524 338156
rect 667572 338104 667624 338156
rect 46204 336744 46256 336796
rect 62120 336744 62172 336796
rect 651472 324300 651524 324352
rect 667020 324300 667072 324352
rect 53288 322940 53340 322992
rect 62120 322940 62172 322992
rect 54484 310496 54536 310548
rect 62120 310496 62172 310548
rect 651472 310496 651524 310548
rect 667204 310496 667256 310548
rect 45468 298120 45520 298172
rect 62120 298120 62172 298172
rect 675852 298052 675904 298104
rect 678980 298052 679032 298104
rect 676128 297848 676180 297900
rect 681004 297848 681056 297900
rect 41328 285064 41380 285116
rect 41696 285064 41748 285116
rect 32404 284928 32456 284980
rect 41696 284928 41748 284980
rect 651472 284316 651524 284368
rect 667756 284316 667808 284368
rect 522396 276360 522448 276412
rect 526904 276360 526956 276412
rect 522212 276224 522264 276276
rect 530492 276224 530544 276276
rect 524880 276088 524932 276140
rect 88340 275952 88392 276004
rect 143356 275952 143408 276004
rect 156880 275952 156932 276004
rect 193864 275952 193916 276004
rect 201776 275952 201828 276004
rect 222108 275952 222160 276004
rect 389180 275952 389232 276004
rect 393320 275952 393372 276004
rect 400588 275952 400640 276004
rect 415768 275952 415820 276004
rect 427820 275952 427872 276004
rect 443000 275952 443052 276004
rect 443736 275952 443788 276004
rect 453580 275952 453632 276004
rect 456984 275952 457036 276004
rect 486700 275952 486752 276004
rect 486884 275952 486936 276004
rect 495164 275952 495216 276004
rect 495440 275952 495492 276004
rect 504548 275952 504600 276004
rect 504916 275952 504968 276004
rect 507032 275952 507084 276004
rect 508044 275952 508096 276004
rect 514024 275952 514076 276004
rect 95424 275816 95476 275868
rect 104808 275816 104860 275868
rect 113180 275816 113232 275868
rect 169944 275816 169996 275868
rect 181720 275816 181772 275868
rect 218888 275816 218940 275868
rect 393596 275816 393648 275868
rect 412272 275816 412324 275868
rect 415308 275816 415360 275868
rect 425244 275816 425296 275868
rect 432972 275816 433024 275868
rect 487896 275816 487948 275868
rect 488908 275816 488960 275868
rect 492588 275816 492640 275868
rect 498200 275816 498252 275868
rect 505652 275816 505704 275868
rect 507216 275816 507268 275868
rect 512736 275816 512788 275868
rect 512920 275816 512972 275868
rect 519820 275952 519872 276004
rect 520004 275952 520056 276004
rect 515496 275816 515548 275868
rect 81256 275680 81308 275732
rect 88984 275680 89036 275732
rect 103704 275680 103756 275732
rect 160100 275680 160152 275732
rect 178132 275680 178184 275732
rect 216864 275680 216916 275732
rect 299940 275680 299992 275732
rect 300768 275680 300820 275732
rect 370504 275680 370556 275732
rect 388628 275680 388680 275732
rect 410064 275680 410116 275732
rect 428832 275680 428884 275732
rect 429200 275680 429252 275732
rect 446496 275680 446548 275732
rect 446772 275680 446824 275732
rect 502064 275680 502116 275732
rect 76472 275544 76524 275596
rect 86868 275544 86920 275596
rect 96620 275544 96672 275596
rect 156604 275544 156656 275596
rect 163964 275544 164016 275596
rect 202144 275544 202196 275596
rect 221924 275544 221976 275596
rect 233884 275544 233936 275596
rect 236092 275544 236144 275596
rect 251088 275544 251140 275596
rect 350724 275544 350776 275596
rect 361396 275544 361448 275596
rect 362224 275544 362276 275596
rect 385040 275544 385092 275596
rect 388168 275544 388220 275596
rect 418160 275544 418212 275596
rect 418344 275544 418396 275596
rect 435916 275544 435968 275596
rect 449164 275544 449216 275596
rect 509148 275680 509200 275732
rect 512184 275680 512236 275732
rect 516232 275680 516284 275732
rect 516784 275816 516836 275868
rect 604920 275952 604972 276004
rect 524880 275816 524932 275868
rect 612004 275816 612056 275868
rect 519176 275680 519228 275732
rect 519360 275680 519412 275732
rect 522212 275680 522264 275732
rect 530308 275680 530360 275732
rect 85948 275408 86000 275460
rect 146760 275408 146812 275460
rect 160468 275408 160520 275460
rect 167736 275408 167788 275460
rect 171048 275408 171100 275460
rect 210792 275408 210844 275460
rect 218336 275408 218388 275460
rect 237472 275408 237524 275460
rect 244372 275408 244424 275460
rect 254584 275408 254636 275460
rect 260932 275408 260984 275460
rect 273536 275408 273588 275460
rect 273904 275408 273956 275460
rect 282920 275408 282972 275460
rect 326436 275408 326488 275460
rect 335360 275408 335412 275460
rect 341524 275408 341576 275460
rect 354312 275408 354364 275460
rect 298744 275340 298796 275392
rect 300032 275340 300084 275392
rect 70584 275272 70636 275324
rect 140136 275272 140188 275324
rect 142712 275272 142764 275324
rect 183468 275272 183520 275324
rect 186412 275272 186464 275324
rect 187792 275272 187844 275324
rect 188804 275272 188856 275324
rect 222844 275272 222896 275324
rect 225420 275272 225472 275324
rect 245108 275272 245160 275324
rect 250260 275272 250312 275324
rect 266360 275272 266412 275324
rect 266820 275272 266872 275324
rect 276664 275272 276716 275324
rect 284576 275272 284628 275324
rect 290096 275272 290148 275324
rect 329472 275272 329524 275324
rect 338948 275272 339000 275324
rect 74080 275136 74132 275188
rect 77208 275136 77260 275188
rect 110788 275136 110840 275188
rect 162124 275136 162176 275188
rect 338948 275136 339000 275188
rect 353116 275272 353168 275324
rect 353944 275272 353996 275324
rect 360200 275408 360252 275460
rect 363052 275408 363104 275460
rect 367284 275408 367336 275460
rect 369124 275408 369176 275460
rect 377956 275408 378008 275460
rect 382004 275408 382056 275460
rect 414572 275408 414624 275460
rect 416412 275408 416464 275460
rect 463056 275408 463108 275460
rect 467656 275408 467708 275460
rect 519544 275544 519596 275596
rect 519728 275544 519780 275596
rect 522396 275544 522448 275596
rect 530860 275680 530912 275732
rect 619088 275680 619140 275732
rect 536840 275544 536892 275596
rect 537024 275544 537076 275596
rect 537760 275544 537812 275596
rect 537944 275544 537996 275596
rect 626172 275544 626224 275596
rect 504548 275408 504600 275460
rect 538220 275408 538272 275460
rect 356336 275272 356388 275324
rect 368480 275272 368532 275324
rect 375104 275272 375156 275324
rect 403992 275272 404044 275324
rect 411260 275272 411312 275324
rect 455972 275272 456024 275324
rect 420920 275136 420972 275188
rect 434720 275136 434772 275188
rect 437480 275136 437532 275188
rect 450084 275136 450136 275188
rect 455880 275136 455932 275188
rect 512184 275272 512236 275324
rect 456800 275136 456852 275188
rect 467840 275136 467892 275188
rect 468208 275136 468260 275188
rect 494980 275136 495032 275188
rect 495164 275136 495216 275188
rect 519360 275272 519412 275324
rect 519544 275272 519596 275324
rect 537576 275272 537628 275324
rect 537760 275272 537812 275324
rect 540980 275408 541032 275460
rect 541164 275408 541216 275460
rect 544660 275408 544712 275460
rect 544844 275408 544896 275460
rect 546040 275408 546092 275460
rect 546224 275408 546276 275460
rect 641628 275408 641680 275460
rect 538680 275272 538732 275324
rect 633348 275272 633400 275324
rect 224224 275068 224276 275120
rect 226156 275068 226208 275120
rect 294052 275068 294104 275120
rect 295156 275068 295208 275120
rect 135628 275000 135680 275052
rect 182088 275000 182140 275052
rect 449900 275000 449952 275052
rect 460664 275000 460716 275052
rect 494704 275000 494756 275052
rect 498568 275000 498620 275052
rect 505100 275000 505152 275052
rect 506848 275000 506900 275052
rect 507032 275000 507084 275052
rect 590752 275136 590804 275188
rect 611360 275136 611412 275188
rect 616788 275136 616840 275188
rect 619180 275136 619232 275188
rect 623872 275136 623924 275188
rect 514024 275000 514076 275052
rect 583668 275000 583720 275052
rect 71780 274932 71832 274984
rect 73804 274932 73856 274984
rect 277492 274932 277544 274984
rect 284300 274932 284352 274984
rect 129648 274864 129700 274916
rect 136548 274864 136600 274916
rect 149796 274864 149848 274916
rect 185584 274864 185636 274916
rect 289268 274864 289320 274916
rect 293408 274864 293460 274916
rect 470968 274864 471020 274916
rect 523132 274864 523184 274916
rect 523316 274864 523368 274916
rect 597836 274864 597888 274916
rect 283380 274796 283432 274848
rect 289084 274796 289136 274848
rect 403992 274796 404044 274848
rect 407488 274796 407540 274848
rect 426256 274796 426308 274848
rect 432328 274796 432380 274848
rect 106004 274728 106056 274780
rect 110420 274728 110472 274780
rect 140320 274728 140372 274780
rect 144644 274728 144696 274780
rect 146208 274728 146260 274780
rect 149888 274728 149940 274780
rect 435640 274728 435692 274780
rect 439412 274728 439464 274780
rect 453948 274728 454000 274780
rect 457168 274728 457220 274780
rect 464160 274728 464212 274780
rect 471336 274728 471388 274780
rect 482928 274728 482980 274780
rect 538312 274728 538364 274780
rect 538496 274728 538548 274780
rect 545856 274728 545908 274780
rect 546040 274728 546092 274780
rect 558828 274728 558880 274780
rect 66996 274660 67048 274712
rect 71044 274660 71096 274712
rect 90640 274660 90692 274712
rect 95884 274660 95936 274712
rect 161572 274660 161624 274712
rect 163136 274660 163188 274712
rect 170128 274660 170180 274712
rect 173072 274660 173124 274712
rect 185216 274660 185268 274712
rect 187148 274660 187200 274712
rect 238484 274660 238536 274712
rect 239772 274660 239824 274712
rect 285772 274660 285824 274712
rect 286968 274660 287020 274712
rect 290464 274660 290516 274712
rect 294144 274660 294196 274712
rect 296352 274660 296404 274712
rect 298376 274660 298428 274712
rect 360292 274660 360344 274712
rect 363788 274660 363840 274712
rect 367100 274660 367152 274712
rect 369676 274660 369728 274712
rect 386052 274660 386104 274712
rect 389732 274660 389784 274712
rect 407120 274660 407172 274712
rect 411076 274660 411128 274712
rect 104808 274592 104860 274644
rect 157616 274592 157668 274644
rect 195888 274592 195940 274644
rect 206284 274592 206336 274644
rect 424968 274592 425020 274644
rect 474924 274592 474976 274644
rect 475384 274592 475436 274644
rect 490564 274592 490616 274644
rect 490748 274592 490800 274644
rect 496176 274592 496228 274644
rect 121368 274456 121420 274508
rect 176752 274456 176804 274508
rect 182916 274456 182968 274508
rect 199660 274456 199712 274508
rect 210056 274456 210108 274508
rect 237840 274456 237892 274508
rect 392584 274456 392636 274508
rect 402796 274456 402848 274508
rect 406844 274456 406896 274508
rect 437480 274456 437532 274508
rect 440884 274456 440936 274508
rect 488448 274456 488500 274508
rect 101312 274320 101364 274372
rect 160928 274320 160980 274372
rect 187792 274320 187844 274372
rect 220912 274320 220964 274372
rect 362868 274320 362920 274372
rect 386236 274320 386288 274372
rect 395896 274320 395948 274372
rect 420920 274320 420972 274372
rect 471244 274320 471296 274372
rect 491024 274456 491076 274508
rect 491208 274456 491260 274508
rect 570696 274592 570748 274644
rect 570880 274592 570932 274644
rect 587164 274592 587216 274644
rect 501972 274456 502024 274508
rect 490564 274320 490616 274372
rect 504732 274456 504784 274508
rect 577780 274456 577832 274508
rect 585784 274456 585836 274508
rect 82360 274184 82412 274236
rect 145564 274184 145616 274236
rect 160100 274184 160152 274236
rect 164240 274184 164292 274236
rect 176936 274184 176988 274236
rect 214656 274184 214708 274236
rect 220544 274184 220596 274236
rect 240600 274184 240652 274236
rect 342904 274184 342956 274236
rect 347228 274184 347280 274236
rect 366916 274184 366968 274236
rect 389180 274184 389232 274236
rect 390284 274184 390336 274236
rect 426440 274184 426492 274236
rect 438768 274184 438820 274236
rect 490748 274184 490800 274236
rect 490932 274184 490984 274236
rect 493784 274184 493836 274236
rect 496268 274184 496320 274236
rect 504180 274184 504232 274236
rect 586060 274320 586112 274372
rect 601424 274320 601476 274372
rect 84752 274048 84804 274100
rect 148324 274048 148376 274100
rect 158076 274048 158128 274100
rect 200672 274048 200724 274100
rect 206560 274048 206612 274100
rect 235448 274048 235500 274100
rect 239588 274048 239640 274100
rect 258632 274048 258684 274100
rect 360108 274048 360160 274100
rect 383844 274048 383896 274100
rect 384948 274048 385000 274100
rect 419356 274048 419408 274100
rect 421564 274048 421616 274100
rect 458364 274048 458416 274100
rect 459376 274048 459428 274100
rect 516600 274048 516652 274100
rect 518440 274184 518492 274236
rect 602528 274184 602580 274236
rect 613384 274184 613436 274236
rect 615592 274184 615644 274236
rect 527824 274048 527876 274100
rect 528008 274048 528060 274100
rect 619180 274048 619232 274100
rect 77208 273912 77260 273964
rect 143540 273912 143592 273964
rect 145012 273912 145064 273964
rect 192484 273912 192536 273964
rect 193496 273912 193548 273964
rect 226340 273912 226392 273964
rect 234896 273912 234948 273964
rect 255504 273912 255556 273964
rect 256148 273912 256200 273964
rect 270592 273912 270644 273964
rect 271512 273912 271564 273964
rect 280804 273912 280856 273964
rect 346308 273912 346360 273964
rect 362592 273912 362644 273964
rect 377772 273912 377824 273964
rect 408684 273912 408736 273964
rect 413928 273912 413980 273964
rect 449900 273912 449952 273964
rect 451096 273912 451148 273964
rect 513840 273912 513892 273964
rect 519728 273912 519780 273964
rect 524236 273912 524288 273964
rect 524420 273912 524472 273964
rect 613200 273912 613252 273964
rect 123760 273776 123812 273828
rect 177488 273776 177540 273828
rect 426900 273776 426952 273828
rect 477224 273776 477276 273828
rect 488448 273776 488500 273828
rect 490932 273776 490984 273828
rect 492036 273776 492088 273828
rect 571800 273776 571852 273828
rect 280988 273708 281040 273760
rect 287520 273708 287572 273760
rect 134432 273640 134484 273692
rect 185032 273640 185084 273692
rect 460020 273640 460072 273692
rect 484308 273640 484360 273692
rect 487988 273640 488040 273692
rect 565912 273640 565964 273692
rect 144644 273504 144696 273556
rect 187792 273504 187844 273556
rect 429016 273504 429068 273556
rect 482008 273504 482060 273556
rect 487068 273504 487120 273556
rect 563520 273504 563572 273556
rect 481364 273368 481416 273420
rect 556436 273368 556488 273420
rect 347044 273232 347096 273284
rect 349620 273232 349672 273284
rect 350264 273232 350316 273284
rect 356336 273232 356388 273284
rect 409144 273232 409196 273284
rect 409880 273232 409932 273284
rect 114284 273164 114336 273216
rect 169024 273164 169076 273216
rect 104992 273028 105044 273080
rect 163320 273028 163372 273080
rect 167552 273028 167604 273080
rect 184204 273028 184256 273080
rect 187608 273028 187660 273080
rect 211988 273164 212040 273216
rect 419172 273164 419224 273216
rect 456800 273164 456852 273216
rect 463148 273164 463200 273216
rect 486884 273164 486936 273216
rect 493692 273164 493744 273216
rect 574192 273164 574244 273216
rect 578884 273164 578936 273216
rect 594340 273164 594392 273216
rect 211252 273028 211304 273080
rect 220084 273028 220136 273080
rect 382924 273028 382976 273080
rect 392124 273028 392176 273080
rect 404176 273028 404228 273080
rect 429200 273028 429252 273080
rect 434628 273028 434680 273080
rect 488724 273028 488776 273080
rect 496636 273028 496688 273080
rect 578516 273028 578568 273080
rect 580264 273028 580316 273080
rect 640432 273028 640484 273080
rect 78864 272892 78916 272944
rect 138664 272892 138716 272944
rect 141792 272892 141844 272944
rect 189816 272892 189868 272944
rect 191196 272892 191248 272944
rect 224868 272892 224920 272944
rect 288072 272892 288124 272944
rect 290464 272892 290516 272944
rect 373264 272892 373316 272944
rect 382648 272892 382700 272944
rect 94228 272756 94280 272808
rect 156052 272756 156104 272808
rect 180524 272756 180576 272808
rect 217232 272756 217284 272808
rect 228824 272756 228876 272808
rect 249064 272756 249116 272808
rect 352932 272756 352984 272808
rect 372988 272756 373040 272808
rect 380716 272756 380768 272808
rect 388628 272892 388680 272944
rect 391848 272892 391900 272944
rect 410064 272892 410116 272944
rect 412456 272892 412508 272944
rect 453948 272892 454000 272944
rect 458088 272892 458140 272944
rect 521844 272892 521896 272944
rect 87144 272620 87196 272672
rect 152004 272620 152056 272672
rect 168656 272620 168708 272672
rect 208492 272620 208544 272672
rect 217416 272620 217468 272672
rect 242164 272620 242216 272672
rect 242348 272620 242400 272672
rect 259552 272620 259604 272672
rect 331036 272620 331088 272672
rect 342444 272620 342496 272672
rect 368388 272620 368440 272672
rect 394516 272756 394568 272808
rect 397276 272756 397328 272808
rect 418344 272756 418396 272808
rect 426072 272756 426124 272808
rect 478420 272756 478472 272808
rect 482744 272756 482796 272808
rect 524374 272892 524426 272944
rect 524512 272892 524564 272944
rect 611360 272892 611412 272944
rect 388628 272620 388680 272672
rect 393596 272620 393648 272672
rect 393964 272620 394016 272672
rect 406292 272620 406344 272672
rect 408408 272620 408460 272672
rect 452476 272620 452528 272672
rect 453856 272620 453908 272672
rect 516416 272620 516468 272672
rect 516600 272620 516652 272672
rect 606116 272756 606168 272808
rect 524328 272620 524380 272672
rect 524512 272620 524564 272672
rect 524880 272620 524932 272672
rect 614396 272620 614448 272672
rect 77668 272484 77720 272536
rect 145104 272484 145156 272536
rect 152188 272484 152240 272536
rect 197544 272484 197596 272536
rect 199476 272484 199528 272536
rect 230572 272484 230624 272536
rect 231400 272484 231452 272536
rect 252744 272484 252796 272536
rect 252928 272484 252980 272536
rect 267740 272484 267792 272536
rect 268016 272484 268068 272536
rect 278780 272484 278832 272536
rect 279792 272484 279844 272536
rect 287152 272484 287204 272536
rect 338028 272484 338080 272536
rect 351920 272484 351972 272536
rect 358636 272484 358688 272536
rect 380348 272484 380400 272536
rect 380532 272484 380584 272536
rect 413376 272484 413428 272536
rect 415124 272484 415176 272536
rect 461860 272484 461912 272536
rect 463516 272484 463568 272536
rect 524604 272484 524656 272536
rect 525064 272484 525116 272536
rect 533988 272484 534040 272536
rect 534172 272484 534224 272536
rect 632152 272484 632204 272536
rect 127348 272348 127400 272400
rect 179880 272348 179932 272400
rect 439320 272348 439372 272400
rect 473728 272348 473780 272400
rect 474648 272348 474700 272400
rect 495440 272348 495492 272400
rect 501604 272348 501656 272400
rect 581276 272348 581328 272400
rect 139124 272212 139176 272264
rect 141608 272212 141660 272264
rect 143908 272212 143960 272264
rect 190736 272212 190788 272264
rect 451740 272212 451792 272264
rect 480812 272212 480864 272264
rect 488356 272212 488408 272264
rect 567108 272212 567160 272264
rect 153292 272076 153344 272128
rect 171784 272076 171836 272128
rect 473084 272076 473136 272128
rect 482928 272076 482980 272128
rect 483756 272076 483808 272128
rect 560024 272076 560076 272128
rect 478696 271940 478748 271992
rect 552480 271940 552532 271992
rect 552848 271940 552900 271992
rect 580080 271940 580132 271992
rect 110420 271804 110472 271856
rect 164976 271804 165028 271856
rect 175832 271804 175884 271856
rect 207664 271804 207716 271856
rect 214840 271804 214892 271856
rect 221464 271804 221516 271856
rect 222108 271804 222160 271856
rect 232136 271804 232188 271856
rect 356520 271804 356572 271856
rect 359004 271804 359056 271856
rect 394332 271804 394384 271856
rect 426256 271804 426308 271856
rect 427084 271804 427136 271856
rect 433524 271804 433576 271856
rect 447784 271804 447836 271856
rect 503996 271804 504048 271856
rect 504732 271804 504784 271856
rect 589556 271804 589608 271856
rect 318616 271736 318668 271788
rect 324780 271736 324832 271788
rect 93032 271668 93084 271720
rect 120724 271668 120776 271720
rect 120908 271668 120960 271720
rect 175280 271668 175332 271720
rect 192300 271668 192352 271720
rect 225512 271668 225564 271720
rect 237472 271668 237524 271720
rect 243728 271668 243780 271720
rect 355324 271668 355376 271720
rect 374368 271668 374420 271720
rect 387708 271668 387760 271720
rect 421380 271668 421432 271720
rect 421748 271668 421800 271720
rect 438216 271668 438268 271720
rect 442908 271668 442960 271720
rect 500500 271668 500552 271720
rect 500868 271668 500920 271720
rect 508044 271668 508096 271720
rect 508964 271668 509016 271720
rect 596640 271804 596692 271856
rect 591488 271668 591540 271720
rect 603724 271668 603776 271720
rect 111984 271532 112036 271584
rect 168380 271532 168432 271584
rect 173440 271532 173492 271584
rect 212632 271532 212684 271584
rect 226156 271532 226208 271584
rect 247132 271532 247184 271584
rect 259736 271532 259788 271584
rect 272616 271532 272668 271584
rect 372528 271532 372580 271584
rect 400404 271532 400456 271584
rect 409788 271532 409840 271584
rect 443736 271532 443788 271584
rect 453304 271532 453356 271584
rect 511540 271532 511592 271584
rect 511908 271532 511960 271584
rect 600228 271532 600280 271584
rect 607864 271532 607916 271584
rect 643928 271532 643980 271584
rect 89720 271396 89772 271448
rect 152648 271396 152700 271448
rect 165160 271396 165212 271448
rect 205732 271396 205784 271448
rect 223580 271396 223632 271448
rect 247316 271396 247368 271448
rect 247868 271396 247920 271448
rect 264336 271396 264388 271448
rect 334624 271396 334676 271448
rect 341340 271396 341392 271448
rect 342168 271396 342220 271448
rect 356704 271396 356756 271448
rect 360844 271396 360896 271448
rect 381544 271396 381596 271448
rect 398104 271396 398156 271448
rect 427084 271396 427136 271448
rect 427268 271396 427320 271448
rect 68192 271260 68244 271312
rect 138480 271260 138532 271312
rect 150992 271260 151044 271312
rect 195980 271260 196032 271312
rect 215944 271260 215996 271312
rect 242072 271260 242124 271312
rect 243176 271260 243228 271312
rect 261024 271260 261076 271312
rect 275100 271260 275152 271312
rect 283472 271260 283524 271312
rect 315764 271260 315816 271312
rect 319996 271260 320048 271312
rect 325516 271260 325568 271312
rect 334164 271260 334216 271312
rect 340604 271260 340656 271312
rect 355508 271260 355560 271312
rect 364156 271260 364208 271312
rect 386052 271260 386104 271312
rect 400128 271260 400180 271312
rect 435640 271260 435692 271312
rect 436928 271396 436980 271448
rect 454776 271396 454828 271448
rect 457444 271396 457496 271448
rect 511724 271396 511776 271448
rect 448888 271260 448940 271312
rect 454684 271260 454736 271312
rect 515128 271396 515180 271448
rect 515312 271396 515364 271448
rect 518624 271396 518676 271448
rect 520096 271396 520148 271448
rect 523960 271396 524012 271448
rect 524144 271396 524196 271448
rect 514484 271260 514536 271312
rect 529020 271260 529072 271312
rect 529388 271396 529440 271448
rect 610808 271396 610860 271448
rect 617984 271260 618036 271312
rect 72976 271124 73028 271176
rect 142160 271124 142212 271176
rect 148600 271124 148652 271176
rect 194784 271124 194836 271176
rect 208860 271124 208912 271176
rect 237472 271124 237524 271176
rect 240784 271124 240836 271176
rect 259828 271124 259880 271176
rect 262128 271124 262180 271176
rect 274640 271124 274692 271176
rect 276296 271124 276348 271176
rect 284484 271124 284536 271176
rect 333888 271124 333940 271176
rect 344468 271124 344520 271176
rect 344652 271124 344704 271176
rect 350724 271124 350776 271176
rect 351828 271124 351880 271176
rect 372068 271124 372120 271176
rect 379428 271124 379480 271176
rect 407120 271124 407172 271176
rect 416596 271124 416648 271176
rect 463976 271124 464028 271176
rect 464528 271124 464580 271176
rect 524604 271124 524656 271176
rect 524788 271124 524840 271176
rect 529388 271124 529440 271176
rect 529572 271124 529624 271176
rect 532792 271124 532844 271176
rect 533160 271124 533212 271176
rect 621480 271124 621532 271176
rect 621664 271124 621716 271176
rect 636844 271124 636896 271176
rect 128544 270988 128596 271040
rect 181352 270988 181404 271040
rect 190000 270988 190052 271040
rect 216128 270988 216180 271040
rect 381544 270988 381596 271040
rect 399208 270988 399260 271040
rect 401324 270988 401376 271040
rect 130844 270852 130896 270904
rect 182456 270852 182508 270904
rect 200488 270852 200540 270904
rect 224224 270852 224276 270904
rect 389088 270852 389140 270904
rect 415308 270852 415360 270904
rect 425704 270988 425756 271040
rect 427268 270988 427320 271040
rect 431684 270988 431736 271040
rect 485504 270988 485556 271040
rect 488540 270988 488592 271040
rect 551744 270988 551796 271040
rect 552664 270988 552716 271040
rect 591488 270988 591540 271040
rect 427820 270852 427872 270904
rect 435364 270852 435416 270904
rect 436928 270852 436980 270904
rect 445024 270852 445076 270904
rect 497372 270852 497424 270904
rect 507676 270852 507728 270904
rect 523960 270852 524012 270904
rect 524880 270852 524932 270904
rect 593144 270852 593196 270904
rect 137928 270716 137980 270768
rect 187884 270716 187936 270768
rect 433156 270716 433208 270768
rect 456984 270716 457036 270768
rect 465724 270716 465776 270768
rect 526260 270716 526312 270768
rect 526444 270716 526496 270768
rect 528652 270716 528704 270768
rect 529020 270716 529072 270768
rect 116676 270580 116728 270632
rect 151084 270580 151136 270632
rect 237288 270580 237340 270632
rect 115848 270444 115900 270496
rect 171232 270444 171284 270496
rect 172428 270444 172480 270496
rect 208676 270444 208728 270496
rect 210792 270444 210844 270496
rect 211804 270444 211856 270496
rect 233148 270444 233200 270496
rect 237288 270444 237340 270496
rect 428464 270580 428516 270632
rect 466644 270580 466696 270632
rect 478144 270580 478196 270632
rect 538864 270580 538916 270632
rect 540520 270716 540572 270768
rect 543556 270716 543608 270768
rect 543694 270716 543746 270768
rect 607312 270716 607364 270768
rect 552664 270580 552716 270632
rect 252008 270444 252060 270496
rect 292856 270444 292908 270496
rect 296260 270444 296312 270496
rect 359004 270444 359056 270496
rect 376760 270444 376812 270496
rect 377588 270444 377640 270496
rect 394700 270444 394752 270496
rect 396264 270444 396316 270496
rect 423680 270444 423732 270496
rect 424600 270444 424652 270496
rect 476304 270444 476356 270496
rect 479248 270444 479300 270496
rect 552204 270444 552256 270496
rect 552388 270444 552440 270496
rect 564440 270444 564492 270496
rect 110236 270308 110288 270360
rect 167920 270308 167972 270360
rect 173072 270308 173124 270360
rect 210148 270308 210200 270360
rect 212448 270308 212500 270360
rect 239956 270308 240008 270360
rect 253848 270308 253900 270360
rect 265072 270308 265124 270360
rect 291660 270308 291712 270360
rect 295524 270308 295576 270360
rect 356704 270308 356756 270360
rect 378140 270308 378192 270360
rect 385684 270308 385736 270360
rect 419540 270308 419592 270360
rect 429568 270308 429620 270360
rect 483112 270308 483164 270360
rect 486700 270308 486752 270360
rect 494336 270308 494388 270360
rect 494520 270308 494572 270360
rect 560300 270308 560352 270360
rect 316960 270240 317012 270292
rect 321560 270240 321612 270292
rect 97908 270172 97960 270224
rect 158812 270172 158864 270224
rect 166908 270172 166960 270224
rect 207388 270172 207440 270224
rect 213828 270172 213880 270224
rect 240508 270172 240560 270224
rect 249616 270172 249668 270224
rect 263324 270172 263376 270224
rect 269212 270172 269264 270224
rect 279700 270172 279752 270224
rect 321928 270172 321980 270224
rect 328460 270172 328512 270224
rect 348424 270172 348476 270224
rect 363052 270172 363104 270224
rect 364984 270172 365036 270224
rect 390560 270172 390612 270224
rect 392308 270172 392360 270224
rect 429384 270172 429436 270224
rect 446956 270172 447008 270224
rect 504180 270172 504232 270224
rect 504364 270172 504416 270224
rect 528468 270172 528520 270224
rect 309784 270104 309836 270156
rect 311348 270104 311400 270156
rect 339316 270104 339368 270156
rect 341524 270104 341576 270156
rect 80060 270036 80112 270088
rect 146392 270036 146444 270088
rect 146760 270036 146812 270088
rect 151360 270036 151412 270088
rect 75828 269900 75880 269952
rect 142620 269900 142672 269952
rect 143356 269900 143408 269952
rect 153844 270036 153896 270088
rect 159916 270036 159968 270088
rect 202696 270036 202748 270088
rect 205548 270036 205600 270088
rect 234988 270036 235040 270088
rect 239772 270036 239824 270088
rect 253204 270036 253256 270088
rect 266176 270036 266228 270088
rect 277216 270036 277268 270088
rect 323584 270036 323636 270088
rect 331220 270036 331272 270088
rect 332324 270036 332376 270088
rect 336740 270036 336792 270088
rect 341800 270036 341852 270088
rect 357440 270036 357492 270088
rect 369400 270036 369452 270088
rect 396080 270036 396132 270088
rect 403072 270036 403124 270088
rect 444380 270036 444432 270088
rect 466000 270036 466052 270088
rect 533896 270172 533948 270224
rect 534034 270172 534086 270224
rect 626540 270172 626592 270224
rect 529020 270036 529072 270088
rect 538864 270036 538916 270088
rect 540980 270036 541032 270088
rect 541808 270036 541860 270088
rect 541992 270036 542044 270088
rect 633624 270036 633676 270088
rect 154488 269900 154540 269952
rect 198188 269900 198240 269952
rect 198648 269900 198700 269952
rect 230020 269900 230072 269952
rect 230388 269900 230440 269952
rect 252376 269900 252428 269952
rect 258448 269900 258500 269952
rect 272248 269900 272300 269952
rect 273076 269900 273128 269952
rect 282184 269900 282236 269952
rect 286784 269900 286836 269952
rect 292120 269900 292172 269952
rect 326896 269900 326948 269952
rect 335912 269900 335964 269952
rect 336832 269900 336884 269952
rect 350540 269900 350592 269952
rect 354220 269900 354272 269952
rect 375380 269900 375432 269952
rect 376576 269900 376628 269952
rect 403992 269900 404044 269952
rect 413008 269900 413060 269952
rect 459560 269900 459612 269952
rect 461860 269900 461912 269952
rect 529204 269900 529256 269952
rect 529756 269900 529808 269952
rect 530308 269900 530360 269952
rect 530584 269900 530636 269952
rect 532884 269900 532936 269952
rect 533068 269900 533120 269952
rect 630680 269900 630732 269952
rect 69388 269764 69440 269816
rect 139768 269764 139820 269816
rect 139952 269764 140004 269816
rect 181168 269764 181220 269816
rect 182088 269764 182140 269816
rect 186964 269764 187016 269816
rect 187332 269764 187384 269816
rect 191932 269764 191984 269816
rect 194600 269764 194652 269816
rect 227260 269764 227312 269816
rect 84108 269628 84160 269680
rect 119804 269628 119856 269680
rect 119068 269492 119120 269544
rect 173716 269628 173768 269680
rect 184756 269628 184808 269680
rect 213828 269628 213880 269680
rect 226616 269628 226668 269680
rect 249892 269764 249944 269816
rect 251456 269764 251508 269816
rect 267280 269764 267332 269816
rect 270316 269764 270368 269816
rect 280528 269764 280580 269816
rect 314476 269764 314528 269816
rect 318984 269764 319036 269816
rect 329656 269764 329708 269816
rect 339500 269764 339552 269816
rect 347596 269764 347648 269816
rect 365720 269764 365772 269816
rect 372344 269764 372396 269816
rect 401784 269764 401836 269816
rect 457720 269764 457772 269816
rect 470968 269764 471020 269816
rect 471612 269764 471664 269816
rect 537944 269764 537996 269816
rect 538864 269764 538916 269816
rect 552296 269764 552348 269816
rect 552480 269764 552532 269816
rect 641904 269764 641956 269816
rect 253204 269628 253256 269680
rect 258172 269628 258224 269680
rect 351644 269628 351696 269680
rect 364340 269628 364392 269680
rect 384028 269628 384080 269680
rect 388168 269628 388220 269680
rect 404360 269628 404412 269680
rect 426624 269628 426676 269680
rect 427360 269628 427412 269680
rect 478880 269628 478932 269680
rect 484216 269628 484268 269680
rect 494520 269628 494572 269680
rect 494888 269628 494940 269680
rect 504364 269628 504416 269680
rect 504548 269628 504600 269680
rect 553032 269628 553084 269680
rect 558920 269628 558972 269680
rect 572720 269628 572772 269680
rect 126888 269492 126940 269544
rect 178684 269492 178736 269544
rect 183468 269492 183520 269544
rect 187332 269492 187384 269544
rect 208308 269492 208360 269544
rect 230756 269492 230808 269544
rect 394700 269492 394752 269544
rect 416780 269492 416832 269544
rect 419632 269492 419684 269544
rect 468024 269492 468076 269544
rect 474280 269492 474332 269544
rect 335636 269424 335688 269476
rect 343824 269424 343876 269476
rect 118608 269356 118660 269408
rect 166908 269356 166960 269408
rect 401600 269356 401652 269408
rect 430580 269356 430632 269408
rect 449900 269356 449952 269408
rect 471980 269356 472032 269408
rect 476764 269356 476816 269408
rect 537944 269492 537996 269544
rect 540980 269492 541032 269544
rect 541348 269492 541400 269544
rect 552388 269492 552440 269544
rect 568580 269492 568632 269544
rect 136824 269220 136876 269272
rect 182180 269220 182232 269272
rect 264888 269220 264940 269272
rect 269120 269220 269172 269272
rect 321100 269220 321152 269272
rect 327908 269220 327960 269272
rect 417148 269220 417200 269272
rect 465080 269220 465132 269272
rect 468760 269220 468812 269272
rect 537024 269220 537076 269272
rect 546224 269356 546276 269408
rect 546408 269356 546460 269408
rect 551928 269356 551980 269408
rect 549444 269220 549496 269272
rect 549628 269220 549680 269272
rect 553032 269356 553084 269408
rect 557540 269356 557592 269408
rect 552296 269220 552348 269272
rect 607588 269220 607640 269272
rect 282736 269084 282788 269136
rect 288808 269084 288860 269136
rect 295340 269084 295392 269136
rect 297548 269084 297600 269136
rect 319444 269084 319496 269136
rect 325700 269084 325752 269136
rect 434444 269084 434496 269136
rect 490196 269084 490248 269136
rect 108948 269016 109000 269068
rect 166264 269016 166316 269068
rect 185584 269016 185636 269068
rect 196900 269016 196952 269068
rect 251088 269016 251140 269068
rect 256516 269016 256568 269068
rect 86868 268880 86920 268932
rect 144736 268880 144788 268932
rect 179328 268880 179380 268932
rect 215944 268880 215996 268932
rect 382372 268880 382424 268932
rect 400588 268880 400640 268932
rect 102508 268744 102560 268796
rect 162952 268744 163004 268796
rect 163136 268744 163188 268796
rect 203524 268744 203576 268796
rect 203892 268744 203944 268796
rect 227720 268744 227772 268796
rect 227904 268744 227956 268796
rect 250720 268744 250772 268796
rect 387340 268744 387392 268796
rect 422300 269016 422352 269068
rect 499120 269016 499172 269068
rect 582380 269016 582432 269068
rect 590660 269016 590712 269068
rect 418988 268880 419040 268932
rect 440240 268880 440292 268932
rect 443644 268880 443696 268932
rect 502524 268880 502576 268932
rect 503076 268880 503128 268932
rect 505100 268880 505152 268932
rect 508228 268880 508280 268932
rect 594800 268880 594852 268932
rect 422300 268744 422352 268796
rect 436100 268744 436152 268796
rect 441160 268744 441212 268796
rect 499580 268744 499632 268796
rect 504088 268744 504140 268796
rect 509332 268744 509384 268796
rect 510712 268744 510764 268796
rect 514300 268744 514352 268796
rect 581644 268744 581696 268796
rect 581828 268744 581880 268796
rect 598848 268744 598900 268796
rect 99288 268608 99340 268660
rect 160468 268608 160520 268660
rect 162768 268608 162820 268660
rect 205180 268608 205232 268660
rect 219532 268608 219584 268660
rect 244924 268608 244976 268660
rect 363052 268608 363104 268660
rect 386420 268608 386472 268660
rect 402244 268608 402296 268660
rect 443276 268608 443328 268660
rect 446128 268608 446180 268660
rect 503076 268608 503128 268660
rect 503260 268608 503312 268660
rect 513748 268608 513800 268660
rect 590660 268608 590712 268660
rect 608692 268608 608744 268660
rect 92388 268472 92440 268524
rect 155500 268472 155552 268524
rect 155868 268472 155920 268524
rect 200212 268472 200264 268524
rect 202972 268472 203024 268524
rect 233332 268472 233384 268524
rect 245568 268472 245620 268524
rect 263140 268472 263192 268524
rect 263508 268472 263560 268524
rect 275560 268472 275612 268524
rect 333520 268472 333572 268524
rect 345112 268472 345164 268524
rect 345940 268472 345992 268524
rect 360292 268472 360344 268524
rect 361028 268472 361080 268524
rect 369860 268472 369912 268524
rect 370320 268472 370372 268524
rect 397460 268472 397512 268524
rect 400588 268472 400640 268524
rect 441620 268472 441672 268524
rect 442724 268472 442776 268524
rect 446772 268472 446824 268524
rect 448612 268472 448664 268524
rect 504088 268472 504140 268524
rect 504272 268472 504324 268524
rect 66260 268336 66312 268388
rect 137284 268336 137336 268388
rect 147588 268336 147640 268388
rect 193588 268336 193640 268388
rect 197268 268336 197320 268388
rect 229192 268336 229244 268388
rect 233700 268336 233752 268388
rect 254860 268336 254912 268388
rect 255320 268336 255372 268388
rect 269764 268336 269816 268388
rect 322756 268336 322808 268388
rect 329840 268336 329892 268388
rect 335176 268336 335228 268388
rect 347780 268336 347832 268388
rect 350080 268336 350132 268388
rect 367100 268336 367152 268388
rect 374920 268336 374972 268388
rect 404544 268336 404596 268388
rect 407212 268336 407264 268388
rect 451464 268336 451516 268388
rect 461032 268336 461084 268388
rect 518808 268336 518860 268388
rect 519360 268472 519412 268524
rect 533896 268472 533948 268524
rect 534034 268472 534086 268524
rect 619640 268472 619692 268524
rect 520280 268336 520332 268388
rect 520464 268336 520516 268388
rect 526996 268336 527048 268388
rect 527180 268336 527232 268388
rect 547512 268336 547564 268388
rect 547696 268336 547748 268388
rect 638960 268336 639012 268388
rect 122748 268200 122800 268252
rect 176200 268200 176252 268252
rect 436192 268200 436244 268252
rect 488908 268200 488960 268252
rect 133788 268064 133840 268116
rect 183652 268064 183704 268116
rect 420460 268064 420512 268116
rect 469036 268064 469088 268116
rect 469220 268064 469272 268116
rect 504272 268200 504324 268252
rect 505744 268200 505796 268252
rect 591028 268200 591080 268252
rect 492772 268064 492824 268116
rect 498200 268064 498252 268116
rect 500684 268064 500736 268116
rect 580448 268064 580500 268116
rect 581644 268064 581696 268116
rect 587900 268064 587952 268116
rect 125508 267928 125560 267980
rect 147588 267928 147640 267980
rect 437848 267928 437900 267980
rect 468208 267928 468260 267980
rect 431960 267792 432012 267844
rect 447140 267792 447192 267844
rect 533896 267928 533948 267980
rect 534034 267928 534086 267980
rect 581828 267928 581880 267980
rect 88984 267656 89036 267708
rect 144552 267656 144604 267708
rect 144920 267656 144972 267708
rect 150532 267656 150584 267708
rect 171784 267656 171836 267708
rect 199384 267656 199436 267708
rect 207664 267656 207716 267708
rect 213460 267656 213512 267708
rect 368204 267656 368256 267708
rect 377588 267656 377640 267708
rect 383200 267656 383252 267708
rect 394700 267656 394752 267708
rect 398472 267656 398524 267708
rect 421748 267656 421800 267708
rect 435640 267656 435692 267708
rect 465540 267656 465592 267708
rect 466828 267656 466880 267708
rect 477592 267656 477644 267708
rect 488540 267792 488592 267844
rect 489184 267792 489236 267844
rect 567292 267792 567344 267844
rect 580448 267792 580500 267844
rect 584036 267792 584088 267844
rect 95884 267520 95936 267572
rect 154672 267520 154724 267572
rect 162124 267520 162176 267572
rect 169576 267520 169628 267572
rect 187148 267520 187200 267572
rect 221740 267520 221792 267572
rect 227720 267520 227772 267572
rect 234160 267520 234212 267572
rect 370780 267520 370832 267572
rect 381544 267520 381596 267572
rect 390652 267520 390704 267572
rect 404360 267520 404412 267572
rect 409604 267520 409656 267572
rect 435364 267520 435416 267572
rect 445300 267520 445352 267572
rect 492772 267656 492824 267708
rect 492956 267656 493008 267708
rect 558920 267656 558972 267708
rect 485228 267520 485280 267572
rect 502340 267520 502392 267572
rect 502800 267520 502852 267572
rect 506204 267520 506256 267572
rect 506480 267520 506532 267572
rect 507216 267520 507268 267572
rect 507400 267520 507452 267572
rect 578884 267520 578936 267572
rect 107568 267384 107620 267436
rect 167092 267384 167144 267436
rect 167736 267384 167788 267436
rect 204352 267384 204404 267436
rect 211988 267384 212040 267436
rect 222568 267384 222620 267436
rect 224224 267384 224276 267436
rect 231676 267384 231728 267436
rect 233884 267384 233936 267436
rect 246580 267384 246632 267436
rect 313648 267384 313700 267436
rect 317788 267384 317840 267436
rect 334348 267384 334400 267436
rect 342904 267384 342956 267436
rect 350908 267384 350960 267436
rect 361028 267384 361080 267436
rect 365812 267384 365864 267436
rect 382924 267384 382976 267436
rect 397092 267384 397144 267436
rect 422300 267384 422352 267436
rect 440332 267384 440384 267436
rect 494704 267384 494756 267436
rect 497464 267384 497516 267436
rect 552848 267384 552900 267436
rect 553032 267384 553084 267436
rect 570880 267384 570932 267436
rect 100668 267248 100720 267300
rect 162124 267248 162176 267300
rect 166908 267248 166960 267300
rect 174544 267248 174596 267300
rect 175096 267248 175148 267300
rect 214288 267248 214340 267300
rect 220084 267248 220136 267300
rect 239128 267248 239180 267300
rect 254584 267248 254636 267300
rect 262312 267248 262364 267300
rect 312820 267248 312872 267300
rect 316040 267248 316092 267300
rect 343456 267248 343508 267300
rect 353944 267248 353996 267300
rect 359188 267248 359240 267300
rect 373264 267248 373316 267300
rect 375748 267248 375800 267300
rect 393964 267248 394016 267300
rect 399760 267248 399812 267300
rect 418988 267248 419040 267300
rect 421288 267248 421340 267300
rect 464160 267248 464212 267300
rect 465540 267248 465592 267300
rect 471244 267248 471296 267300
rect 471796 267248 471848 267300
rect 475384 267248 475436 267300
rect 475936 267248 475988 267300
rect 518900 267248 518952 267300
rect 519176 267248 519228 267300
rect 521660 267248 521712 267300
rect 522948 267248 523000 267300
rect 73804 267112 73856 267164
rect 141424 267112 141476 267164
rect 144552 267112 144604 267164
rect 147404 267112 147456 267164
rect 147588 267112 147640 267164
rect 149060 267112 149112 267164
rect 149888 267112 149940 267164
rect 194416 267112 194468 267164
rect 199660 267112 199712 267164
rect 218428 267112 218480 267164
rect 221464 267112 221516 267164
rect 241612 267112 241664 267164
rect 246856 267112 246908 267164
rect 263968 267112 264020 267164
rect 342628 267112 342680 267164
rect 356520 267112 356572 267164
rect 363328 267112 363380 267164
rect 370504 267112 370556 267164
rect 373264 267112 373316 267164
rect 392584 267112 392636 267164
rect 404728 267112 404780 267164
rect 431960 267112 432012 267164
rect 71044 266976 71096 267028
rect 138112 266976 138164 267028
rect 141608 266976 141660 267028
rect 184020 266976 184072 267028
rect 184204 266976 184256 267028
rect 132408 266840 132460 266892
rect 184480 266840 184532 266892
rect 193864 266976 193916 267028
rect 201868 266976 201920 267028
rect 206284 266976 206336 267028
rect 228364 266976 228416 267028
rect 237288 266976 237340 267028
rect 254032 266976 254084 267028
rect 271420 266976 271472 267028
rect 276664 266976 276716 267028
rect 278044 266976 278096 267028
rect 286968 266976 287020 267028
rect 291292 266976 291344 267028
rect 295156 266976 295208 267028
rect 297088 266976 297140 267028
rect 324412 266976 324464 267028
rect 332508 266976 332560 267028
rect 353392 266976 353444 267028
rect 355324 266976 355376 267028
rect 355876 266976 355928 267028
rect 369124 266976 369176 267028
rect 378232 266976 378284 267028
rect 409144 266976 409196 267028
rect 422116 266976 422168 267028
rect 449900 267112 449952 267164
rect 450268 267112 450320 267164
rect 499764 267112 499816 267164
rect 499948 267112 500000 267164
rect 500868 267112 500920 267164
rect 501052 267112 501104 267164
rect 506388 267112 506440 267164
rect 506572 267112 506624 267164
rect 507676 267112 507728 267164
rect 507860 267112 507912 267164
rect 523592 267112 523644 267164
rect 523960 267248 524012 267300
rect 543556 267248 543608 267300
rect 543694 267248 543746 267300
rect 621664 267248 621716 267300
rect 585784 267112 585836 267164
rect 446404 266976 446456 267028
rect 451740 266976 451792 267028
rect 451924 266976 451976 267028
rect 460020 266976 460072 267028
rect 465172 266976 465224 267028
rect 519176 266976 519228 267028
rect 519360 266976 519412 267028
rect 520096 266976 520148 267028
rect 520280 266976 520332 267028
rect 522948 266976 523000 267028
rect 523132 266976 523184 267028
rect 524328 266976 524380 267028
rect 524788 266976 524840 267028
rect 525708 266976 525760 267028
rect 525892 266976 525944 267028
rect 533896 266976 533948 267028
rect 534034 266976 534086 267028
rect 622400 266976 622452 267028
rect 209320 266840 209372 266892
rect 216128 266840 216180 266892
rect 223396 266840 223448 266892
rect 249064 266840 249116 266892
rect 251548 266840 251600 266892
rect 257988 266840 258040 266892
rect 316132 266840 316184 266892
rect 320180 266840 320232 266892
rect 331864 266840 331916 266892
rect 335636 266840 335688 266892
rect 336004 266840 336056 266892
rect 347044 266840 347096 266892
rect 393136 266840 393188 266892
rect 401600 266840 401652 266892
rect 405556 266840 405608 266892
rect 425704 266840 425756 266892
rect 265072 266772 265124 266824
rect 268936 266772 268988 266824
rect 120724 266704 120776 266756
rect 156420 266704 156472 266756
rect 156604 266704 156656 266756
rect 159640 266704 159692 266756
rect 169024 266704 169076 266756
rect 172060 266704 172112 266756
rect 184020 266704 184072 266756
rect 189448 266704 189500 266756
rect 245108 266704 245160 266756
rect 249064 266704 249116 266756
rect 320272 266704 320324 266756
rect 327448 266704 327500 266756
rect 358360 266704 358412 266756
rect 360844 266704 360896 266756
rect 388168 266704 388220 266756
rect 396264 266704 396316 266756
rect 412180 266704 412232 266756
rect 330208 266636 330260 266688
rect 334624 266636 334676 266688
rect 138664 266568 138716 266620
rect 119804 266432 119856 266484
rect 144920 266432 144972 266484
rect 149060 266568 149112 266620
rect 179512 266568 179564 266620
rect 208676 266568 208728 266620
rect 210976 266568 211028 266620
rect 213828 266568 213880 266620
rect 220084 266568 220136 266620
rect 360844 266568 360896 266620
rect 362224 266568 362276 266620
rect 417976 266704 418028 266756
rect 428464 266704 428516 266756
rect 430396 266704 430448 266756
rect 451234 266840 451286 266892
rect 456432 266840 456484 266892
rect 469220 266840 469272 266892
rect 470140 266840 470192 266892
rect 432052 266704 432104 266756
rect 446404 266704 446456 266756
rect 449440 266704 449492 266756
rect 453304 266772 453356 266824
rect 455236 266772 455288 266824
rect 512920 266704 512972 266756
rect 513380 266704 513432 266756
rect 515496 266704 515548 266756
rect 516508 266704 516560 266756
rect 518716 266704 518768 266756
rect 519176 266840 519228 266892
rect 533988 266840 534040 266892
rect 534172 266840 534224 266892
rect 537208 266840 537260 266892
rect 537392 266840 537444 266892
rect 539508 266840 539560 266892
rect 539692 266840 539744 266892
rect 580264 266840 580316 266892
rect 524374 266704 524426 266756
rect 524512 266704 524564 266756
rect 613384 266704 613436 266756
rect 452752 266636 452804 266688
rect 455788 266636 455840 266688
rect 421564 266568 421616 266620
rect 422944 266568 422996 266620
rect 439320 266568 439372 266620
rect 439504 266568 439556 266620
rect 145564 266500 145616 266552
rect 148876 266500 148928 266552
rect 240692 266500 240744 266552
rect 245752 266500 245804 266552
rect 308680 266500 308732 266552
rect 310888 266500 310940 266552
rect 311164 266500 311216 266552
rect 313280 266500 313332 266552
rect 327724 266500 327776 266552
rect 332324 266500 332376 266552
rect 346768 266500 346820 266552
rect 351644 266500 351696 266552
rect 355048 266500 355100 266552
rect 359004 266500 359056 266552
rect 394792 266500 394844 266552
rect 398104 266500 398156 266552
rect 151084 266432 151136 266484
rect 172888 266432 172940 266484
rect 361672 266432 361724 266484
rect 362776 266432 362828 266484
rect 427912 266432 427964 266484
rect 147220 266364 147272 266416
rect 148324 266364 148376 266416
rect 149704 266364 149756 266416
rect 182180 266364 182232 266416
rect 186136 266364 186188 266416
rect 202144 266364 202196 266416
rect 206836 266364 206888 266416
rect 222844 266364 222896 266416
rect 224224 266364 224276 266416
rect 230756 266364 230808 266416
rect 236644 266364 236696 266416
rect 242256 266364 242308 266416
rect 243268 266364 243320 266416
rect 252008 266364 252060 266416
rect 257344 266364 257396 266416
rect 263324 266364 263376 266416
rect 265624 266364 265676 266416
rect 269120 266364 269172 266416
rect 276388 266364 276440 266416
rect 278596 266364 278648 266416
rect 286324 266364 286376 266416
rect 290464 266364 290516 266416
rect 292948 266364 293000 266416
rect 297916 266364 297968 266416
rect 299572 266364 299624 266416
rect 301044 266364 301096 266416
rect 302056 266364 302108 266416
rect 307852 266364 307904 266416
rect 309508 266364 309560 266416
rect 310336 266364 310388 266416
rect 311900 266364 311952 266416
rect 312360 266364 312412 266416
rect 314660 266364 314712 266416
rect 317788 266364 317840 266416
rect 323124 266364 323176 266416
rect 328552 266364 328604 266416
rect 329472 266364 329524 266416
rect 332692 266364 332744 266416
rect 333888 266364 333940 266416
rect 340972 266364 341024 266416
rect 342168 266364 342220 266416
rect 345112 266364 345164 266416
rect 346308 266364 346360 266416
rect 349252 266364 349304 266416
rect 350264 266364 350316 266416
rect 357532 266364 357584 266416
rect 358636 266364 358688 266416
rect 367468 266364 367520 266416
rect 368388 266364 368440 266416
rect 371608 266364 371660 266416
rect 372528 266364 372580 266416
rect 374092 266364 374144 266416
rect 375104 266364 375156 266416
rect 379888 266364 379940 266416
rect 380716 266364 380768 266416
rect 386512 266364 386564 266416
rect 387708 266364 387760 266416
rect 396448 266364 396500 266416
rect 397276 266364 397328 266416
rect 398932 266364 398984 266416
rect 400128 266364 400180 266416
rect 408868 266364 408920 266416
rect 409788 266364 409840 266416
rect 411352 266364 411404 266416
rect 412456 266364 412508 266416
rect 415492 266364 415544 266416
rect 416412 266364 416464 266416
rect 423772 266364 423824 266416
rect 424968 266364 425020 266416
rect 425428 266364 425480 266416
rect 426900 266364 426952 266416
rect 432052 266364 432104 266416
rect 432328 266364 432380 266416
rect 433156 266364 433208 266416
rect 433708 266364 433760 266416
rect 434628 266364 434680 266416
rect 437020 266364 437072 266416
rect 440884 266364 440936 266416
rect 441988 266364 442040 266416
rect 442908 266364 442960 266416
rect 459192 266568 459244 266620
rect 464160 266568 464212 266620
rect 464344 266568 464396 266620
rect 465724 266568 465776 266620
rect 469312 266568 469364 266620
rect 473268 266568 473320 266620
rect 473452 266568 473504 266620
rect 474648 266568 474700 266620
rect 474832 266568 474884 266620
rect 478144 266568 478196 266620
rect 481732 266568 481784 266620
rect 485228 266568 485280 266620
rect 485872 266568 485924 266620
rect 487068 266568 487120 266620
rect 490012 266568 490064 266620
rect 444472 266500 444524 266552
rect 447784 266500 447836 266552
rect 454408 266500 454460 266552
rect 457444 266500 457496 266552
rect 543694 266568 543746 266620
rect 553032 266568 553084 266620
rect 460204 266432 460256 266484
rect 445024 266364 445076 266416
rect 447784 266364 447836 266416
rect 449164 266364 449216 266416
rect 451924 266364 451976 266416
rect 454684 266364 454736 266416
rect 456892 266364 456944 266416
rect 458088 266364 458140 266416
rect 458548 266364 458600 266416
rect 459376 266364 459428 266416
rect 498568 266296 498620 266348
rect 501604 266296 501656 266348
rect 517336 266432 517388 266484
rect 512368 266364 512420 266416
rect 513380 266228 513432 266280
rect 514852 266364 514904 266416
rect 516784 266364 516836 266416
rect 549628 266432 549680 266484
rect 520280 266296 520332 266348
rect 522672 266296 522724 266348
rect 524512 266296 524564 266348
rect 546408 266296 546460 266348
rect 475108 266024 475160 266076
rect 547880 266024 547932 266076
rect 485044 265888 485096 265940
rect 561680 265888 561732 265940
rect 494980 265752 495032 265804
rect 575572 265752 575624 265804
rect 187700 265616 187752 265668
rect 188252 265616 188304 265668
rect 247132 265616 247184 265668
rect 247868 265616 247920 265668
rect 259552 265616 259604 265668
rect 260380 265616 260432 265668
rect 284300 265616 284352 265668
rect 285220 265616 285272 265668
rect 480076 265616 480128 265668
rect 554780 265616 554832 265668
rect 558184 265616 558236 265668
rect 647240 265616 647292 265668
rect 570604 261468 570656 261520
rect 645860 261468 645912 261520
rect 554412 260856 554464 260908
rect 568580 260856 568632 260908
rect 554320 259428 554372 259480
rect 567844 259428 567896 259480
rect 35808 256708 35860 256760
rect 40684 256708 40736 256760
rect 553952 256708 554004 256760
rect 562324 256708 562376 256760
rect 554504 253376 554556 253428
rect 559564 253376 559616 253428
rect 35624 252832 35676 252884
rect 41696 252832 41748 252884
rect 35808 252696 35860 252748
rect 40684 252696 40736 252748
rect 35440 252560 35492 252612
rect 41696 252560 41748 252612
rect 675852 252220 675904 252272
rect 678244 252220 678296 252272
rect 675852 251540 675904 251592
rect 678428 251540 678480 251592
rect 35808 251200 35860 251252
rect 36544 251200 36596 251252
rect 553492 251200 553544 251252
rect 555424 251200 555476 251252
rect 553676 249024 553728 249076
rect 571340 249024 571392 249076
rect 553860 246304 553912 246356
rect 632704 246304 632756 246356
rect 554412 245624 554464 245676
rect 591304 245624 591356 245676
rect 554504 244264 554556 244316
rect 624424 244264 624476 244316
rect 36544 242836 36596 242888
rect 41696 242836 41748 242888
rect 576124 242156 576176 242208
rect 648620 242156 648672 242208
rect 553952 241476 554004 241528
rect 628564 241476 628616 241528
rect 553860 240116 553912 240168
rect 577504 240116 577556 240168
rect 554320 238688 554372 238740
rect 576124 238688 576176 238740
rect 672172 238008 672224 238060
rect 671252 237600 671304 237652
rect 668768 237396 668820 237448
rect 671436 237124 671488 237176
rect 673304 237056 673356 237108
rect 671620 236920 671672 236972
rect 673414 236852 673466 236904
rect 673528 236648 673580 236700
rect 673414 236444 673466 236496
rect 673752 236240 673804 236292
rect 672632 236104 672684 236156
rect 554504 236036 554556 236088
rect 558184 236036 558236 236088
rect 671068 235832 671120 235884
rect 673000 235696 673052 235748
rect 669780 235492 669832 235544
rect 668124 235288 668176 235340
rect 591304 235220 591356 235272
rect 633624 235220 633676 235272
rect 674426 234744 674478 234796
rect 672540 234608 672592 234660
rect 554412 234540 554464 234592
rect 570604 234540 570656 234592
rect 675852 234540 675904 234592
rect 679624 234540 679676 234592
rect 669596 234200 669648 234252
rect 674564 234200 674616 234252
rect 675852 234336 675904 234388
rect 679992 234336 680044 234388
rect 674886 234268 674938 234320
rect 675852 234200 675904 234252
rect 679808 234200 679860 234252
rect 674978 234064 675030 234116
rect 670792 233996 670844 234048
rect 671804 233996 671856 234048
rect 675096 233860 675148 233912
rect 669136 233588 669188 233640
rect 675852 233656 675904 233708
rect 677784 233656 677836 233708
rect 671804 233316 671856 233368
rect 676036 233384 676088 233436
rect 683488 233384 683540 233436
rect 671160 232976 671212 233028
rect 674748 232976 674800 233028
rect 670884 232772 670936 232824
rect 675024 232772 675076 232824
rect 652024 232500 652076 232552
rect 675484 232500 675536 232552
rect 675852 232500 675904 232552
rect 680176 232500 680228 232552
rect 662328 232364 662380 232416
rect 675346 232296 675398 232348
rect 665088 232160 665140 232212
rect 673920 232024 673972 232076
rect 674564 232024 674616 232076
rect 675346 232024 675398 232076
rect 675180 231752 675232 231804
rect 675070 231548 675122 231600
rect 674956 231276 675008 231328
rect 675852 231208 675904 231260
rect 677600 231208 677652 231260
rect 674840 231140 674892 231192
rect 673552 231004 673604 231056
rect 674564 231004 674616 231056
rect 674732 230868 674784 230920
rect 673460 230800 673512 230852
rect 144644 230528 144696 230580
rect 150532 230528 150584 230580
rect 150900 230528 150952 230580
rect 158260 230664 158312 230716
rect 90364 230392 90416 230444
rect 165436 230528 165488 230580
rect 172060 230528 172112 230580
rect 176108 230528 176160 230580
rect 181076 230528 181128 230580
rect 439320 230528 439372 230580
rect 161112 230392 161164 230444
rect 161296 230392 161348 230444
rect 215208 230392 215260 230444
rect 223396 230392 223448 230444
rect 271880 230392 271932 230444
rect 274180 230392 274232 230444
rect 307944 230392 307996 230444
rect 312544 230392 312596 230444
rect 315672 230392 315724 230444
rect 377404 230392 377456 230444
rect 378784 230392 378836 230444
rect 674012 230528 674064 230580
rect 440700 230392 440752 230444
rect 441896 230392 441948 230444
rect 443460 230392 443512 230444
rect 468300 230392 468352 230444
rect 469036 230392 469088 230444
rect 534632 230392 534684 230444
rect 544200 230392 544252 230444
rect 669320 230392 669372 230444
rect 673920 230392 673972 230444
rect 674518 230460 674570 230512
rect 404268 230324 404320 230376
rect 412272 230324 412324 230376
rect 436100 230324 436152 230376
rect 436744 230324 436796 230376
rect 438676 230324 438728 230376
rect 439320 230324 439372 230376
rect 443828 230324 443880 230376
rect 444840 230324 444892 230376
rect 446404 230324 446456 230376
rect 449164 230324 449216 230376
rect 449624 230324 449676 230376
rect 450544 230324 450596 230376
rect 452844 230324 452896 230376
rect 454316 230324 454368 230376
rect 455420 230324 455472 230376
rect 457168 230324 457220 230376
rect 463792 230324 463844 230376
rect 465724 230324 465776 230376
rect 475384 230324 475436 230376
rect 478328 230324 478380 230376
rect 480536 230324 480588 230376
rect 481548 230324 481600 230376
rect 492772 230324 492824 230376
rect 493968 230324 494020 230376
rect 494704 230324 494756 230376
rect 496360 230324 496412 230376
rect 499856 230324 499908 230376
rect 501144 230324 501196 230376
rect 503720 230324 503772 230376
rect 506940 230324 506992 230376
rect 516600 230324 516652 230376
rect 517428 230324 517480 230376
rect 520464 230324 520516 230376
rect 521568 230324 521620 230376
rect 526904 230324 526956 230376
rect 527824 230324 527876 230376
rect 118424 230256 118476 230308
rect 189448 230256 189500 230308
rect 190920 230256 190972 230308
rect 202328 230256 202380 230308
rect 203708 230256 203760 230308
rect 256424 230256 256476 230308
rect 261392 230256 261444 230308
rect 297640 230256 297692 230308
rect 302884 230256 302936 230308
rect 305368 230256 305420 230308
rect 307852 230256 307904 230308
rect 323400 230256 323452 230308
rect 497924 230256 497976 230308
rect 499672 230256 499724 230308
rect 408868 230188 408920 230240
rect 410984 230188 411036 230240
rect 447048 230188 447100 230240
rect 449900 230188 449952 230240
rect 451556 230188 451608 230240
rect 453304 230188 453356 230240
rect 454132 230188 454184 230240
rect 455236 230188 455288 230240
rect 470876 230188 470928 230240
rect 471888 230188 471940 230240
rect 493416 230188 493468 230240
rect 495164 230188 495216 230240
rect 513380 230188 513432 230240
rect 515404 230188 515456 230240
rect 517244 230188 517296 230240
rect 529204 230256 529256 230308
rect 541624 230256 541676 230308
rect 667940 230256 667992 230308
rect 673828 230256 673880 230308
rect 522304 230188 522356 230240
rect 111064 230120 111116 230172
rect 184296 230120 184348 230172
rect 88248 229984 88300 230036
rect 166264 229984 166316 230036
rect 166448 229984 166500 230036
rect 181720 229984 181772 230036
rect 184204 229984 184256 230036
rect 191564 230120 191616 230172
rect 196992 230120 197044 230172
rect 251272 230120 251324 230172
rect 276848 230120 276900 230172
rect 313096 230120 313148 230172
rect 315304 230120 315356 230172
rect 340144 230120 340196 230172
rect 476672 230120 476724 230172
rect 479708 230120 479760 230172
rect 345664 230052 345716 230104
rect 353024 230052 353076 230104
rect 444472 230052 444524 230104
rect 447600 230052 447652 230104
rect 490840 230052 490892 230104
rect 493784 230052 493836 230104
rect 494336 230052 494388 230104
rect 503260 230120 503312 230172
rect 515680 230052 515732 230104
rect 189724 229984 189776 230036
rect 246120 229984 246172 230036
rect 251732 229984 251784 230036
rect 292488 229984 292540 230036
rect 296904 229984 296956 230036
rect 302516 229984 302568 230036
rect 305644 229984 305696 230036
rect 334992 229984 335044 230036
rect 380440 229984 380492 230036
rect 389088 229984 389140 230036
rect 468852 229984 468904 230036
rect 475384 229984 475436 230036
rect 476028 229984 476080 230036
rect 479524 229984 479576 230036
rect 483112 229984 483164 230036
rect 484308 229984 484360 230036
rect 484768 229984 484820 230036
rect 490656 229984 490708 230036
rect 499672 229984 499724 230036
rect 504364 229984 504416 230036
rect 511448 229916 511500 229968
rect 516784 229916 516836 229968
rect 74448 229848 74500 229900
rect 155960 229848 156012 229900
rect 156328 229848 156380 229900
rect 176568 229848 176620 229900
rect 177580 229848 177632 229900
rect 67548 229712 67600 229764
rect 144644 229712 144696 229764
rect 144828 229712 144880 229764
rect 140044 229576 140096 229628
rect 146944 229576 146996 229628
rect 148600 229712 148652 229764
rect 150900 229712 150952 229764
rect 151360 229712 151412 229764
rect 190920 229712 190972 229764
rect 191564 229848 191616 229900
rect 240968 229848 241020 229900
rect 245660 229848 245712 229900
rect 287336 229848 287388 229900
rect 300124 229848 300176 229900
rect 329840 229848 329892 229900
rect 334256 229848 334308 229900
rect 345296 229848 345348 229900
rect 352564 229848 352616 229900
rect 358176 229848 358228 229900
rect 364156 229848 364208 229900
rect 381360 229848 381412 229900
rect 384304 229848 384356 229900
rect 394240 229848 394292 229900
rect 412456 229848 412508 229900
rect 419356 229848 419408 229900
rect 467012 229848 467064 229900
rect 474004 229848 474056 229900
rect 481824 229848 481876 229900
rect 489920 229848 489972 229900
rect 495992 229848 496044 229900
rect 509240 229848 509292 229900
rect 519176 230052 519228 230104
rect 529020 230188 529072 230240
rect 674058 230188 674110 230240
rect 530768 230120 530820 230172
rect 523040 229984 523092 230036
rect 534724 229984 534776 230036
rect 536564 230120 536616 230172
rect 549260 230120 549312 230172
rect 673644 230052 673696 230104
rect 547144 229984 547196 230036
rect 555424 229984 555476 230036
rect 569960 229984 570012 230036
rect 673948 229916 674000 229968
rect 525524 229848 525576 229900
rect 538496 229848 538548 229900
rect 556804 229848 556856 229900
rect 433524 229780 433576 229832
rect 434168 229780 434220 229832
rect 675852 229848 675904 229900
rect 676956 229848 677008 229900
rect 235816 229712 235868 229764
rect 236920 229712 236972 229764
rect 282184 229712 282236 229764
rect 285312 229712 285364 229764
rect 318248 229712 318300 229764
rect 324044 229712 324096 229764
rect 350448 229712 350500 229764
rect 210056 229576 210108 229628
rect 210240 229576 210292 229628
rect 261576 229576 261628 229628
rect 350540 229576 350592 229628
rect 371056 229712 371108 229764
rect 370964 229576 371016 229628
rect 386512 229712 386564 229764
rect 386972 229712 387024 229764
rect 396816 229712 396868 229764
rect 399852 229712 399904 229764
rect 409696 229712 409748 229764
rect 411168 229712 411220 229764
rect 417424 229712 417476 229764
rect 457352 229712 457404 229764
rect 463884 229712 463936 229764
rect 465448 229712 465500 229764
rect 467472 229712 467524 229764
rect 469588 229712 469640 229764
rect 476764 229712 476816 229764
rect 479248 229712 479300 229764
rect 484124 229712 484176 229764
rect 486332 229712 486384 229764
rect 500224 229712 500276 229764
rect 505652 229712 505704 229764
rect 516048 229712 516100 229764
rect 518900 229712 518952 229764
rect 521108 229712 521160 229764
rect 529940 229712 529992 229764
rect 532700 229712 532752 229764
rect 555608 229712 555660 229764
rect 490656 229576 490708 229628
rect 497464 229576 497516 229628
rect 509516 229576 509568 229628
rect 666836 229644 666888 229696
rect 524972 229576 525024 229628
rect 532424 229576 532476 229628
rect 675852 229576 675904 229628
rect 677140 229576 677192 229628
rect 131120 229440 131172 229492
rect 197176 229440 197228 229492
rect 200212 229440 200264 229492
rect 200764 229440 200816 229492
rect 231124 229440 231176 229492
rect 277032 229440 277084 229492
rect 673828 229440 673880 229492
rect 448980 229372 449032 229424
rect 451372 229372 451424 229424
rect 122932 229304 122984 229356
rect 179144 229304 179196 229356
rect 181352 229304 181404 229356
rect 230664 229304 230716 229356
rect 453488 229304 453540 229356
rect 455788 229304 455840 229356
rect 673460 229304 673512 229356
rect 358084 229236 358136 229288
rect 360752 229236 360804 229288
rect 360936 229236 360988 229288
rect 363328 229236 363380 229288
rect 419448 229236 419500 229288
rect 424508 229236 424560 229288
rect 450268 229236 450320 229288
rect 451832 229236 451884 229288
rect 479892 229236 479944 229288
rect 482284 229236 482336 229288
rect 483756 229236 483808 229288
rect 486792 229236 486844 229288
rect 501788 229236 501840 229288
rect 507124 229236 507176 229288
rect 675852 229304 675904 229356
rect 677324 229304 677376 229356
rect 92480 229168 92532 229220
rect 146300 229168 146352 229220
rect 146944 229168 146996 229220
rect 153384 229168 153436 229220
rect 153844 229168 153896 229220
rect 163688 229168 163740 229220
rect 163872 229168 163924 229220
rect 166448 229168 166500 229220
rect 166908 229168 166960 229220
rect 172244 229168 172296 229220
rect 172428 229168 172480 229220
rect 220360 229168 220412 229220
rect 378968 229100 379020 229152
rect 383936 229100 383988 229152
rect 97908 229032 97960 229084
rect 107292 229032 107344 229084
rect 107476 229032 107528 229084
rect 102048 228896 102100 228948
rect 166908 228896 166960 228948
rect 82084 228624 82136 228676
rect 107108 228760 107160 228812
rect 107292 228760 107344 228812
rect 166448 228760 166500 228812
rect 96252 228624 96304 228676
rect 165436 228624 165488 228676
rect 168196 229032 168248 229084
rect 173992 229032 174044 229084
rect 174820 229032 174872 229084
rect 172244 228896 172296 228948
rect 175280 228896 175332 228948
rect 175648 228896 175700 228948
rect 168012 228760 168064 228812
rect 181260 228692 181312 228744
rect 179788 228624 179840 228676
rect 181720 229032 181772 229084
rect 192668 229032 192720 229084
rect 192852 229032 192904 229084
rect 194600 229032 194652 229084
rect 195612 229032 195664 229084
rect 250628 229032 250680 229084
rect 259276 229032 259328 229084
rect 298284 229032 298336 229084
rect 413836 229032 413888 229084
rect 420000 229100 420052 229152
rect 420184 229100 420236 229152
rect 421932 229100 421984 229152
rect 424324 229100 424376 229152
rect 427728 229100 427780 229152
rect 441252 229100 441304 229152
rect 442080 229100 442132 229152
rect 450912 229100 450964 229152
rect 452752 229100 452804 229152
rect 507584 229100 507636 229152
rect 511264 229100 511316 229152
rect 517888 229032 517940 229084
rect 540520 229032 540572 229084
rect 673598 229032 673650 229084
rect 675852 229032 675904 229084
rect 676404 229032 676456 229084
rect 181904 228896 181956 228948
rect 237104 228896 237156 228948
rect 251088 228896 251140 228948
rect 291200 228896 291252 228948
rect 319812 228896 319864 228948
rect 345940 228896 345992 228948
rect 350172 228896 350224 228948
rect 369124 228896 369176 228948
rect 507124 228896 507176 228948
rect 520096 228896 520148 228948
rect 526260 228896 526312 228948
rect 551560 228896 551612 228948
rect 673506 228828 673558 228880
rect 190552 228760 190604 228812
rect 190736 228760 190788 228812
rect 241612 228760 241664 228812
rect 246304 228760 246356 228812
rect 253848 228760 253900 228812
rect 255136 228760 255188 228812
rect 295708 228760 295760 228812
rect 317972 228760 318024 228812
rect 344652 228760 344704 228812
rect 346216 228760 346268 228812
rect 366548 228760 366600 228812
rect 376576 228760 376628 228812
rect 389732 228760 389784 228812
rect 401416 228760 401468 228812
rect 408408 228760 408460 228812
rect 493784 228760 493836 228812
rect 506020 228760 506072 228812
rect 519820 228760 519872 228812
rect 543188 228760 543240 228812
rect 675852 228760 675904 228812
rect 676220 228760 676272 228812
rect 231308 228624 231360 228676
rect 239404 228624 239456 228676
rect 284116 228624 284168 228676
rect 292396 228624 292448 228676
rect 326620 228624 326672 228676
rect 333244 228624 333296 228676
rect 355600 228624 355652 228676
rect 62764 228488 62816 228540
rect 140780 228488 140832 228540
rect 140964 228488 141016 228540
rect 66168 228352 66220 228404
rect 147634 228352 147686 228404
rect 153292 228488 153344 228540
rect 200580 228488 200632 228540
rect 200764 228488 200816 228540
rect 219348 228488 219400 228540
rect 267372 228488 267424 228540
rect 267556 228488 267608 228540
rect 307300 228488 307352 228540
rect 307668 228488 307720 228540
rect 335636 228488 335688 228540
rect 336648 228488 336700 228540
rect 358820 228488 358872 228540
rect 157432 228352 157484 228404
rect 157800 228352 157852 228404
rect 212172 228352 212224 228404
rect 226156 228352 226208 228404
rect 226340 228352 226392 228404
rect 273812 228352 273864 228404
rect 284116 228352 284168 228404
rect 320180 228352 320232 228404
rect 326896 228352 326948 228404
rect 351092 228352 351144 228404
rect 355232 228352 355284 228404
rect 369768 228624 369820 228676
rect 373816 228624 373868 228676
rect 387248 228624 387300 228676
rect 390284 228624 390336 228676
rect 400036 228624 400088 228676
rect 410892 228624 410944 228676
rect 416136 228624 416188 228676
rect 478788 228624 478840 228676
rect 483572 228624 483624 228676
rect 484124 228624 484176 228676
rect 490564 228624 490616 228676
rect 495348 228624 495400 228676
rect 511816 228624 511868 228676
rect 512092 228624 512144 228676
rect 533528 228624 533580 228676
rect 533988 228624 534040 228676
rect 561588 228624 561640 228676
rect 366916 228488 366968 228540
rect 382004 228488 382056 228540
rect 362868 228352 362920 228404
rect 379428 228352 379480 228404
rect 381728 228352 381780 228404
rect 392952 228488 393004 228540
rect 393228 228488 393280 228540
rect 391848 228352 391900 228404
rect 400128 228488 400180 228540
rect 407764 228488 407816 228540
rect 482468 228488 482520 228540
rect 494612 228488 494664 228540
rect 502432 228488 502484 228540
rect 520924 228488 520976 228540
rect 531412 228488 531464 228540
rect 558184 228488 558236 228540
rect 673388 228488 673440 228540
rect 671804 228420 671856 228472
rect 107108 228216 107160 228268
rect 140964 228216 141016 228268
rect 141148 228216 141200 228268
rect 190920 228216 190972 228268
rect 106188 228080 106240 228132
rect 107476 228080 107528 228132
rect 112996 228080 113048 228132
rect 122748 227944 122800 227996
rect 181076 227944 181128 227996
rect 181904 228080 181956 228132
rect 200764 228216 200816 228268
rect 201408 228216 201460 228268
rect 252560 228216 252612 228268
rect 277216 228216 277268 228268
rect 311808 228216 311860 228268
rect 402612 228352 402664 228404
rect 409788 228352 409840 228404
rect 415492 228352 415544 228404
rect 487620 228352 487672 228404
rect 501512 228352 501564 228404
rect 506296 228352 506348 228404
rect 525892 228352 525944 228404
rect 537852 228352 537904 228404
rect 566372 228352 566424 228404
rect 403900 228216 403952 228268
rect 479708 228216 479760 228268
rect 487804 228216 487856 228268
rect 671068 228216 671120 228268
rect 197912 228080 197964 228132
rect 204904 228080 204956 228132
rect 205364 228080 205416 228132
rect 257068 228080 257120 228132
rect 288164 228080 288216 228132
rect 321468 228080 321520 228132
rect 184940 227944 184992 227996
rect 186136 227944 186188 227996
rect 190736 227944 190788 227996
rect 190920 227944 190972 227996
rect 200212 227944 200264 227996
rect 200580 227944 200632 227996
rect 210700 227944 210752 227996
rect 212172 227944 212224 227996
rect 218428 227944 218480 227996
rect 226156 227944 226208 227996
rect 272524 227944 272576 227996
rect 369124 227876 369176 227928
rect 375564 227876 375616 227928
rect 407764 227876 407816 227928
rect 411628 227876 411680 227928
rect 471520 227876 471572 227928
rect 479340 227876 479392 227928
rect 673046 227876 673098 227928
rect 133788 227808 133840 227860
rect 200396 227808 200448 227860
rect 225696 227808 225748 227860
rect 226340 227808 226392 227860
rect 671804 227808 671856 227860
rect 242716 227740 242768 227792
rect 245660 227740 245712 227792
rect 255964 227740 256016 227792
rect 259000 227740 259052 227792
rect 366364 227740 366416 227792
rect 372988 227740 373040 227792
rect 393964 227740 394016 227792
rect 395528 227740 395580 227792
rect 396632 227740 396684 227792
rect 397460 227740 397512 227792
rect 402244 227740 402296 227792
rect 403256 227740 403308 227792
rect 404084 227740 404136 227792
rect 408868 227740 408920 227792
rect 409052 227740 409104 227792
rect 410340 227740 410392 227792
rect 411904 227740 411956 227792
rect 413560 227740 413612 227792
rect 416688 227740 416740 227792
rect 420644 227740 420696 227792
rect 475016 227740 475068 227792
rect 482928 227740 482980 227792
rect 110144 227672 110196 227724
rect 182364 227672 182416 227724
rect 185492 227672 185544 227724
rect 187516 227672 187568 227724
rect 191564 227672 191616 227724
rect 270132 227672 270184 227724
rect 306656 227672 306708 227724
rect 321376 227672 321428 227724
rect 346584 227672 346636 227724
rect 525524 227672 525576 227724
rect 537484 227672 537536 227724
rect 248052 227604 248104 227656
rect 465908 227604 465960 227656
rect 469864 227604 469916 227656
rect 672604 227604 672656 227656
rect 100668 227536 100720 227588
rect 174636 227536 174688 227588
rect 179052 227536 179104 227588
rect 236460 227536 236512 227588
rect 252468 227536 252520 227588
rect 293132 227536 293184 227588
rect 299296 227536 299348 227588
rect 328552 227536 328604 227588
rect 359372 227536 359424 227588
rect 374920 227536 374972 227588
rect 515864 227536 515916 227588
rect 538956 227536 539008 227588
rect 89628 227400 89680 227452
rect 159640 227400 159692 227452
rect 160008 227400 160060 227452
rect 166816 227400 166868 227452
rect 175188 227400 175240 227452
rect 231952 227400 232004 227452
rect 248236 227400 248288 227452
rect 291844 227400 291896 227452
rect 293776 227400 293828 227452
rect 325332 227400 325384 227452
rect 340604 227400 340656 227452
rect 361396 227400 361448 227452
rect 369768 227400 369820 227452
rect 385868 227400 385920 227452
rect 524328 227400 524380 227452
rect 547880 227400 547932 227452
rect 672448 227400 672500 227452
rect 676404 227332 676456 227384
rect 677048 227332 677100 227384
rect 86868 227264 86920 227316
rect 151912 227264 151964 227316
rect 152924 227264 152976 227316
rect 164332 227264 164384 227316
rect 165436 227264 165488 227316
rect 227444 227264 227496 227316
rect 75828 227128 75880 227180
rect 150164 227128 150216 227180
rect 150348 227128 150400 227180
rect 57888 226992 57940 227044
rect 134984 226992 135036 227044
rect 135444 226992 135496 227044
rect 151912 226992 151964 227044
rect 152280 227128 152332 227180
rect 168840 227128 168892 227180
rect 169576 227128 169628 227180
rect 228732 227128 228784 227180
rect 213276 226992 213328 227044
rect 226892 226992 226944 227044
rect 233240 227264 233292 227316
rect 234528 227264 234580 227316
rect 278320 227264 278372 227316
rect 280712 227264 280764 227316
rect 312084 227264 312136 227316
rect 326344 227264 326396 227316
rect 352380 227264 352432 227316
rect 355508 227264 355560 227316
rect 372344 227264 372396 227316
rect 235908 227128 235960 227180
rect 280252 227128 280304 227180
rect 296444 227128 296496 227180
rect 329196 227128 329248 227180
rect 329748 227128 329800 227180
rect 353668 227128 353720 227180
rect 354588 227128 354640 227180
rect 373632 227264 373684 227316
rect 382924 227264 382976 227316
rect 391664 227264 391716 227316
rect 395988 227264 396040 227316
rect 406476 227264 406528 227316
rect 485044 227264 485096 227316
rect 498752 227264 498804 227316
rect 501144 227264 501196 227316
rect 517796 227264 517848 227316
rect 521752 227264 521804 227316
rect 545120 227264 545172 227316
rect 373264 227128 373316 227180
rect 383292 227128 383344 227180
rect 386328 227128 386380 227180
rect 398748 227128 398800 227180
rect 481180 227128 481232 227180
rect 492956 227128 493008 227180
rect 498568 227128 498620 227180
rect 515864 227128 515916 227180
rect 516048 227128 516100 227180
rect 525064 227128 525116 227180
rect 535920 227128 535972 227180
rect 563888 227128 563940 227180
rect 672604 227060 672656 227112
rect 229054 226992 229106 227044
rect 271236 226992 271288 227044
rect 271788 226992 271840 227044
rect 308588 226992 308640 227044
rect 308772 226992 308824 227044
rect 336280 226992 336332 227044
rect 336464 226992 336516 227044
rect 360108 226992 360160 227044
rect 361212 226992 361264 227044
rect 377220 226992 377272 227044
rect 381912 226992 381964 227044
rect 396172 226992 396224 227044
rect 398472 226992 398524 227044
rect 408684 226992 408736 227044
rect 472164 226992 472216 227044
rect 481180 226992 481232 227044
rect 497280 226992 497332 227044
rect 106924 226856 106976 226908
rect 125784 226856 125836 226908
rect 121092 226720 121144 226772
rect 191104 226856 191156 226908
rect 200028 226856 200080 226908
rect 251916 226856 251968 226908
rect 272432 226856 272484 226908
rect 284760 226856 284812 226908
rect 514024 226992 514076 227044
rect 535644 226992 535696 227044
rect 537208 226992 537260 227044
rect 565636 226992 565688 227044
rect 514300 226856 514352 226908
rect 672494 226856 672546 226908
rect 119988 226584 120040 226636
rect 190092 226720 190144 226772
rect 195796 226720 195848 226772
rect 199476 226720 199528 226772
rect 212172 226720 212224 226772
rect 262220 226720 262272 226772
rect 672380 226720 672432 226772
rect 125784 226448 125836 226500
rect 135444 226584 135496 226636
rect 135628 226584 135680 226636
rect 129372 226448 129424 226500
rect 137192 226448 137244 226500
rect 137560 226584 137612 226636
rect 197452 226584 197504 226636
rect 222016 226584 222068 226636
rect 269948 226584 270000 226636
rect 668308 226584 668360 226636
rect 142114 226448 142166 226500
rect 142252 226448 142304 226500
rect 205548 226448 205600 226500
rect 213184 226448 213236 226500
rect 217784 226448 217836 226500
rect 221832 226448 221884 226500
rect 229008 226448 229060 226500
rect 232504 226448 232556 226500
rect 266728 226448 266780 226500
rect 666652 226448 666704 226500
rect 291844 226380 291896 226432
rect 295064 226380 295116 226432
rect 83464 226244 83516 226296
rect 69572 226108 69624 226160
rect 137468 226108 137520 226160
rect 137652 226108 137704 226160
rect 141516 226108 141568 226160
rect 141700 226108 141752 226160
rect 146760 226108 146812 226160
rect 166816 226312 166868 226364
rect 221004 226312 221056 226364
rect 152832 226244 152884 226296
rect 161940 226244 161992 226296
rect 162308 226244 162360 226296
rect 166632 226244 166684 226296
rect 222476 226244 222528 226296
rect 225512 226244 225564 226296
rect 228732 226244 228784 226296
rect 275100 226244 275152 226296
rect 278504 226244 278556 226296
rect 315028 226244 315080 226296
rect 317328 226244 317380 226296
rect 334256 226244 334308 226296
rect 503260 226244 503312 226296
rect 510160 226244 510212 226296
rect 529940 226244 529992 226296
rect 544936 226244 544988 226296
rect 562324 226244 562376 226296
rect 567568 226244 567620 226296
rect 672034 226244 672086 226296
rect 157432 226108 157484 226160
rect 157616 226108 157668 226160
rect 215852 226108 215904 226160
rect 216496 226108 216548 226160
rect 264796 226108 264848 226160
rect 266268 226108 266320 226160
rect 303436 226108 303488 226160
rect 325424 226108 325476 226160
rect 349160 226108 349212 226160
rect 510804 226108 510856 226160
rect 531688 226108 531740 226160
rect 666008 226040 666060 226092
rect 93768 225972 93820 226024
rect 166816 225972 166868 226024
rect 166954 225972 167006 226024
rect 176476 225972 176528 226024
rect 178684 225972 178736 226024
rect 187148 225972 187200 226024
rect 187332 225972 187384 226024
rect 224224 225972 224276 226024
rect 95148 225836 95200 225888
rect 161204 225836 161256 225888
rect 161940 225836 161992 225888
rect 176108 225836 176160 225888
rect 177212 225836 177264 225888
rect 233884 225972 233936 226024
rect 243452 225972 243504 226024
rect 248696 225972 248748 226024
rect 267694 225972 267746 226024
rect 304080 225972 304132 226024
rect 313096 225972 313148 226024
rect 340788 225972 340840 226024
rect 64788 225700 64840 225752
rect 92480 225700 92532 225752
rect 108304 225700 108356 225752
rect 176476 225700 176528 225752
rect 176660 225700 176712 225752
rect 185676 225700 185728 225752
rect 187516 225700 187568 225752
rect 239036 225836 239088 225888
rect 249708 225836 249760 225888
rect 290556 225836 290608 225888
rect 294972 225836 295024 225888
rect 325976 225836 326028 225888
rect 340144 225836 340196 225888
rect 347872 225972 347924 226024
rect 349068 225972 349120 226024
rect 367192 225972 367244 226024
rect 518532 225972 518584 226024
rect 541440 225972 541492 226024
rect 544200 225972 544252 226024
rect 562692 225972 562744 226024
rect 347044 225836 347096 225888
rect 365904 225836 365956 225888
rect 367652 225836 367704 225888
rect 380072 225836 380124 225888
rect 488908 225836 488960 225888
rect 502984 225836 503036 225888
rect 528192 225836 528244 225888
rect 554044 225836 554096 225888
rect 458640 225768 458692 225820
rect 462964 225768 463016 225820
rect 61292 225564 61344 225616
rect 136824 225564 136876 225616
rect 137008 225564 137060 225616
rect 146944 225564 146996 225616
rect 147128 225564 147180 225616
rect 201040 225564 201092 225616
rect 222476 225564 222528 225616
rect 224224 225564 224276 225616
rect 242900 225700 242952 225752
rect 257712 225700 257764 225752
rect 299572 225700 299624 225752
rect 304908 225700 304960 225752
rect 333704 225700 333756 225752
rect 335268 225700 335320 225752
rect 356888 225700 356940 225752
rect 379336 225700 379388 225752
rect 393596 225700 393648 225752
rect 394608 225700 394660 225752
rect 404544 225700 404596 225752
rect 491484 225700 491536 225752
rect 506848 225700 506900 225752
rect 507308 225700 507360 225752
rect 526720 225700 526772 225752
rect 527548 225700 527600 225752
rect 553216 225700 553268 225752
rect 671820 225700 671872 225752
rect 234344 225564 234396 225616
rect 281540 225564 281592 225616
rect 285496 225564 285548 225616
rect 318892 225564 318944 225616
rect 322848 225564 322900 225616
rect 349804 225564 349856 225616
rect 351184 225564 351236 225616
rect 370412 225564 370464 225616
rect 372528 225564 372580 225616
rect 388076 225564 388128 225616
rect 388444 225564 388496 225616
rect 399392 225564 399444 225616
rect 467656 225564 467708 225616
rect 476580 225564 476632 225616
rect 477316 225564 477368 225616
rect 489184 225564 489236 225616
rect 495164 225564 495216 225616
rect 509700 225564 509752 225616
rect 510344 225564 510396 225616
rect 530492 225564 530544 225616
rect 532056 225564 532108 225616
rect 559012 225564 559064 225616
rect 103428 225428 103480 225480
rect 108304 225428 108356 225480
rect 106004 225292 106056 225344
rect 127440 225428 127492 225480
rect 117228 225292 117280 225344
rect 185492 225428 185544 225480
rect 187332 225428 187384 225480
rect 195796 225428 195848 225480
rect 199384 225428 199436 225480
rect 200488 225428 200540 225480
rect 127440 225156 127492 225208
rect 137008 225292 137060 225344
rect 128268 225156 128320 225208
rect 146944 225292 146996 225344
rect 147128 225292 147180 225344
rect 671712 225496 671764 225548
rect 201040 225428 201092 225480
rect 242256 225428 242308 225480
rect 669412 225428 669464 225480
rect 463148 225360 463200 225412
rect 467288 225360 467340 225412
rect 126888 225020 126940 225072
rect 185676 225156 185728 225208
rect 187332 225156 187384 225208
rect 200580 225156 200632 225208
rect 207756 225292 207808 225344
rect 208032 225292 208084 225344
rect 260932 225292 260984 225344
rect 671068 225224 671120 225276
rect 202512 225156 202564 225208
rect 202696 225156 202748 225208
rect 254492 225156 254544 225208
rect 137468 225020 137520 225072
rect 143540 225020 143592 225072
rect 146944 225020 146996 225072
rect 162308 225020 162360 225072
rect 162492 225020 162544 225072
rect 166448 225020 166500 225072
rect 166816 225020 166868 225072
rect 167000 225020 167052 225072
rect 167368 225020 167420 225072
rect 185676 225020 185728 225072
rect 187056 225020 187108 225072
rect 223580 225020 223632 225072
rect 224868 225020 224920 225072
rect 270592 225020 270644 225072
rect 668308 225020 668360 225072
rect 275836 224952 275888 225004
rect 276848 224952 276900 225004
rect 282736 224952 282788 225004
rect 285312 224952 285364 225004
rect 489920 224952 489972 225004
rect 494796 224952 494848 225004
rect 509240 224952 509292 225004
rect 512644 224952 512696 225004
rect 122564 224884 122616 224936
rect 193956 224884 194008 224936
rect 194508 224884 194560 224936
rect 247408 224884 247460 224936
rect 264152 224884 264204 224936
rect 269304 224884 269356 224936
rect 285680 224884 285732 224936
rect 316316 224884 316368 224936
rect 406752 224884 406804 224936
rect 414848 224884 414900 224936
rect 516784 224884 516836 224936
rect 531320 224884 531372 224936
rect 667940 224884 667992 224936
rect 668308 224884 668360 224936
rect 671068 224884 671120 224936
rect 115848 224748 115900 224800
rect 116768 224612 116820 224664
rect 118148 224612 118200 224664
rect 118792 224748 118844 224800
rect 191380 224748 191432 224800
rect 192484 224748 192536 224800
rect 246764 224748 246816 224800
rect 247592 224748 247644 224800
rect 289268 224748 289320 224800
rect 315856 224748 315908 224800
rect 341432 224748 341484 224800
rect 532424 224748 532476 224800
rect 549904 224748 549956 224800
rect 460572 224680 460624 224732
rect 463148 224680 463200 224732
rect 188804 224612 188856 224664
rect 195612 224612 195664 224664
rect 248880 224612 248932 224664
rect 249064 224612 249116 224664
rect 263876 224612 263928 224664
rect 271604 224612 271656 224664
rect 309876 224612 309928 224664
rect 319996 224612 320048 224664
rect 347228 224612 347280 224664
rect 514668 224612 514720 224664
rect 536656 224612 536708 224664
rect 667940 224612 667992 224664
rect 456064 224544 456116 224596
rect 459652 224544 459704 224596
rect 60648 224476 60700 224528
rect 103612 224476 103664 224528
rect 108672 224476 108724 224528
rect 118608 224476 118660 224528
rect 126704 224476 126756 224528
rect 131120 224476 131172 224528
rect 131304 224476 131356 224528
rect 196532 224476 196584 224528
rect 201224 224476 201276 224528
rect 255780 224476 255832 224528
rect 261852 224476 261904 224528
rect 300860 224476 300912 224528
rect 303252 224476 303304 224528
rect 333060 224476 333112 224528
rect 333888 224476 333940 224528
rect 356244 224476 356296 224528
rect 357348 224476 357400 224528
rect 374276 224476 374328 224528
rect 479524 224476 479576 224528
rect 486608 224476 486660 224528
rect 508228 224476 508280 224528
rect 528376 224476 528428 224528
rect 530124 224476 530176 224528
rect 556528 224476 556580 224528
rect 671022 224408 671074 224460
rect 82728 224340 82780 224392
rect 157294 224340 157346 224392
rect 157432 224340 157484 224392
rect 170956 224340 171008 224392
rect 171094 224340 171146 224392
rect 186872 224340 186924 224392
rect 188988 224340 189040 224392
rect 243820 224340 243872 224392
rect 246948 224340 247000 224392
rect 288624 224340 288676 224392
rect 289636 224340 289688 224392
rect 307852 224340 307904 224392
rect 308956 224340 309008 224392
rect 339500 224340 339552 224392
rect 344652 224340 344704 224392
rect 364616 224340 364668 224392
rect 375288 224340 375340 224392
rect 387800 224340 387852 224392
rect 462504 224340 462556 224392
rect 469312 224340 469364 224392
rect 470232 224340 470284 224392
rect 479708 224340 479760 224392
rect 486792 224340 486844 224392
rect 496912 224340 496964 224392
rect 499212 224340 499264 224392
rect 516784 224340 516836 224392
rect 525708 224340 525760 224392
rect 550640 224340 550692 224392
rect 58992 224204 59044 224256
rect 116768 224204 116820 224256
rect 116952 224204 117004 224256
rect 118424 224204 118476 224256
rect 118608 224204 118660 224256
rect 183836 224204 183888 224256
rect 184664 224204 184716 224256
rect 239680 224204 239732 224256
rect 241980 224204 242032 224256
rect 104808 224068 104860 224120
rect 117964 224068 118016 224120
rect 118148 224068 118200 224120
rect 76564 223932 76616 223984
rect 142160 223932 142212 223984
rect 142620 224068 142672 224120
rect 209412 224068 209464 224120
rect 209688 224068 209740 224120
rect 259644 224068 259696 224120
rect 282552 224204 282604 224256
rect 285680 224204 285732 224256
rect 288348 224204 288400 224256
rect 322388 224204 322440 224256
rect 342076 224204 342128 224256
rect 364800 224204 364852 224256
rect 364984 224204 365036 224256
rect 378140 224204 378192 224256
rect 389088 224204 389140 224256
rect 400956 224204 401008 224256
rect 416504 224204 416556 224256
rect 422208 224204 422260 224256
rect 423312 224204 423364 224256
rect 424324 224204 424376 224256
rect 451372 224204 451424 224256
rect 452200 224204 452252 224256
rect 474740 224204 474792 224256
rect 484584 224204 484636 224256
rect 485688 224204 485740 224256
rect 499396 224204 499448 224256
rect 508872 224204 508924 224256
rect 529388 224204 529440 224256
rect 535276 224204 535328 224256
rect 563796 224204 563848 224256
rect 567844 224204 567896 224256
rect 568948 224204 569000 224256
rect 669412 224136 669464 224188
rect 285036 224068 285088 224120
rect 286692 224068 286744 224120
rect 319536 224068 319588 224120
rect 145196 223932 145248 223984
rect 147680 223932 147732 223984
rect 154580 223932 154632 223984
rect 156880 223932 156932 223984
rect 217140 223932 217192 223984
rect 217324 223932 217376 223984
rect 228088 223932 228140 223984
rect 231308 223932 231360 223984
rect 278964 223932 279016 223984
rect 117964 223796 118016 223848
rect 122932 223796 122984 223848
rect 125232 223796 125284 223848
rect 131304 223796 131356 223848
rect 134984 223796 135036 223848
rect 204260 223796 204312 223848
rect 205272 223796 205324 223848
rect 212632 223796 212684 223848
rect 215944 223796 215996 223848
rect 222936 223796 222988 223848
rect 238668 223796 238720 223848
rect 282368 223796 282420 223848
rect 132408 223660 132460 223712
rect 201684 223660 201736 223712
rect 85488 223524 85540 223576
rect 161940 223524 161992 223576
rect 162124 223524 162176 223576
rect 167828 223524 167880 223576
rect 168288 223524 168340 223576
rect 226708 223524 226760 223576
rect 269028 223524 269080 223576
rect 298008 223524 298060 223576
rect 300124 223524 300176 223576
rect 426440 223592 426492 223644
rect 426992 223592 427044 223644
rect 306012 223524 306064 223576
rect 329104 223524 329156 223576
rect 342720 223524 342772 223576
rect 457996 223524 458048 223576
rect 460204 223524 460256 223576
rect 473452 223524 473504 223576
rect 475568 223524 475620 223576
rect 679256 223524 679308 223576
rect 680176 223524 680228 223576
rect 112812 223388 112864 223440
rect 185860 223388 185912 223440
rect 203892 223388 203944 223440
rect 254860 223388 254912 223440
rect 260104 223388 260156 223440
rect 298928 223388 298980 223440
rect 302148 223388 302200 223440
rect 331128 223388 331180 223440
rect 518900 223388 518952 223440
rect 530032 223388 530084 223440
rect 81348 223252 81400 223304
rect 156880 223252 156932 223304
rect 157432 223252 157484 223304
rect 159824 223252 159876 223304
rect 160928 223252 160980 223304
rect 164516 223252 164568 223304
rect 78588 223116 78640 223168
rect 157064 223116 157116 223168
rect 157248 223116 157300 223168
rect 161204 223116 161256 223168
rect 161388 223116 161440 223168
rect 89444 222980 89496 223032
rect 162124 222980 162176 223032
rect 164148 223116 164200 223168
rect 224040 223252 224092 223304
rect 264796 223252 264848 223304
rect 304724 223252 304776 223304
rect 306288 223252 306340 223304
rect 336924 223252 336976 223304
rect 343548 223252 343600 223304
rect 363972 223252 364024 223304
rect 489552 223252 489604 223304
rect 504364 223252 504416 223304
rect 505100 223252 505152 223304
rect 523960 223252 524012 223304
rect 529020 223252 529072 223304
rect 543648 223252 543700 223304
rect 165068 223116 165120 223168
rect 222292 223116 222344 223168
rect 224224 223116 224276 223168
rect 238392 223116 238444 223168
rect 245292 223116 245344 223168
rect 287612 223116 287664 223168
rect 290832 223116 290884 223168
rect 323676 223116 323728 223168
rect 330484 223116 330536 223168
rect 354956 223116 355008 223168
rect 357072 223116 357124 223168
rect 376208 223116 376260 223168
rect 490196 223116 490248 223168
rect 505652 223116 505704 223168
rect 513104 223116 513156 223168
rect 534448 223116 534500 223168
rect 534724 223116 534776 223168
rect 547420 223116 547472 223168
rect 92112 222844 92164 222896
rect 166448 222844 166500 222896
rect 166954 222980 167006 223032
rect 176108 222980 176160 223032
rect 176292 222980 176344 223032
rect 234804 222980 234856 223032
rect 235172 222980 235224 223032
rect 243268 222980 243320 223032
rect 250904 222980 250956 223032
rect 294420 222980 294472 223032
rect 300308 222980 300360 223032
rect 331312 222980 331364 223032
rect 337936 222980 337988 223032
rect 359188 222980 359240 223032
rect 370504 222980 370556 223032
rect 384580 222980 384632 223032
rect 387708 222980 387760 223032
rect 398104 222980 398156 223032
rect 501788 222980 501840 223032
rect 519268 222980 519320 223032
rect 523684 222980 523736 223032
rect 548064 222980 548116 223032
rect 549260 222980 549312 223032
rect 564808 222980 564860 223032
rect 566832 222912 566884 222964
rect 576400 222912 576452 222964
rect 221648 222844 221700 222896
rect 231952 222844 232004 222896
rect 277676 222844 277728 222896
rect 283380 222844 283432 222896
rect 316960 222844 317012 222896
rect 317144 222844 317196 222896
rect 343364 222844 343416 222896
rect 347596 222844 347648 222896
rect 368480 222844 368532 222896
rect 375104 222844 375156 222896
rect 391020 222844 391072 222896
rect 397368 222844 397420 222896
rect 407120 222844 407172 222896
rect 408408 222844 408460 222896
rect 416872 222844 416924 222896
rect 420828 222844 420880 222896
rect 425152 222844 425204 222896
rect 459928 222844 459980 222896
rect 467104 222844 467156 222896
rect 467472 222844 467524 222896
rect 473728 222844 473780 222896
rect 478328 222844 478380 222896
rect 486148 222844 486200 222896
rect 486976 222844 487028 222896
rect 501052 222844 501104 222896
rect 504640 222844 504692 222896
rect 523776 222844 523828 222896
rect 533712 222844 533764 222896
rect 560668 222844 560720 222896
rect 563796 222776 563848 222828
rect 569960 222776 570012 222828
rect 87972 222708 88024 222760
rect 160928 222708 160980 222760
rect 161204 222708 161256 222760
rect 99288 222572 99340 222624
rect 175464 222572 175516 222624
rect 176108 222708 176160 222760
rect 192024 222708 192076 222760
rect 192300 222708 192352 222760
rect 207480 222708 207532 222760
rect 209504 222708 209556 222760
rect 210240 222708 210292 222760
rect 213828 222708 213880 222760
rect 262864 222708 262916 222760
rect 263508 222708 263560 222760
rect 296904 222708 296956 222760
rect 562508 222640 562560 222692
rect 564624 222640 564676 222692
rect 564808 222640 564860 222692
rect 574100 222640 574152 222692
rect 56508 222436 56560 222488
rect 133512 222436 133564 222488
rect 142988 222436 143040 222488
rect 143356 222436 143408 222488
rect 144828 222436 144880 222488
rect 145012 222436 145064 222488
rect 151360 222436 151412 222488
rect 154212 222436 154264 222488
rect 214380 222436 214432 222488
rect 214748 222572 214800 222624
rect 260288 222572 260340 222624
rect 219716 222436 219768 222488
rect 220084 222436 220136 222488
rect 268660 222436 268712 222488
rect 142344 222300 142396 222352
rect 144276 222300 144328 222352
rect 208768 222300 208820 222352
rect 210976 222300 211028 222352
rect 214748 222300 214800 222352
rect 220452 222300 220504 222352
rect 268016 222300 268068 222352
rect 214932 222232 214984 222284
rect 216220 222232 216272 222284
rect 107844 222096 107896 222148
rect 171048 222096 171100 222148
rect 104532 221960 104584 222012
rect 174912 222164 174964 222216
rect 176292 222164 176344 222216
rect 482928 222164 482980 222216
rect 562508 222232 562560 222284
rect 571708 222504 571760 222556
rect 567384 222368 567436 222420
rect 572812 222504 572864 222556
rect 564624 222232 564676 222284
rect 593972 222368 594024 222420
rect 178224 222096 178276 222148
rect 176108 222028 176160 222080
rect 71412 221824 71464 221876
rect 68100 221688 68152 221740
rect 142114 221688 142166 221740
rect 142344 221688 142396 221740
rect 144460 221688 144512 221740
rect 146208 221688 146260 221740
rect 149244 221824 149296 221876
rect 61476 221552 61528 221604
rect 137284 221552 137336 221604
rect 137468 221552 137520 221604
rect 152096 221688 152148 221740
rect 162124 221824 162176 221876
rect 172980 221960 173032 222012
rect 176292 221960 176344 222012
rect 180616 221960 180668 222012
rect 181628 222096 181680 222148
rect 240140 222096 240192 222148
rect 261024 222096 261076 222148
rect 301688 222096 301740 222148
rect 331404 222096 331456 222148
rect 353944 222096 353996 222148
rect 424968 222096 425020 222148
rect 429292 222096 429344 222148
rect 462136 222096 462188 222148
rect 468760 222096 468812 222148
rect 471888 222096 471940 222148
rect 477868 222096 477920 222148
rect 553584 222096 553636 222148
rect 563704 222096 563756 222148
rect 597560 222232 597612 222284
rect 593236 222096 593288 222148
rect 607496 222096 607548 222148
rect 237564 221960 237616 222012
rect 243636 221960 243688 222012
rect 285864 221960 285916 222012
rect 309876 221960 309928 222012
rect 338396 221960 338448 222012
rect 529756 221960 529808 222012
rect 555792 221960 555844 222012
rect 556804 221960 556856 222012
rect 562692 221960 562744 222012
rect 563428 221960 563480 222012
rect 569316 221960 569368 222012
rect 569592 221960 569644 222012
rect 596456 221960 596508 222012
rect 596640 221960 596692 222012
rect 171508 221824 171560 221876
rect 229652 221824 229704 221876
rect 230388 221824 230440 221876
rect 258724 221824 258776 221876
rect 267832 221824 267884 221876
rect 273996 221824 274048 221876
rect 303712 221824 303764 221876
rect 334072 221824 334124 221876
rect 496176 221824 496228 221876
rect 513380 221824 513432 221876
rect 515404 221824 515456 221876
rect 535000 221824 535052 221876
rect 545120 221824 545172 221876
rect 596824 221824 596876 221876
rect 597192 221960 597244 222012
rect 607312 221960 607364 222012
rect 606024 221824 606076 221876
rect 162308 221688 162360 221740
rect 162676 221688 162728 221740
rect 224500 221688 224552 221740
rect 227076 221688 227128 221740
rect 272708 221688 272760 221740
rect 275100 221688 275152 221740
rect 310888 221688 310940 221740
rect 311532 221688 311584 221740
rect 338580 221688 338632 221740
rect 64604 221416 64656 221468
rect 142114 221416 142166 221468
rect 142252 221416 142304 221468
rect 144000 221416 144052 221468
rect 144460 221416 144512 221468
rect 146668 221416 146720 221468
rect 204904 221552 204956 221604
rect 205088 221552 205140 221604
rect 214196 221552 214248 221604
rect 214656 221552 214708 221604
rect 258540 221552 258592 221604
rect 258724 221552 258776 221604
rect 275284 221552 275336 221604
rect 278320 221552 278372 221604
rect 313280 221552 313332 221604
rect 314476 221552 314528 221604
rect 341616 221688 341668 221740
rect 359556 221688 359608 221740
rect 376852 221688 376904 221740
rect 500040 221688 500092 221740
rect 518440 221688 518492 221740
rect 522856 221688 522908 221740
rect 546592 221688 546644 221740
rect 547144 221688 547196 221740
rect 556712 221688 556764 221740
rect 557816 221688 557868 221740
rect 558276 221688 558328 221740
rect 562876 221688 562928 221740
rect 563060 221688 563112 221740
rect 566648 221688 566700 221740
rect 567384 221688 567436 221740
rect 567752 221688 567804 221740
rect 569592 221688 569644 221740
rect 569960 221688 570012 221740
rect 610532 221688 610584 221740
rect 341340 221552 341392 221604
rect 361580 221552 361632 221604
rect 162124 221416 162176 221468
rect 162308 221416 162360 221468
rect 95424 221280 95476 221332
rect 114468 221280 114520 221332
rect 185124 221280 185176 221332
rect 185768 221416 185820 221468
rect 232136 221416 232188 221468
rect 241152 221416 241204 221468
rect 285864 221416 285916 221468
rect 286048 221416 286100 221468
rect 289820 221416 289872 221468
rect 290004 221416 290056 221468
rect 321744 221416 321796 221468
rect 338856 221416 338908 221468
rect 362224 221552 362276 221604
rect 377772 221552 377824 221604
rect 390008 221552 390060 221604
rect 456708 221552 456760 221604
rect 462136 221552 462188 221604
rect 484308 221552 484360 221604
rect 496084 221552 496136 221604
rect 503444 221552 503496 221604
rect 521752 221552 521804 221604
rect 525892 221552 525944 221604
rect 601516 221552 601568 221604
rect 362040 221416 362092 221468
rect 379888 221416 379940 221468
rect 391020 221416 391072 221468
rect 400404 221416 400456 221468
rect 405096 221416 405148 221468
rect 414204 221416 414256 221468
rect 452568 221416 452620 221468
rect 456708 221416 456760 221468
rect 483756 221416 483808 221468
rect 538680 221416 538732 221468
rect 543280 221416 543332 221468
rect 596640 221416 596692 221468
rect 596824 221416 596876 221468
rect 606668 221552 606720 221604
rect 655704 221552 655756 221604
rect 659292 221552 659344 221604
rect 654232 221416 654284 221468
rect 655520 221416 655572 221468
rect 195244 221280 195296 221332
rect 195428 221280 195480 221332
rect 245108 221280 245160 221332
rect 258540 221280 258592 221332
rect 265716 221280 265768 221332
rect 273444 221280 273496 221332
rect 309232 221280 309284 221332
rect 542912 221212 542964 221264
rect 550364 221212 550416 221264
rect 550640 221212 550692 221264
rect 551284 221212 551336 221264
rect 569132 221212 569184 221264
rect 569316 221212 569368 221264
rect 610072 221212 610124 221264
rect 137100 221144 137152 221196
rect 137284 221144 137336 221196
rect 142114 221144 142166 221196
rect 142252 221144 142304 221196
rect 203248 221144 203300 221196
rect 117780 221008 117832 221060
rect 180754 221008 180806 221060
rect 180892 221008 180944 221060
rect 185768 221008 185820 221060
rect 185952 221008 186004 221060
rect 187884 221008 187936 221060
rect 188160 221008 188212 221060
rect 128544 220872 128596 220924
rect 195244 221008 195296 221060
rect 205088 221144 205140 221196
rect 206008 221144 206060 221196
rect 258356 221144 258408 221196
rect 548064 221076 548116 221128
rect 593236 221076 593288 221128
rect 596456 221076 596508 221128
rect 204904 221008 204956 221060
rect 211620 221008 211672 221060
rect 237104 221008 237156 221060
rect 280436 221008 280488 221060
rect 415032 221008 415084 221060
rect 420184 221008 420236 221060
rect 545120 221008 545172 221060
rect 545764 221008 545816 221060
rect 552848 220940 552900 220992
rect 553216 220940 553268 220992
rect 567752 220940 567804 220992
rect 569132 220940 569184 220992
rect 597192 220940 597244 220992
rect 597560 221076 597612 221128
rect 608692 221076 608744 221128
rect 608876 220940 608928 220992
rect 91284 220736 91336 220788
rect 97724 220600 97776 220652
rect 162308 220736 162360 220788
rect 172704 220736 172756 220788
rect 173348 220736 173400 220788
rect 182640 220736 182692 220788
rect 183100 220736 183152 220788
rect 184204 220736 184256 220788
rect 190460 220736 190512 220788
rect 194784 220736 194836 220788
rect 195428 220872 195480 220924
rect 198924 220872 198976 220924
rect 203248 220872 203300 220924
rect 206376 220872 206428 220924
rect 256056 220872 256108 220924
rect 261392 220872 261444 220924
rect 420644 220804 420696 220856
rect 423772 220804 423824 220856
rect 466092 220804 466144 220856
rect 470600 220804 470652 220856
rect 518440 220804 518492 220856
rect 591948 220804 592000 220856
rect 196072 220736 196124 220788
rect 197728 220736 197780 220788
rect 198096 220736 198148 220788
rect 252744 220736 252796 220788
rect 253572 220736 253624 220788
rect 293316 220736 293368 220788
rect 293592 220736 293644 220788
rect 299940 220736 299992 220788
rect 306748 220736 306800 220788
rect 320364 220736 320416 220788
rect 329564 220736 329616 220788
rect 331956 220736 332008 220788
rect 414204 220736 414256 220788
rect 418252 220736 418304 220788
rect 455236 220736 455288 220788
rect 458824 220736 458876 220788
rect 475384 220736 475436 220788
rect 476212 220736 476264 220788
rect 476764 220736 476816 220788
rect 478696 220736 478748 220788
rect 504180 220736 504232 220788
rect 515772 220736 515824 220788
rect 592132 220736 592184 220788
rect 620284 220736 620336 220788
rect 465724 220668 465776 220720
rect 469588 220668 469640 220720
rect 676036 220668 676088 220720
rect 677416 220668 677468 220720
rect 83004 220464 83056 220516
rect 157340 220464 157392 220516
rect 157524 220464 157576 220516
rect 167184 220600 167236 220652
rect 170772 220600 170824 220652
rect 76380 220328 76432 220380
rect 150716 220328 150768 220380
rect 150900 220328 150952 220380
rect 161756 220328 161808 220380
rect 162308 220464 162360 220516
rect 162860 220464 162912 220516
rect 173532 220464 173584 220516
rect 177396 220600 177448 220652
rect 234068 220600 234120 220652
rect 254400 220600 254452 220652
rect 296720 220600 296772 220652
rect 299940 220600 299992 220652
rect 330024 220600 330076 220652
rect 474004 220600 474056 220652
rect 475384 220600 475436 220652
rect 511264 220600 511316 220652
rect 527548 220600 527600 220652
rect 542728 220600 542780 220652
rect 543648 220600 543700 220652
rect 545948 220600 546000 220652
rect 546132 220600 546184 220652
rect 550272 220600 550324 220652
rect 550548 220600 550600 220652
rect 553768 220600 553820 220652
rect 555608 220600 555660 220652
rect 559840 220600 559892 220652
rect 626632 220600 626684 220652
rect 229284 220464 229336 220516
rect 240324 220464 240376 220516
rect 283012 220464 283064 220516
rect 296628 220464 296680 220516
rect 327540 220464 327592 220516
rect 328092 220464 328144 220516
rect 351368 220464 351420 220516
rect 371148 220464 371200 220516
rect 385224 220464 385276 220516
rect 482284 220464 482336 220516
rect 491944 220464 491996 220516
rect 493968 220464 494020 220516
rect 508504 220464 508556 220516
rect 522304 220464 522356 220516
rect 540060 220464 540112 220516
rect 622676 220464 622728 220516
rect 218612 220328 218664 220380
rect 229744 220328 229796 220380
rect 276112 220328 276164 220380
rect 280068 220328 280120 220380
rect 313924 220328 313976 220380
rect 323124 220328 323176 220380
rect 348148 220328 348200 220380
rect 352932 220328 352984 220380
rect 371424 220328 371476 220380
rect 481548 220328 481600 220380
rect 492772 220328 492824 220380
rect 496360 220328 496412 220380
rect 510988 220328 511040 220380
rect 517428 220328 517480 220380
rect 539140 220328 539192 220380
rect 541716 220328 541768 220380
rect 554964 220328 555016 220380
rect 66444 220192 66496 220244
rect 142114 220192 142166 220244
rect 142252 220192 142304 220244
rect 205732 220192 205784 220244
rect 211344 220192 211396 220244
rect 263048 220192 263100 220244
rect 263324 220192 263376 220244
rect 301044 220192 301096 220244
rect 311808 220192 311860 220244
rect 327264 220192 327316 220244
rect 332232 220192 332284 220244
rect 357532 220192 357584 220244
rect 360384 220192 360436 220244
rect 377404 220192 377456 220244
rect 390100 220192 390152 220244
rect 401692 220192 401744 220244
rect 432236 220192 432288 220244
rect 434812 220192 434864 220244
rect 459468 220192 459520 220244
rect 465448 220192 465500 220244
rect 469036 220192 469088 220244
rect 474556 220192 474608 220244
rect 478512 220192 478564 220244
rect 489460 220192 489512 220244
rect 492312 220192 492364 220244
rect 507676 220192 507728 220244
rect 521568 220192 521620 220244
rect 544200 220192 544252 220244
rect 63132 220056 63184 220108
rect 146484 220056 146536 220108
rect 147588 220056 147640 220108
rect 204536 220056 204588 220108
rect 204720 220056 204772 220108
rect 214012 220056 214064 220108
rect 217140 220056 217192 220108
rect 265164 220056 265216 220108
rect 280896 220056 280948 220108
rect 317512 220056 317564 220108
rect 318156 220056 318208 220108
rect 343732 220056 343784 220108
rect 345480 220056 345532 220108
rect 367376 220056 367428 220108
rect 367836 220056 367888 220108
rect 382464 220056 382516 220108
rect 382740 220056 382792 220108
rect 394792 220056 394844 220108
rect 397644 220056 397696 220108
rect 405832 220056 405884 220108
rect 421656 220056 421708 220108
rect 426808 220056 426860 220108
rect 427912 220056 427964 220108
rect 428740 220056 428792 220108
rect 472992 220056 473044 220108
rect 482008 220056 482060 220108
rect 488264 220056 488316 220108
rect 502708 220056 502760 220108
rect 507032 220056 507084 220108
rect 522580 220056 522632 220108
rect 527824 220056 527876 220108
rect 552480 220192 552532 220244
rect 559564 220328 559616 220380
rect 567200 220328 567252 220380
rect 567384 220328 567436 220380
rect 572352 220328 572404 220380
rect 572812 220328 572864 220380
rect 582196 220328 582248 220380
rect 582380 220328 582432 220380
rect 591856 220328 591908 220380
rect 591994 220328 592046 220380
rect 628196 220328 628248 220380
rect 562692 220192 562744 220244
rect 563060 220192 563112 220244
rect 620100 220192 620152 220244
rect 620284 220192 620336 220244
rect 628012 220192 628064 220244
rect 625528 220056 625580 220108
rect 647240 220056 647292 220108
rect 652760 220056 652812 220108
rect 553216 219988 553268 220040
rect 553584 219988 553636 220040
rect 553768 219988 553820 220040
rect 558000 219988 558052 220040
rect 111248 219920 111300 219972
rect 173348 219920 173400 219972
rect 173532 219920 173584 219972
rect 124404 219784 124456 219836
rect 193312 219784 193364 219836
rect 195428 219920 195480 219972
rect 244464 219920 244516 219972
rect 256884 219920 256936 219972
rect 295892 219920 295944 219972
rect 296812 219920 296864 219972
rect 310704 219920 310756 219972
rect 540796 219852 540848 219904
rect 548892 219852 548944 219904
rect 550088 219852 550140 219904
rect 625344 219852 625396 219904
rect 204720 219784 204772 219836
rect 131028 219648 131080 219700
rect 190460 219648 190512 219700
rect 190644 219648 190696 219700
rect 195428 219648 195480 219700
rect 197268 219648 197320 219700
rect 249892 219784 249944 219836
rect 531320 219716 531372 219768
rect 532608 219716 532660 219768
rect 621020 219716 621072 219768
rect 207204 219648 207256 219700
rect 257252 219648 257304 219700
rect 520096 219648 520148 219700
rect 464988 219580 465040 219632
rect 472072 219580 472124 219632
rect 618260 219580 618312 219632
rect 620100 219580 620152 219632
rect 626816 219580 626868 219632
rect 137652 219512 137704 219564
rect 140780 219512 140832 219564
rect 140964 219512 141016 219564
rect 141976 219512 142028 219564
rect 142160 219512 142212 219564
rect 203432 219512 203484 219564
rect 204536 219512 204588 219564
rect 211160 219512 211212 219564
rect 105820 219444 105872 219496
rect 63960 219376 64012 219428
rect 64880 219376 64932 219428
rect 72240 219376 72292 219428
rect 73160 219376 73212 219428
rect 80520 219376 80572 219428
rect 90272 219376 90324 219428
rect 90456 219376 90508 219428
rect 106924 219240 106976 219292
rect 117964 219376 118016 219428
rect 123484 219376 123536 219428
rect 126060 219376 126112 219428
rect 126980 219376 127032 219428
rect 130200 219376 130252 219428
rect 134156 219376 134208 219428
rect 134340 219376 134392 219428
rect 135260 219376 135312 219428
rect 135812 219376 135864 219428
rect 139952 219376 140004 219428
rect 140136 219376 140188 219428
rect 145748 219376 145800 219428
rect 146484 219376 146536 219428
rect 197912 219376 197964 219428
rect 199752 219376 199804 219428
rect 203340 219376 203392 219428
rect 208860 219376 208912 219428
rect 209780 219376 209832 219428
rect 148370 219240 148422 219292
rect 149244 219240 149296 219292
rect 150348 219240 150400 219292
rect 152556 219240 152608 219292
rect 153108 219240 153160 219292
rect 153384 219240 153436 219292
rect 162308 219240 162360 219292
rect 162860 219240 162912 219292
rect 163964 219240 164016 219292
rect 164976 219240 165028 219292
rect 165436 219240 165488 219292
rect 165804 219240 165856 219292
rect 166448 219240 166500 219292
rect 85304 219104 85356 219156
rect 117964 219104 118016 219156
rect 123576 219104 123628 219156
rect 128728 219104 128780 219156
rect 131856 219104 131908 219156
rect 132408 219104 132460 219156
rect 70584 218968 70636 219020
rect 132776 218968 132828 219020
rect 133788 218968 133840 219020
rect 134156 219104 134208 219156
rect 135812 218968 135864 219020
rect 135996 218968 136048 219020
rect 136548 218968 136600 219020
rect 136916 219104 136968 219156
rect 146484 219104 146536 219156
rect 146944 219104 146996 219156
rect 152280 219104 152332 219156
rect 168932 219240 168984 219292
rect 169116 219240 169168 219292
rect 167092 219104 167144 219156
rect 185768 219104 185820 219156
rect 193128 219240 193180 219292
rect 195428 219240 195480 219292
rect 196072 219240 196124 219292
rect 199384 219240 199436 219292
rect 225420 219376 225472 219428
rect 226156 219376 226208 219428
rect 228548 219376 228600 219428
rect 232504 219376 232556 219428
rect 233700 219376 233752 219428
rect 234620 219376 234672 219428
rect 234804 219376 234856 219428
rect 279240 219444 279292 219496
rect 405924 219444 405976 219496
rect 412732 219444 412784 219496
rect 285864 219376 285916 219428
rect 301504 219376 301556 219428
rect 325608 219376 325660 219428
rect 326344 219376 326396 219428
rect 343824 219376 343876 219428
rect 347044 219376 347096 219428
rect 352104 219376 352156 219428
rect 366364 219376 366416 219428
rect 374460 219376 374512 219428
rect 375380 219376 375432 219428
rect 380256 219376 380308 219428
rect 384304 219376 384356 219428
rect 399300 219376 399352 219428
rect 400220 219376 400272 219428
rect 403440 219376 403492 219428
rect 404360 219376 404412 219428
rect 415860 219376 415912 219428
rect 416780 219376 416832 219428
rect 417516 219376 417568 219428
rect 421012 219444 421064 219496
rect 432052 219512 432104 219564
rect 515220 219512 515272 219564
rect 515772 219512 515824 219564
rect 667940 219512 667992 219564
rect 669320 219512 669372 219564
rect 428280 219376 428332 219428
rect 488724 219376 488776 219428
rect 489184 219376 489236 219428
rect 518808 219376 518860 219428
rect 519820 219376 519872 219428
rect 567844 219376 567896 219428
rect 568120 219376 568172 219428
rect 617248 219444 617300 219496
rect 504640 219308 504692 219360
rect 505284 219308 505336 219360
rect 195060 219104 195112 219156
rect 195244 219104 195296 219156
rect 226892 219240 226944 219292
rect 229376 219240 229428 219292
rect 235172 219240 235224 219292
rect 237840 219240 237892 219292
rect 239404 219240 239456 219292
rect 246120 219240 246172 219292
rect 286048 219240 286100 219292
rect 327264 219240 327316 219292
rect 152740 218968 152792 219020
rect 200580 218968 200632 219020
rect 201500 218968 201552 219020
rect 203340 219104 203392 219156
rect 246304 219104 246356 219156
rect 258540 219104 258592 219156
rect 259276 219104 259328 219156
rect 259460 219104 259512 219156
rect 291844 219104 291896 219156
rect 294144 219104 294196 219156
rect 311808 219104 311860 219156
rect 315672 219104 315724 219156
rect 317972 219104 318024 219156
rect 320640 219104 320692 219156
rect 340144 219104 340196 219156
rect 383568 219240 383620 219292
rect 387064 219240 387116 219292
rect 419172 219240 419224 219292
rect 422668 219240 422720 219292
rect 450728 219240 450780 219292
rect 453856 219240 453908 219292
rect 479708 219240 479760 219292
rect 480352 219240 480404 219292
rect 507124 219172 507176 219224
rect 516600 219308 516652 219360
rect 535000 219308 535052 219360
rect 543832 219308 543884 219360
rect 544016 219308 544068 219360
rect 553216 219240 553268 219292
rect 345664 219104 345716 219156
rect 204904 218968 204956 219020
rect 206376 218968 206428 219020
rect 255872 218968 255924 219020
rect 259276 218968 259328 219020
rect 293592 218968 293644 219020
rect 301504 218968 301556 219020
rect 306748 218968 306800 219020
rect 62304 218832 62356 218884
rect 76564 218832 76616 218884
rect 83832 218832 83884 218884
rect 148232 218832 148284 218884
rect 148416 218832 148468 218884
rect 148968 218832 149020 218884
rect 149888 218832 149940 218884
rect 152096 218832 152148 218884
rect 152280 218832 152332 218884
rect 166080 218832 166132 218884
rect 166954 218832 167006 218884
rect 215944 218832 215996 218884
rect 217968 218832 218020 218884
rect 220084 218832 220136 218884
rect 77208 218696 77260 218748
rect 142252 218696 142304 218748
rect 59820 218560 59872 218612
rect 69572 218560 69624 218612
rect 92940 218560 92992 218612
rect 93768 218560 93820 218612
rect 145564 218696 145616 218748
rect 145748 218696 145800 218748
rect 146944 218696 146996 218748
rect 93768 218424 93820 218476
rect 142620 218560 142672 218612
rect 143172 218560 143224 218612
rect 145104 218560 145156 218612
rect 146208 218560 146260 218612
rect 146760 218560 146812 218612
rect 152740 218696 152792 218748
rect 152924 218696 152976 218748
rect 156328 218696 156380 218748
rect 156696 218696 156748 218748
rect 107016 218424 107068 218476
rect 157984 218560 158036 218612
rect 159180 218560 159232 218612
rect 160008 218560 160060 218612
rect 160836 218560 160888 218612
rect 161388 218560 161440 218612
rect 162308 218696 162360 218748
rect 213184 218696 213236 218748
rect 213552 218696 213604 218748
rect 217324 218696 217376 218748
rect 218796 218696 218848 218748
rect 219348 218696 219400 218748
rect 219624 218696 219676 218748
rect 220912 218696 220964 218748
rect 228548 218696 228600 218748
rect 229928 218832 229980 218884
rect 264152 218696 264204 218748
rect 167276 218560 167328 218612
rect 169944 218560 169996 218612
rect 177580 218560 177632 218612
rect 185584 218560 185636 218612
rect 195244 218560 195296 218612
rect 195428 218560 195480 218612
rect 243452 218560 243504 218612
rect 252744 218560 252796 218612
rect 259460 218560 259512 218612
rect 274272 218832 274324 218884
rect 280712 218832 280764 218884
rect 281080 218832 281132 218884
rect 312544 218832 312596 218884
rect 265992 218696 266044 218748
rect 267832 218560 267884 218612
rect 272616 218560 272668 218612
rect 296812 218560 296864 218612
rect 300768 218696 300820 218748
rect 329564 218968 329616 219020
rect 333704 218968 333756 219020
rect 352564 219104 352616 219156
rect 354404 219104 354456 219156
rect 355508 219104 355560 219156
rect 358728 219104 358780 219156
rect 364984 219104 365036 219156
rect 483572 219104 483624 219156
rect 490288 219104 490340 219156
rect 502984 219104 503036 219156
rect 503536 219104 503588 219156
rect 524420 219104 524472 219156
rect 533896 219104 533948 219156
rect 538864 219104 538916 219156
rect 544016 219104 544068 219156
rect 568028 219240 568080 219292
rect 351368 218968 351420 219020
rect 355232 218968 355284 219020
rect 355416 218968 355468 219020
rect 369124 218968 369176 219020
rect 373632 218968 373684 219020
rect 380072 218968 380124 219020
rect 384396 218968 384448 219020
rect 393964 218968 394016 219020
rect 401784 218968 401836 219020
rect 407764 218968 407816 219020
rect 502524 218968 502576 219020
rect 507308 218968 507360 219020
rect 515036 218968 515088 219020
rect 542544 218968 542596 219020
rect 543832 218968 543884 219020
rect 553492 219104 553544 219156
rect 558552 219104 558604 219156
rect 558736 219104 558788 219156
rect 563014 219104 563066 219156
rect 572168 219240 572220 219292
rect 572352 219240 572404 219292
rect 573732 219240 573784 219292
rect 574100 219240 574152 219292
rect 577872 219240 577924 219292
rect 568396 219104 568448 219156
rect 572352 219104 572404 219156
rect 314016 218832 314068 218884
rect 329104 218832 329156 218884
rect 337200 218832 337252 218884
rect 357716 218832 357768 218884
rect 366732 218832 366784 218884
rect 378784 218832 378836 218884
rect 386052 218832 386104 218884
rect 396632 218832 396684 218884
rect 402612 218832 402664 218884
rect 409052 218832 409104 218884
rect 411720 218832 411772 218884
rect 412456 218832 412508 218884
rect 510160 218832 510212 218884
rect 514760 218832 514812 218884
rect 524144 218832 524196 218884
rect 524604 218832 524656 218884
rect 525064 218832 525116 218884
rect 529572 218832 529624 218884
rect 534264 218832 534316 218884
rect 545304 218832 545356 218884
rect 547420 218832 547472 218884
rect 548248 218832 548300 218884
rect 562876 218968 562928 219020
rect 563152 218968 563204 219020
rect 563336 218968 563388 219020
rect 566924 218968 566976 219020
rect 567200 218968 567252 219020
rect 570972 218968 571024 219020
rect 571156 218968 571208 219020
rect 576032 219104 576084 219156
rect 592132 219104 592184 219156
rect 599216 219104 599268 219156
rect 302884 218560 302936 218612
rect 307392 218560 307444 218612
rect 337016 218696 337068 218748
rect 340512 218696 340564 218748
rect 360844 218696 360896 218748
rect 379152 218696 379204 218748
rect 392124 218696 392176 218748
rect 395804 218696 395856 218748
rect 404544 218696 404596 218748
rect 412548 218696 412600 218748
rect 417148 218696 417200 218748
rect 429936 218696 429988 218748
rect 432696 218696 432748 218748
rect 460204 218696 460256 218748
rect 461308 218696 461360 218748
rect 482928 218696 482980 218748
rect 485320 218696 485372 218748
rect 519728 218696 519780 218748
rect 530308 218696 530360 218748
rect 534080 218696 534132 218748
rect 534632 218696 534684 218748
rect 537484 218696 537536 218748
rect 548892 218832 548944 218884
rect 553584 218832 553636 218884
rect 567200 218832 567252 218884
rect 576216 218968 576268 219020
rect 469864 218560 469916 218612
rect 471244 218560 471296 218612
rect 475568 218560 475620 218612
rect 482836 218560 482888 218612
rect 518808 218628 518860 218680
rect 148232 218424 148284 218476
rect 149888 218424 149940 218476
rect 150072 218424 150124 218476
rect 157248 218424 157300 218476
rect 157708 218424 157760 218476
rect 160652 218424 160704 218476
rect 161664 218424 161716 218476
rect 162676 218424 162728 218476
rect 163320 218424 163372 218476
rect 166264 218424 166316 218476
rect 167000 218424 167052 218476
rect 213552 218424 213604 218476
rect 216312 218424 216364 218476
rect 220912 218424 220964 218476
rect 221096 218424 221148 218476
rect 224224 218424 224276 218476
rect 224592 218424 224644 218476
rect 225696 218424 225748 218476
rect 226248 218424 226300 218476
rect 229928 218424 229980 218476
rect 239496 218424 239548 218476
rect 272432 218424 272484 218476
rect 279240 218424 279292 218476
rect 281080 218424 281132 218476
rect 291660 218424 291712 218476
rect 324596 218424 324648 218476
rect 501052 218424 501104 218476
rect 529204 218560 529256 218612
rect 557264 218696 557316 218748
rect 562876 218696 562928 218748
rect 563336 218696 563388 218748
rect 573088 218832 573140 218884
rect 575434 218832 575486 218884
rect 575572 218832 575624 218884
rect 567660 218696 567712 218748
rect 568120 218696 568172 218748
rect 572720 218696 572772 218748
rect 572904 218696 572956 218748
rect 575572 218696 575624 218748
rect 575848 218696 575900 218748
rect 582932 218696 582984 218748
rect 514760 218424 514812 218476
rect 538864 218424 538916 218476
rect 542360 218424 542412 218476
rect 543648 218424 543700 218476
rect 545948 218424 546000 218476
rect 571156 218560 571208 218612
rect 571984 218560 572036 218612
rect 572536 218560 572588 218612
rect 591948 218696 592000 218748
rect 592132 218696 592184 218748
rect 675852 218628 675904 218680
rect 677048 218628 677100 218680
rect 548800 218424 548852 218476
rect 567384 218424 567436 218476
rect 567568 218424 567620 218476
rect 596824 218560 596876 218612
rect 75552 218288 75604 218340
rect 83464 218288 83516 218340
rect 100392 218288 100444 218340
rect 105820 218288 105872 218340
rect 113640 218288 113692 218340
rect 56324 218152 56376 218204
rect 62764 218152 62816 218204
rect 79692 218152 79744 218204
rect 82084 218152 82136 218204
rect 120264 218152 120316 218204
rect 55680 218016 55732 218068
rect 56508 218016 56560 218068
rect 57336 218016 57388 218068
rect 57888 218016 57940 218068
rect 58164 218016 58216 218068
rect 61292 218016 61344 218068
rect 65616 218016 65668 218068
rect 66168 218016 66220 218068
rect 73896 218016 73948 218068
rect 74448 218016 74500 218068
rect 74724 218016 74776 218068
rect 75828 218016 75880 218068
rect 78036 218016 78088 218068
rect 78588 218016 78640 218068
rect 78864 218016 78916 218068
rect 79968 218016 80020 218068
rect 82176 218016 82228 218068
rect 82728 218016 82780 218068
rect 84660 218016 84712 218068
rect 85488 218016 85540 218068
rect 86316 218016 86368 218068
rect 86868 218016 86920 218068
rect 87144 218016 87196 218068
rect 88248 218016 88300 218068
rect 88800 218016 88852 218068
rect 89444 218016 89496 218068
rect 94596 218016 94648 218068
rect 95148 218016 95200 218068
rect 97080 218016 97132 218068
rect 98000 218016 98052 218068
rect 98736 218016 98788 218068
rect 99288 218016 99340 218068
rect 99564 218016 99616 218068
rect 100668 218016 100720 218068
rect 101220 218016 101272 218068
rect 102140 218016 102192 218068
rect 102876 218016 102928 218068
rect 103428 218016 103480 218068
rect 103704 218016 103756 218068
rect 104808 218016 104860 218068
rect 105360 218016 105412 218068
rect 106004 218016 106056 218068
rect 109500 218016 109552 218068
rect 110144 218016 110196 218068
rect 110328 218016 110380 218068
rect 110972 218016 111024 218068
rect 111984 218016 112036 218068
rect 112812 218016 112864 218068
rect 115296 218016 115348 218068
rect 115848 218016 115900 218068
rect 116124 218016 116176 218068
rect 117228 218016 117280 218068
rect 119436 218016 119488 218068
rect 119988 218016 120040 218068
rect 121920 218016 121972 218068
rect 122564 218016 122616 218068
rect 127716 218152 127768 218204
rect 128268 218152 128320 218204
rect 128728 218288 128780 218340
rect 174544 218288 174596 218340
rect 159640 218152 159692 218204
rect 166448 218152 166500 218204
rect 166632 218152 166684 218204
rect 167000 218152 167052 218204
rect 168104 218152 168156 218204
rect 171048 218152 171100 218204
rect 171600 218152 171652 218204
rect 176292 218288 176344 218340
rect 175740 218152 175792 218204
rect 176476 218152 176528 218204
rect 160008 218016 160060 218068
rect 166816 218016 166868 218068
rect 167460 218016 167512 218068
rect 168288 218016 168340 218068
rect 169116 218016 169168 218068
rect 169576 218016 169628 218068
rect 173256 218016 173308 218068
rect 174084 218016 174136 218068
rect 175188 218016 175240 218068
rect 176568 218016 176620 218068
rect 177212 218016 177264 218068
rect 185584 218288 185636 218340
rect 185768 218288 185820 218340
rect 192300 218288 192352 218340
rect 193772 218288 193824 218340
rect 229376 218288 229428 218340
rect 229560 218288 229612 218340
rect 231124 218288 231176 218340
rect 232872 218288 232924 218340
rect 234804 218288 234856 218340
rect 365352 218288 365404 218340
rect 373264 218288 373316 218340
rect 426624 218288 426676 218340
rect 429568 218288 429620 218340
rect 434904 218288 434956 218340
rect 436652 218288 436704 218340
rect 500040 218288 500092 218340
rect 507124 218288 507176 218340
rect 507676 218288 507728 218340
rect 529204 218288 529256 218340
rect 529572 218288 529624 218340
rect 571156 218288 571208 218340
rect 179880 218152 179932 218204
rect 221096 218152 221148 218204
rect 221280 218152 221332 218204
rect 221832 218152 221884 218204
rect 222936 218152 222988 218204
rect 223396 218152 223448 218204
rect 223764 218152 223816 218204
rect 224868 218152 224920 218204
rect 227904 218152 227956 218204
rect 229744 218152 229796 218204
rect 235356 218152 235408 218204
rect 235908 218152 235960 218204
rect 236184 218152 236236 218204
rect 236920 218152 236972 218204
rect 177580 218016 177632 218068
rect 181352 218016 181404 218068
rect 182364 218016 182416 218068
rect 183284 218016 183336 218068
rect 184020 218016 184072 218068
rect 184664 218016 184716 218068
rect 185676 218016 185728 218068
rect 186136 218016 186188 218068
rect 186504 218016 186556 218068
rect 189816 218016 189868 218068
rect 190276 218016 190328 218068
rect 193772 218016 193824 218068
rect 193956 218016 194008 218068
rect 194508 218016 194560 218068
rect 194784 218016 194836 218068
rect 195888 218016 195940 218068
rect 196440 218016 196492 218068
rect 197084 218016 197136 218068
rect 198924 218016 198976 218068
rect 200028 218016 200080 218068
rect 202236 218016 202288 218068
rect 202696 218016 202748 218068
rect 203064 218016 203116 218068
rect 203708 218016 203760 218068
rect 204720 218016 204772 218068
rect 206008 218016 206060 218068
rect 210516 218016 210568 218068
rect 210976 218016 211028 218068
rect 213000 218016 213052 218068
rect 215484 218016 215536 218068
rect 216496 218016 216548 218068
rect 249064 218152 249116 218204
rect 249432 218152 249484 218204
rect 251732 218152 251784 218204
rect 269304 218152 269356 218204
rect 273904 218152 273956 218204
rect 299112 218152 299164 218204
rect 300308 218152 300360 218204
rect 304080 218152 304132 218204
rect 305644 218152 305696 218204
rect 310704 218152 310756 218204
rect 315304 218152 315356 218204
rect 330668 218152 330720 218204
rect 333244 218152 333296 218204
rect 348792 218152 348844 218204
rect 351184 218152 351236 218204
rect 364524 218152 364576 218204
rect 367652 218152 367704 218204
rect 369492 218152 369544 218204
rect 370504 218152 370556 218204
rect 376944 218152 376996 218204
rect 382924 218152 382976 218204
rect 386880 218152 386932 218204
rect 388444 218152 388496 218204
rect 394332 218152 394384 218204
rect 402244 218152 402296 218204
rect 407580 218152 407632 218204
rect 411904 218152 411956 218204
rect 422484 218152 422536 218204
rect 425428 218152 425480 218204
rect 425796 218152 425848 218204
rect 428464 218152 428516 218204
rect 433248 218152 433300 218204
rect 435272 218152 435324 218204
rect 455052 218152 455104 218204
rect 460480 218152 460532 218204
rect 461952 218152 462004 218204
rect 466276 218152 466328 218204
rect 494612 218152 494664 218204
rect 495256 218152 495308 218204
rect 519728 218152 519780 218204
rect 519912 218152 519964 218204
rect 524604 218152 524656 218204
rect 527548 218152 527600 218204
rect 572536 218288 572588 218340
rect 572720 218288 572772 218340
rect 574836 218288 574888 218340
rect 575756 218424 575808 218476
rect 576584 218424 576636 218476
rect 607128 218424 607180 218476
rect 604460 218288 604512 218340
rect 571616 218152 571668 218204
rect 581920 218152 581972 218204
rect 582104 218152 582156 218204
rect 582564 218152 582616 218204
rect 582748 218152 582800 218204
rect 592316 218152 592368 218204
rect 676404 218084 676456 218136
rect 677600 218084 677652 218136
rect 244464 218016 244516 218068
rect 247592 218016 247644 218068
rect 247776 218016 247828 218068
rect 248236 218016 248288 218068
rect 248604 218016 248656 218068
rect 249708 218016 249760 218068
rect 250260 218016 250312 218068
rect 251180 218016 251232 218068
rect 251916 218016 251968 218068
rect 252468 218016 252520 218068
rect 262680 218016 262732 218068
rect 263600 218016 263652 218068
rect 264336 218016 264388 218068
rect 264796 218016 264848 218068
rect 265164 218016 265216 218068
rect 266268 218016 266320 218068
rect 266820 218016 266872 218068
rect 267694 218016 267746 218068
rect 268476 218016 268528 218068
rect 269028 218016 269080 218068
rect 270960 218016 271012 218068
rect 271604 218016 271656 218068
rect 276756 218016 276808 218068
rect 277216 218016 277268 218068
rect 277584 218016 277636 218068
rect 278504 218016 278556 218068
rect 281724 218016 281776 218068
rect 282552 218016 282604 218068
rect 285036 218016 285088 218068
rect 285496 218016 285548 218068
rect 287520 218016 287572 218068
rect 288440 218016 288492 218068
rect 289176 218016 289228 218068
rect 289636 218016 289688 218068
rect 293316 218016 293368 218068
rect 293776 218016 293828 218068
rect 295800 218016 295852 218068
rect 296444 218016 296496 218068
rect 297456 218016 297508 218068
rect 298008 218016 298060 218068
rect 298284 218016 298336 218068
rect 299296 218016 299348 218068
rect 301596 218016 301648 218068
rect 302148 218016 302200 218068
rect 302424 218016 302476 218068
rect 303712 218016 303764 218068
rect 305736 218016 305788 218068
rect 306288 218016 306340 218068
rect 306564 218016 306616 218068
rect 307668 218016 307720 218068
rect 308220 218016 308272 218068
rect 308772 218016 308824 218068
rect 312360 218016 312412 218068
rect 314476 218016 314528 218068
rect 314844 218016 314896 218068
rect 315856 218016 315908 218068
rect 316500 218016 316552 218068
rect 317144 218016 317196 218068
rect 318984 218016 319036 218068
rect 319996 218016 320048 218068
rect 322296 218016 322348 218068
rect 322848 218016 322900 218068
rect 324780 218016 324832 218068
rect 325424 218016 325476 218068
rect 326436 218016 326488 218068
rect 326896 218016 326948 218068
rect 328920 218016 328972 218068
rect 330484 218016 330536 218068
rect 333060 218016 333112 218068
rect 333888 218016 333940 218068
rect 334716 218016 334768 218068
rect 335268 218016 335320 218068
rect 335544 218016 335596 218068
rect 336372 218016 336424 218068
rect 339684 218016 339736 218068
rect 340696 218016 340748 218068
rect 342996 218016 343048 218068
rect 343548 218016 343600 218068
rect 347136 218016 347188 218068
rect 347596 218016 347648 218068
rect 347964 218016 348016 218068
rect 349068 218016 349120 218068
rect 349620 218016 349672 218068
rect 350172 218016 350224 218068
rect 353760 218016 353812 218068
rect 354588 218016 354640 218068
rect 356244 218016 356296 218068
rect 357348 218016 357400 218068
rect 357900 218016 357952 218068
rect 359372 218016 359424 218068
rect 363696 218016 363748 218068
rect 364156 218016 364208 218068
rect 366180 218016 366232 218068
rect 366916 218016 366968 218068
rect 368664 218016 368716 218068
rect 369768 218016 369820 218068
rect 370320 218016 370372 218068
rect 370964 218016 371016 218068
rect 371976 218016 372028 218068
rect 372528 218016 372580 218068
rect 372804 218016 372856 218068
rect 373816 218016 373868 218068
rect 376116 218016 376168 218068
rect 376576 218016 376628 218068
rect 378600 218016 378652 218068
rect 379336 218016 379388 218068
rect 381084 218016 381136 218068
rect 381728 218016 381780 218068
rect 385224 218016 385276 218068
rect 386328 218016 386380 218068
rect 388536 218016 388588 218068
rect 389088 218016 389140 218068
rect 389364 218016 389416 218068
rect 390284 218016 390336 218068
rect 392676 218016 392728 218068
rect 393228 218016 393280 218068
rect 393504 218016 393556 218068
rect 394608 218016 394660 218068
rect 395160 218016 395212 218068
rect 395988 218016 396040 218068
rect 396816 218016 396868 218068
rect 397368 218016 397420 218068
rect 400956 218016 401008 218068
rect 401416 218016 401468 218068
rect 409236 218016 409288 218068
rect 409788 218016 409840 218068
rect 410064 218016 410116 218068
rect 411168 218016 411220 218068
rect 413376 218016 413428 218068
rect 413836 218016 413888 218068
rect 418344 218016 418396 218068
rect 419448 218016 419500 218068
rect 420000 218016 420052 218068
rect 420920 218016 420972 218068
rect 424140 218016 424192 218068
rect 426992 218016 427044 218068
rect 427452 218016 427504 218068
rect 427912 218016 427964 218068
rect 429108 218016 429160 218068
rect 430580 218016 430632 218068
rect 432420 218016 432472 218068
rect 433800 218016 433852 218068
rect 435732 218016 435784 218068
rect 436284 218016 436336 218068
rect 436560 218016 436612 218068
rect 437480 218016 437532 218068
rect 438216 218016 438268 218068
rect 438860 218016 438912 218068
rect 439872 218016 439924 218068
rect 440332 218016 440384 218068
rect 453304 218016 453356 218068
rect 455512 218016 455564 218068
rect 456708 218016 456760 218068
rect 457168 218016 457220 218068
rect 463148 218016 463200 218068
rect 464620 218016 464672 218068
rect 467288 218016 467340 218068
rect 467932 218016 467984 218068
rect 470600 218016 470652 218068
rect 472900 218016 472952 218068
rect 488724 218016 488776 218068
rect 497556 218016 497608 218068
rect 505284 218016 505336 218068
rect 505652 218016 505704 218068
rect 613844 218016 613896 218068
rect 505468 217812 505520 217864
rect 514668 217812 514720 217864
rect 528376 217812 528428 217864
rect 602896 217812 602948 217864
rect 603080 217812 603132 217864
rect 612280 217812 612332 217864
rect 514484 217676 514536 217728
rect 519912 217676 519964 217728
rect 533436 217676 533488 217728
rect 542176 217676 542228 217728
rect 542360 217676 542412 217728
rect 551008 217744 551060 217796
rect 551192 217676 551244 217728
rect 603448 217676 603500 217728
rect 604460 217676 604512 217728
rect 615684 217676 615736 217728
rect 523776 217540 523828 217592
rect 524604 217540 524656 217592
rect 533712 217540 533764 217592
rect 534264 217540 534316 217592
rect 538404 217540 538456 217592
rect 542912 217540 542964 217592
rect 543464 217540 543516 217592
rect 543694 217540 543746 217592
rect 543832 217540 543884 217592
rect 557264 217540 557316 217592
rect 557540 217540 557592 217592
rect 572720 217540 572772 217592
rect 575204 217540 575256 217592
rect 576032 217540 576084 217592
rect 593512 217540 593564 217592
rect 596824 217540 596876 217592
rect 623320 217540 623372 217592
rect 524420 217404 524472 217456
rect 541992 217404 542044 217456
rect 542176 217404 542228 217456
rect 549076 217404 549128 217456
rect 549260 217404 549312 217456
rect 551744 217404 551796 217456
rect 553492 217404 553544 217456
rect 564164 217404 564216 217456
rect 564348 217404 564400 217456
rect 571800 217404 571852 217456
rect 571984 217404 572036 217456
rect 572536 217404 572588 217456
rect 572720 217404 572772 217456
rect 573272 217404 573324 217456
rect 609060 217404 609112 217456
rect 436100 217200 436152 217252
rect 437342 217200 437394 217252
rect 447140 217200 447192 217252
rect 448106 217200 448158 217252
rect 448612 217200 448664 217252
rect 449762 217200 449814 217252
rect 469312 217200 469364 217252
rect 470462 217200 470514 217252
rect 530492 217200 530544 217252
rect 530906 217200 530958 217252
rect 542360 217268 542412 217320
rect 535874 217132 535926 217184
rect 548432 217268 548484 217320
rect 550272 217268 550324 217320
rect 551008 217268 551060 217320
rect 557540 217268 557592 217320
rect 558368 217268 558420 217320
rect 562876 217268 562928 217320
rect 563428 217268 563480 217320
rect 570788 217268 570840 217320
rect 571156 217268 571208 217320
rect 547880 217132 547932 217184
rect 520970 217064 521022 217116
rect 546132 217064 546184 217116
rect 549122 217064 549174 217116
rect 549444 217064 549496 217116
rect 550364 217064 550416 217116
rect 550916 217132 550968 217184
rect 551376 217132 551428 217184
rect 551744 217132 551796 217184
rect 571984 217132 572036 217184
rect 572444 217064 572496 217116
rect 573272 217268 573324 217320
rect 604552 217268 604604 217320
rect 607128 217268 607180 217320
rect 616144 217268 616196 217320
rect 573088 217132 573140 217184
rect 574192 217132 574244 217184
rect 575204 217132 575256 217184
rect 604000 217132 604052 217184
rect 582656 216996 582708 217048
rect 590292 216996 590344 217048
rect 591764 216996 591816 217048
rect 592224 216996 592276 217048
rect 592592 216996 592644 217048
rect 614120 216996 614172 217048
rect 582472 216860 582524 216912
rect 590752 216860 590804 216912
rect 593512 216860 593564 216912
rect 605104 216860 605156 216912
rect 605840 216724 605892 216776
rect 574652 216588 574704 216640
rect 582564 216588 582616 216640
rect 591764 216588 591816 216640
rect 595904 216588 595956 216640
rect 576860 216452 576912 216504
rect 582748 216452 582800 216504
rect 592040 216452 592092 216504
rect 596824 216452 596876 216504
rect 582380 216248 582432 216300
rect 592224 216248 592276 216300
rect 590108 216112 590160 216164
rect 597928 216112 597980 216164
rect 590752 215976 590804 216028
rect 596364 215976 596416 216028
rect 599216 215908 599268 215960
rect 613384 215908 613436 215960
rect 652852 215908 652904 215960
rect 654784 215908 654836 215960
rect 590292 215568 590344 215620
rect 598480 215568 598532 215620
rect 613844 215364 613896 215416
rect 615040 215364 615092 215416
rect 636660 215296 636712 215348
rect 639604 215296 639656 215348
rect 575572 215228 575624 215280
rect 621664 215228 621716 215280
rect 574376 215092 574428 215144
rect 619640 215092 619692 215144
rect 675944 215092 675996 215144
rect 677232 215092 677284 215144
rect 577688 214956 577740 215008
rect 626080 214956 626132 215008
rect 576400 214820 576452 214872
rect 622400 214820 622452 214872
rect 574836 214684 574888 214736
rect 616696 214684 616748 214736
rect 616880 214684 616932 214736
rect 617800 214684 617852 214736
rect 624424 214684 624476 214736
rect 633808 214684 633860 214736
rect 577872 214548 577924 214600
rect 575756 214412 575808 214464
rect 620008 214412 620060 214464
rect 626632 214548 626684 214600
rect 627184 214548 627236 214600
rect 628012 214548 628064 214600
rect 628840 214548 628892 214600
rect 630772 214548 630824 214600
rect 631600 214548 631652 214600
rect 628380 214412 628432 214464
rect 600412 214276 600464 214328
rect 600780 214276 600832 214328
rect 607312 214276 607364 214328
rect 607864 214276 607916 214328
rect 608692 214276 608744 214328
rect 609520 214276 609572 214328
rect 616696 214276 616748 214328
rect 624424 214276 624476 214328
rect 658740 214140 658792 214192
rect 661684 214140 661736 214192
rect 662052 214004 662104 214056
rect 665824 214004 665876 214056
rect 35808 213936 35860 213988
rect 40684 213936 40736 213988
rect 675852 213936 675904 213988
rect 676496 213936 676548 213988
rect 626448 213868 626500 213920
rect 629392 213868 629444 213920
rect 638316 213868 638368 213920
rect 640064 213868 640116 213920
rect 648528 213868 648580 213920
rect 650644 213868 650696 213920
rect 655704 213868 655756 213920
rect 656808 213868 656860 213920
rect 660396 213868 660448 213920
rect 660948 213868 661000 213920
rect 651840 213732 651892 213784
rect 658004 213732 658056 213784
rect 660948 213732 661000 213784
rect 662972 213732 663024 213784
rect 663156 213732 663208 213784
rect 664444 213732 664496 213784
rect 576216 213596 576268 213648
rect 601792 213596 601844 213648
rect 645492 213596 645544 213648
rect 659476 213596 659528 213648
rect 574192 213460 574244 213512
rect 601240 213460 601292 213512
rect 639972 213460 640024 213512
rect 642088 213460 642140 213512
rect 650460 213460 650512 213512
rect 575664 213324 575716 213376
rect 612832 213324 612884 213376
rect 635556 213324 635608 213376
rect 652024 213324 652076 213376
rect 666008 213324 666060 213376
rect 575388 213188 575440 213240
rect 623872 213188 623924 213240
rect 641628 213188 641680 213240
rect 658924 213188 658976 213240
rect 654048 212984 654100 213036
rect 654784 212984 654836 213036
rect 664260 212984 664312 213036
rect 665088 212984 665140 213036
rect 632704 212848 632756 212900
rect 634360 212848 634412 212900
rect 628564 212712 628616 212764
rect 632704 212712 632756 212764
rect 637212 212712 637264 212764
rect 641444 212712 641496 212764
rect 578516 211624 578568 211676
rect 580448 211624 580500 211676
rect 35808 211148 35860 211200
rect 41696 211148 41748 211200
rect 579252 209788 579304 209840
rect 581736 209788 581788 209840
rect 581552 208564 581604 208616
rect 632152 209516 632204 209568
rect 652208 209516 652260 209568
rect 666836 209040 666888 209092
rect 35808 208360 35860 208412
rect 40040 208360 40092 208412
rect 578884 208292 578936 208344
rect 589464 208292 589516 208344
rect 580448 207612 580500 207664
rect 589464 207612 589516 207664
rect 581736 206252 581788 206304
rect 589648 206252 589700 206304
rect 579528 205776 579580 205828
rect 581000 205776 581052 205828
rect 579712 204212 579764 204264
rect 589464 204212 589516 204264
rect 35808 202852 35860 202904
rect 37924 202852 37976 202904
rect 578332 202852 578384 202904
rect 580264 202852 580316 202904
rect 581000 202784 581052 202836
rect 589464 202784 589516 202836
rect 578792 200132 578844 200184
rect 590384 200132 590436 200184
rect 580264 199996 580316 200048
rect 589464 199996 589516 200048
rect 669136 199316 669188 199368
rect 670792 199316 670844 199368
rect 579528 198704 579580 198756
rect 589464 198704 589516 198756
rect 578516 195984 578568 196036
rect 589280 195984 589332 196036
rect 579528 194556 579580 194608
rect 589464 194556 589516 194608
rect 669136 194284 669188 194336
rect 670792 194284 670844 194336
rect 579528 191836 579580 191888
rect 589464 191836 589516 191888
rect 579528 190476 579580 190528
rect 590568 190476 590620 190528
rect 667940 189388 667992 189440
rect 670792 189388 670844 189440
rect 579528 187688 579580 187740
rect 589464 187688 589516 187740
rect 579528 186260 579580 186312
rect 589648 186260 589700 186312
rect 579528 184832 579580 184884
rect 589464 184832 589516 184884
rect 579528 182112 579580 182164
rect 589464 182112 589516 182164
rect 578792 180752 578844 180804
rect 590568 180752 590620 180804
rect 578792 178032 578844 178084
rect 589464 178032 589516 178084
rect 579528 177896 579580 177948
rect 589648 177896 589700 177948
rect 579988 175244 580040 175296
rect 589464 175312 589516 175364
rect 667940 174700 667992 174752
rect 669780 174700 669832 174752
rect 578424 174496 578476 174548
rect 589648 174496 589700 174548
rect 578240 172864 578292 172916
rect 579988 172864 580040 172916
rect 580908 172524 580960 172576
rect 589464 172524 589516 172576
rect 579896 171096 579948 171148
rect 589464 171096 589516 171148
rect 578700 169736 578752 169788
rect 580908 169736 580960 169788
rect 582380 169736 582432 169788
rect 589464 169736 589516 169788
rect 668032 169668 668084 169720
rect 670332 169668 670384 169720
rect 579712 168376 579764 168428
rect 589464 168376 589516 168428
rect 583760 167016 583812 167068
rect 589464 167016 589516 167068
rect 578884 165520 578936 165572
rect 582380 165520 582432 165572
rect 667940 164908 667992 164960
rect 670148 164908 670200 164960
rect 582472 164228 582524 164280
rect 589464 164228 589516 164280
rect 580908 162868 580960 162920
rect 589464 162868 589516 162920
rect 676128 162800 676180 162852
rect 678244 162800 678296 162852
rect 578424 162664 578476 162716
rect 582472 162664 582524 162716
rect 675944 162596 675996 162648
rect 679624 162596 679676 162648
rect 578240 162528 578292 162580
rect 583760 162528 583812 162580
rect 675852 161712 675904 161764
rect 681004 161712 681056 161764
rect 580540 161440 580592 161492
rect 589464 161440 589516 161492
rect 580724 160080 580776 160132
rect 589464 160080 589516 160132
rect 578884 158720 578936 158772
rect 580908 158720 580960 158772
rect 587164 158720 587216 158772
rect 589832 158720 589884 158772
rect 585784 157360 585836 157412
rect 589464 157360 589516 157412
rect 578332 154640 578384 154692
rect 580540 154640 580592 154692
rect 584404 154572 584456 154624
rect 589464 154572 589516 154624
rect 583024 153212 583076 153264
rect 589464 153212 589516 153264
rect 578240 152736 578292 152788
rect 580724 152736 580776 152788
rect 580448 151784 580500 151836
rect 589464 151784 589516 151836
rect 578332 151036 578384 151088
rect 587164 151036 587216 151088
rect 578884 149064 578936 149116
rect 589464 149064 589516 149116
rect 578700 147228 578752 147280
rect 585784 147228 585836 147280
rect 668584 145528 668636 145580
rect 670792 145528 670844 145580
rect 585968 144916 586020 144968
rect 589464 144916 589516 144968
rect 579252 144644 579304 144696
rect 584404 144644 584456 144696
rect 584588 143556 584640 143608
rect 589464 143556 589516 143608
rect 579528 143420 579580 143472
rect 583024 143420 583076 143472
rect 587164 142400 587216 142452
rect 589832 142400 589884 142452
rect 583024 140768 583076 140820
rect 589464 140768 589516 140820
rect 578608 140700 578660 140752
rect 580448 140700 580500 140752
rect 580264 139408 580316 139460
rect 589464 139408 589516 139460
rect 578608 139272 578660 139324
rect 589924 139272 589976 139324
rect 578700 137232 578752 137284
rect 588544 137232 588596 137284
rect 579068 137096 579120 137148
rect 585968 137096 586020 137148
rect 585784 136620 585836 136672
rect 589464 136620 589516 136672
rect 667940 136348 667992 136400
rect 669964 136348 670016 136400
rect 584404 135260 584456 135312
rect 589464 135260 589516 135312
rect 675852 133900 675904 133952
rect 676496 133900 676548 133952
rect 580632 131724 580684 131776
rect 590292 131724 590344 131776
rect 578884 131248 578936 131300
rect 589464 131248 589516 131300
rect 579068 131112 579120 131164
rect 584588 131112 584640 131164
rect 579160 128256 579212 128308
rect 587164 128256 587216 128308
rect 587624 127168 587676 127220
rect 589464 127168 589516 127220
rect 579068 126216 579120 126268
rect 587624 126216 587676 126268
rect 667940 125536 667992 125588
rect 669780 125536 669832 125588
rect 579528 125332 579580 125384
rect 583024 125332 583076 125384
rect 583208 124856 583260 124908
rect 589648 124856 589700 124908
rect 578332 124108 578384 124160
rect 580264 124108 580316 124160
rect 580448 122816 580500 122868
rect 589464 122816 589516 122868
rect 581828 122068 581880 122120
rect 590108 122068 590160 122120
rect 587348 121456 587400 121508
rect 589280 121456 589332 121508
rect 579528 121388 579580 121440
rect 585784 121388 585836 121440
rect 584588 118668 584640 118720
rect 589464 118668 589516 118720
rect 578700 118532 578752 118584
rect 584404 118532 584456 118584
rect 668032 118464 668084 118516
rect 670332 118464 670384 118516
rect 585968 117308 586020 117360
rect 589464 117308 589516 117360
rect 675852 117240 675904 117292
rect 682384 117240 682436 117292
rect 578700 117172 578752 117224
rect 580632 117172 580684 117224
rect 585784 115948 585836 116000
rect 589464 115948 589516 116000
rect 579252 114452 579304 114504
rect 581644 114452 581696 114504
rect 668124 114112 668176 114164
rect 669964 114112 670016 114164
rect 584404 113160 584456 113212
rect 589464 113160 589516 113212
rect 579160 113024 579212 113076
rect 588728 113024 588780 113076
rect 581644 111052 581696 111104
rect 589924 111052 589976 111104
rect 583024 109692 583076 109744
rect 589372 109692 589424 109744
rect 578884 108944 578936 108996
rect 581828 108944 581880 108996
rect 578884 107584 578936 107636
rect 589464 107652 589516 107704
rect 581828 106292 581880 106344
rect 589464 106292 589516 106344
rect 668400 106156 668452 106208
rect 670792 106156 670844 106208
rect 580264 104864 580316 104916
rect 589464 104864 589516 104916
rect 578332 103300 578384 103352
rect 583208 103300 583260 103352
rect 578516 102076 578568 102128
rect 580448 102076 580500 102128
rect 587164 100716 587216 100768
rect 589556 100716 589608 100768
rect 624792 100104 624844 100156
rect 668124 100104 668176 100156
rect 580448 99968 580500 100020
rect 590108 99968 590160 100020
rect 614856 99900 614908 99952
rect 667940 99968 667992 100020
rect 622308 99288 622360 99340
rect 630772 99288 630824 99340
rect 579252 99220 579304 99272
rect 581644 99220 581696 99272
rect 623688 99152 623740 99204
rect 633440 99152 633492 99204
rect 577504 99084 577556 99136
rect 595260 99084 595312 99136
rect 625068 99016 625120 99068
rect 636292 99016 636344 99068
rect 629024 98880 629076 98932
rect 643652 98880 643704 98932
rect 629760 98744 629812 98796
rect 645124 98744 645176 98796
rect 630496 98608 630548 98660
rect 646596 98608 646648 98660
rect 578332 97928 578384 97980
rect 587348 97928 587400 97980
rect 605472 97928 605524 97980
rect 606484 97928 606536 97980
rect 618720 97928 618772 97980
rect 625804 97928 625856 97980
rect 628288 97928 628340 97980
rect 642180 98132 642232 98184
rect 627552 97792 627604 97844
rect 640708 97996 640760 98048
rect 634176 97792 634228 97844
rect 650736 97928 650788 97980
rect 655428 97928 655480 97980
rect 662512 97928 662564 97980
rect 647148 97792 647200 97844
rect 659016 97792 659068 97844
rect 659200 97792 659252 97844
rect 663892 97792 663944 97844
rect 621664 97656 621716 97708
rect 629300 97656 629352 97708
rect 631968 97656 632020 97708
rect 648620 97656 648672 97708
rect 653956 97656 654008 97708
rect 655060 97656 655112 97708
rect 659936 97656 659988 97708
rect 665364 97656 665416 97708
rect 626080 97520 626132 97572
rect 637764 97520 637816 97572
rect 639052 97520 639104 97572
rect 613568 97384 613620 97436
rect 618904 97384 618956 97436
rect 620192 97384 620244 97436
rect 625988 97384 626040 97436
rect 631232 97384 631284 97436
rect 639788 97384 639840 97436
rect 643008 97520 643060 97572
rect 659752 97588 659804 97640
rect 658188 97452 658240 97504
rect 663064 97452 663116 97504
rect 647056 97384 647108 97436
rect 651104 97384 651156 97436
rect 654600 97384 654652 97436
rect 656808 97316 656860 97368
rect 661408 97316 661460 97368
rect 623136 97248 623188 97300
rect 632060 97248 632112 97300
rect 632704 97248 632756 97300
rect 650552 97248 650604 97300
rect 651840 97248 651892 97300
rect 654324 97248 654376 97300
rect 626816 97112 626868 97164
rect 639236 97112 639288 97164
rect 644296 97112 644348 97164
rect 658832 97180 658884 97232
rect 659016 97180 659068 97232
rect 661960 97180 662012 97232
rect 612648 97044 612700 97096
rect 621664 97044 621716 97096
rect 624608 96976 624660 97028
rect 635004 96976 635056 97028
rect 635556 96976 635608 97028
rect 639052 96976 639104 97028
rect 639420 96976 639472 97028
rect 647516 96976 647568 97028
rect 650368 96976 650420 97028
rect 658280 97044 658332 97096
rect 596180 96908 596232 96960
rect 596732 96908 596784 96960
rect 615776 96908 615828 96960
rect 616788 96908 616840 96960
rect 654784 96908 654836 96960
rect 655428 96908 655480 96960
rect 660672 96908 660724 96960
rect 663248 96908 663300 96960
rect 612096 96840 612148 96892
rect 612648 96840 612700 96892
rect 617248 96840 617300 96892
rect 618168 96840 618220 96892
rect 633256 96840 633308 96892
rect 606208 96704 606260 96756
rect 612004 96704 612056 96756
rect 634728 96704 634780 96756
rect 639420 96704 639472 96756
rect 639788 96840 639840 96892
rect 647332 96840 647384 96892
rect 654324 96772 654376 96824
rect 659568 96772 659620 96824
rect 650184 96704 650236 96756
rect 638592 96568 638644 96620
rect 639604 96432 639656 96484
rect 642640 96432 642692 96484
rect 645768 96568 645820 96620
rect 652024 96568 652076 96620
rect 652576 96568 652628 96620
rect 664352 96568 664404 96620
rect 652208 96432 652260 96484
rect 653312 96432 653364 96484
rect 665180 96432 665232 96484
rect 640064 96296 640116 96348
rect 647884 96296 647936 96348
rect 648896 96296 648948 96348
rect 664168 96296 664220 96348
rect 637580 96160 637632 96212
rect 660672 96160 660724 96212
rect 610624 96024 610676 96076
rect 623044 96024 623096 96076
rect 641536 96024 641588 96076
rect 663708 96024 663760 96076
rect 577504 95888 577556 95940
rect 601884 95888 601936 95940
rect 607680 95888 607732 95940
rect 622308 95888 622360 95940
rect 645308 95888 645360 95940
rect 649448 95888 649500 95940
rect 649954 95888 650006 95940
rect 664536 95888 664588 95940
rect 642640 95684 642692 95736
rect 651840 95684 651892 95736
rect 641996 95548 642048 95600
rect 646228 95548 646280 95600
rect 646412 95548 646464 95600
rect 640524 95412 640576 95464
rect 643468 95412 643520 95464
rect 649264 95412 649316 95464
rect 620928 95140 620980 95192
rect 626448 95140 626500 95192
rect 647056 95140 647108 95192
rect 648896 95140 648948 95192
rect 653404 95276 653456 95328
rect 649908 95140 649960 95192
rect 579436 95004 579488 95056
rect 584588 95004 584640 95056
rect 649448 94800 649500 94852
rect 656164 94800 656216 94852
rect 609152 94460 609204 94512
rect 620284 94460 620336 94512
rect 648160 93848 648212 93900
rect 654416 93848 654468 93900
rect 619548 93780 619600 93832
rect 626448 93780 626500 93832
rect 579528 93372 579580 93424
rect 585968 93372 586020 93424
rect 611268 93100 611320 93152
rect 619548 93100 619600 93152
rect 647700 92760 647752 92812
rect 655428 92760 655480 92812
rect 607128 92556 607180 92608
rect 610072 92556 610124 92608
rect 617984 92420 618036 92472
rect 626448 92420 626500 92472
rect 652208 92420 652260 92472
rect 655244 92420 655296 92472
rect 579344 91944 579396 91996
rect 585784 91944 585836 91996
rect 579528 91740 579580 91792
rect 588544 91740 588596 91792
rect 616604 91740 616656 91792
rect 626264 91740 626316 91792
rect 618168 90992 618220 91044
rect 626448 90992 626500 91044
rect 622308 89632 622360 89684
rect 626448 89632 626500 89684
rect 581644 88952 581696 89004
rect 600320 88952 600372 89004
rect 649724 88748 649776 88800
rect 658556 88748 658608 88800
rect 662328 88748 662380 88800
rect 663892 88748 663944 88800
rect 610072 88272 610124 88324
rect 626448 88272 626500 88324
rect 655060 88272 655112 88324
rect 658464 88272 658516 88324
rect 619548 88136 619600 88188
rect 626264 88136 626316 88188
rect 578332 86912 578384 86964
rect 580448 86912 580500 86964
rect 659568 86912 659620 86964
rect 663248 86912 663300 86964
rect 652024 86844 652076 86896
rect 657728 86844 657780 86896
rect 649264 86708 649316 86760
rect 661408 86708 661460 86760
rect 647884 86572 647936 86624
rect 660120 86572 660172 86624
rect 656164 86436 656216 86488
rect 660672 86436 660724 86488
rect 623044 86300 623096 86352
rect 626448 86300 626500 86352
rect 654416 86300 654468 86352
rect 662512 86300 662564 86352
rect 653404 86164 653456 86216
rect 657176 86164 657228 86216
rect 609888 85484 609940 85536
rect 626448 85484 626500 85536
rect 578424 85416 578476 85468
rect 581828 85416 581880 85468
rect 620284 85348 620336 85400
rect 625252 85348 625304 85400
rect 608508 84124 608560 84176
rect 625804 84124 625856 84176
rect 579528 83988 579580 84040
rect 583024 83988 583076 84040
rect 579436 82424 579488 82476
rect 584404 82424 584456 82476
rect 628748 81064 628800 81116
rect 642456 81064 642508 81116
rect 618904 80928 618956 80980
rect 649080 80928 649132 80980
rect 614028 80792 614080 80844
rect 646044 80792 646096 80844
rect 595444 80656 595496 80708
rect 636108 80656 636160 80708
rect 585784 79432 585836 79484
rect 589924 79432 589976 79484
rect 629208 79432 629260 79484
rect 645308 79432 645360 79484
rect 579068 79296 579120 79348
rect 598940 79296 598992 79348
rect 615408 79296 615460 79348
rect 646228 79296 646280 79348
rect 631048 78072 631100 78124
rect 643100 78072 643152 78124
rect 621664 77936 621716 77988
rect 648712 77936 648764 77988
rect 578332 77664 578384 77716
rect 580264 77664 580316 77716
rect 584404 77256 584456 77308
rect 631048 77392 631100 77444
rect 628472 77256 628524 77308
rect 632796 77256 632848 77308
rect 616788 76644 616840 76696
rect 646780 76644 646832 76696
rect 606484 76508 606536 76560
rect 662420 76508 662472 76560
rect 588544 75896 588596 75948
rect 628472 75896 628524 75948
rect 612648 75420 612700 75472
rect 646596 75420 646648 75472
rect 612004 75284 612056 75336
rect 646412 75284 646464 75336
rect 578884 75148 578936 75200
rect 666560 75148 666612 75200
rect 579528 73108 579580 73160
rect 587164 73108 587216 73160
rect 579528 71204 579580 71256
rect 585784 71204 585836 71256
rect 585784 68280 585836 68332
rect 601884 68280 601936 68332
rect 579528 66240 579580 66292
rect 623044 66240 623096 66292
rect 579528 64812 579580 64864
rect 614856 64812 614908 64864
rect 578516 62024 578568 62076
rect 613384 62024 613436 62076
rect 580264 58624 580316 58676
rect 600504 58624 600556 58676
rect 579528 57876 579580 57928
rect 624424 57876 624476 57928
rect 576860 57196 576912 57248
rect 603080 57196 603132 57248
rect 579528 56516 579580 56568
rect 588544 56516 588596 56568
rect 574560 56108 574612 56160
rect 596456 56108 596508 56160
rect 574928 55972 574980 56024
rect 596180 55972 596232 56024
rect 574744 55836 574796 55888
rect 599124 55836 599176 55888
rect 462228 53592 462280 53644
rect 581644 55156 581696 55208
rect 459468 53456 459520 53508
rect 579068 55020 579120 55072
rect 584404 54884 584456 54936
rect 589924 54748 589976 54800
rect 597652 54612 597704 54664
rect 597928 54476 597980 54528
rect 583024 54340 583076 54392
rect 580264 54204 580316 54256
rect 574744 54068 574796 54120
rect 574560 53932 574612 53984
rect 462780 53592 462832 53644
rect 463608 53592 463660 53644
rect 464344 53592 464396 53644
rect 472716 53592 472768 53644
rect 473176 53592 473228 53644
rect 476764 53592 476816 53644
rect 477868 53592 477920 53644
rect 481732 53592 481784 53644
rect 482284 53592 482336 53644
rect 485228 53592 485280 53644
rect 463148 53456 463200 53508
rect 472532 53524 472584 53576
rect 477132 53456 477184 53508
rect 482100 53456 482152 53508
rect 482468 53456 482520 53508
rect 574928 53796 574980 53848
rect 50344 53320 50396 53372
rect 130384 53320 130436 53372
rect 460388 53320 460440 53372
rect 462780 53320 462832 53372
rect 465448 53320 465500 53372
rect 477868 53320 477920 53372
rect 47768 53184 47820 53236
rect 130568 53184 130620 53236
rect 463424 53184 463476 53236
rect 476764 53184 476816 53236
rect 312360 53116 312412 53168
rect 313740 53116 313792 53168
rect 316316 53116 316368 53168
rect 317696 53116 317748 53168
rect 46204 53048 46256 53100
rect 129004 53048 129056 53100
rect 464528 53048 464580 53100
rect 473176 53048 473228 53100
rect 464068 52912 464120 52964
rect 477132 52912 477184 52964
rect 464666 52776 464718 52828
rect 485228 52776 485280 52828
rect 460986 52708 461038 52760
rect 463608 52708 463660 52760
rect 465908 52640 465960 52692
rect 472716 52640 472768 52692
rect 145380 52436 145432 52488
rect 306012 52436 306064 52488
rect 49148 51960 49200 52012
rect 126428 51960 126480 52012
rect 48964 51824 49016 51876
rect 129464 51824 129516 51876
rect 46388 51688 46440 51740
rect 130752 51688 130804 51740
rect 126428 50736 126480 50788
rect 129280 50736 129332 50788
rect 50528 50464 50580 50516
rect 128636 50464 128688 50516
rect 318340 50464 318392 50516
rect 458364 50464 458416 50516
rect 45468 50328 45520 50380
rect 129004 50328 129056 50380
rect 314016 50328 314068 50380
rect 458180 50328 458232 50380
rect 51724 49104 51776 49156
rect 128452 49104 128504 49156
rect 47584 48968 47636 49020
rect 129648 48968 129700 49020
rect 128636 48084 128688 48136
rect 132132 48084 132184 48136
rect 129188 47676 129240 47728
rect 131856 47676 131908 47728
rect 623044 46452 623096 46504
rect 661592 46452 661644 46504
rect 129556 45024 129608 45076
rect 129740 44888 129792 44940
rect 128452 44616 128504 44668
rect 129372 44480 129424 44532
rect 131856 44548 131908 44600
rect 132132 44448 132184 44500
rect 132408 44412 132460 44464
rect 130752 44276 130804 44328
rect 129004 44140 129056 44192
rect 132224 44140 132276 44192
rect 130384 44004 130436 44056
rect 130568 43868 130620 43920
rect 43444 42780 43496 42832
rect 187332 43528 187384 43580
rect 431224 43596 431276 43648
rect 310428 42712 310480 42764
rect 364892 42712 364944 42764
rect 431224 42712 431276 42764
rect 456064 42712 456116 42764
rect 463884 42712 463936 42764
rect 427084 42576 427136 42628
rect 455420 42440 455472 42492
rect 462964 42440 463016 42492
rect 404452 42304 404504 42356
rect 405188 42304 405240 42356
rect 420736 42304 420788 42356
rect 426900 42304 426952 42356
rect 663800 42173 663852 42225
rect 427084 42032 427136 42084
rect 431224 42032 431276 42084
rect 456064 42032 456116 42084
rect 455420 41896 455472 41948
rect 404452 41420 404504 41472
rect 420736 41420 420788 41472
rect 426900 41420 426952 41472
rect 459192 41420 459244 41472
<< metal2 >>
rect 110170 1029098 110262 1029126
rect 212934 1029098 213026 1029126
rect 264362 1029098 264454 1029126
rect 315974 1029098 316066 1029126
rect 366390 1029098 366482 1029126
rect 433734 1029098 433826 1029126
rect 510738 1029098 510830 1029126
rect 562166 1029098 562258 1029126
rect 110170 1028622 110262 1028650
rect 212934 1028622 213026 1028650
rect 264362 1028622 264454 1028650
rect 315974 1028622 316066 1028650
rect 366390 1028622 366482 1028650
rect 433734 1028622 433826 1028650
rect 510738 1028622 510830 1028650
rect 562166 1028622 562258 1028650
rect 110170 1028177 110262 1028205
rect 212934 1028177 213026 1028205
rect 264362 1028177 264454 1028205
rect 315974 1028177 316066 1028205
rect 366390 1028177 366482 1028205
rect 433734 1028177 433826 1028205
rect 510738 1028177 510830 1028205
rect 562166 1028177 562258 1028205
rect 366180 1027880 366232 1027886
rect 366180 1027822 366232 1027828
rect 366548 1027880 366600 1027886
rect 366548 1027822 366600 1027828
rect 110170 1027738 110262 1027766
rect 212934 1027738 213026 1027766
rect 264362 1027738 264454 1027766
rect 315974 1027738 316066 1027766
rect 366192 1027752 366220 1027822
rect 366560 1027752 366588 1027822
rect 433734 1027738 433826 1027766
rect 510738 1027738 510830 1027766
rect 562166 1027738 562258 1027766
rect 110170 1027262 110262 1027290
rect 212934 1027262 213026 1027290
rect 264362 1027262 264454 1027290
rect 315974 1027262 316066 1027290
rect 366390 1027262 366482 1027290
rect 433734 1027262 433826 1027290
rect 510738 1027262 510830 1027290
rect 562166 1027262 562258 1027290
rect 110170 1026786 110262 1026814
rect 212934 1026786 213026 1026814
rect 264362 1026786 264454 1026814
rect 315974 1026786 316066 1026814
rect 366390 1026786 366482 1026814
rect 433734 1026786 433826 1026814
rect 510738 1026786 510830 1026814
rect 562166 1026786 562258 1026814
rect 110170 1026310 110262 1026338
rect 212934 1026310 213026 1026338
rect 264362 1026310 264454 1026338
rect 315974 1026310 316066 1026338
rect 366284 1026202 366312 1026324
rect 366468 1026202 366496 1026324
rect 433734 1026310 433826 1026338
rect 510738 1026310 510830 1026338
rect 562166 1026310 562258 1026338
rect 366284 1026174 366496 1026202
rect 366284 1026038 366496 1026066
rect 110170 1025902 110262 1025930
rect 212934 1025902 213026 1025930
rect 264362 1025902 264454 1025930
rect 315974 1025902 316066 1025930
rect 366284 1025916 366312 1026038
rect 366468 1025916 366496 1026038
rect 433734 1025902 433826 1025930
rect 510738 1025902 510830 1025930
rect 562166 1025902 562258 1025930
rect 110170 1025426 110262 1025454
rect 212934 1025426 213026 1025454
rect 264362 1025426 264454 1025454
rect 315974 1025426 316066 1025454
rect 366390 1025426 366482 1025454
rect 433734 1025426 433826 1025454
rect 510738 1025426 510830 1025454
rect 562166 1025426 562258 1025454
rect 110170 1024950 110262 1024978
rect 212934 1024950 213026 1024978
rect 264362 1024950 264454 1024978
rect 315974 1024950 316066 1024978
rect 366390 1024950 366482 1024978
rect 433734 1024950 433826 1024978
rect 510738 1024950 510830 1024978
rect 562166 1024950 562258 1024978
rect 110170 1024474 110262 1024502
rect 212934 1024474 213026 1024502
rect 264362 1024474 264454 1024502
rect 315974 1024474 316066 1024502
rect 366192 1024418 366220 1024488
rect 366560 1024418 366588 1024488
rect 433734 1024474 433826 1024502
rect 510738 1024474 510830 1024502
rect 562166 1024474 562258 1024502
rect 366180 1024412 366232 1024418
rect 366180 1024354 366232 1024360
rect 366548 1024412 366600 1024418
rect 366548 1024354 366600 1024360
rect 110170 1024037 110262 1024065
rect 212934 1024037 213026 1024065
rect 264362 1024037 264454 1024065
rect 315974 1024037 316066 1024065
rect 366390 1024037 366482 1024065
rect 433734 1024037 433826 1024065
rect 510738 1024037 510830 1024065
rect 562166 1024037 562258 1024065
rect 110170 1023590 110262 1023618
rect 212934 1023590 213026 1023618
rect 264362 1023590 264454 1023618
rect 315974 1023590 316066 1023618
rect 366390 1023590 366482 1023618
rect 433734 1023590 433826 1023618
rect 510738 1023590 510830 1023618
rect 562166 1023590 562258 1023618
rect 426346 1007176 426402 1007185
rect 426346 1007111 426348 1007120
rect 426400 1007111 426402 1007120
rect 437480 1007140 437532 1007146
rect 426348 1007082 426400 1007088
rect 437480 1007082 437532 1007088
rect 358542 1007040 358598 1007049
rect 358542 1006975 358544 1006984
rect 358596 1006975 358598 1006984
rect 373264 1007004 373316 1007010
rect 358544 1006946 358596 1006952
rect 373264 1006946 373316 1006952
rect 359370 1006904 359426 1006913
rect 359370 1006839 359372 1006848
rect 359424 1006839 359426 1006848
rect 359372 1006810 359424 1006816
rect 360198 1006768 360254 1006777
rect 144184 1006732 144236 1006738
rect 144184 1006674 144236 1006680
rect 150256 1006732 150308 1006738
rect 150256 1006674 150308 1006680
rect 161940 1006732 161992 1006738
rect 161940 1006674 161992 1006680
rect 164884 1006732 164936 1006738
rect 360198 1006703 360200 1006712
rect 164884 1006674 164936 1006680
rect 360252 1006703 360254 1006712
rect 360200 1006674 360252 1006680
rect 101954 1006632 102010 1006641
rect 94504 1006596 94556 1006602
rect 101954 1006567 101956 1006576
rect 94504 1006538 94556 1006544
rect 102008 1006567 102010 1006576
rect 101956 1006538 102008 1006544
rect 93124 1006460 93176 1006466
rect 93124 1006402 93176 1006408
rect 92480 1006188 92532 1006194
rect 92480 1006130 92532 1006136
rect 92492 1003354 92520 1006130
rect 92308 1003326 92520 1003354
rect 92308 998578 92336 1003326
rect 92296 998572 92348 998578
rect 92296 998514 92348 998520
rect 92848 998572 92900 998578
rect 92848 998514 92900 998520
rect 92296 998436 92348 998442
rect 92296 998378 92348 998384
rect 82266 995752 82322 995761
rect 82018 995710 82266 995738
rect 86498 995752 86554 995761
rect 86342 995710 86498 995738
rect 82266 995687 82322 995696
rect 88982 995752 89038 995761
rect 88734 995710 88982 995738
rect 86498 995687 86554 995696
rect 89626 995752 89682 995761
rect 89378 995710 89626 995738
rect 88982 995687 89038 995696
rect 90270 995752 90326 995761
rect 90022 995710 90270 995738
rect 89626 995687 89682 995696
rect 90270 995687 90326 995696
rect 84658 995480 84714 995489
rect 77036 995081 77064 995452
rect 77022 995072 77078 995081
rect 77022 995007 77078 995016
rect 77680 994702 77708 995452
rect 78338 995438 78628 995466
rect 78600 995058 78628 995438
rect 78600 995030 78720 995058
rect 78692 994809 78720 995030
rect 80164 994838 80192 995452
rect 80152 994832 80204 994838
rect 78678 994800 78734 994809
rect 80152 994774 80204 994780
rect 78678 994735 78734 994744
rect 77668 994696 77720 994702
rect 77668 994638 77720 994644
rect 80716 994430 80744 995452
rect 81360 994566 81388 995452
rect 84502 995438 84658 995466
rect 84658 995415 84714 995424
rect 81348 994560 81400 994566
rect 81348 994502 81400 994508
rect 80704 994424 80756 994430
rect 80704 994366 80756 994372
rect 85040 994265 85068 995452
rect 85698 995438 86080 995466
rect 87538 995438 87920 995466
rect 91218 995438 91692 995466
rect 86052 994537 86080 995438
rect 86038 994528 86094 994537
rect 86038 994463 86094 994472
rect 85026 994256 85082 994265
rect 85026 994191 85082 994200
rect 87892 993993 87920 995438
rect 91664 995330 91692 995438
rect 92308 995330 92336 998378
rect 92664 997824 92716 997830
rect 92664 997766 92716 997772
rect 92480 997688 92532 997694
rect 92480 997630 92532 997636
rect 92492 996985 92520 997630
rect 92478 996976 92534 996985
rect 92478 996911 92534 996920
rect 92676 996033 92704 997766
rect 92662 996024 92718 996033
rect 92662 995959 92718 995968
rect 92664 995852 92716 995858
rect 92664 995794 92716 995800
rect 92480 995580 92532 995586
rect 92480 995522 92532 995528
rect 91664 995302 92336 995330
rect 92492 994537 92520 995522
rect 92478 994528 92534 994537
rect 92478 994463 92534 994472
rect 92676 994265 92704 995794
rect 92860 995489 92888 998514
rect 93136 995761 93164 1006402
rect 93308 999796 93360 999802
rect 93308 999738 93360 999744
rect 93122 995752 93178 995761
rect 93122 995687 93178 995696
rect 92846 995480 92902 995489
rect 92846 995415 92902 995424
rect 92662 994256 92718 994265
rect 92662 994191 92718 994200
rect 93320 993993 93348 999738
rect 94516 994430 94544 1006538
rect 98274 1006496 98330 1006505
rect 98274 1006431 98276 1006440
rect 98328 1006431 98330 1006440
rect 98276 1006402 98328 1006408
rect 103978 1006360 104034 1006369
rect 101404 1006324 101456 1006330
rect 103978 1006295 103980 1006304
rect 101404 1006266 101456 1006272
rect 104032 1006295 104034 1006304
rect 108486 1006360 108542 1006369
rect 108486 1006295 108488 1006304
rect 103980 1006266 104032 1006272
rect 108540 1006295 108542 1006304
rect 126244 1006324 126296 1006330
rect 108488 1006266 108540 1006272
rect 126244 1006266 126296 1006272
rect 99470 1006088 99526 1006097
rect 94688 1006052 94740 1006058
rect 99470 1006023 99472 1006032
rect 94688 1005994 94740 1006000
rect 99524 1006023 99526 1006032
rect 99472 1005994 99524 1006000
rect 94700 997257 94728 1005994
rect 100298 1002688 100354 1002697
rect 97264 1002652 97316 1002658
rect 100298 1002623 100300 1002632
rect 97264 1002594 97316 1002600
rect 100352 1002623 100354 1002632
rect 100300 1002594 100352 1002600
rect 96068 1002108 96120 1002114
rect 96068 1002050 96120 1002056
rect 95884 1001972 95936 1001978
rect 95884 1001914 95936 1001920
rect 94686 997248 94742 997257
rect 94686 997183 94742 997192
rect 94504 994424 94556 994430
rect 94504 994366 94556 994372
rect 87878 993984 87934 993993
rect 87878 993919 87934 993928
rect 93306 993984 93362 993993
rect 93306 993919 93362 993928
rect 50344 993200 50396 993206
rect 50344 993142 50396 993148
rect 44824 993064 44876 993070
rect 44824 993006 44876 993012
rect 43444 975724 43496 975730
rect 43444 975666 43496 975672
rect 42168 969218 42196 969272
rect 42260 969258 42564 969286
rect 42260 969218 42288 969258
rect 42168 969190 42288 969218
rect 42536 969218 42564 969258
rect 42536 969190 42840 969218
rect 42182 968034 42564 968062
rect 41800 967201 41828 967405
rect 41786 967192 41842 967201
rect 41786 967127 41842 967136
rect 42338 966784 42394 966793
rect 42182 966742 42338 966770
rect 42338 966719 42394 966728
rect 42536 966014 42564 968034
rect 42536 965986 42656 966014
rect 42182 965551 42472 965579
rect 42444 964753 42472 965551
rect 42430 964744 42486 964753
rect 42430 964679 42486 964688
rect 42182 964362 42472 964390
rect 42182 963711 42288 963739
rect 42076 962826 42104 963084
rect 42260 962985 42288 963711
rect 42444 963393 42472 964362
rect 42430 963384 42486 963393
rect 42430 963319 42486 963328
rect 42246 962976 42302 962985
rect 42246 962911 42302 962920
rect 42076 962798 42288 962826
rect 41800 962169 41828 962540
rect 41786 962160 41842 962169
rect 41786 962095 41842 962104
rect 42260 962033 42288 962798
rect 42246 962024 42302 962033
rect 42246 961959 42302 961968
rect 41800 959857 41828 960024
rect 41786 959848 41842 959857
rect 41786 959783 41842 959792
rect 41800 959177 41828 959412
rect 41786 959168 41842 959177
rect 41786 959103 41842 959112
rect 42168 958854 42288 958882
rect 42168 958732 42196 958854
rect 42260 958746 42288 958854
rect 42430 958760 42486 958769
rect 42260 958718 42430 958746
rect 42430 958695 42486 958704
rect 41800 957817 41828 958188
rect 41786 957808 41842 957817
rect 41786 957743 41842 957752
rect 42182 956338 42288 956366
rect 41800 955505 41828 955740
rect 41786 955496 41842 955505
rect 41786 955431 41842 955440
rect 41800 954689 41828 955060
rect 41786 954680 41842 954689
rect 41786 954615 41842 954624
rect 41786 954408 41842 954417
rect 41786 954343 41842 954352
rect 35162 952912 35218 952921
rect 35162 952847 35218 952856
rect 33784 951516 33836 951522
rect 33784 951458 33836 951464
rect 31758 946656 31814 946665
rect 31758 946591 31814 946600
rect 31772 945334 31800 946591
rect 28724 945328 28776 945334
rect 28724 945270 28776 945276
rect 31760 945328 31812 945334
rect 31760 945270 31812 945276
rect 8588 944180 8616 944316
rect 9048 944180 9076 944316
rect 9508 944180 9536 944316
rect 9968 944180 9996 944316
rect 10428 944180 10456 944316
rect 10888 944180 10916 944316
rect 11348 944180 11376 944316
rect 11808 944180 11836 944316
rect 12268 944180 12296 944316
rect 12728 944180 12756 944316
rect 13188 944180 13216 944316
rect 13648 944180 13676 944316
rect 14108 944180 14136 944316
rect 28736 942721 28764 945270
rect 28722 942712 28778 942721
rect 28722 942647 28778 942656
rect 33796 938233 33824 951458
rect 33782 938224 33838 938233
rect 33782 938159 33838 938168
rect 35176 937825 35204 952847
rect 41800 952626 41828 954343
rect 41524 952598 41828 952626
rect 37922 952504 37978 952513
rect 37922 952439 37978 952448
rect 36544 952400 36596 952406
rect 36544 952342 36596 952348
rect 35806 943120 35862 943129
rect 35806 943055 35862 943064
rect 35820 942614 35848 943055
rect 35808 942608 35860 942614
rect 35808 942550 35860 942556
rect 35806 941896 35862 941905
rect 35806 941831 35862 941840
rect 35820 941254 35848 941831
rect 35808 941248 35860 941254
rect 35808 941190 35860 941196
rect 35806 940264 35862 940273
rect 35806 940199 35862 940208
rect 35820 939826 35848 940199
rect 35808 939820 35860 939826
rect 35808 939762 35860 939768
rect 36556 939049 36584 952342
rect 36542 939040 36598 939049
rect 36542 938975 36598 938984
rect 37936 938641 37964 952439
rect 39302 952232 39358 952241
rect 39302 952167 39358 952176
rect 37922 938632 37978 938641
rect 37922 938567 37978 938576
rect 35162 937816 35218 937825
rect 35162 937751 35218 937760
rect 39316 937417 39344 952167
rect 40038 951688 40094 951697
rect 40038 951623 40094 951632
rect 39762 943800 39818 943809
rect 39762 943735 39818 943744
rect 39302 937408 39358 937417
rect 39302 937343 39358 937352
rect 39776 935785 39804 943735
rect 39762 935776 39818 935785
rect 39762 935711 39818 935720
rect 40052 934561 40080 951623
rect 41524 951522 41552 952598
rect 42260 952490 42288 956338
rect 41708 952462 42288 952490
rect 41708 952406 41736 952462
rect 41696 952400 41748 952406
rect 41696 952342 41748 952348
rect 41512 951516 41564 951522
rect 41512 951458 41564 951464
rect 42628 949454 42656 965986
rect 42536 949426 42656 949454
rect 41696 942608 41748 942614
rect 41748 942556 41828 942562
rect 41696 942550 41828 942556
rect 41708 942534 41828 942550
rect 41420 941248 41472 941254
rect 41420 941190 41472 941196
rect 40038 934552 40094 934561
rect 40038 934487 40094 934496
rect 41432 911713 41460 941190
rect 41604 939820 41656 939826
rect 41604 939762 41656 939768
rect 41616 911985 41644 939762
rect 41800 935626 41828 942534
rect 42062 940672 42118 940681
rect 42062 940607 42118 940616
rect 42076 939865 42104 940607
rect 42062 939856 42118 939865
rect 42062 939791 42118 939800
rect 42536 939794 42564 949426
rect 42352 939766 42564 939794
rect 41970 935640 42026 935649
rect 41800 935598 41970 935626
rect 41970 935575 42026 935584
rect 42352 932929 42380 939766
rect 42812 937009 42840 969190
rect 43456 966793 43484 975666
rect 43442 966784 43498 966793
rect 43442 966719 43498 966728
rect 43258 964744 43314 964753
rect 43258 964679 43314 964688
rect 42982 963384 43038 963393
rect 42982 963319 43038 963328
rect 42798 937000 42854 937009
rect 42798 936935 42854 936944
rect 42996 933745 43024 963319
rect 43272 935377 43300 964679
rect 43442 962976 43498 962985
rect 43442 962911 43498 962920
rect 43258 935368 43314 935377
rect 43258 935303 43314 935312
rect 43456 934969 43484 962911
rect 44270 962024 44326 962033
rect 44270 961959 44326 961968
rect 43442 934960 43498 934969
rect 43442 934895 43498 934904
rect 44284 934153 44312 961959
rect 44454 958760 44510 958769
rect 44454 958695 44510 958704
rect 44468 936193 44496 958695
rect 44836 941497 44864 993006
rect 47584 991772 47636 991778
rect 47584 991714 47636 991720
rect 46204 961920 46256 961926
rect 46204 961862 46256 961868
rect 46216 946665 46244 961862
rect 46202 946656 46258 946665
rect 46202 946591 46258 946600
rect 45560 946008 45612 946014
rect 45560 945950 45612 945956
rect 45572 943537 45600 945950
rect 45558 943528 45614 943537
rect 45558 943463 45614 943472
rect 44822 941488 44878 941497
rect 44822 941423 44878 941432
rect 44638 941080 44694 941089
rect 44638 941015 44694 941024
rect 44454 936184 44510 936193
rect 44454 936119 44510 936128
rect 44270 934144 44326 934153
rect 44270 934079 44326 934088
rect 42982 933736 43038 933745
rect 42982 933671 43038 933680
rect 43350 933328 43406 933337
rect 43350 933263 43406 933272
rect 42338 932920 42394 932929
rect 42338 932855 42394 932864
rect 41602 911976 41658 911985
rect 41602 911911 41658 911920
rect 41418 911704 41474 911713
rect 41418 911639 41474 911648
rect 43074 892800 43130 892809
rect 43074 892735 43130 892744
rect 42844 892528 42900 892537
rect 42844 892463 42846 892472
rect 42898 892463 42900 892472
rect 42846 892434 42898 892440
rect 43088 892362 43116 892735
rect 43076 892356 43128 892362
rect 43076 892298 43128 892304
rect 42936 892256 42992 892265
rect 42936 892191 42992 892200
rect 41602 885456 41658 885465
rect 41602 885391 41658 885400
rect 41418 885184 41474 885193
rect 41418 885119 41474 885128
rect 8588 818380 8616 818516
rect 9048 818380 9076 818516
rect 9508 818380 9536 818516
rect 9968 818380 9996 818516
rect 10428 818380 10456 818516
rect 10888 818380 10916 818516
rect 11348 818380 11376 818516
rect 11808 818380 11836 818516
rect 12268 818380 12296 818516
rect 12728 818380 12756 818516
rect 13188 818380 13216 818516
rect 13648 818380 13676 818516
rect 14108 818380 14136 818516
rect 35806 817320 35862 817329
rect 35806 817255 35862 817264
rect 35820 817086 35848 817255
rect 35808 817080 35860 817086
rect 35808 817022 35860 817028
rect 35806 816504 35862 816513
rect 35806 816439 35862 816448
rect 35820 815658 35848 816439
rect 41432 815658 41460 885119
rect 41616 823874 41644 885391
rect 42062 884640 42118 884649
rect 42062 884575 42118 884584
rect 42076 823874 42104 884575
rect 41524 823846 41644 823874
rect 41708 823846 42104 823874
rect 41524 815810 41552 823846
rect 41708 817086 41736 823846
rect 41696 817080 41748 817086
rect 41696 817022 41748 817028
rect 41524 815782 41644 815810
rect 35808 815652 35860 815658
rect 35808 815594 35860 815600
rect 41420 815652 41472 815658
rect 41420 815594 41472 815600
rect 35806 814872 35862 814881
rect 35806 814807 35862 814816
rect 35820 814298 35848 814807
rect 41616 814298 41644 815782
rect 35808 814292 35860 814298
rect 35808 814234 35860 814240
rect 41604 814292 41656 814298
rect 41604 814234 41656 814240
rect 41326 812832 41382 812841
rect 41326 812767 41382 812776
rect 40958 812424 41014 812433
rect 40958 812359 41014 812368
rect 35162 811608 35218 811617
rect 35162 811543 35218 811552
rect 35176 802466 35204 811543
rect 35898 811200 35954 811209
rect 35898 811135 35954 811144
rect 35164 802460 35216 802466
rect 35164 802402 35216 802408
rect 35912 802330 35940 811135
rect 40774 808344 40830 808353
rect 40592 808308 40644 808314
rect 40774 808279 40830 808288
rect 40592 808250 40644 808256
rect 40604 805225 40632 808250
rect 40590 805216 40646 805225
rect 40590 805151 40646 805160
rect 40788 805089 40816 808279
rect 40774 805080 40830 805089
rect 40774 805015 40830 805024
rect 40972 804817 41000 812359
rect 41142 812016 41198 812025
rect 41142 811951 41198 811960
rect 40958 804808 41014 804817
rect 40958 804743 41014 804752
rect 41156 804545 41184 811951
rect 41340 811510 41368 812767
rect 41328 811504 41380 811510
rect 41328 811446 41380 811452
rect 41696 811504 41748 811510
rect 41748 811452 42012 811458
rect 41696 811446 42012 811452
rect 41708 811430 42012 811446
rect 41786 808752 41842 808761
rect 41616 808710 41786 808738
rect 41616 808314 41644 808710
rect 41786 808687 41842 808696
rect 41604 808308 41656 808314
rect 41604 808250 41656 808256
rect 41984 804554 42012 811430
rect 43166 810792 43222 810801
rect 43166 810727 43222 810736
rect 42798 809976 42854 809985
rect 42798 809911 42854 809920
rect 42338 806712 42394 806721
rect 42338 806647 42394 806656
rect 41142 804536 41198 804545
rect 41984 804526 42288 804554
rect 41142 804471 41198 804480
rect 41694 802496 41750 802505
rect 41694 802431 41696 802440
rect 41748 802431 41750 802440
rect 41696 802402 41748 802408
rect 35900 802324 35952 802330
rect 35900 802266 35952 802272
rect 41696 802324 41748 802330
rect 41696 802266 41748 802272
rect 41708 802210 41736 802266
rect 41708 802182 41828 802210
rect 41800 800329 41828 802182
rect 41786 800320 41842 800329
rect 41786 800255 41842 800264
rect 41786 799912 41842 799921
rect 41786 799847 41842 799856
rect 41800 799445 41828 799847
rect 42260 798969 42288 804526
rect 42352 801794 42380 806647
rect 42614 802496 42670 802505
rect 42614 802431 42670 802440
rect 42352 801766 42472 801794
rect 42246 798960 42302 798969
rect 42246 798895 42302 798904
rect 42444 798402 42472 801766
rect 42168 798374 42472 798402
rect 42168 798252 42196 798374
rect 42430 798144 42486 798153
rect 42430 798079 42486 798088
rect 42154 797872 42210 797881
rect 42154 797807 42210 797816
rect 42168 797605 42196 797807
rect 42444 797450 42472 798079
rect 42168 797422 42472 797450
rect 42168 796960 42196 797422
rect 42338 797192 42394 797201
rect 42338 797127 42394 797136
rect 42352 796906 42380 797127
rect 42260 796878 42380 796906
rect 42260 795779 42288 796878
rect 42430 796784 42486 796793
rect 42430 796719 42486 796728
rect 42182 795751 42288 795779
rect 42444 795002 42472 796719
rect 42168 794974 42472 795002
rect 42168 794580 42196 794974
rect 42430 794880 42486 794889
rect 42430 794815 42486 794824
rect 41786 794200 41842 794209
rect 41786 794135 41842 794144
rect 41800 793900 41828 794135
rect 42444 793302 42472 794815
rect 42182 793274 42472 793302
rect 42628 792826 42656 802431
rect 42536 792798 42656 792826
rect 42536 792758 42564 792798
rect 42182 792730 42564 792758
rect 42246 792568 42302 792577
rect 42246 792503 42302 792512
rect 42260 790650 42288 792503
rect 42812 792146 42840 809911
rect 42982 807528 43038 807537
rect 42982 807463 43038 807472
rect 42720 792134 42840 792146
rect 42168 790622 42288 790650
rect 42352 792118 42840 792134
rect 42352 792106 42748 792118
rect 42168 790228 42196 790622
rect 42352 789630 42380 792106
rect 42182 789602 42380 789630
rect 42154 789304 42210 789313
rect 42154 789239 42210 789248
rect 42168 788936 42196 789239
rect 42706 789032 42762 789041
rect 42536 788990 42706 789018
rect 41786 788624 41842 788633
rect 41786 788559 41842 788568
rect 41800 788392 41828 788559
rect 42246 788216 42302 788225
rect 42246 788151 42302 788160
rect 41786 786856 41842 786865
rect 41786 786791 41842 786800
rect 41800 786556 41828 786791
rect 42260 786162 42288 788151
rect 42076 786134 42288 786162
rect 42076 785944 42104 786134
rect 42536 785278 42564 788990
rect 42706 788967 42762 788976
rect 42798 788624 42854 788633
rect 42798 788559 42854 788568
rect 42182 785250 42564 785278
rect 42812 782474 42840 788559
rect 42628 782446 42840 782474
rect 42628 779714 42656 782446
rect 41708 779686 42656 779714
rect 8588 775132 8616 775268
rect 9048 775132 9076 775268
rect 9508 775132 9536 775268
rect 9968 775132 9996 775268
rect 10428 775132 10456 775268
rect 10888 775132 10916 775268
rect 11348 775132 11376 775268
rect 11808 775132 11836 775268
rect 12268 775132 12296 775268
rect 12728 775132 12756 775268
rect 13188 775132 13216 775268
rect 13648 775132 13676 775268
rect 14108 775132 14136 775268
rect 35806 773528 35862 773537
rect 35806 773463 35862 773472
rect 35820 772886 35848 773463
rect 41708 772886 41736 779686
rect 35808 772880 35860 772886
rect 35808 772822 35860 772828
rect 41696 772880 41748 772886
rect 41696 772822 41748 772828
rect 35622 769448 35678 769457
rect 35622 769383 35678 769392
rect 35438 769040 35494 769049
rect 35438 768975 35494 768984
rect 35452 768738 35480 768975
rect 35636 768874 35664 769383
rect 35806 769040 35862 769049
rect 35806 768975 35808 768984
rect 35860 768975 35862 768984
rect 41328 769004 41380 769010
rect 35808 768946 35860 768952
rect 41328 768946 41380 768952
rect 35624 768868 35676 768874
rect 35624 768810 35676 768816
rect 35440 768732 35492 768738
rect 35440 768674 35492 768680
rect 40040 768732 40092 768738
rect 40040 768674 40092 768680
rect 31022 768224 31078 768233
rect 31022 768159 31078 768168
rect 31036 758334 31064 768159
rect 35806 767816 35862 767825
rect 35806 767751 35862 767760
rect 35820 767582 35848 767751
rect 35808 767576 35860 767582
rect 35808 767518 35860 767524
rect 37924 767508 37976 767514
rect 37924 767450 37976 767456
rect 35806 767408 35862 767417
rect 35806 767343 35808 767352
rect 35860 767343 35862 767352
rect 36544 767372 36596 767378
rect 35808 767314 35860 767320
rect 36544 767314 36596 767320
rect 35162 767000 35218 767009
rect 35162 766935 35218 766944
rect 35176 759014 35204 766935
rect 35164 759008 35216 759014
rect 35164 758950 35216 758956
rect 31024 758328 31076 758334
rect 31024 758270 31076 758276
rect 36556 757761 36584 767314
rect 37094 763328 37150 763337
rect 37094 763263 37096 763272
rect 37148 763263 37150 763272
rect 37096 763234 37148 763240
rect 37936 759150 37964 767450
rect 40052 764561 40080 768674
rect 41340 765785 41368 768946
rect 41696 768868 41748 768874
rect 41696 768810 41748 768816
rect 41708 765914 41736 768810
rect 41708 765886 42104 765914
rect 41326 765776 41382 765785
rect 41326 765711 41382 765720
rect 40038 764552 40094 764561
rect 40038 764487 40094 764496
rect 39304 763292 39356 763298
rect 39304 763234 39356 763240
rect 37924 759144 37976 759150
rect 39316 759121 39344 763234
rect 40868 759144 40920 759150
rect 37924 759086 37976 759092
rect 39302 759112 39358 759121
rect 40868 759086 40920 759092
rect 39302 759047 39358 759056
rect 40316 759008 40368 759014
rect 40316 758950 40368 758956
rect 36542 757752 36598 757761
rect 36542 757687 36598 757696
rect 40328 757353 40356 758950
rect 40592 758328 40644 758334
rect 40590 758296 40592 758305
rect 40644 758296 40646 758305
rect 40590 758231 40646 758240
rect 40880 757353 40908 759086
rect 42076 758713 42104 765886
rect 42246 765776 42302 765785
rect 42246 765711 42302 765720
rect 42260 763154 42288 765711
rect 42260 763126 42932 763154
rect 42338 759112 42394 759121
rect 42338 759047 42394 759056
rect 42062 758704 42118 758713
rect 42062 758639 42118 758648
rect 42352 758146 42380 759047
rect 42522 758296 42578 758305
rect 42522 758231 42578 758240
rect 42352 758118 42472 758146
rect 40314 757344 40370 757353
rect 40314 757279 40370 757288
rect 40866 757344 40922 757353
rect 40866 757279 40922 757288
rect 41786 756664 41842 756673
rect 41786 756599 41842 756608
rect 41800 756228 41828 756599
rect 42444 755086 42472 758118
rect 42536 757772 42564 758231
rect 42536 757744 42656 757772
rect 42628 757466 42656 757744
rect 42168 755018 42196 755072
rect 42260 755058 42472 755086
rect 42536 757438 42656 757466
rect 42260 755018 42288 755058
rect 42168 754990 42288 755018
rect 42338 754896 42394 754905
rect 42338 754831 42394 754840
rect 42352 754406 42380 754831
rect 42182 754378 42380 754406
rect 42062 754080 42118 754089
rect 42062 754015 42118 754024
rect 42076 753780 42104 754015
rect 42338 753672 42394 753681
rect 42338 753607 42394 753616
rect 42062 752992 42118 753001
rect 42062 752927 42118 752936
rect 42076 752556 42104 752927
rect 42168 751346 42196 751369
rect 42352 751346 42380 753607
rect 42536 753494 42564 757438
rect 42904 754746 42932 763126
rect 42168 751318 42380 751346
rect 42444 753466 42564 753494
rect 42628 754718 42932 754746
rect 41970 751088 42026 751097
rect 41970 751023 42026 751032
rect 41984 750720 42012 751023
rect 42444 750802 42472 753466
rect 42352 750774 42472 750802
rect 41786 750408 41842 750417
rect 41786 750343 41842 750352
rect 41800 750108 41828 750343
rect 42352 749714 42380 750774
rect 42260 749686 42380 749714
rect 42260 749543 42288 749686
rect 42182 749515 42288 749543
rect 41786 747416 41842 747425
rect 41786 747351 41842 747360
rect 41800 747048 41828 747351
rect 42154 746736 42210 746745
rect 42154 746671 42210 746680
rect 42168 746401 42196 746671
rect 42628 746594 42656 754718
rect 42798 754624 42854 754633
rect 42798 754559 42854 754568
rect 42812 753250 42840 754559
rect 42444 746566 42656 746594
rect 42720 753222 42840 753250
rect 42154 746056 42210 746065
rect 42154 745991 42210 746000
rect 42168 745756 42196 745991
rect 42444 745906 42472 746566
rect 42720 746065 42748 753222
rect 42706 746056 42762 746065
rect 42706 745991 42762 746000
rect 42260 745878 42472 745906
rect 42260 745498 42288 745878
rect 42076 745470 42288 745498
rect 42076 745212 42104 745470
rect 42246 745376 42302 745385
rect 42246 745311 42302 745320
rect 42260 744274 42288 745311
rect 42614 744424 42670 744433
rect 42444 744382 42614 744410
rect 42260 744246 42380 744274
rect 41786 743744 41842 743753
rect 41786 743679 41842 743688
rect 41800 743376 41828 743679
rect 42168 742750 42288 742778
rect 42168 742696 42196 742750
rect 42260 742710 42288 742750
rect 42352 742710 42380 744246
rect 42260 742682 42380 742710
rect 42444 742098 42472 744382
rect 42614 744359 42670 744368
rect 42614 743064 42670 743073
rect 42614 742999 42670 743008
rect 42182 742070 42472 742098
rect 42628 741826 42656 742999
rect 42260 741798 42656 741826
rect 8588 731884 8616 732020
rect 9048 731884 9076 732020
rect 9508 731884 9536 732020
rect 9968 731884 9996 732020
rect 10428 731884 10456 732020
rect 10888 731884 10916 732020
rect 11348 731884 11376 732020
rect 11808 731884 11836 732020
rect 12268 731884 12296 732020
rect 12728 731884 12756 732020
rect 13188 731884 13216 732020
rect 13648 731884 13676 732020
rect 14108 731884 14136 732020
rect 42260 731414 42288 741798
rect 42430 741704 42486 741713
rect 42430 741639 42486 741648
rect 42444 731414 42472 741639
rect 41524 731386 42288 731414
rect 42352 731386 42472 731414
rect 35622 731368 35678 731377
rect 35622 731303 35678 731312
rect 35636 730250 35664 731303
rect 35806 730960 35862 730969
rect 35806 730895 35862 730904
rect 35624 730244 35676 730250
rect 35624 730186 35676 730192
rect 35820 730114 35848 730895
rect 41524 730114 41552 731386
rect 42352 730266 42380 731386
rect 41708 730250 42380 730266
rect 41696 730244 42380 730250
rect 41748 730238 42380 730244
rect 41696 730186 41748 730192
rect 35808 730108 35860 730114
rect 35808 730050 35860 730056
rect 41512 730108 41564 730114
rect 41512 730050 41564 730056
rect 41326 726472 41382 726481
rect 41326 726407 41382 726416
rect 41340 726102 41368 726407
rect 41328 726096 41380 726102
rect 41142 726064 41198 726073
rect 41328 726038 41380 726044
rect 41696 726096 41748 726102
rect 41748 726044 42196 726050
rect 41696 726038 42196 726044
rect 41708 726022 42196 726038
rect 41142 725999 41198 726008
rect 31022 725248 31078 725257
rect 31022 725183 31078 725192
rect 31036 716922 31064 725183
rect 36542 724840 36598 724849
rect 36542 724775 36598 724784
rect 33046 724024 33102 724033
rect 33046 723959 33102 723968
rect 31024 716916 31076 716922
rect 31024 716858 31076 716864
rect 33060 715562 33088 723959
rect 33782 723208 33838 723217
rect 33782 723143 33838 723152
rect 33796 715698 33824 723143
rect 33784 715692 33836 715698
rect 33784 715634 33836 715640
rect 33048 715556 33100 715562
rect 33048 715498 33100 715504
rect 36556 715358 36584 724775
rect 40682 724432 40738 724441
rect 40682 724367 40738 724376
rect 40038 720352 40094 720361
rect 40038 720287 40094 720296
rect 39856 715692 39908 715698
rect 39856 715634 39908 715640
rect 36544 715352 36596 715358
rect 36544 715294 36596 715300
rect 39868 715193 39896 715634
rect 39854 715184 39910 715193
rect 39854 715119 39910 715128
rect 40052 714513 40080 720287
rect 40222 715592 40278 715601
rect 40222 715527 40224 715536
rect 40276 715527 40278 715536
rect 40224 715498 40276 715504
rect 40696 714785 40724 724367
rect 41156 721777 41184 725999
rect 41326 725656 41382 725665
rect 41326 725591 41382 725600
rect 41340 724538 41368 725591
rect 41328 724532 41380 724538
rect 41328 724474 41380 724480
rect 41696 724532 41748 724538
rect 41696 724474 41748 724480
rect 41142 721768 41198 721777
rect 41142 721703 41198 721712
rect 41708 719273 41736 724474
rect 41878 722392 41934 722401
rect 41878 722327 41934 722336
rect 41694 719264 41750 719273
rect 41694 719199 41750 719208
rect 41892 718593 41920 722327
rect 41878 718584 41934 718593
rect 41878 718519 41934 718528
rect 42168 718321 42196 726022
rect 42522 719264 42578 719273
rect 42522 719199 42578 719208
rect 42154 718312 42210 718321
rect 42154 718247 42210 718256
rect 41512 716916 41564 716922
rect 41512 716858 41564 716864
rect 40682 714776 40738 714785
rect 40682 714711 40738 714720
rect 40038 714504 40094 714513
rect 40038 714439 40094 714448
rect 41524 714241 41552 716858
rect 41696 715352 41748 715358
rect 41696 715294 41748 715300
rect 41708 715034 41736 715294
rect 42338 715184 42394 715193
rect 42338 715119 42394 715128
rect 41708 715006 41920 715034
rect 41892 714762 41920 715006
rect 42062 714776 42118 714785
rect 41892 714734 42062 714762
rect 42062 714711 42118 714720
rect 42062 714504 42118 714513
rect 42062 714439 42118 714448
rect 41510 714232 41566 714241
rect 42076 714218 42104 714439
rect 42076 714190 42288 714218
rect 41510 714167 41566 714176
rect 41970 713416 42026 713425
rect 41970 713351 42026 713360
rect 41984 713048 42012 713351
rect 42260 712314 42288 714190
rect 42352 713474 42380 715119
rect 42352 713446 42472 713474
rect 42168 712286 42288 712314
rect 42168 711824 42196 712286
rect 42444 711906 42472 713446
rect 42352 711878 42472 711906
rect 42154 711648 42210 711657
rect 42154 711583 42210 711592
rect 42168 711212 42196 711583
rect 42154 710832 42210 710841
rect 42154 710767 42210 710776
rect 42168 710561 42196 710767
rect 42352 709390 42380 711878
rect 42182 709362 42380 709390
rect 42246 709200 42302 709209
rect 42302 709158 42472 709186
rect 42246 709135 42302 709144
rect 42154 708520 42210 708529
rect 42154 708455 42210 708464
rect 42168 708152 42196 708455
rect 42062 707704 42118 707713
rect 42062 707639 42118 707648
rect 42076 707540 42104 707639
rect 41786 707432 41842 707441
rect 41786 707367 41842 707376
rect 41800 706860 41828 707367
rect 42062 706616 42118 706625
rect 42062 706551 42118 706560
rect 42076 706316 42104 706551
rect 42246 705256 42302 705265
rect 42246 705191 42302 705200
rect 42260 704041 42288 705191
rect 42246 704032 42302 704041
rect 42246 703967 42302 703976
rect 42444 703882 42472 709158
rect 42168 703746 42196 703868
rect 42260 703854 42472 703882
rect 42260 703746 42288 703854
rect 42168 703718 42288 703746
rect 42246 703624 42302 703633
rect 42246 703559 42302 703568
rect 42260 703202 42288 703559
rect 42182 703174 42288 703202
rect 42062 703080 42118 703089
rect 42062 703015 42118 703024
rect 42076 702576 42104 703015
rect 42536 702434 42564 719199
rect 42706 715592 42762 715601
rect 42706 715527 42762 715536
rect 42720 712094 42748 715527
rect 42720 712066 42840 712094
rect 42812 703089 42840 712066
rect 42798 703080 42854 703089
rect 42798 703015 42854 703024
rect 42536 702406 42748 702434
rect 42720 702250 42748 702406
rect 42352 702222 42748 702250
rect 42168 701978 42196 702032
rect 42352 701978 42380 702222
rect 42614 702128 42670 702137
rect 42614 702063 42670 702072
rect 42168 701950 42380 701978
rect 42246 701856 42302 701865
rect 42246 701791 42302 701800
rect 42260 700179 42288 701791
rect 42430 701584 42486 701593
rect 42430 701519 42486 701528
rect 42182 700151 42288 700179
rect 42444 699530 42472 701519
rect 42182 699502 42472 699530
rect 42628 698918 42656 702063
rect 42168 698850 42196 698904
rect 42260 698890 42656 698918
rect 42260 698850 42288 698890
rect 42168 698822 42288 698850
rect 41694 697912 41750 697921
rect 41694 697847 41750 697856
rect 35622 691384 35678 691393
rect 35622 691319 35678 691328
rect 8588 688772 8616 688908
rect 9048 688772 9076 688908
rect 9508 688772 9536 688908
rect 9968 688772 9996 688908
rect 10428 688772 10456 688908
rect 10888 688772 10916 688908
rect 11348 688772 11376 688908
rect 11808 688772 11836 688908
rect 12268 688772 12296 688908
rect 12728 688772 12756 688908
rect 13188 688772 13216 688908
rect 13648 688772 13676 688908
rect 14108 688772 14136 688908
rect 35636 687313 35664 691319
rect 35806 687712 35862 687721
rect 35806 687647 35862 687656
rect 35622 687304 35678 687313
rect 35820 687274 35848 687647
rect 41708 687274 41736 697847
rect 35622 687239 35678 687248
rect 35808 687268 35860 687274
rect 35808 687210 35860 687216
rect 41696 687268 41748 687274
rect 41696 687210 41748 687216
rect 35806 683224 35862 683233
rect 35806 683159 35808 683168
rect 35860 683159 35862 683168
rect 41696 683188 41748 683194
rect 35808 683130 35860 683136
rect 41696 683130 41748 683136
rect 35438 682816 35494 682825
rect 35438 682751 35494 682760
rect 35452 681086 35480 682751
rect 35622 682408 35678 682417
rect 35622 682343 35678 682352
rect 35636 681902 35664 682343
rect 35806 682000 35862 682009
rect 41708 681986 41736 683130
rect 41708 681958 42656 681986
rect 35806 681935 35862 681944
rect 35624 681896 35676 681902
rect 35624 681838 35676 681844
rect 35820 681766 35848 681935
rect 41696 681896 41748 681902
rect 41748 681844 42472 681850
rect 41696 681838 42472 681844
rect 41708 681822 42472 681838
rect 35808 681760 35860 681766
rect 35808 681702 35860 681708
rect 41328 681760 41380 681766
rect 41328 681702 41380 681708
rect 35622 681592 35678 681601
rect 35622 681527 35678 681536
rect 35440 681080 35492 681086
rect 35440 681022 35492 681028
rect 35162 680776 35218 680785
rect 35162 680711 35218 680720
rect 35176 672790 35204 680711
rect 35636 680678 35664 681527
rect 35806 681184 35862 681193
rect 35806 681119 35862 681128
rect 35624 680672 35676 680678
rect 35624 680614 35676 680620
rect 35820 680406 35848 681119
rect 36544 680672 36596 680678
rect 36544 680614 36596 680620
rect 35808 680400 35860 680406
rect 35808 680342 35860 680348
rect 35164 672784 35216 672790
rect 35164 672726 35216 672732
rect 36556 672110 36584 680614
rect 37924 680400 37976 680406
rect 37924 680342 37976 680348
rect 36544 672104 36596 672110
rect 36544 672046 36596 672052
rect 37936 670993 37964 680342
rect 41340 678858 41368 681702
rect 41604 681080 41656 681086
rect 41786 681048 41842 681057
rect 41656 681028 41786 681034
rect 41604 681022 41786 681028
rect 41616 681006 41786 681022
rect 41786 680983 41842 680992
rect 42444 678974 42472 681822
rect 42352 678946 42472 678974
rect 42628 678974 42656 681958
rect 42798 679960 42854 679969
rect 42798 679895 42854 679904
rect 42628 678946 42748 678974
rect 41340 678830 41552 678858
rect 39946 677104 40002 677113
rect 39946 677039 40002 677048
rect 38936 672784 38988 672790
rect 38936 672726 38988 672732
rect 38948 672217 38976 672726
rect 39960 672489 39988 677039
rect 39946 672480 40002 672489
rect 39946 672415 40002 672424
rect 38934 672208 38990 672217
rect 38934 672143 38990 672152
rect 39580 672104 39632 672110
rect 39580 672046 39632 672052
rect 39592 671265 39620 672046
rect 41524 671265 41552 678830
rect 42352 674834 42380 678946
rect 42720 676214 42748 678946
rect 42628 676186 42748 676214
rect 42352 674806 42472 674834
rect 42444 672489 42472 674806
rect 42628 674257 42656 676186
rect 42614 674248 42670 674257
rect 42614 674183 42670 674192
rect 42246 672480 42302 672489
rect 42246 672415 42302 672424
rect 42430 672480 42486 672489
rect 42430 672415 42486 672424
rect 39578 671256 39634 671265
rect 39578 671191 39634 671200
rect 41510 671256 41566 671265
rect 41510 671191 41566 671200
rect 37922 670984 37978 670993
rect 37922 670919 37978 670928
rect 41786 670304 41842 670313
rect 41786 670239 41842 670248
rect 41800 669868 41828 670239
rect 42260 668658 42288 672415
rect 42812 672330 42840 679895
rect 42182 668630 42288 668658
rect 42352 672302 42840 672330
rect 41970 668536 42026 668545
rect 41970 668471 42026 668480
rect 41984 668032 42012 668471
rect 41878 667720 41934 667729
rect 41878 667655 41934 667664
rect 41892 667352 41920 667655
rect 42352 666618 42380 672302
rect 42522 672208 42578 672217
rect 42522 672143 42578 672152
rect 42798 672208 42854 672217
rect 42798 672143 42854 672152
rect 42536 671922 42564 672143
rect 42168 666590 42380 666618
rect 42444 671894 42564 671922
rect 42168 666165 42196 666590
rect 42154 665408 42210 665417
rect 42154 665343 42210 665352
rect 42168 665174 42196 665343
rect 42168 665146 42288 665174
rect 42260 664986 42288 665146
rect 42182 664958 42288 664986
rect 42154 664864 42210 664873
rect 42154 664799 42210 664808
rect 42168 664325 42196 664799
rect 41786 664184 41842 664193
rect 41786 664119 41842 664128
rect 41800 663680 41828 664119
rect 42246 664048 42302 664057
rect 42246 663983 42302 663992
rect 42260 663150 42288 663983
rect 42182 663122 42288 663150
rect 42062 662824 42118 662833
rect 42118 662782 42380 662810
rect 42062 662759 42118 662768
rect 42062 661056 42118 661065
rect 42062 660991 42118 661000
rect 42076 660620 42104 660991
rect 42352 660022 42380 662782
rect 42182 659994 42380 660022
rect 42444 659818 42472 671894
rect 42812 667570 42840 672143
rect 42260 659790 42472 659818
rect 42536 667542 42840 667570
rect 42260 659371 42288 659790
rect 42536 659654 42564 667542
rect 42798 667312 42854 667321
rect 42628 667270 42798 667298
rect 42628 664034 42656 667270
rect 42798 667247 42854 667256
rect 42798 664048 42854 664057
rect 42628 664006 42798 664034
rect 42798 663983 42854 663992
rect 42706 663776 42762 663785
rect 42706 663711 42762 663720
rect 42720 661065 42748 663711
rect 42706 661056 42762 661065
rect 42706 660991 42762 661000
rect 42706 660784 42762 660793
rect 42706 660719 42762 660728
rect 42720 659654 42748 660719
rect 42182 659343 42288 659371
rect 42444 659626 42564 659654
rect 42628 659626 42748 659654
rect 42168 658838 42288 658866
rect 42168 658784 42196 658838
rect 42260 658798 42288 658838
rect 42444 658798 42472 659626
rect 42260 658770 42472 658798
rect 42430 658608 42486 658617
rect 42430 658543 42486 658552
rect 42246 658336 42302 658345
rect 42246 658271 42302 658280
rect 42062 657384 42118 657393
rect 42062 657319 42118 657328
rect 42076 656948 42104 657319
rect 42260 656350 42288 658271
rect 42182 656322 42288 656350
rect 42168 655710 42288 655738
rect 42168 655656 42196 655710
rect 42260 655670 42288 655710
rect 42444 655670 42472 658543
rect 42628 657393 42656 659626
rect 42614 657384 42670 657393
rect 42614 657319 42670 657328
rect 42260 655642 42472 655670
rect 35806 646776 35862 646785
rect 35806 646711 35862 646720
rect 8588 645524 8616 645660
rect 9048 645524 9076 645660
rect 9508 645524 9536 645660
rect 9968 645524 9996 645660
rect 10428 645524 10456 645660
rect 10888 645524 10916 645660
rect 11348 645524 11376 645660
rect 11808 645524 11836 645660
rect 12268 645524 12296 645660
rect 12728 645524 12756 645660
rect 13188 645524 13216 645660
rect 13648 645524 13676 645660
rect 14108 645524 14136 645660
rect 35820 644745 35848 646711
rect 35806 644736 35862 644745
rect 35806 644671 35862 644680
rect 41786 641676 41842 641685
rect 41786 641611 41842 641620
rect 41800 641209 41828 641611
rect 41786 641200 41842 641209
rect 41786 641135 41842 641144
rect 35806 639840 35862 639849
rect 35806 639775 35862 639784
rect 35820 639198 35848 639775
rect 35808 639192 35860 639198
rect 35808 639134 35860 639140
rect 41696 639124 41748 639130
rect 41696 639066 41748 639072
rect 35806 639024 35862 639033
rect 41708 639010 41736 639066
rect 35806 638959 35808 638968
rect 35860 638959 35862 638968
rect 40040 638988 40092 638994
rect 35808 638930 35860 638936
rect 41708 638982 42564 639010
rect 40040 638930 40092 638936
rect 35806 638616 35862 638625
rect 35806 638551 35862 638560
rect 32402 638208 32458 638217
rect 32402 638143 32458 638152
rect 32416 629950 32444 638143
rect 35820 637634 35848 638551
rect 35808 637628 35860 637634
rect 35808 637570 35860 637576
rect 40052 637401 40080 638930
rect 41970 638072 42026 638081
rect 41970 638007 42026 638016
rect 41328 637628 41380 637634
rect 41984 637605 42012 638007
rect 41328 637570 41380 637576
rect 41970 637596 42026 637605
rect 40038 637392 40094 637401
rect 40038 637327 40094 637336
rect 41340 634814 41368 637570
rect 41970 637531 42026 637540
rect 41340 634786 41460 634814
rect 32404 629944 32456 629950
rect 32404 629886 32456 629892
rect 41432 627745 41460 634786
rect 42338 633856 42394 633865
rect 42338 633791 42394 633800
rect 41696 629944 41748 629950
rect 41748 629892 42288 629898
rect 41696 629886 42288 629892
rect 41708 629870 42288 629886
rect 41418 627736 41474 627745
rect 41418 627671 41474 627680
rect 42260 627178 42288 629870
rect 42168 627150 42288 627178
rect 42168 626620 42196 627150
rect 42352 625682 42380 633791
rect 42536 626226 42564 638982
rect 42706 627328 42762 627337
rect 42706 627263 42762 627272
rect 42720 626226 42748 627263
rect 42168 625654 42380 625682
rect 42444 626198 42564 626226
rect 42628 626198 42748 626226
rect 42168 625464 42196 625654
rect 42444 625002 42472 626198
rect 42628 626090 42656 626198
rect 42168 624974 42472 625002
rect 42536 626062 42656 626090
rect 42168 624784 42196 624974
rect 42536 624730 42564 626062
rect 42260 624702 42564 624730
rect 42260 624186 42288 624702
rect 42430 624608 42486 624617
rect 42430 624543 42486 624552
rect 42182 624158 42288 624186
rect 42246 623792 42302 623801
rect 42246 623727 42302 623736
rect 42062 623384 42118 623393
rect 42062 623319 42118 623328
rect 42076 622948 42104 623319
rect 42168 621738 42196 621792
rect 42260 621738 42288 623727
rect 42168 621710 42288 621738
rect 42444 621126 42472 624543
rect 42182 621098 42472 621126
rect 42062 620936 42118 620945
rect 42062 620871 42118 620880
rect 42076 620500 42104 620871
rect 42246 620664 42302 620673
rect 42246 620599 42302 620608
rect 41786 620256 41842 620265
rect 41786 620191 41842 620200
rect 41800 619956 41828 620191
rect 42260 617454 42288 620599
rect 42430 620392 42486 620401
rect 42430 620327 42486 620336
rect 42444 619154 42472 620327
rect 42706 619984 42762 619993
rect 42706 619919 42762 619928
rect 42444 619126 42656 619154
rect 42430 619032 42486 619041
rect 42430 618967 42486 618976
rect 42182 617426 42288 617454
rect 42444 616842 42472 618967
rect 42628 618254 42656 619126
rect 42168 616706 42196 616828
rect 42260 616814 42472 616842
rect 42536 618226 42656 618254
rect 42260 616706 42288 616814
rect 42168 616678 42288 616706
rect 42536 616434 42564 618226
rect 42168 616406 42564 616434
rect 42168 616148 42196 616406
rect 42062 615904 42118 615913
rect 42062 615839 42118 615848
rect 42076 615604 42104 615839
rect 42430 615496 42486 615505
rect 42430 615431 42486 615440
rect 42062 615224 42118 615233
rect 42118 615182 42380 615210
rect 42062 615159 42118 615168
rect 41878 614136 41934 614145
rect 41878 614071 41934 614080
rect 41892 613768 41920 614071
rect 42352 613135 42380 615182
rect 42182 613107 42380 613135
rect 42444 612490 42472 615431
rect 42182 612462 42472 612490
rect 42720 611017 42748 619919
rect 42996 612377 43024 807463
rect 43180 788225 43208 810727
rect 43166 788216 43222 788225
rect 43166 788151 43222 788160
rect 43166 766320 43222 766329
rect 43166 766255 43222 766264
rect 43180 753001 43208 766255
rect 43166 752992 43222 753001
rect 43166 752927 43222 752936
rect 43166 723616 43222 723625
rect 43166 723551 43222 723560
rect 43180 705265 43208 723551
rect 43166 705256 43222 705265
rect 43166 705191 43222 705200
rect 43166 679144 43222 679153
rect 43166 679079 43222 679088
rect 43180 663785 43208 679079
rect 43166 663776 43222 663785
rect 43166 663711 43222 663720
rect 43166 636304 43222 636313
rect 43166 636239 43222 636248
rect 43180 624617 43208 636239
rect 43166 624608 43222 624617
rect 43166 624543 43222 624552
rect 43364 613034 43392 933263
rect 43534 932104 43590 932113
rect 43534 932039 43590 932048
rect 43364 613006 43411 613034
rect 43383 612746 43411 613006
rect 43548 612950 43576 932039
rect 44086 891984 44142 891993
rect 44086 891919 44088 891928
rect 44140 891919 44142 891928
rect 44088 891890 44140 891896
rect 44362 816096 44418 816105
rect 44362 816031 44418 816040
rect 44178 814464 44234 814473
rect 44178 814399 44234 814408
rect 43902 809568 43958 809577
rect 43902 809503 43958 809512
rect 43718 806304 43774 806313
rect 43718 806239 43774 806248
rect 43536 612944 43588 612950
rect 43536 612886 43588 612892
rect 43371 612740 43423 612746
rect 43371 612682 43423 612688
rect 43732 612542 43760 806239
rect 43916 797745 43944 809503
rect 43902 797736 43958 797745
rect 43902 797671 43958 797680
rect 44192 773106 44220 814399
rect 44376 773265 44404 816031
rect 44652 815697 44680 941015
rect 47596 891993 47624 991714
rect 48964 990140 49016 990146
rect 48964 990082 49016 990088
rect 48976 940137 49004 990082
rect 48962 940128 49018 940137
rect 48962 940063 49018 940072
rect 50356 939865 50384 993142
rect 54484 992928 54536 992934
rect 54484 992870 54536 992876
rect 51724 991636 51776 991642
rect 51724 991578 51776 991584
rect 51736 942313 51764 991578
rect 53288 990276 53340 990282
rect 53288 990218 53340 990224
rect 51722 942304 51778 942313
rect 51722 942239 51778 942248
rect 50342 939856 50398 939865
rect 50342 939791 50398 939800
rect 53104 923296 53156 923302
rect 53104 923238 53156 923244
rect 50344 909492 50396 909498
rect 50344 909434 50396 909440
rect 47768 897048 47820 897054
rect 47768 896990 47820 896996
rect 47582 891984 47638 891993
rect 47582 891919 47638 891928
rect 46204 870868 46256 870874
rect 46204 870810 46256 870816
rect 44638 815688 44694 815697
rect 44638 815623 44694 815632
rect 44822 815280 44878 815289
rect 44822 815215 44878 815224
rect 44546 810384 44602 810393
rect 44546 810319 44602 810328
rect 44560 789313 44588 810319
rect 44546 789304 44602 789313
rect 44546 789239 44602 789248
rect 44362 773256 44418 773265
rect 44362 773191 44418 773200
rect 44192 773078 44404 773106
rect 44178 772032 44234 772041
rect 44178 771967 44234 771976
rect 44192 729337 44220 771967
rect 44376 771633 44404 773078
rect 44638 772848 44694 772857
rect 44638 772783 44694 772792
rect 44362 771624 44418 771633
rect 44362 771559 44418 771568
rect 44362 771216 44418 771225
rect 44362 771151 44418 771160
rect 44178 729328 44234 729337
rect 44178 729263 44234 729272
rect 44376 728521 44404 771151
rect 44652 730153 44680 772783
rect 44836 772449 44864 815215
rect 45006 813648 45062 813657
rect 45006 813583 45062 813592
rect 44822 772440 44878 772449
rect 44822 772375 44878 772384
rect 45020 770817 45048 813583
rect 45190 807936 45246 807945
rect 45190 807871 45246 807880
rect 45204 796793 45232 807871
rect 45190 796784 45246 796793
rect 45190 796719 45246 796728
rect 45006 770808 45062 770817
rect 45006 770743 45062 770752
rect 45098 770400 45154 770409
rect 45098 770335 45154 770344
rect 44822 766728 44878 766737
rect 44822 766663 44878 766672
rect 44836 746745 44864 766663
rect 44822 746736 44878 746745
rect 44822 746671 44878 746680
rect 44638 730144 44694 730153
rect 44638 730079 44694 730088
rect 44546 729736 44602 729745
rect 44546 729671 44602 729680
rect 44362 728512 44418 728521
rect 44362 728447 44418 728456
rect 44270 727288 44326 727297
rect 44270 727223 44326 727232
rect 43902 721576 43958 721585
rect 43902 721511 43958 721520
rect 43916 708529 43944 721511
rect 43902 708520 43958 708529
rect 43902 708455 43958 708464
rect 44284 684457 44312 727223
rect 44560 686905 44588 729671
rect 44914 728920 44970 728929
rect 44914 728855 44970 728864
rect 44730 721168 44786 721177
rect 44730 721103 44786 721112
rect 44546 686896 44602 686905
rect 44546 686831 44602 686840
rect 44546 686488 44602 686497
rect 44546 686423 44602 686432
rect 44560 685098 44588 686423
rect 44548 685092 44600 685098
rect 44548 685034 44600 685040
rect 44270 684448 44326 684457
rect 44270 684383 44326 684392
rect 44362 684040 44418 684049
rect 44362 683975 44418 683984
rect 44178 680368 44234 680377
rect 44178 680303 44234 680312
rect 44192 662833 44220 680303
rect 44178 662824 44234 662833
rect 44178 662759 44234 662768
rect 44376 641481 44404 683975
rect 44744 669314 44772 721103
rect 44928 686089 44956 728855
rect 45112 727705 45140 770335
rect 45282 764824 45338 764833
rect 45282 764759 45338 764768
rect 45296 753681 45324 764759
rect 45558 764280 45614 764289
rect 45558 764215 45614 764224
rect 45282 753672 45338 753681
rect 45282 753607 45338 753616
rect 45282 728104 45338 728113
rect 45282 728039 45338 728048
rect 45098 727696 45154 727705
rect 45098 727631 45154 727640
rect 45098 722800 45154 722809
rect 45098 722735 45154 722744
rect 45112 707713 45140 722735
rect 45098 707704 45154 707713
rect 45098 707639 45154 707648
rect 45296 692774 45324 728039
rect 45296 692746 45416 692774
rect 44914 686080 44970 686089
rect 44914 686015 44970 686024
rect 45098 685672 45154 685681
rect 45098 685607 45154 685616
rect 44914 684856 44970 684865
rect 44914 684791 44970 684800
rect 44928 683114 44956 684791
rect 45112 683114 45140 685607
rect 45388 685386 45416 692746
rect 45296 685358 45416 685386
rect 45296 685273 45324 685358
rect 45282 685264 45338 685273
rect 45282 685199 45338 685208
rect 45376 685092 45428 685098
rect 45376 685034 45428 685040
rect 44836 683086 44956 683114
rect 45020 683086 45140 683114
rect 44836 678974 44864 683086
rect 45020 678974 45048 683086
rect 45190 679552 45246 679561
rect 45190 679487 45246 679496
rect 44836 678946 44956 678974
rect 45020 678946 45140 678974
rect 44928 669314 44956 678946
rect 45112 669314 45140 678946
rect 44652 669286 44772 669314
rect 44836 669286 44956 669314
rect 45020 669286 45140 669314
rect 44652 659654 44680 669286
rect 44836 659654 44864 669286
rect 45020 659654 45048 669286
rect 45204 664873 45232 679487
rect 45190 664864 45246 664873
rect 45190 664799 45246 664808
rect 44652 659626 44772 659654
rect 44836 659626 44956 659654
rect 45020 659626 45140 659654
rect 44744 653177 44772 659626
rect 44730 653168 44786 653177
rect 44730 653103 44786 653112
rect 44546 643376 44602 643385
rect 44546 643311 44602 643320
rect 44362 641472 44418 641481
rect 44362 641407 44418 641416
rect 44178 636576 44234 636585
rect 44234 636534 44404 636562
rect 44178 636511 44234 636520
rect 44376 635610 44404 636534
rect 44284 635582 44404 635610
rect 43902 635352 43958 635361
rect 43902 635287 43958 635296
rect 43916 620945 43944 635287
rect 44088 626136 44140 626142
rect 44088 626078 44140 626084
rect 43902 620936 43958 620945
rect 43902 620871 43958 620880
rect 44100 620673 44128 626078
rect 44284 623393 44312 635582
rect 44560 627914 44588 643311
rect 44730 642560 44786 642569
rect 44730 642495 44786 642504
rect 44468 627886 44588 627914
rect 44270 623384 44326 623393
rect 44270 623319 44326 623328
rect 44086 620664 44142 620673
rect 44086 620599 44142 620608
rect 44468 618254 44496 627886
rect 44744 623098 44772 642495
rect 44928 642297 44956 659626
rect 45112 643113 45140 659626
rect 45388 643657 45416 685034
rect 45374 643648 45430 643657
rect 45374 643583 45430 643592
rect 45098 643104 45154 643113
rect 45098 643039 45154 643048
rect 44914 642288 44970 642297
rect 44914 642223 44970 642232
rect 45282 641200 45338 641209
rect 45282 641135 45338 641144
rect 44914 640928 44970 640937
rect 44914 640863 44970 640872
rect 44928 636002 44956 640863
rect 44916 635996 44968 636002
rect 44916 635938 44968 635944
rect 44914 635760 44970 635769
rect 44914 635695 44970 635704
rect 45100 635724 45152 635730
rect 44928 626142 44956 635695
rect 45100 635666 45152 635672
rect 44916 626136 44968 626142
rect 44916 626078 44968 626084
rect 44744 623070 44956 623098
rect 44928 618254 44956 623070
rect 45112 618254 45140 635666
rect 45296 635474 45324 641135
rect 44468 618226 44680 618254
rect 44178 614136 44234 614145
rect 44178 614071 44234 614080
rect 43720 612536 43772 612542
rect 43720 612478 43772 612484
rect 42982 612368 43038 612377
rect 42982 612303 43038 612312
rect 43580 612368 43636 612377
rect 43580 612303 43582 612312
rect 43634 612303 43636 612312
rect 43582 612274 43634 612280
rect 44192 611590 44220 614071
rect 44180 611584 44232 611590
rect 44180 611526 44232 611532
rect 42706 611008 42762 611017
rect 42706 610943 42762 610952
rect 44270 611008 44326 611017
rect 44270 610943 44326 610952
rect 44284 610586 44312 610943
rect 44502 610632 44554 610638
rect 44284 610580 44502 610586
rect 44284 610574 44554 610580
rect 44284 610558 44542 610574
rect 44652 605834 44680 618226
rect 44560 605806 44680 605834
rect 44836 618226 44956 618254
rect 45020 618226 45140 618254
rect 45204 635446 45324 635474
rect 8588 602276 8616 602412
rect 9048 602276 9076 602412
rect 9508 602276 9536 602412
rect 9968 602276 9996 602412
rect 10428 602276 10456 602412
rect 10888 602276 10916 602412
rect 11348 602276 11376 602412
rect 11808 602276 11836 602412
rect 12268 602276 12296 602412
rect 12728 602276 12756 602412
rect 13188 602276 13216 602412
rect 13648 602276 13676 602412
rect 14108 602276 14136 602412
rect 44560 600545 44588 605806
rect 44546 600536 44602 600545
rect 44546 600471 44602 600480
rect 44638 600128 44694 600137
rect 44638 600063 44694 600072
rect 40314 597272 40370 597281
rect 40314 597207 40370 597216
rect 40328 596222 40356 597207
rect 42982 597000 43038 597009
rect 42982 596935 43038 596944
rect 42614 596864 42670 596873
rect 42614 596799 42670 596808
rect 40316 596216 40368 596222
rect 40316 596158 40368 596164
rect 40866 596218 40922 596227
rect 40866 596153 40922 596162
rect 41142 596218 41198 596227
rect 41142 596153 41198 596162
rect 41696 596216 41748 596222
rect 41748 596164 41828 596174
rect 41696 596158 41828 596164
rect 40880 596086 40908 596153
rect 40868 596080 40920 596086
rect 40868 596022 40920 596028
rect 32402 595640 32458 595649
rect 32402 595575 32458 595584
rect 32416 585818 32444 595575
rect 36542 595232 36598 595241
rect 36542 595167 36598 595176
rect 35162 594416 35218 594425
rect 35162 594351 35218 594360
rect 35176 585954 35204 594351
rect 35164 585948 35216 585954
rect 35164 585890 35216 585896
rect 32404 585812 32456 585818
rect 32404 585754 32456 585760
rect 36556 585206 36584 595167
rect 37922 594824 37978 594833
rect 37922 594759 37978 594768
rect 36544 585200 36596 585206
rect 37936 585177 37964 594759
rect 41156 594674 41184 596153
rect 41708 596146 41828 596158
rect 41328 596080 41380 596086
rect 41800 596057 41828 596146
rect 41328 596022 41380 596028
rect 41786 596048 41842 596057
rect 41340 594946 41368 596022
rect 41786 595983 41842 595992
rect 41694 594960 41750 594969
rect 41340 594918 41694 594946
rect 41694 594895 41750 594904
rect 41156 594646 41460 594674
rect 40684 593292 40736 593298
rect 40684 593234 40736 593240
rect 39946 590744 40002 590753
rect 39946 590679 40002 590688
rect 39960 585993 39988 590679
rect 39946 585984 40002 585993
rect 39946 585919 40002 585928
rect 40500 585948 40552 585954
rect 40500 585890 40552 585896
rect 39488 585812 39540 585818
rect 39488 585754 39540 585760
rect 36544 585142 36596 585148
rect 37922 585168 37978 585177
rect 37922 585103 37978 585112
rect 39500 584905 39528 585754
rect 40512 585721 40540 585890
rect 40498 585712 40554 585721
rect 40498 585647 40554 585656
rect 39486 584896 39542 584905
rect 39486 584831 39542 584840
rect 40696 584633 40724 593234
rect 40960 593088 41012 593094
rect 40960 593030 41012 593036
rect 40972 589665 41000 593030
rect 40958 589656 41014 589665
rect 40958 589591 41014 589600
rect 41432 585449 41460 594646
rect 41786 593600 41842 593609
rect 41616 593558 41786 593586
rect 41616 593298 41644 593558
rect 41786 593535 41842 593544
rect 42628 593314 42656 596799
rect 42798 594008 42854 594017
rect 42798 593943 42854 593952
rect 41604 593292 41656 593298
rect 42628 593286 42748 593314
rect 41604 593234 41656 593240
rect 41786 593192 41842 593201
rect 41616 593150 41786 593178
rect 41616 593094 41644 593150
rect 41786 593127 41842 593136
rect 41604 593088 41656 593094
rect 41604 593030 41656 593036
rect 41786 592784 41842 592793
rect 41786 592719 41842 592728
rect 41800 589393 41828 592719
rect 41786 589384 41842 589393
rect 41786 589319 41842 589328
rect 42720 586129 42748 593286
rect 42812 589274 42840 593943
rect 42812 589246 42932 589274
rect 42706 586120 42762 586129
rect 42706 586055 42762 586064
rect 42246 585984 42302 585993
rect 42246 585919 42302 585928
rect 41418 585440 41474 585449
rect 41418 585375 41474 585384
rect 42260 585290 42288 585919
rect 42614 585712 42670 585721
rect 42670 585670 42840 585698
rect 42614 585647 42670 585656
rect 42430 585440 42486 585449
rect 42430 585375 42486 585384
rect 42260 585262 42380 585290
rect 41420 585200 41472 585206
rect 41420 585142 41472 585148
rect 40682 584624 40738 584633
rect 40682 584559 40738 584568
rect 41432 584474 41460 585142
rect 41432 584446 42288 584474
rect 42260 583454 42288 584446
rect 42182 583426 42288 583454
rect 42352 582263 42380 585262
rect 42444 582298 42472 585375
rect 42444 582270 42656 582298
rect 42182 582235 42380 582263
rect 42338 581904 42394 581913
rect 42338 581839 42394 581848
rect 42352 581618 42380 581839
rect 42182 581590 42380 581618
rect 42246 581496 42302 581505
rect 42302 581454 42472 581482
rect 42246 581431 42302 581440
rect 42062 581224 42118 581233
rect 42062 581159 42118 581168
rect 42076 580961 42104 581159
rect 42246 580816 42302 580825
rect 42246 580751 42302 580760
rect 41786 580272 41842 580281
rect 41786 580207 41842 580216
rect 41800 579768 41828 580207
rect 42260 578626 42288 580751
rect 42168 578598 42288 578626
rect 42168 578544 42196 578598
rect 41786 578232 41842 578241
rect 41786 578167 41842 578176
rect 41800 577932 41828 578167
rect 41786 577552 41842 577561
rect 41786 577487 41842 577496
rect 41800 577281 41828 577487
rect 42444 577266 42472 581454
rect 42628 579614 42656 582270
rect 42812 579614 42840 585670
rect 42260 577238 42472 577266
rect 42536 579586 42656 579614
rect 42720 579586 42840 579614
rect 42260 576994 42288 577238
rect 42076 576966 42288 576994
rect 42076 576708 42104 576966
rect 42246 576872 42302 576881
rect 42246 576807 42302 576816
rect 42260 574274 42288 576807
rect 42536 576201 42564 579586
rect 42522 576192 42578 576201
rect 42522 576127 42578 576136
rect 42182 574246 42288 574274
rect 42720 573866 42748 579586
rect 42628 573838 42748 573866
rect 42076 573345 42104 573580
rect 42628 573458 42656 573838
rect 42536 573430 42656 573458
rect 42062 573336 42118 573345
rect 42062 573271 42118 573280
rect 42536 572982 42564 573430
rect 42706 573336 42762 573345
rect 42904 573322 42932 589246
rect 42762 573294 42932 573322
rect 42706 573271 42762 573280
rect 42182 572954 42564 572982
rect 41970 572656 42026 572665
rect 41970 572591 42026 572600
rect 41984 572424 42012 572591
rect 42246 572248 42302 572257
rect 42246 572183 42302 572192
rect 42062 571024 42118 571033
rect 42062 570959 42118 570968
rect 42076 570588 42104 570959
rect 42260 569922 42288 572183
rect 42614 571976 42670 571985
rect 42614 571911 42670 571920
rect 42182 569894 42288 569922
rect 42628 569514 42656 571911
rect 42076 569486 42656 569514
rect 42076 569296 42104 569486
rect 42338 569256 42394 569265
rect 42338 569191 42394 569200
rect 42352 567194 42380 569191
rect 41524 567166 42380 567194
rect 8588 559164 8616 559300
rect 9048 559164 9076 559300
rect 9508 559164 9536 559300
rect 9968 559164 9996 559300
rect 10428 559164 10456 559300
rect 10888 559164 10916 559300
rect 11348 559164 11376 559300
rect 11808 559164 11836 559300
rect 12268 559164 12296 559300
rect 12728 559164 12756 559300
rect 13188 559164 13216 559300
rect 13648 559164 13676 559300
rect 14108 559164 14136 559300
rect 35806 558104 35862 558113
rect 35806 558039 35862 558048
rect 35820 557598 35848 558039
rect 41524 557598 41552 567166
rect 42062 558512 42118 558521
rect 42062 558447 42118 558456
rect 35808 557592 35860 557598
rect 35808 557534 35860 557540
rect 41512 557592 41564 557598
rect 42076 557569 42104 558447
rect 41512 557534 41564 557540
rect 42062 557560 42118 557569
rect 42996 557534 43024 596935
rect 44454 591968 44510 591977
rect 44454 591903 44510 591912
rect 43442 590336 43498 590345
rect 43442 590271 43498 590280
rect 42062 557495 42118 557504
rect 42812 557506 43024 557534
rect 35806 554840 35862 554849
rect 42812 554826 42840 557506
rect 41708 554810 42840 554826
rect 35806 554775 35808 554784
rect 35860 554775 35862 554784
rect 41696 554804 42840 554810
rect 35808 554746 35860 554752
rect 41748 554798 42840 554804
rect 41696 554746 41748 554752
rect 35622 554024 35678 554033
rect 35622 553959 35678 553968
rect 35636 553450 35664 553959
rect 35806 553616 35862 553625
rect 35806 553551 35808 553560
rect 35860 553551 35862 553560
rect 41420 553580 41472 553586
rect 35808 553522 35860 553528
rect 41420 553522 41472 553528
rect 35624 553444 35676 553450
rect 35624 553386 35676 553392
rect 41432 553394 41460 553522
rect 41696 553444 41748 553450
rect 41432 553366 41552 553394
rect 41748 553392 41828 553394
rect 41696 553386 41828 553392
rect 41708 553366 41828 553386
rect 40866 553208 40922 553217
rect 40866 553143 40922 553152
rect 33782 551984 33838 551993
rect 33782 551919 33838 551928
rect 31758 547496 31814 547505
rect 31758 547431 31760 547440
rect 31812 547431 31814 547440
rect 31760 547402 31812 547408
rect 33796 543046 33824 551919
rect 40880 549794 40908 553143
rect 41050 552800 41106 552809
rect 41050 552735 41106 552744
rect 41064 552158 41092 552735
rect 41052 552152 41104 552158
rect 41052 552094 41104 552100
rect 41234 551168 41290 551177
rect 41234 551103 41290 551112
rect 41248 550662 41276 551103
rect 41236 550656 41288 550662
rect 41236 550598 41288 550604
rect 40880 549766 41184 549794
rect 41156 547754 41184 549766
rect 41326 548312 41382 548321
rect 41326 548247 41382 548256
rect 41340 547942 41368 548247
rect 41328 547936 41380 547942
rect 41328 547878 41380 547884
rect 41156 547726 41368 547754
rect 37096 547460 37148 547466
rect 37096 547402 37148 547408
rect 33784 543040 33836 543046
rect 33784 542982 33836 542988
rect 37108 542366 37136 547402
rect 41340 546417 41368 547726
rect 41326 546408 41382 546417
rect 41326 546343 41382 546352
rect 41524 543734 41552 553366
rect 41800 553217 41828 553366
rect 41786 553208 41842 553217
rect 41786 553143 41842 553152
rect 42982 552392 43038 552401
rect 42982 552327 43038 552336
rect 41708 552090 41920 552106
rect 41696 552084 41920 552090
rect 41748 552078 41920 552084
rect 41696 552026 41748 552032
rect 41892 551993 41920 552078
rect 41878 551984 41934 551993
rect 41878 551919 41934 551928
rect 41696 550656 41748 550662
rect 41748 550616 42840 550644
rect 41696 550598 41748 550604
rect 42062 550352 42118 550361
rect 42062 550287 42118 550296
rect 41696 547936 41748 547942
rect 41696 547878 41748 547884
rect 41708 547777 41736 547878
rect 41694 547768 41750 547777
rect 41694 547703 41750 547712
rect 42076 545737 42104 550287
rect 42062 545728 42118 545737
rect 42062 545663 42118 545672
rect 41524 543706 42472 543734
rect 41512 543040 41564 543046
rect 41512 542982 41564 542988
rect 37096 542360 37148 542366
rect 37096 542302 37148 542308
rect 41524 542178 41552 542982
rect 41696 542360 41748 542366
rect 41748 542308 42288 542314
rect 41696 542302 42288 542308
rect 41708 542286 42288 542302
rect 41524 542150 41828 542178
rect 41800 541113 41828 542150
rect 41786 541104 41842 541113
rect 41786 541039 41842 541048
rect 42260 540818 42288 542286
rect 42260 540790 42380 540818
rect 41786 540696 41842 540705
rect 41786 540631 41842 540640
rect 41800 540260 41828 540631
rect 42352 539050 42380 540790
rect 42182 539022 42380 539050
rect 42444 538778 42472 543706
rect 42614 540288 42670 540297
rect 42614 540223 42670 540232
rect 42076 538750 42472 538778
rect 42076 538424 42104 538750
rect 42338 538656 42394 538665
rect 42338 538591 42394 538600
rect 42352 538506 42380 538591
rect 42352 538478 42472 538506
rect 42246 538248 42302 538257
rect 42246 538183 42302 538192
rect 42260 538098 42288 538183
rect 42260 538070 42380 538098
rect 42062 537976 42118 537985
rect 42062 537911 42118 537920
rect 42076 537744 42104 537911
rect 42352 537758 42380 538070
rect 42444 537826 42472 538478
rect 42628 537985 42656 540223
rect 42614 537976 42670 537985
rect 42614 537911 42670 537920
rect 42444 537798 42564 537826
rect 42260 537730 42380 537758
rect 42168 536466 42196 536588
rect 42260 536466 42288 537730
rect 42536 537690 42564 537798
rect 42168 536438 42288 536466
rect 42444 537662 42564 537690
rect 42246 536344 42302 536353
rect 42246 536279 42302 536288
rect 42260 535378 42288 536279
rect 42182 535350 42288 535378
rect 42444 534766 42472 537662
rect 42614 537160 42670 537169
rect 42614 537095 42670 537104
rect 42168 534698 42196 534752
rect 42260 534738 42472 534766
rect 42260 534698 42288 534738
rect 42168 534670 42288 534698
rect 42628 534086 42656 537095
rect 42182 534058 42656 534086
rect 42154 533896 42210 533905
rect 42154 533831 42210 533840
rect 42168 533528 42196 533831
rect 42246 533216 42302 533225
rect 42246 533151 42302 533160
rect 42260 531162 42288 533151
rect 42522 532808 42578 532817
rect 42522 532743 42578 532752
rect 42168 531134 42288 531162
rect 42168 531045 42196 531134
rect 42536 530890 42564 532743
rect 42812 531314 42840 550616
rect 42996 533905 43024 552327
rect 43166 549536 43222 549545
rect 43166 549471 43222 549480
rect 42982 533896 43038 533905
rect 42982 533831 43038 533840
rect 43180 533225 43208 549471
rect 43166 533216 43222 533225
rect 43166 533151 43222 533160
rect 42352 530862 42564 530890
rect 42720 531286 42840 531314
rect 42352 530754 42380 530862
rect 42260 530726 42380 530754
rect 42260 530414 42288 530726
rect 42522 530632 42578 530641
rect 42182 530386 42288 530414
rect 42352 530590 42522 530618
rect 42154 530088 42210 530097
rect 42154 530023 42210 530032
rect 42168 529757 42196 530023
rect 41878 529408 41934 529417
rect 41878 529343 41934 529352
rect 41892 529205 41920 529343
rect 42352 527626 42380 530590
rect 42522 530567 42578 530576
rect 42720 530097 42748 531286
rect 42706 530088 42762 530097
rect 42706 530023 42762 530032
rect 42614 529680 42670 529689
rect 42614 529615 42670 529624
rect 42168 527598 42380 527626
rect 42168 527340 42196 527598
rect 42628 526742 42656 529615
rect 42890 529136 42946 529145
rect 42182 526714 42656 526742
rect 42720 529094 42890 529122
rect 42720 526091 42748 529094
rect 42890 529071 42946 529080
rect 42182 526063 42748 526091
rect 8588 431596 8616 431664
rect 9048 431596 9076 431664
rect 9508 431596 9536 431664
rect 9968 431596 9996 431664
rect 10428 431596 10456 431664
rect 10888 431596 10916 431664
rect 11348 431596 11376 431664
rect 11808 431596 11836 431664
rect 12268 431596 12296 431664
rect 12728 431596 12756 431664
rect 13188 431596 13216 431664
rect 13648 431596 13676 431664
rect 14108 431596 14136 431664
rect 41326 426048 41382 426057
rect 41326 425983 41382 425992
rect 40958 425640 41014 425649
rect 40958 425575 41014 425584
rect 36542 424416 36598 424425
rect 36542 424351 36598 424360
rect 36556 415410 36584 424351
rect 40972 422226 41000 425575
rect 41340 425054 41368 425983
rect 41340 425026 41552 425054
rect 41326 424008 41382 424017
rect 41326 423943 41382 423952
rect 41340 423706 41368 423943
rect 41328 423700 41380 423706
rect 41328 423642 41380 423648
rect 40972 422198 41184 422226
rect 41156 418849 41184 422198
rect 41142 418840 41198 418849
rect 41142 418775 41198 418784
rect 41524 418577 41552 425026
rect 41696 423700 41748 423706
rect 41748 423660 42840 423688
rect 41696 423642 41748 423648
rect 41878 422784 41934 422793
rect 41878 422719 41934 422728
rect 41510 418568 41566 418577
rect 41510 418503 41566 418512
rect 41892 417897 41920 422719
rect 42062 421968 42118 421977
rect 42062 421903 42118 421912
rect 41878 417888 41934 417897
rect 41878 417823 41934 417832
rect 42076 417625 42104 421903
rect 42430 419928 42486 419937
rect 42430 419863 42486 419872
rect 42246 418568 42302 418577
rect 42246 418503 42302 418512
rect 42062 417616 42118 417625
rect 42062 417551 42118 417560
rect 36544 415404 36596 415410
rect 36544 415346 36596 415352
rect 41696 415404 41748 415410
rect 42260 415394 42288 418503
rect 42444 415394 42472 419863
rect 42260 415366 42380 415394
rect 42444 415366 42564 415394
rect 41696 415346 41748 415352
rect 41708 415290 41736 415346
rect 41708 415262 42288 415290
rect 42260 413114 42288 415262
rect 42168 413086 42288 413114
rect 42168 412624 42196 413086
rect 42352 412026 42380 415366
rect 42260 411998 42380 412026
rect 42062 411904 42118 411913
rect 42062 411839 42118 411848
rect 42076 411468 42104 411839
rect 42260 411074 42288 411998
rect 42536 411913 42564 415366
rect 42522 411904 42578 411913
rect 42522 411839 42578 411848
rect 42168 411046 42288 411074
rect 42168 410788 42196 411046
rect 42182 410162 42472 410190
rect 41786 409456 41842 409465
rect 41786 409391 41842 409400
rect 41800 408952 41828 409391
rect 42444 408513 42472 410162
rect 42430 408504 42486 408513
rect 42430 408439 42486 408448
rect 42430 407824 42486 407833
rect 42168 407674 42196 407796
rect 42260 407782 42430 407810
rect 42260 407674 42288 407782
rect 42430 407759 42486 407768
rect 42168 407646 42288 407674
rect 42182 407102 42656 407130
rect 42430 407008 42486 407017
rect 42430 406943 42486 406952
rect 42444 406518 42472 406943
rect 42168 406450 42196 406504
rect 42260 406490 42472 406518
rect 42260 406450 42288 406490
rect 42168 406422 42288 406450
rect 41786 406328 41842 406337
rect 41786 406263 41842 406272
rect 41800 405929 41828 406263
rect 42628 405657 42656 407102
rect 42614 405648 42670 405657
rect 42614 405583 42670 405592
rect 41786 403880 41842 403889
rect 41786 403815 41842 403824
rect 41800 403444 41828 403815
rect 42338 402928 42394 402937
rect 42168 402886 42338 402914
rect 42168 402801 42196 402886
rect 42338 402863 42394 402872
rect 42182 402138 42472 402166
rect 41786 401840 41842 401849
rect 41786 401775 41842 401784
rect 41800 401608 41828 401775
rect 42444 400217 42472 402138
rect 42430 400208 42486 400217
rect 42430 400143 42486 400152
rect 42430 399800 42486 399809
rect 42182 399758 42430 399786
rect 42430 399735 42486 399744
rect 42812 399135 42840 423660
rect 43074 423192 43130 423201
rect 43074 423127 43130 423136
rect 43088 402937 43116 423127
rect 43258 421152 43314 421161
rect 43258 421087 43314 421096
rect 43272 407833 43300 421087
rect 43258 407824 43314 407833
rect 43258 407759 43314 407768
rect 43074 402928 43130 402937
rect 43074 402863 43130 402872
rect 42182 399107 42840 399135
rect 41786 398848 41842 398857
rect 41786 398783 41842 398792
rect 41800 398480 41828 398783
rect 8588 388348 8616 388484
rect 9048 388348 9076 388484
rect 9508 388348 9536 388484
rect 9968 388348 9996 388484
rect 10428 388348 10456 388484
rect 10888 388348 10916 388484
rect 11348 388348 11376 388484
rect 11808 388348 11836 388484
rect 12268 388348 12296 388484
rect 12728 388348 12756 388484
rect 13188 388348 13216 388484
rect 13648 388348 13676 388484
rect 14108 388348 14136 388484
rect 41340 387654 41552 387682
rect 41142 387152 41198 387161
rect 41142 387087 41144 387096
rect 41196 387087 41198 387096
rect 41144 387058 41196 387064
rect 41340 386753 41368 387654
rect 41524 386753 41552 387654
rect 41708 387122 41920 387138
rect 41696 387116 41920 387122
rect 41748 387110 41920 387116
rect 41696 387058 41748 387064
rect 41892 387025 41920 387110
rect 41878 387016 41934 387025
rect 41878 386951 41934 386960
rect 41326 386744 41382 386753
rect 41326 386679 41382 386688
rect 41510 386744 41566 386753
rect 41510 386679 41566 386688
rect 41326 382664 41382 382673
rect 41326 382599 41382 382608
rect 41340 382430 41368 382599
rect 41328 382424 41380 382430
rect 41328 382366 41380 382372
rect 41512 382424 41564 382430
rect 41512 382366 41564 382372
rect 40038 382256 40094 382265
rect 40038 382191 40094 382200
rect 37922 381440 37978 381449
rect 37922 381375 37978 381384
rect 33782 380216 33838 380225
rect 33782 380151 33838 380160
rect 28538 376544 28594 376553
rect 28538 376479 28594 376488
rect 28552 373289 28580 376479
rect 28538 373280 28594 373289
rect 28538 373215 28594 373224
rect 33796 371929 33824 380151
rect 35808 379568 35860 379574
rect 35808 379510 35860 379516
rect 35820 379409 35848 379510
rect 35806 379400 35862 379409
rect 35806 379335 35862 379344
rect 35806 376136 35862 376145
rect 35806 376071 35862 376080
rect 35820 375426 35848 376071
rect 35808 375420 35860 375426
rect 35808 375362 35860 375368
rect 37936 372638 37964 381375
rect 40052 376961 40080 382191
rect 40222 381032 40278 381041
rect 40222 380967 40278 380976
rect 40236 378554 40264 380967
rect 41524 379250 41552 382366
rect 41696 379568 41748 379574
rect 41748 379516 42840 379522
rect 41696 379510 42840 379516
rect 41708 379494 42840 379510
rect 41524 379222 42472 379250
rect 40224 378548 40276 378554
rect 40224 378490 40276 378496
rect 41696 378548 41748 378554
rect 41696 378490 41748 378496
rect 41708 378434 41736 378490
rect 41708 378406 42380 378434
rect 40038 376952 40094 376961
rect 40038 376887 40094 376896
rect 41694 375456 41750 375465
rect 41694 375391 41696 375400
rect 41748 375391 41750 375400
rect 41696 375362 41748 375368
rect 37924 372632 37976 372638
rect 41696 372632 41748 372638
rect 37924 372574 37976 372580
rect 41694 372600 41696 372609
rect 41748 372600 41750 372609
rect 41694 372535 41750 372544
rect 33782 371920 33838 371929
rect 33782 371855 33838 371864
rect 42352 370002 42380 378406
rect 42168 369974 42380 370002
rect 42168 369444 42196 369974
rect 42444 369854 42472 379222
rect 42614 372600 42670 372609
rect 42614 372535 42670 372544
rect 42352 369826 42472 369854
rect 41786 368520 41842 368529
rect 41786 368455 41842 368464
rect 41800 368249 41828 368455
rect 42352 367622 42380 369826
rect 42182 367594 42380 367622
rect 42430 367024 42486 367033
rect 42182 366968 42430 366975
rect 42182 366959 42486 366968
rect 42182 366947 42472 366959
rect 42628 365922 42656 372535
rect 42536 365894 42656 365922
rect 42338 365800 42394 365809
rect 42182 365758 42338 365786
rect 42338 365735 42394 365744
rect 42154 364984 42210 364993
rect 42154 364919 42210 364928
rect 42168 364548 42196 364919
rect 42536 364426 42564 365894
rect 42812 365809 42840 379494
rect 43456 379514 43484 590271
rect 44468 581097 44496 591903
rect 44454 581088 44510 581097
rect 44454 581023 44510 581032
rect 44652 557297 44680 600063
rect 44836 599729 44864 618226
rect 44822 599720 44878 599729
rect 44822 599655 44878 599664
rect 44822 599312 44878 599321
rect 44822 599247 44878 599256
rect 44638 557288 44694 557297
rect 44638 557223 44694 557232
rect 44836 556481 44864 599247
rect 45020 598097 45048 618226
rect 45204 598913 45232 635446
rect 45374 633448 45430 633457
rect 45374 633383 45430 633392
rect 45388 610910 45416 633383
rect 45572 612202 45600 764215
rect 46216 754089 46244 870810
rect 47584 818372 47636 818378
rect 47584 818314 47636 818320
rect 46386 763056 46442 763065
rect 46386 762991 46442 763000
rect 46202 754080 46258 754089
rect 46202 754015 46258 754024
rect 45742 676696 45798 676705
rect 45742 676631 45798 676640
rect 45560 612196 45612 612202
rect 45560 612138 45612 612144
rect 45756 611318 45784 676631
rect 46018 637800 46074 637809
rect 46018 637735 46074 637744
rect 46032 615641 46060 637735
rect 46202 636984 46258 636993
rect 46202 636919 46258 636928
rect 46216 619041 46244 636919
rect 46202 619032 46258 619041
rect 46202 618967 46258 618976
rect 46018 615632 46074 615641
rect 46018 615567 46074 615576
rect 46400 612406 46428 762991
rect 46938 719944 46994 719953
rect 46938 719879 46994 719888
rect 46388 612400 46440 612406
rect 46388 612342 46440 612348
rect 46952 611726 46980 719879
rect 47596 710841 47624 818314
rect 47780 817737 47808 896990
rect 47766 817728 47822 817737
rect 47766 817663 47822 817672
rect 50356 816921 50384 909434
rect 50342 816912 50398 816921
rect 50342 816847 50398 816856
rect 50344 805996 50396 806002
rect 50344 805938 50396 805944
rect 48964 767372 49016 767378
rect 48964 767314 49016 767320
rect 47582 710832 47638 710841
rect 47582 710767 47638 710776
rect 47214 677920 47270 677929
rect 47214 677855 47270 677864
rect 46940 611720 46992 611726
rect 46940 611662 46992 611668
rect 45744 611312 45796 611318
rect 45744 611254 45796 611260
rect 47228 611114 47256 677855
rect 48976 669361 49004 767314
rect 50356 730561 50384 805938
rect 53116 799241 53144 923238
rect 53300 892809 53328 990218
rect 53286 892800 53342 892809
rect 53286 892735 53342 892744
rect 54496 892265 54524 992870
rect 55864 991500 55916 991506
rect 55864 991442 55916 991448
rect 55876 892265 55904 991442
rect 95896 990282 95924 1001914
rect 96080 991778 96108 1002050
rect 97276 996169 97304 1002594
rect 98644 1002516 98696 1002522
rect 98644 1002458 98696 1002464
rect 97448 1002380 97500 1002386
rect 97448 1002322 97500 1002328
rect 97262 996160 97318 996169
rect 97262 996095 97318 996104
rect 97460 995858 97488 1002322
rect 98274 1002008 98330 1002017
rect 98274 1001943 98276 1001952
rect 98328 1001943 98330 1001952
rect 98276 1001914 98328 1001920
rect 97448 995852 97500 995858
rect 97448 995794 97500 995800
rect 98656 994566 98684 1002458
rect 100298 1002416 100354 1002425
rect 100298 1002351 100300 1002360
rect 100352 1002351 100354 1002360
rect 100484 1002380 100536 1002386
rect 100300 1002322 100352 1002328
rect 100484 1002322 100536 1002328
rect 98828 1002244 98880 1002250
rect 98828 1002186 98880 1002192
rect 98840 995586 98868 1002186
rect 99102 1002144 99158 1002153
rect 99102 1002079 99104 1002088
rect 99156 1002079 99158 1002088
rect 100024 1002108 100076 1002114
rect 99104 1002050 99156 1002056
rect 100024 1002050 100076 1002056
rect 99012 1001972 99064 1001978
rect 99012 1001914 99064 1001920
rect 99024 999802 99052 1001914
rect 99012 999796 99064 999802
rect 99012 999738 99064 999744
rect 98828 995580 98880 995586
rect 98828 995522 98880 995528
rect 100036 994702 100064 1002050
rect 100496 998442 100524 1002322
rect 101126 1002280 101182 1002289
rect 101126 1002215 101128 1002224
rect 101180 1002215 101182 1002224
rect 101128 1002186 101180 1002192
rect 101126 1002008 101182 1002017
rect 101126 1001943 101128 1001952
rect 101180 1001943 101182 1001952
rect 101128 1001914 101180 1001920
rect 100484 998436 100536 998442
rect 100484 998378 100536 998384
rect 101416 995081 101444 1006266
rect 104806 1006224 104862 1006233
rect 101588 1006188 101640 1006194
rect 104806 1006159 104808 1006168
rect 101588 1006130 101640 1006136
rect 104860 1006159 104862 1006168
rect 106830 1006224 106886 1006233
rect 106830 1006159 106832 1006168
rect 104808 1006130 104860 1006136
rect 106884 1006159 106886 1006168
rect 113824 1006188 113876 1006194
rect 106832 1006130 106884 1006136
rect 113824 1006130 113876 1006136
rect 101600 997694 101628 1006130
rect 103150 1006088 103206 1006097
rect 103150 1006023 103152 1006032
rect 103204 1006023 103206 1006032
rect 106002 1006088 106058 1006097
rect 106002 1006023 106004 1006032
rect 103152 1005994 103204 1006000
rect 106056 1006023 106058 1006032
rect 106004 1005994 106056 1006000
rect 102784 1005304 102836 1005310
rect 108856 1005304 108908 1005310
rect 102784 1005246 102836 1005252
rect 108854 1005272 108856 1005281
rect 108908 1005272 108910 1005281
rect 101954 1002552 102010 1002561
rect 101954 1002487 101956 1002496
rect 102008 1002487 102010 1002496
rect 101956 1002458 102008 1002464
rect 102322 1002144 102378 1002153
rect 102322 1002079 102324 1002088
rect 102376 1002079 102378 1002088
rect 102324 1002050 102376 1002056
rect 101588 997688 101640 997694
rect 101588 997630 101640 997636
rect 101402 995072 101458 995081
rect 101402 995007 101458 995016
rect 100024 994696 100076 994702
rect 100024 994638 100076 994644
rect 98644 994560 98696 994566
rect 98644 994502 98696 994508
rect 96068 991772 96120 991778
rect 96068 991714 96120 991720
rect 95884 990276 95936 990282
rect 95884 990218 95936 990224
rect 89628 986128 89680 986134
rect 89628 986070 89680 986076
rect 73436 985992 73488 985998
rect 73436 985934 73488 985940
rect 73448 983620 73476 985934
rect 89640 983620 89668 986070
rect 102796 985998 102824 1005246
rect 108854 1005207 108910 1005216
rect 108486 1004728 108542 1004737
rect 106188 1004692 106240 1004698
rect 108486 1004663 108488 1004672
rect 106188 1004634 106240 1004640
rect 108540 1004663 108542 1004672
rect 108488 1004634 108540 1004640
rect 103150 1002416 103206 1002425
rect 103150 1002351 103152 1002360
rect 103204 1002351 103206 1002360
rect 103152 1002322 103204 1002328
rect 105634 1002280 105690 1002289
rect 105634 1002215 105636 1002224
rect 105688 1002215 105690 1002224
rect 105636 1002186 105688 1002192
rect 103978 1002144 104034 1002153
rect 103978 1002079 103980 1002088
rect 104032 1002079 104034 1002088
rect 103980 1002050 104032 1002056
rect 104806 1002008 104862 1002017
rect 104176 1001966 104806 1001994
rect 104176 994809 104204 1001966
rect 104806 1001943 104862 1001952
rect 106002 1002008 106058 1002017
rect 106002 1001943 106004 1001952
rect 106056 1001943 106058 1001952
rect 106004 1001914 106056 1001920
rect 104162 994800 104218 994809
rect 104162 994735 104218 994744
rect 102784 985992 102836 985998
rect 102784 985934 102836 985940
rect 106200 983634 106228 1004634
rect 107658 1002416 107714 1002425
rect 107658 1002351 107660 1002360
rect 107712 1002351 107714 1002360
rect 109500 1002380 109552 1002386
rect 107660 1002322 107712 1002328
rect 109500 1002322 109552 1002328
rect 108026 1002280 108082 1002289
rect 107844 1002244 107896 1002250
rect 108026 1002215 108028 1002224
rect 107844 1002186 107896 1002192
rect 108080 1002215 108082 1002224
rect 108028 1002186 108080 1002192
rect 106830 1002144 106886 1002153
rect 106464 1002108 106516 1002114
rect 107856 1002130 107884 1002186
rect 107856 1002102 108160 1002130
rect 106830 1002079 106832 1002088
rect 106464 1002050 106516 1002056
rect 106884 1002079 106886 1002088
rect 106832 1002050 106884 1002056
rect 106476 994838 106504 1002050
rect 107752 1001972 107804 1001978
rect 107752 1001914 107804 1001920
rect 106464 994832 106516 994838
rect 106464 994774 106516 994780
rect 107764 993206 107792 1001914
rect 107752 993200 107804 993206
rect 107752 993142 107804 993148
rect 108132 990146 108160 1002102
rect 109040 1002108 109092 1002114
rect 109040 1002050 109092 1002056
rect 109052 993070 109080 1002050
rect 109512 997694 109540 1002322
rect 110420 1002244 110472 1002250
rect 110420 1002186 110472 1002192
rect 109682 1002144 109738 1002153
rect 109682 1002079 109684 1002088
rect 109736 1002079 109738 1002088
rect 109684 1002050 109736 1002056
rect 109500 997688 109552 997694
rect 109500 997630 109552 997636
rect 109040 993064 109092 993070
rect 109040 993006 109092 993012
rect 110432 991642 110460 1002186
rect 111800 1002108 111852 1002114
rect 111800 1002050 111852 1002056
rect 110420 991636 110472 991642
rect 110420 991578 110472 991584
rect 108120 990140 108172 990146
rect 108120 990082 108172 990088
rect 111812 986134 111840 1002050
rect 113836 997558 113864 1006130
rect 124864 1006052 124916 1006058
rect 124864 1005994 124916 1006000
rect 121736 997824 121788 997830
rect 121736 997766 121788 997772
rect 117228 997688 117280 997694
rect 117228 997630 117280 997636
rect 113824 997552 113876 997558
rect 113824 997494 113876 997500
rect 116952 997552 117004 997558
rect 116952 997494 117004 997500
rect 116964 996985 116992 997494
rect 117240 997257 117268 997630
rect 117226 997248 117282 997257
rect 117226 997183 117282 997192
rect 116950 996976 117006 996985
rect 116950 996911 117006 996920
rect 111800 986128 111852 986134
rect 111800 986070 111852 986076
rect 105846 983606 106228 983634
rect 121748 983634 121776 997766
rect 124876 995081 124904 1005994
rect 126256 996305 126284 1006266
rect 144000 998436 144052 998442
rect 144000 998378 144052 998384
rect 143816 997756 143868 997762
rect 143816 997698 143868 997704
rect 143828 997257 143856 997698
rect 143814 997248 143870 997257
rect 143814 997183 143870 997192
rect 143724 996396 143776 996402
rect 143724 996338 143776 996344
rect 126242 996296 126298 996305
rect 126242 996231 126298 996240
rect 140792 995858 140820 995860
rect 140780 995852 140832 995858
rect 140780 995794 140832 995800
rect 131854 995752 131910 995761
rect 131606 995710 131854 995738
rect 131854 995687 131910 995696
rect 132958 995752 133014 995761
rect 136730 995752 136786 995761
rect 133014 995710 133446 995738
rect 136482 995710 136730 995738
rect 132958 995687 133014 995696
rect 137374 995752 137430 995761
rect 137126 995710 137374 995738
rect 136730 995687 136786 995696
rect 140410 995752 140466 995761
rect 140162 995710 140410 995738
rect 137374 995687 137430 995696
rect 143736 995738 143764 996338
rect 144012 995858 144040 998378
rect 144196 996169 144224 1006674
rect 145748 1006596 145800 1006602
rect 145748 1006538 145800 1006544
rect 145564 1006460 145616 1006466
rect 145564 1006402 145616 1006408
rect 144368 1006256 144420 1006262
rect 144368 1006198 144420 1006204
rect 144380 996441 144408 1006198
rect 144828 997620 144880 997626
rect 144828 997562 144880 997568
rect 144644 997076 144696 997082
rect 144644 997018 144696 997024
rect 144366 996432 144422 996441
rect 144366 996367 144422 996376
rect 144182 996160 144238 996169
rect 144182 996095 144238 996104
rect 144000 995852 144052 995858
rect 144000 995794 144052 995800
rect 140410 995687 140466 995696
rect 143460 995710 143764 995738
rect 141790 995616 141846 995625
rect 141450 995574 141790 995602
rect 141790 995551 141846 995560
rect 124862 995072 124918 995081
rect 124862 995007 124918 995016
rect 128464 994430 128492 995452
rect 129108 994702 129136 995452
rect 129752 994838 129780 995452
rect 129740 994832 129792 994838
rect 132144 994809 132172 995452
rect 132802 995438 133184 995466
rect 132406 995344 132462 995353
rect 132406 995279 132462 995288
rect 129740 994774 129792 994780
rect 132130 994800 132186 994809
rect 132130 994735 132186 994744
rect 129096 994696 129148 994702
rect 129096 994638 129148 994644
rect 132420 994566 132448 995279
rect 132408 994560 132460 994566
rect 133156 994537 133184 995438
rect 135916 994809 135944 995452
rect 137100 994832 137152 994838
rect 135902 994800 135958 994809
rect 137100 994774 137152 994780
rect 137284 994832 137336 994838
rect 137284 994774 137336 994780
rect 135902 994735 135958 994744
rect 132408 994502 132460 994508
rect 133142 994528 133198 994537
rect 133142 994463 133198 994472
rect 128452 994424 128504 994430
rect 128452 994366 128504 994372
rect 137112 994294 137140 994774
rect 137296 994430 137324 994774
rect 137284 994424 137336 994430
rect 137284 994366 137336 994372
rect 137100 994288 137152 994294
rect 137100 994230 137152 994236
rect 137756 993721 137784 995452
rect 138966 995438 139348 995466
rect 142646 995438 143028 995466
rect 139320 995058 139348 995438
rect 143000 995330 143028 995438
rect 143460 995330 143488 995710
rect 143724 995580 143776 995586
rect 143724 995522 143776 995528
rect 143000 995302 143488 995330
rect 139320 995030 139440 995058
rect 139216 994152 139268 994158
rect 139216 994094 139268 994100
rect 139228 993993 139256 994094
rect 139412 993993 139440 995030
rect 141882 994800 141938 994809
rect 141882 994735 141938 994744
rect 142066 994800 142122 994809
rect 142066 994735 142122 994744
rect 141896 994022 141924 994735
rect 142080 994158 142108 994735
rect 143736 994265 143764 995522
rect 144656 994294 144684 997018
rect 144840 996985 144868 997562
rect 144826 996976 144882 996985
rect 144826 996911 144882 996920
rect 144644 994288 144696 994294
rect 143722 994256 143778 994265
rect 143722 994191 143778 994200
rect 143906 994256 143962 994265
rect 144644 994230 144696 994236
rect 143906 994191 143962 994200
rect 142068 994152 142120 994158
rect 142068 994094 142120 994100
rect 141884 994016 141936 994022
rect 139214 993984 139270 993993
rect 139214 993919 139270 993928
rect 139398 993984 139454 993993
rect 141884 993958 141936 993964
rect 142344 994016 142396 994022
rect 142344 993958 142396 993964
rect 139398 993919 139454 993928
rect 142160 993744 142212 993750
rect 137742 993712 137798 993721
rect 137742 993647 137798 993656
rect 142158 993712 142160 993721
rect 142356 993721 142384 993958
rect 143920 993750 143948 994191
rect 145576 993993 145604 1006402
rect 145760 995586 145788 1006538
rect 150268 1006126 150296 1006674
rect 153750 1006632 153806 1006641
rect 153750 1006567 153752 1006576
rect 153804 1006567 153806 1006576
rect 157430 1006632 157486 1006641
rect 157430 1006567 157432 1006576
rect 153752 1006538 153804 1006544
rect 157484 1006567 157486 1006576
rect 157432 1006538 157484 1006544
rect 152922 1006496 152978 1006505
rect 152922 1006431 152924 1006440
rect 152976 1006431 152978 1006440
rect 160282 1006496 160338 1006505
rect 161952 1006466 161980 1006674
rect 160282 1006431 160284 1006440
rect 152924 1006402 152976 1006408
rect 160336 1006431 160338 1006440
rect 161940 1006460 161992 1006466
rect 160284 1006402 160336 1006408
rect 161940 1006402 161992 1006408
rect 162768 1006460 162820 1006466
rect 162768 1006402 162820 1006408
rect 152094 1006360 152150 1006369
rect 152094 1006295 152096 1006304
rect 152148 1006295 152150 1006304
rect 158258 1006360 158314 1006369
rect 158258 1006295 158260 1006304
rect 152096 1006266 152148 1006272
rect 158312 1006295 158314 1006304
rect 158260 1006266 158312 1006272
rect 151268 1006256 151320 1006262
rect 151266 1006224 151268 1006233
rect 151320 1006224 151322 1006233
rect 151266 1006159 151322 1006168
rect 158626 1006224 158682 1006233
rect 162780 1006194 162808 1006402
rect 158626 1006159 158628 1006168
rect 158680 1006159 158682 1006168
rect 162768 1006188 162820 1006194
rect 158628 1006130 158680 1006136
rect 162768 1006130 162820 1006136
rect 148876 1006120 148928 1006126
rect 147126 1006088 147182 1006097
rect 147126 1006023 147182 1006032
rect 148874 1006088 148876 1006097
rect 150072 1006120 150124 1006126
rect 148928 1006088 148930 1006097
rect 148874 1006023 148930 1006032
rect 150070 1006088 150072 1006097
rect 150256 1006120 150308 1006126
rect 150124 1006088 150126 1006097
rect 150256 1006062 150308 1006068
rect 158258 1006088 158314 1006097
rect 150070 1006023 150126 1006032
rect 153936 1006052 153988 1006058
rect 146944 1001972 146996 1001978
rect 146944 1001914 146996 1001920
rect 145748 995580 145800 995586
rect 145748 995522 145800 995528
rect 145562 993984 145618 993993
rect 145562 993919 145618 993928
rect 143908 993744 143960 993750
rect 142212 993712 142214 993721
rect 142158 993647 142214 993656
rect 142342 993712 142398 993721
rect 143908 993686 143960 993692
rect 142342 993647 142398 993656
rect 138296 991636 138348 991642
rect 138296 991578 138348 991584
rect 121748 983606 122130 983634
rect 138308 983620 138336 991578
rect 146956 991506 146984 1001914
rect 147140 995625 147168 1006023
rect 158258 1006023 158260 1006032
rect 153936 1005994 153988 1006000
rect 158312 1006023 158314 1006032
rect 159454 1006088 159510 1006097
rect 159454 1006023 159456 1006032
rect 158260 1005994 158312 1006000
rect 159508 1006023 159510 1006032
rect 159456 1005994 159508 1006000
rect 153750 1005136 153806 1005145
rect 151084 1005100 151136 1005106
rect 153750 1005071 153752 1005080
rect 151084 1005042 151136 1005048
rect 153804 1005071 153806 1005080
rect 153752 1005042 153804 1005048
rect 149704 1004964 149756 1004970
rect 149704 1004906 149756 1004912
rect 148508 1002380 148560 1002386
rect 148508 1002322 148560 1002328
rect 148324 1002108 148376 1002114
rect 148324 1002050 148376 1002056
rect 147126 995616 147182 995625
rect 147126 995551 147182 995560
rect 148336 992934 148364 1002050
rect 148520 994265 148548 1002322
rect 149242 1002008 149298 1002017
rect 149242 1001943 149244 1001952
rect 149296 1001943 149298 1001952
rect 149244 1001914 149296 1001920
rect 149716 994537 149744 1004906
rect 149888 1004692 149940 1004698
rect 149888 1004634 149940 1004640
rect 149900 994566 149928 1004634
rect 150898 1002416 150954 1002425
rect 150898 1002351 150900 1002360
rect 150952 1002351 150954 1002360
rect 150900 1002322 150952 1002328
rect 150898 1002144 150954 1002153
rect 150898 1002079 150900 1002088
rect 150952 1002079 150954 1002088
rect 150900 1002050 150952 1002056
rect 151096 994702 151124 1005042
rect 152922 1005000 152978 1005009
rect 152922 1004935 152924 1004944
rect 152976 1004935 152978 1004944
rect 152924 1004906 152976 1004912
rect 151268 1004828 151320 1004834
rect 151268 1004770 151320 1004776
rect 151280 996402 151308 1004770
rect 151726 1004728 151782 1004737
rect 151726 1004663 151728 1004672
rect 151780 1004663 151782 1004672
rect 151728 1004634 151780 1004640
rect 152464 1002108 152516 1002114
rect 152464 1002050 152516 1002056
rect 151268 996396 151320 996402
rect 151268 996338 151320 996344
rect 151084 994696 151136 994702
rect 151084 994638 151136 994644
rect 149888 994560 149940 994566
rect 149702 994528 149758 994537
rect 149888 994502 149940 994508
rect 149702 994463 149758 994472
rect 148506 994256 148562 994265
rect 148506 994191 148562 994200
rect 152476 993721 152504 1002050
rect 153948 997762 153976 1005994
rect 154118 1004864 154174 1004873
rect 154118 1004799 154120 1004808
rect 154172 1004799 154174 1004808
rect 160650 1004864 160706 1004873
rect 160650 1004799 160652 1004808
rect 154120 1004770 154172 1004776
rect 160704 1004799 160706 1004808
rect 163136 1004828 163188 1004834
rect 160652 1004770 160704 1004776
rect 163136 1004770 163188 1004776
rect 161110 1004728 161166 1004737
rect 161110 1004663 161112 1004672
rect 161164 1004663 161166 1004672
rect 162952 1004692 163004 1004698
rect 161112 1004634 161164 1004640
rect 162952 1004634 163004 1004640
rect 155774 1002280 155830 1002289
rect 155774 1002215 155776 1002224
rect 155828 1002215 155830 1002224
rect 157340 1002244 157392 1002250
rect 155776 1002186 155828 1002192
rect 157340 1002186 157392 1002192
rect 154578 1002144 154634 1002153
rect 154578 1002079 154580 1002088
rect 154632 1002079 154634 1002088
rect 154580 1002050 154632 1002056
rect 154946 1002008 155002 1002017
rect 154592 1001966 154946 1001994
rect 153936 997756 153988 997762
rect 153936 997698 153988 997704
rect 154302 995752 154358 995761
rect 154302 995687 154358 995696
rect 154316 995081 154344 995687
rect 154302 995072 154358 995081
rect 154302 995007 154358 995016
rect 154592 994537 154620 1001966
rect 154946 1001943 155002 1001952
rect 155774 1002008 155830 1002017
rect 156602 1002008 156658 1002017
rect 155830 1001966 156000 1001994
rect 155774 1001943 155830 1001952
rect 155972 998442 156000 1001966
rect 156602 1001943 156604 1001952
rect 156656 1001943 156658 1001952
rect 156604 1001914 156656 1001920
rect 155960 998436 156012 998442
rect 155960 998378 156012 998384
rect 157352 994702 157380 1002186
rect 157798 1002144 157854 1002153
rect 157798 1002079 157800 1002088
rect 157852 1002079 157854 1002088
rect 160100 1002108 160152 1002114
rect 157800 1002050 157852 1002056
rect 160100 1002050 160152 1002056
rect 158720 1001972 158772 1001978
rect 158720 1001914 158772 1001920
rect 158732 997082 158760 1001914
rect 160112 997626 160140 1002050
rect 160100 997620 160152 997626
rect 160100 997562 160152 997568
rect 162964 997218 162992 1004634
rect 160744 997212 160796 997218
rect 160744 997154 160796 997160
rect 162952 997212 163004 997218
rect 162952 997154 163004 997160
rect 158720 997076 158772 997082
rect 158720 997018 158772 997024
rect 157340 994696 157392 994702
rect 157340 994638 157392 994644
rect 154578 994528 154634 994537
rect 154578 994463 154634 994472
rect 152462 993712 152518 993721
rect 152462 993647 152518 993656
rect 148324 992928 148376 992934
rect 148324 992870 148376 992876
rect 146944 991500 146996 991506
rect 146944 991442 146996 991448
rect 160756 985726 160784 997154
rect 163148 991642 163176 1004770
rect 163136 991636 163188 991642
rect 163136 991578 163188 991584
rect 164896 990894 164924 1006674
rect 166264 1006596 166316 1006602
rect 166264 1006538 166316 1006544
rect 173164 1006596 173216 1006602
rect 173164 1006538 173216 1006544
rect 364892 1006596 364944 1006602
rect 364892 1006538 364944 1006544
rect 371884 1006596 371936 1006602
rect 371884 1006538 371936 1006544
rect 166276 1006194 166304 1006538
rect 171784 1006324 171836 1006330
rect 171784 1006266 171836 1006272
rect 166264 1006188 166316 1006194
rect 166264 1006130 166316 1006136
rect 171796 996130 171824 1006266
rect 171784 996124 171836 996130
rect 171784 996066 171836 996072
rect 170680 995988 170732 995994
rect 170680 995930 170732 995936
rect 171232 995988 171284 995994
rect 171232 995930 171284 995936
rect 169392 995852 169444 995858
rect 169392 995794 169444 995800
rect 169404 994158 169432 995794
rect 170496 994764 170548 994770
rect 170496 994706 170548 994712
rect 169392 994152 169444 994158
rect 169392 994094 169444 994100
rect 170508 993682 170536 994706
rect 170692 994634 170720 995930
rect 171048 995580 171100 995586
rect 171048 995522 171100 995528
rect 170862 995344 170918 995353
rect 170862 995279 170918 995288
rect 170680 994628 170732 994634
rect 170680 994570 170732 994576
rect 170876 994498 170904 995279
rect 171060 994770 171088 995522
rect 171244 995111 171272 995930
rect 171508 995852 171560 995858
rect 171508 995794 171560 995800
rect 171520 995223 171548 995794
rect 171690 995344 171746 995353
rect 171690 995279 171692 995288
rect 171744 995279 171746 995288
rect 171692 995271 171744 995277
rect 171508 995217 171560 995223
rect 171508 995159 171560 995165
rect 171232 995105 171284 995111
rect 173176 995081 173204 1006538
rect 256146 1006496 256202 1006505
rect 247684 1006460 247736 1006466
rect 256146 1006431 256148 1006440
rect 247684 1006402 247736 1006408
rect 256200 1006431 256202 1006440
rect 354862 1006496 354918 1006505
rect 354862 1006431 354864 1006440
rect 256148 1006402 256200 1006408
rect 354916 1006431 354918 1006440
rect 363604 1006460 363656 1006466
rect 354864 1006402 354916 1006408
rect 363604 1006402 363656 1006408
rect 210422 1006224 210478 1006233
rect 175924 1006188 175976 1006194
rect 210422 1006159 210424 1006168
rect 175924 1006130 175976 1006136
rect 210476 1006159 210478 1006168
rect 228364 1006188 228416 1006194
rect 210424 1006130 210476 1006136
rect 228364 1006130 228416 1006136
rect 175936 995897 175964 1006130
rect 201038 1006088 201094 1006097
rect 177304 1006052 177356 1006058
rect 177304 1005994 177356 1006000
rect 195152 1006052 195204 1006058
rect 201038 1006023 201040 1006032
rect 195152 1005994 195204 1006000
rect 201092 1006023 201094 1006032
rect 208398 1006088 208454 1006097
rect 208398 1006023 208400 1006032
rect 201040 1005994 201092 1006000
rect 208452 1006023 208454 1006032
rect 208400 1005994 208452 1006000
rect 175922 995888 175978 995897
rect 175922 995823 175978 995832
rect 177316 995625 177344 1005994
rect 195164 1004654 195192 1005994
rect 204904 1005304 204956 1005310
rect 212080 1005304 212132 1005310
rect 204904 1005246 204956 1005252
rect 212078 1005272 212080 1005281
rect 212132 1005272 212134 1005281
rect 195164 1004626 195468 1004654
rect 195152 1001768 195204 1001774
rect 195152 1001710 195204 1001716
rect 195164 997754 195192 1001710
rect 195164 997726 195284 997754
rect 195058 995888 195114 995897
rect 195058 995823 195114 995832
rect 192482 995786 192538 995795
rect 192188 995730 192482 995738
rect 192188 995721 192538 995730
rect 192188 995710 192524 995721
rect 177302 995616 177358 995625
rect 177302 995551 177358 995560
rect 194876 995512 194928 995518
rect 179860 995438 180196 995466
rect 180504 995438 180748 995466
rect 181148 995438 181484 995466
rect 180168 995110 180196 995438
rect 180720 995382 180748 995438
rect 180708 995376 180760 995382
rect 180708 995318 180760 995324
rect 180156 995104 180208 995110
rect 171232 995047 171284 995053
rect 173162 995072 173218 995081
rect 180156 995046 180208 995052
rect 173162 995007 173218 995016
rect 181456 994974 181484 995438
rect 182974 995246 183002 995452
rect 183540 995438 183876 995466
rect 184184 995438 184520 995466
rect 184828 995438 184888 995466
rect 187312 995438 187648 995466
rect 187864 995438 188200 995466
rect 188508 995438 188844 995466
rect 189152 995438 189488 995466
rect 190348 995438 190408 995466
rect 191544 995438 191788 995466
rect 192832 995438 193168 995466
rect 194028 995438 194456 995466
rect 194876 995454 194928 995460
rect 183848 995353 183876 995438
rect 183834 995344 183890 995353
rect 183834 995279 183890 995288
rect 182962 995240 183014 995246
rect 182962 995182 183014 995188
rect 181444 994968 181496 994974
rect 181444 994910 181496 994916
rect 171232 994881 171284 994887
rect 171232 994823 171284 994829
rect 171048 994764 171100 994770
rect 171048 994706 171100 994712
rect 170864 994492 170916 994498
rect 170864 994434 170916 994440
rect 171244 993818 171272 994823
rect 184492 994362 184520 995438
rect 184480 994356 184532 994362
rect 184480 994298 184532 994304
rect 184860 994265 184888 995438
rect 187620 994809 187648 995438
rect 187606 994800 187662 994809
rect 187606 994735 187662 994744
rect 184846 994256 184902 994265
rect 184846 994191 184902 994200
rect 171232 993812 171284 993818
rect 171232 993754 171284 993760
rect 170496 993676 170548 993682
rect 170496 993618 170548 993624
rect 188172 993546 188200 995438
rect 188816 994537 188844 995438
rect 188802 994528 188858 994537
rect 188802 994463 188858 994472
rect 189460 993993 189488 995438
rect 190380 994537 190408 995438
rect 190366 994528 190422 994537
rect 190366 994463 190422 994472
rect 191760 994362 191788 995438
rect 191104 994356 191156 994362
rect 191104 994298 191156 994304
rect 191748 994356 191800 994362
rect 191748 994298 191800 994304
rect 191116 994022 191144 994298
rect 191104 994016 191156 994022
rect 189446 993984 189502 993993
rect 191104 993958 191156 993964
rect 189446 993919 189502 993928
rect 193140 993721 193168 995438
rect 194428 995330 194456 995438
rect 194888 995330 194916 995454
rect 195072 995353 195100 995823
rect 194428 995302 194916 995330
rect 195058 995344 195114 995353
rect 195058 995279 195114 995288
rect 195256 994809 195284 997726
rect 195242 994800 195298 994809
rect 195242 994735 195298 994744
rect 195440 994004 195468 1004626
rect 202880 1002516 202932 1002522
rect 202880 1002458 202932 1002464
rect 202892 1001978 202920 1002458
rect 202880 1001972 202932 1001978
rect 202880 1001914 202932 1001920
rect 204168 1001972 204220 1001978
rect 204168 1001914 204220 1001920
rect 202694 1001192 202750 1001201
rect 202524 1001150 202694 1001178
rect 200212 998844 200264 998850
rect 200212 998786 200264 998792
rect 196808 998708 196860 998714
rect 196808 998650 196860 998656
rect 196624 998572 196676 998578
rect 196624 998514 196676 998520
rect 195704 998436 195756 998442
rect 195704 998378 195756 998384
rect 195716 997754 195744 998378
rect 196070 997792 196126 997801
rect 195716 997726 195836 997754
rect 196070 997727 196126 997736
rect 195612 996260 195664 996266
rect 195612 996202 195664 996208
rect 195624 995602 195652 996202
rect 195808 996146 195836 997726
rect 195348 993976 195468 994004
rect 195532 995574 195652 995602
rect 195716 996118 195836 996146
rect 195348 993721 195376 993976
rect 195532 993818 195560 995574
rect 195716 995518 195744 996118
rect 195888 995988 195940 995994
rect 195888 995930 195940 995936
rect 195704 995512 195756 995518
rect 195704 995454 195756 995460
rect 195520 993812 195572 993818
rect 195520 993754 195572 993760
rect 193126 993712 193182 993721
rect 193126 993647 193182 993656
rect 195334 993712 195390 993721
rect 195334 993647 195390 993656
rect 195900 993546 195928 995930
rect 196084 994537 196112 997727
rect 196070 994528 196126 994537
rect 196070 994463 196126 994472
rect 196636 994265 196664 998514
rect 196622 994256 196678 994265
rect 196622 994191 196678 994200
rect 196820 994022 196848 998650
rect 199384 998096 199436 998102
rect 199384 998038 199436 998044
rect 197544 997960 197596 997966
rect 197544 997902 197596 997908
rect 197360 997076 197412 997082
rect 197360 997018 197412 997024
rect 197372 994362 197400 997018
rect 197360 994356 197412 994362
rect 197360 994298 197412 994304
rect 196808 994016 196860 994022
rect 196808 993958 196860 993964
rect 197556 993682 197584 997902
rect 199396 993993 199424 998038
rect 200224 997801 200252 998786
rect 200396 998232 200448 998238
rect 200396 998174 200448 998180
rect 200210 997792 200266 997801
rect 200210 997727 200266 997736
rect 200212 997280 200264 997286
rect 200210 997248 200212 997257
rect 200264 997248 200266 997257
rect 200210 997183 200266 997192
rect 200408 996826 200436 998174
rect 201868 997960 201920 997966
rect 201866 997928 201868 997937
rect 202144 997960 202196 997966
rect 201920 997928 201922 997937
rect 202144 997902 202196 997908
rect 201866 997863 201922 997872
rect 200224 996798 200436 996826
rect 200224 996713 200252 996798
rect 200210 996704 200266 996713
rect 200210 996639 200266 996648
rect 200670 996296 200726 996305
rect 200670 996231 200672 996240
rect 200724 996231 200726 996240
rect 200672 996202 200724 996208
rect 202156 995382 202184 997902
rect 202328 997824 202380 997830
rect 202328 997766 202380 997772
rect 202340 995897 202368 997766
rect 202524 995994 202552 1001150
rect 202694 1001127 202750 1001136
rect 203890 998880 203946 998889
rect 203890 998815 203892 998824
rect 203944 998815 203946 998824
rect 203892 998786 203944 998792
rect 203522 998608 203578 998617
rect 203522 998543 203524 998552
rect 203576 998543 203578 998552
rect 203524 998514 203576 998520
rect 204180 998442 204208 1001914
rect 204350 998744 204406 998753
rect 204350 998679 204352 998688
rect 204404 998679 204406 998688
rect 204352 998650 204404 998656
rect 204168 998436 204220 998442
rect 204168 998378 204220 998384
rect 203524 998232 203576 998238
rect 203522 998200 203524 998209
rect 203576 998200 203578 998209
rect 203522 998135 203578 998144
rect 202696 998096 202748 998102
rect 202694 998064 202696 998073
rect 202748 998064 202750 998073
rect 202694 997999 202750 998008
rect 204720 997824 204772 997830
rect 204718 997792 204720 997801
rect 204772 997792 204774 997801
rect 204718 997727 204774 997736
rect 202512 995988 202564 995994
rect 202512 995930 202564 995936
rect 202326 995888 202382 995897
rect 202326 995823 202382 995832
rect 203614 995888 203670 995897
rect 203614 995823 203670 995832
rect 202144 995376 202196 995382
rect 203628 995353 203656 995823
rect 202144 995318 202196 995324
rect 203614 995344 203670 995353
rect 203614 995279 203670 995288
rect 199382 993984 199438 993993
rect 199382 993919 199438 993928
rect 197544 993676 197596 993682
rect 197544 993618 197596 993624
rect 188160 993540 188212 993546
rect 188160 993482 188212 993488
rect 195888 993540 195940 993546
rect 195888 993482 195940 993488
rect 186502 992896 186558 992905
rect 186502 992831 186558 992840
rect 164884 990888 164936 990894
rect 164884 990830 164936 990836
rect 170772 990888 170824 990894
rect 170772 990830 170824 990836
rect 154488 985720 154540 985726
rect 154488 985662 154540 985668
rect 160744 985720 160796 985726
rect 160744 985662 160796 985668
rect 154500 983620 154528 985662
rect 170784 983620 170812 990830
rect 186516 983634 186544 992831
rect 204916 986678 204944 1005246
rect 212078 1005207 212134 1005216
rect 209226 1005000 209282 1005009
rect 209226 1004935 209228 1004944
rect 209280 1004935 209282 1004944
rect 211804 1004964 211856 1004970
rect 209228 1004906 209280 1004912
rect 211804 1004906 211856 1004912
rect 211250 1004864 211306 1004873
rect 211250 1004799 211252 1004808
rect 211304 1004799 211306 1004808
rect 211252 1004770 211304 1004776
rect 209226 1004728 209282 1004737
rect 209226 1004663 209228 1004672
rect 209280 1004663 209282 1004672
rect 211160 1004692 211212 1004698
rect 209228 1004634 209280 1004640
rect 211160 1004634 211212 1004640
rect 206374 1002552 206430 1002561
rect 206374 1002487 206376 1002496
rect 206428 1002487 206430 1002496
rect 206376 1002458 206428 1002464
rect 207202 1002280 207258 1002289
rect 205088 1002244 205140 1002250
rect 207202 1002215 207204 1002224
rect 205088 1002186 205140 1002192
rect 207256 1002215 207258 1002224
rect 207204 1002186 207256 1002192
rect 205100 997286 205128 1002186
rect 206742 1002144 206798 1002153
rect 210882 1002144 210938 1002153
rect 206742 1002079 206744 1002088
rect 206796 1002079 206798 1002088
rect 208584 1002108 208636 1002114
rect 206744 1002050 206796 1002056
rect 210882 1002079 210884 1002088
rect 208584 1002050 208636 1002056
rect 210936 1002079 210938 1002088
rect 210884 1002050 210936 1002056
rect 205546 1002008 205602 1002017
rect 207202 1002008 207258 1002017
rect 205546 1001943 205548 1001952
rect 205600 1001943 205602 1001952
rect 206284 1001972 206336 1001978
rect 205548 1001914 205600 1001920
rect 206284 1001914 206336 1001920
rect 207032 1001966 207202 1001994
rect 205548 997960 205600 997966
rect 205546 997928 205548 997937
rect 205600 997928 205602 997937
rect 205546 997863 205602 997872
rect 205088 997280 205140 997286
rect 205088 997222 205140 997228
rect 206296 994974 206324 1001914
rect 207032 995110 207060 1001966
rect 207202 1001943 207258 1001952
rect 207570 1002008 207626 1002017
rect 207570 1001943 207572 1001952
rect 207624 1001943 207626 1001952
rect 207572 1001914 207624 1001920
rect 208398 995888 208454 995897
rect 208398 995823 208454 995832
rect 207020 995104 207072 995110
rect 208412 995081 208440 995823
rect 208596 995246 208624 1002050
rect 211172 996130 211200 1004634
rect 211160 996124 211212 996130
rect 211160 996066 211212 996072
rect 211816 995858 211844 1004906
rect 215944 1004828 215996 1004834
rect 215944 1004770 215996 1004776
rect 213184 1002108 213236 1002114
rect 213184 1002050 213236 1002056
rect 212538 1002008 212594 1002017
rect 212538 1001943 212540 1001952
rect 212592 1001943 212594 1001952
rect 212540 1001914 212592 1001920
rect 213196 995994 213224 1002050
rect 214564 1001972 214616 1001978
rect 214564 1001914 214616 1001920
rect 213184 995988 213236 995994
rect 213184 995930 213236 995936
rect 211804 995852 211856 995858
rect 211804 995794 211856 995800
rect 208584 995240 208636 995246
rect 208584 995182 208636 995188
rect 207020 995046 207072 995052
rect 208398 995072 208454 995081
rect 208398 995007 208454 995016
rect 206284 994968 206336 994974
rect 206284 994910 206336 994916
rect 214576 991234 214604 1001914
rect 214564 991228 214616 991234
rect 214564 991170 214616 991176
rect 203156 986672 203208 986678
rect 203156 986614 203208 986620
rect 204904 986672 204956 986678
rect 204904 986614 204956 986620
rect 186516 983606 186990 983634
rect 203168 983620 203196 986614
rect 215956 985998 215984 1004770
rect 226340 997076 226392 997082
rect 226340 997018 226392 997024
rect 226352 994294 226380 997018
rect 228376 995081 228404 1006130
rect 229744 1006052 229796 1006058
rect 229744 1005994 229796 1006000
rect 229756 996130 229784 1005994
rect 247132 1003944 247184 1003950
rect 247132 1003886 247184 1003892
rect 246580 1002584 246632 1002590
rect 246580 1002526 246632 1002532
rect 246592 998073 246620 1002526
rect 246948 999796 247000 999802
rect 246948 999738 247000 999744
rect 246764 998368 246816 998374
rect 246764 998310 246816 998316
rect 246578 998064 246634 998073
rect 246578 997999 246634 998008
rect 246776 997754 246804 998310
rect 246776 997726 246896 997754
rect 246672 997688 246724 997694
rect 246672 997630 246724 997636
rect 246684 996441 246712 997630
rect 246670 996432 246726 996441
rect 246670 996367 246726 996376
rect 229744 996124 229796 996130
rect 229744 996066 229796 996072
rect 246670 996024 246726 996033
rect 246868 996010 246896 997726
rect 246726 995982 246896 996010
rect 246670 995959 246726 995968
rect 246960 995761 246988 999738
rect 247144 996713 247172 1003886
rect 247316 998504 247368 998510
rect 247316 998446 247368 998452
rect 247130 996704 247186 996713
rect 247130 996639 247186 996648
rect 238574 995752 238630 995761
rect 239586 995752 239642 995761
rect 238630 995710 238740 995738
rect 239292 995710 239586 995738
rect 238574 995687 238630 995696
rect 240230 995752 240286 995761
rect 239936 995710 240230 995738
rect 239586 995687 239642 995696
rect 240874 995752 240930 995761
rect 240580 995710 240874 995738
rect 240230 995687 240286 995696
rect 243818 995752 243874 995761
rect 243616 995710 243818 995738
rect 240874 995687 240930 995696
rect 243818 995687 243874 995696
rect 244094 995752 244150 995761
rect 245566 995752 245622 995761
rect 244150 995710 244260 995738
rect 245456 995710 245566 995738
rect 244094 995687 244150 995696
rect 245566 995687 245622 995696
rect 246946 995752 247002 995761
rect 246946 995687 247002 995696
rect 247130 995752 247186 995761
rect 247130 995687 247186 995696
rect 247144 995518 247172 995687
rect 246212 995512 246264 995518
rect 231288 995438 231624 995466
rect 231932 995438 232268 995466
rect 232576 995438 232912 995466
rect 231596 995110 231624 995438
rect 231584 995104 231636 995110
rect 228362 995072 228418 995081
rect 231584 995046 231636 995052
rect 228362 995007 228418 995016
rect 226340 994288 226392 994294
rect 226340 994230 226392 994236
rect 232240 994022 232268 995438
rect 232884 994974 232912 995438
rect 234402 995246 234430 995452
rect 234968 995438 235304 995466
rect 235612 995438 235948 995466
rect 236256 995438 236592 995466
rect 241776 995438 242112 995466
rect 242972 995438 243308 995466
rect 246212 995454 246264 995460
rect 247132 995512 247184 995518
rect 247132 995454 247184 995460
rect 234390 995240 234442 995246
rect 234390 995182 234442 995188
rect 232872 994968 232924 994974
rect 232872 994910 232924 994916
rect 235276 994537 235304 995438
rect 235262 994528 235318 994537
rect 235262 994463 235318 994472
rect 235920 994265 235948 995438
rect 236564 995382 236592 995438
rect 236552 995376 236604 995382
rect 242084 995353 242112 995438
rect 236552 995318 236604 995324
rect 242070 995344 242126 995353
rect 242070 995279 242126 995288
rect 243280 994809 243308 995438
rect 245014 995344 245070 995353
rect 246224 995330 246252 995454
rect 245070 995302 246252 995330
rect 245014 995279 245070 995288
rect 247328 994809 247356 998446
rect 243266 994800 243322 994809
rect 243266 994735 243322 994744
rect 247314 994800 247370 994809
rect 247314 994735 247370 994744
rect 247696 994265 247724 1006402
rect 258998 1006360 259054 1006369
rect 255964 1006324 256016 1006330
rect 307758 1006360 307814 1006369
rect 258998 1006295 259000 1006304
rect 255964 1006266 256016 1006272
rect 259052 1006295 259054 1006304
rect 301504 1006324 301556 1006330
rect 259000 1006266 259052 1006272
rect 307758 1006295 307760 1006304
rect 301504 1006266 301556 1006272
rect 307812 1006295 307814 1006304
rect 314658 1006360 314714 1006369
rect 361394 1006360 361450 1006369
rect 314658 1006295 314660 1006304
rect 307760 1006266 307812 1006272
rect 314712 1006295 314714 1006304
rect 320824 1006324 320876 1006330
rect 314660 1006266 314712 1006272
rect 361394 1006295 361396 1006304
rect 320824 1006266 320876 1006272
rect 361448 1006295 361450 1006304
rect 361396 1006266 361448 1006272
rect 249064 1006188 249116 1006194
rect 249064 1006130 249116 1006136
rect 247868 997824 247920 997830
rect 247868 997766 247920 997772
rect 235906 994256 235962 994265
rect 235906 994191 235962 994200
rect 247682 994256 247738 994265
rect 247682 994191 247738 994200
rect 247880 994158 247908 997766
rect 249076 997257 249104 1006130
rect 252466 1006088 252522 1006097
rect 252466 1006023 252522 1006032
rect 251824 1002380 251876 1002386
rect 251824 1002322 251876 1002328
rect 250444 998164 250496 998170
rect 250444 998106 250496 998112
rect 249062 997248 249118 997257
rect 249062 997183 249118 997192
rect 250456 994634 250484 998106
rect 251180 997960 251232 997966
rect 251180 997902 251232 997908
rect 251192 995489 251220 997902
rect 251178 995480 251234 995489
rect 251178 995415 251234 995424
rect 251836 995382 251864 1002322
rect 252480 998374 252508 1006023
rect 255320 1003944 255372 1003950
rect 255318 1003912 255320 1003921
rect 255372 1003912 255374 1003921
rect 255318 1003847 255374 1003856
rect 253112 1002720 253164 1002726
rect 253112 1002662 253164 1002668
rect 252468 998368 252520 998374
rect 252468 998310 252520 998316
rect 252468 997824 252520 997830
rect 252466 997792 252468 997801
rect 252520 997792 252522 997801
rect 252466 997727 252522 997736
rect 251824 995376 251876 995382
rect 251824 995318 251876 995324
rect 250444 994628 250496 994634
rect 250444 994570 250496 994576
rect 253124 994537 253152 1002662
rect 254124 1002584 254176 1002590
rect 254122 1002552 254124 1002561
rect 254176 1002552 254178 1002561
rect 254122 1002487 254178 1002496
rect 254490 1002416 254546 1002425
rect 254490 1002351 254492 1002360
rect 254544 1002351 254546 1002360
rect 254492 1002322 254544 1002328
rect 254584 1002244 254636 1002250
rect 254584 1002186 254636 1002192
rect 253388 1002108 253440 1002114
rect 253388 1002050 253440 1002056
rect 253400 995761 253428 1002050
rect 253662 998200 253718 998209
rect 253662 998135 253664 998144
rect 253716 998135 253718 998144
rect 253664 998106 253716 998112
rect 253664 997960 253716 997966
rect 253662 997928 253664 997937
rect 253716 997928 253718 997937
rect 253662 997863 253718 997872
rect 253386 995752 253442 995761
rect 253386 995687 253442 995696
rect 253110 994528 253166 994537
rect 253110 994463 253166 994472
rect 251456 994288 251508 994294
rect 251456 994230 251508 994236
rect 247868 994152 247920 994158
rect 247868 994094 247920 994100
rect 232228 994016 232280 994022
rect 232228 993958 232280 993964
rect 219440 991228 219492 991234
rect 219440 991170 219492 991176
rect 215944 985992 215996 985998
rect 215944 985934 215996 985940
rect 219452 983620 219480 991170
rect 235632 985992 235684 985998
rect 235632 985934 235684 985940
rect 235644 983620 235672 985934
rect 251468 983634 251496 994230
rect 254596 994022 254624 1002186
rect 255318 1002144 255374 1002153
rect 255318 1002079 255320 1002088
rect 255372 1002079 255374 1002088
rect 255320 1002050 255372 1002056
rect 254768 1001972 254820 1001978
rect 254768 1001914 254820 1001920
rect 254780 999802 254808 1001914
rect 254768 999796 254820 999802
rect 254768 999738 254820 999744
rect 255976 994974 256004 1006266
rect 257342 1006224 257398 1006233
rect 257342 1006159 257344 1006168
rect 257396 1006159 257398 1006168
rect 262678 1006224 262734 1006233
rect 262678 1006159 262680 1006168
rect 257344 1006130 257396 1006136
rect 262732 1006159 262734 1006168
rect 269764 1006188 269816 1006194
rect 262680 1006130 262732 1006136
rect 269764 1006130 269816 1006136
rect 298744 1006188 298796 1006194
rect 298744 1006130 298796 1006136
rect 258170 1006088 258226 1006097
rect 257344 1006052 257396 1006058
rect 258170 1006023 258172 1006032
rect 257344 1005994 257396 1006000
rect 258224 1006023 258226 1006032
rect 261850 1006088 261906 1006097
rect 261850 1006023 261852 1006032
rect 258172 1005994 258224 1006000
rect 261904 1006023 261906 1006032
rect 261852 1005994 261904 1006000
rect 256148 1002720 256200 1002726
rect 256146 1002688 256148 1002697
rect 256200 1002688 256202 1002697
rect 256146 1002623 256202 1002632
rect 256514 1002280 256570 1002289
rect 256514 1002215 256516 1002224
rect 256568 1002215 256570 1002224
rect 256516 1002186 256568 1002192
rect 256974 1002008 257030 1002017
rect 256974 1001943 256976 1001952
rect 257028 1001943 257030 1001952
rect 256976 1001914 257028 1001920
rect 257356 995110 257384 1005994
rect 263046 1005000 263102 1005009
rect 263046 1004935 263048 1004944
rect 263100 1004935 263102 1004944
rect 268384 1004964 268436 1004970
rect 263048 1004906 263100 1004912
rect 268384 1004906 268436 1004912
rect 258170 1004864 258226 1004873
rect 258170 1004799 258172 1004808
rect 258224 1004799 258226 1004808
rect 259460 1004828 259512 1004834
rect 258172 1004770 258224 1004776
rect 259460 1004770 259512 1004776
rect 258998 1002008 259054 1002017
rect 258092 1001966 258998 1001994
rect 258092 997694 258120 1001966
rect 258998 1001943 259054 1001952
rect 258080 997688 258132 997694
rect 258080 997630 258132 997636
rect 259472 995246 259500 1004770
rect 261022 1002416 261078 1002425
rect 261022 1002351 261024 1002360
rect 261076 1002351 261078 1002360
rect 264244 1002380 264296 1002386
rect 261024 1002322 261076 1002328
rect 264244 1002322 264296 1002328
rect 260194 1002280 260250 1002289
rect 260194 1002215 260196 1002224
rect 260248 1002215 260250 1002224
rect 262864 1002244 262916 1002250
rect 260196 1002186 260248 1002192
rect 262864 1002186 262916 1002192
rect 259826 1002144 259882 1002153
rect 259826 1002079 259828 1002088
rect 259880 1002079 259882 1002088
rect 262220 1002108 262272 1002114
rect 259828 1002050 259880 1002056
rect 262220 1002050 262272 1002056
rect 260194 1002008 260250 1002017
rect 261850 1002008 261906 1002017
rect 260194 1001943 260196 1001952
rect 260248 1001943 260250 1001952
rect 260932 1001972 260984 1001978
rect 260196 1001914 260248 1001920
rect 260932 1001914 260984 1001920
rect 261128 1001966 261850 1001994
rect 260944 995858 260972 1001914
rect 261128 995994 261156 1001966
rect 261850 1001943 261906 1001952
rect 262232 996130 262260 1002050
rect 262876 996334 262904 1002186
rect 263874 1002144 263930 1002153
rect 263874 1002079 263876 1002088
rect 263928 1002079 263930 1002088
rect 263876 1002050 263928 1002056
rect 263506 1002008 263562 1002017
rect 263506 1001943 263508 1001952
rect 263560 1001943 263562 1001952
rect 263508 1001914 263560 1001920
rect 262864 996328 262916 996334
rect 262864 996270 262916 996276
rect 262220 996124 262272 996130
rect 262220 996066 262272 996072
rect 264256 995994 264284 1002322
rect 267004 1002108 267056 1002114
rect 267004 1002050 267056 1002056
rect 265624 1001972 265676 1001978
rect 265624 1001914 265676 1001920
rect 261116 995988 261168 995994
rect 261116 995930 261168 995936
rect 264244 995988 264296 995994
rect 264244 995930 264296 995936
rect 260932 995852 260984 995858
rect 260932 995794 260984 995800
rect 259460 995240 259512 995246
rect 259460 995182 259512 995188
rect 257344 995104 257396 995110
rect 257344 995046 257396 995052
rect 255964 994968 256016 994974
rect 255964 994910 256016 994916
rect 254584 994016 254636 994022
rect 254584 993958 254636 993964
rect 265636 990894 265664 1001914
rect 267016 991506 267044 1002050
rect 267004 991500 267056 991506
rect 267004 991442 267056 991448
rect 265624 990888 265676 990894
rect 265624 990830 265676 990836
rect 267648 990888 267700 990894
rect 267648 990830 267700 990836
rect 267660 985334 267688 990830
rect 268396 985998 268424 1004906
rect 269776 996130 269804 1006130
rect 279424 1006052 279476 1006058
rect 279424 1005994 279476 1006000
rect 278228 997824 278280 997830
rect 278228 997766 278280 997772
rect 270408 996328 270460 996334
rect 270408 996270 270460 996276
rect 269764 996124 269816 996130
rect 269764 996066 269816 996072
rect 270420 995081 270448 996270
rect 270406 995072 270462 995081
rect 270406 995007 270462 995016
rect 278240 994294 278268 997766
rect 279436 995353 279464 1005994
rect 298282 1002280 298338 1002289
rect 298282 1002215 298338 1002224
rect 298098 997792 298154 997801
rect 298098 997727 298154 997736
rect 282734 995752 282790 995761
rect 288070 995752 288126 995761
rect 282790 995710 282854 995738
rect 287822 995710 288070 995738
rect 282734 995687 282790 995696
rect 291106 995752 291162 995761
rect 290858 995710 291106 995738
rect 288070 995687 288126 995696
rect 291106 995687 291162 995696
rect 297824 995580 297876 995586
rect 297824 995522 297876 995528
rect 279422 995344 279478 995353
rect 279422 995279 279478 995288
rect 283484 994634 283512 995452
rect 284128 995110 284156 995452
rect 285968 995246 285996 995452
rect 285956 995240 286008 995246
rect 285956 995182 286008 995188
rect 284116 995104 284168 995110
rect 284116 995046 284168 995052
rect 283472 994628 283524 994634
rect 283472 994570 283524 994576
rect 286520 994537 286548 995452
rect 287164 994974 287192 995452
rect 290306 995438 290780 995466
rect 291502 995438 291792 995466
rect 287152 994968 287204 994974
rect 287152 994910 287204 994916
rect 290752 994809 290780 995438
rect 290738 994800 290794 994809
rect 290738 994735 290794 994744
rect 286506 994528 286562 994537
rect 286506 994463 286562 994472
rect 278228 994288 278280 994294
rect 278228 994230 278280 994236
rect 291764 993993 291792 995438
rect 292132 994265 292160 995452
rect 293342 995438 293632 995466
rect 294538 995438 294828 995466
rect 293604 995382 293632 995438
rect 293592 995376 293644 995382
rect 293592 995318 293644 995324
rect 294800 994809 294828 995438
rect 295168 995330 295196 995452
rect 295826 995438 296208 995466
rect 297022 995438 297404 995466
rect 296180 995382 296208 995438
rect 295984 995376 296036 995382
rect 295168 995302 295288 995330
rect 295984 995318 296036 995324
rect 296168 995376 296220 995382
rect 296168 995318 296220 995324
rect 297376 995330 297404 995438
rect 297836 995330 297864 995522
rect 298112 995382 298140 997727
rect 295260 994809 295288 995302
rect 295996 995194 296024 995318
rect 297376 995302 297864 995330
rect 298100 995376 298152 995382
rect 298100 995318 298152 995324
rect 298296 995194 298324 1002215
rect 298756 1001894 298784 1006130
rect 298928 1006052 298980 1006058
rect 298928 1005994 298980 1006000
rect 298664 1001866 298784 1001894
rect 298940 1001894 298968 1005994
rect 300308 1003332 300360 1003338
rect 300308 1003274 300360 1003280
rect 299296 1003196 299348 1003202
rect 299296 1003138 299348 1003144
rect 298940 1001866 299152 1001894
rect 298468 1000544 298520 1000550
rect 298468 1000486 298520 1000492
rect 298480 995586 298508 1000486
rect 298664 997778 298692 1001866
rect 298572 997750 298692 997778
rect 298836 997756 298888 997762
rect 298572 996554 298600 997750
rect 298836 997698 298888 997704
rect 298848 996713 298876 997698
rect 298834 996704 298890 996713
rect 298834 996639 298890 996648
rect 298572 996526 298876 996554
rect 298650 996432 298706 996441
rect 298650 996367 298652 996376
rect 298704 996367 298706 996376
rect 298652 996338 298704 996344
rect 298468 995580 298520 995586
rect 298468 995522 298520 995528
rect 295996 995166 298324 995194
rect 294786 994800 294842 994809
rect 295246 994800 295302 994809
rect 294786 994735 294842 994744
rect 295064 994764 295116 994770
rect 295246 994735 295302 994744
rect 295064 994706 295116 994712
rect 292118 994256 292174 994265
rect 292118 994191 292174 994200
rect 295076 994158 295104 994706
rect 298848 994498 298876 996526
rect 299124 996010 299152 1001866
rect 299308 996985 299336 1003138
rect 300124 1002108 300176 1002114
rect 300124 1002050 300176 1002056
rect 299480 997620 299532 997626
rect 299480 997562 299532 997568
rect 299492 997257 299520 997562
rect 299478 997248 299534 997257
rect 299478 997183 299534 997192
rect 299294 996976 299350 996985
rect 299294 996911 299350 996920
rect 299124 995994 299244 996010
rect 299124 995988 299256 995994
rect 299124 995982 299204 995988
rect 299204 995930 299256 995936
rect 298836 994492 298888 994498
rect 298836 994434 298888 994440
rect 300136 994158 300164 1002050
rect 300320 994265 300348 1003274
rect 301516 994537 301544 1006266
rect 304906 1006224 304962 1006233
rect 304906 1006159 304908 1006168
rect 304960 1006159 304962 1006168
rect 304908 1006130 304960 1006136
rect 301686 1006088 301742 1006097
rect 301686 1006023 301742 1006032
rect 303250 1006088 303306 1006097
rect 303250 1006023 303252 1006032
rect 301700 997801 301728 1006023
rect 303304 1006023 303306 1006032
rect 304078 1006088 304134 1006097
rect 304078 1006023 304080 1006032
rect 303252 1005994 303304 1006000
rect 304132 1006023 304134 1006032
rect 311806 1006088 311862 1006097
rect 311806 1006023 311808 1006032
rect 304080 1005994 304132 1006000
rect 311860 1006023 311862 1006032
rect 314658 1006088 314714 1006097
rect 314658 1006023 314660 1006032
rect 311808 1005994 311860 1006000
rect 314712 1006023 314714 1006032
rect 319444 1006052 319496 1006058
rect 314660 1005994 314712 1006000
rect 319444 1005994 319496 1006000
rect 307298 1005272 307354 1005281
rect 304264 1005236 304316 1005242
rect 307298 1005207 307300 1005216
rect 304264 1005178 304316 1005184
rect 307352 1005207 307354 1005216
rect 307300 1005178 307352 1005184
rect 303620 1004964 303672 1004970
rect 303620 1004906 303672 1004912
rect 303250 1002280 303306 1002289
rect 303068 1002244 303120 1002250
rect 303632 1002266 303660 1004906
rect 303306 1002238 303660 1002266
rect 303250 1002215 303306 1002224
rect 303068 1002186 303120 1002192
rect 302884 1001972 302936 1001978
rect 302884 1001914 302936 1001920
rect 301686 997792 301742 997801
rect 301686 997727 301742 997736
rect 302896 996169 302924 1001914
rect 302882 996160 302938 996169
rect 302882 996095 302938 996104
rect 303080 995897 303108 1002186
rect 304078 1002144 304134 1002153
rect 304078 1002079 304080 1002088
rect 304132 1002079 304134 1002088
rect 304080 1002050 304132 1002056
rect 303066 995888 303122 995897
rect 303066 995823 303122 995832
rect 304276 994974 304304 1005178
rect 306930 1005000 306986 1005009
rect 306930 1004935 306932 1004944
rect 306984 1004935 306986 1004944
rect 306932 1004906 306984 1004912
rect 308954 1004864 309010 1004873
rect 305828 1004828 305880 1004834
rect 308954 1004799 308956 1004808
rect 305828 1004770 305880 1004776
rect 309008 1004799 309010 1004808
rect 313830 1004864 313886 1004873
rect 313830 1004799 313832 1004808
rect 308956 1004770 309008 1004776
rect 313884 1004799 313886 1004808
rect 316040 1004828 316092 1004834
rect 313832 1004770 313884 1004776
rect 316040 1004770 316092 1004776
rect 305644 1004692 305696 1004698
rect 305644 1004634 305696 1004640
rect 305274 1003368 305330 1003377
rect 305274 1003303 305276 1003312
rect 305328 1003303 305330 1003312
rect 305276 1003274 305328 1003280
rect 304264 994968 304316 994974
rect 304264 994910 304316 994916
rect 305656 994634 305684 1004634
rect 305840 1000550 305868 1004770
rect 308126 1004728 308182 1004737
rect 308126 1004663 308128 1004672
rect 308180 1004663 308182 1004672
rect 315486 1004728 315542 1004737
rect 315486 1004663 315488 1004672
rect 308128 1004634 308180 1004640
rect 315540 1004663 315542 1004672
rect 315488 1004634 315540 1004640
rect 308954 1003232 309010 1003241
rect 308954 1003167 308956 1003176
rect 309008 1003167 309010 1003176
rect 308956 1003138 309008 1003144
rect 310610 1002552 310666 1002561
rect 310610 1002487 310666 1002496
rect 310624 1002402 310652 1002487
rect 310440 1002374 310652 1002402
rect 306102 1002280 306158 1002289
rect 306102 1002215 306104 1002224
rect 306156 1002215 306158 1002224
rect 308404 1002244 308456 1002250
rect 306104 1002186 306156 1002192
rect 308404 1002186 308456 1002192
rect 306102 1002008 306158 1002017
rect 306930 1002008 306986 1002017
rect 306102 1001943 306104 1001952
rect 306156 1001943 306158 1001952
rect 306392 1001966 306930 1001994
rect 306104 1001914 306156 1001920
rect 305828 1000544 305880 1000550
rect 305828 1000486 305880 1000492
rect 305644 994628 305696 994634
rect 305644 994570 305696 994576
rect 301502 994528 301558 994537
rect 301502 994463 301558 994472
rect 306392 994265 306420 1001966
rect 306930 1001943 306986 1001952
rect 308416 995110 308444 1002186
rect 309782 1002008 309838 1002017
rect 309152 1001966 309782 1001994
rect 308770 995616 308826 995625
rect 308770 995551 308826 995560
rect 308404 995104 308456 995110
rect 308784 995081 308812 995551
rect 309152 995246 309180 1001966
rect 309782 1001943 309838 1001952
rect 310150 1002008 310206 1002017
rect 310150 1001943 310152 1001952
rect 310204 1001943 310206 1001952
rect 310152 1001914 310204 1001920
rect 310440 1001894 310468 1002374
rect 310610 1002280 310666 1002289
rect 310610 1002215 310612 1002224
rect 310664 1002215 310666 1002224
rect 310612 1002186 310664 1002192
rect 311900 1001972 311952 1001978
rect 311900 1001914 311952 1001920
rect 310440 1001866 310560 1001894
rect 310532 997626 310560 1001866
rect 311912 997762 311940 1001914
rect 311900 997756 311952 997762
rect 311900 997698 311952 997704
rect 310520 997620 310572 997626
rect 310520 997562 310572 997568
rect 316052 996130 316080 1004770
rect 318064 1004692 318116 1004698
rect 318064 1004634 318116 1004640
rect 316040 996124 316092 996130
rect 316040 996066 316092 996072
rect 309140 995240 309192 995246
rect 309140 995182 309192 995188
rect 308404 995046 308456 995052
rect 308770 995072 308826 995081
rect 308770 995007 308826 995016
rect 316408 994288 316460 994294
rect 300306 994256 300362 994265
rect 300306 994191 300362 994200
rect 306378 994256 306434 994265
rect 316408 994230 316460 994236
rect 306378 994191 306434 994200
rect 295064 994152 295116 994158
rect 295064 994094 295116 994100
rect 300124 994152 300176 994158
rect 300124 994094 300176 994100
rect 291750 993984 291806 993993
rect 291750 993919 291806 993928
rect 284300 991500 284352 991506
rect 284300 991442 284352 991448
rect 268384 985992 268436 985998
rect 268384 985934 268436 985940
rect 267660 985306 267780 985334
rect 267752 983634 267780 985306
rect 251468 983606 251850 983634
rect 267752 983606 268134 983634
rect 284312 983620 284340 991442
rect 300492 985992 300544 985998
rect 300492 985934 300544 985940
rect 300504 983620 300532 985934
rect 316420 983634 316448 994230
rect 318076 993070 318104 1004634
rect 318064 993064 318116 993070
rect 318064 993006 318116 993012
rect 319456 992934 319484 1005994
rect 320836 997082 320864 1006266
rect 360566 1006224 360622 1006233
rect 360566 1006159 360568 1006168
rect 360620 1006159 360622 1006168
rect 363418 1006224 363474 1006233
rect 363418 1006159 363420 1006168
rect 360568 1006130 360620 1006136
rect 363472 1006159 363474 1006168
rect 363420 1006130 363472 1006136
rect 358542 1006088 358598 1006097
rect 358542 1006023 358544 1006032
rect 358596 1006023 358598 1006032
rect 362224 1006052 362276 1006058
rect 358544 1005994 358596 1006000
rect 362224 1005994 362276 1006000
rect 360568 1005440 360620 1005446
rect 360566 1005408 360568 1005417
rect 360620 1005408 360622 1005417
rect 360566 1005343 360622 1005352
rect 355692 1005304 355744 1005310
rect 355690 1005272 355692 1005281
rect 355744 1005272 355746 1005281
rect 355690 1005207 355746 1005216
rect 356518 1005000 356574 1005009
rect 354588 1004964 354640 1004970
rect 356518 1004935 356520 1004944
rect 354588 1004906 354640 1004912
rect 356572 1004935 356574 1004944
rect 361394 1005000 361450 1005009
rect 361394 1004935 361396 1004944
rect 356520 1004906 356572 1004912
rect 361448 1004935 361450 1004944
rect 361396 1004906 361448 1004912
rect 353208 1004828 353260 1004834
rect 353208 1004770 353260 1004776
rect 351828 1001972 351880 1001978
rect 351828 1001914 351880 1001920
rect 351840 998714 351868 1001914
rect 353220 1001230 353248 1004770
rect 354034 1002008 354090 1002017
rect 354034 1001943 354036 1001952
rect 354088 1001943 354090 1001952
rect 354036 1001914 354088 1001920
rect 353208 1001224 353260 1001230
rect 353208 1001166 353260 1001172
rect 351828 998708 351880 998714
rect 351828 998650 351880 998656
rect 354600 998442 354628 1004906
rect 355690 1004864 355746 1004873
rect 355690 1004799 355692 1004808
rect 355744 1004799 355746 1004808
rect 355692 1004770 355744 1004776
rect 357714 1002416 357770 1002425
rect 357714 1002351 357716 1002360
rect 357768 1002351 357770 1002360
rect 360844 1002380 360896 1002386
rect 357716 1002322 357768 1002328
rect 360844 1002322 360896 1002328
rect 357714 1002144 357770 1002153
rect 355784 1002108 355836 1002114
rect 357714 1002079 357716 1002088
rect 355784 1002050 355836 1002056
rect 357768 1002079 357770 1002088
rect 357716 1002050 357768 1002056
rect 355796 998578 355824 1002050
rect 356518 1002008 356574 1002017
rect 356072 1001966 356518 1001994
rect 356072 998850 356100 1001966
rect 356518 1001943 356574 1001952
rect 357346 1002008 357402 1002017
rect 359370 1002008 359426 1002017
rect 357402 1001966 358124 1001994
rect 357346 1001943 357402 1001952
rect 356060 998844 356112 998850
rect 356060 998786 356112 998792
rect 355784 998572 355836 998578
rect 355784 998514 355836 998520
rect 354588 998436 354640 998442
rect 354588 998378 354640 998384
rect 320824 997076 320876 997082
rect 320824 997018 320876 997024
rect 332600 997076 332652 997082
rect 332600 997018 332652 997024
rect 319444 992928 319496 992934
rect 319444 992870 319496 992876
rect 332612 983634 332640 997018
rect 358096 995042 358124 1001966
rect 358832 1001966 359370 1001994
rect 358832 997762 358860 1001966
rect 359370 1001943 359426 1001952
rect 358820 997756 358872 997762
rect 358820 997698 358872 997704
rect 360856 995858 360884 1002322
rect 360844 995852 360896 995858
rect 360844 995794 360896 995800
rect 362236 995178 362264 1005994
rect 362590 1004864 362646 1004873
rect 362590 1004799 362592 1004808
rect 362644 1004799 362646 1004808
rect 362592 1004770 362644 1004776
rect 362224 995172 362276 995178
rect 362224 995114 362276 995120
rect 358084 995036 358136 995042
rect 358084 994978 358136 994984
rect 363616 994906 363644 1006402
rect 364904 1006058 364932 1006538
rect 365074 1006088 365130 1006097
rect 364892 1006052 364944 1006058
rect 365074 1006023 365076 1006032
rect 364892 1005994 364944 1006000
rect 365128 1006023 365130 1006032
rect 367744 1006052 367796 1006058
rect 365076 1005994 365128 1006000
rect 367744 1005994 367796 1006000
rect 365074 1005136 365130 1005145
rect 365074 1005071 365076 1005080
rect 365128 1005071 365130 1005080
rect 365076 1005042 365128 1005048
rect 364984 1004964 365036 1004970
rect 364984 1004906 365036 1004912
rect 364246 1004728 364302 1004737
rect 364246 1004663 364248 1004672
rect 364300 1004663 364302 1004672
rect 364248 1004634 364300 1004640
rect 364996 995994 365024 1004906
rect 365168 1004828 365220 1004834
rect 365168 1004770 365220 1004776
rect 365180 997626 365208 1004770
rect 366364 1004692 366416 1004698
rect 366364 1004634 366416 1004640
rect 365902 1002008 365958 1002017
rect 365902 1001943 365904 1001952
rect 365956 1001943 365958 1001952
rect 365904 1001914 365956 1001920
rect 365168 997620 365220 997626
rect 365168 997562 365220 997568
rect 365168 996396 365220 996402
rect 365168 996338 365220 996344
rect 364984 995988 365036 995994
rect 364984 995930 365036 995936
rect 363604 994900 363656 994906
rect 363604 994842 363656 994848
rect 365180 994294 365208 996338
rect 366376 996130 366404 1004634
rect 366364 996124 366416 996130
rect 366364 996066 366416 996072
rect 365168 994288 365220 994294
rect 365168 994230 365220 994236
rect 349160 993064 349212 993070
rect 349160 993006 349212 993012
rect 316420 983606 316802 983634
rect 332612 983606 332994 983634
rect 349172 983620 349200 993006
rect 364984 992928 365036 992934
rect 364984 992870 365036 992876
rect 364996 983634 365024 992870
rect 367756 991506 367784 1005994
rect 370504 1005100 370556 1005106
rect 370504 1005042 370556 1005048
rect 369124 1001972 369176 1001978
rect 369124 1001914 369176 1001920
rect 369136 991642 369164 1001914
rect 369124 991636 369176 991642
rect 369124 991578 369176 991584
rect 367744 991500 367796 991506
rect 367744 991442 367796 991448
rect 370516 985998 370544 1005042
rect 371896 998306 371924 1006538
rect 373276 998850 373304 1006946
rect 380164 1006868 380216 1006874
rect 380164 1006810 380216 1006816
rect 374644 1006460 374696 1006466
rect 374644 1006402 374696 1006408
rect 372160 998844 372212 998850
rect 372160 998786 372212 998792
rect 373264 998844 373316 998850
rect 373264 998786 373316 998792
rect 371884 998300 371936 998306
rect 371884 998242 371936 998248
rect 372172 996010 372200 998786
rect 372988 998300 373040 998306
rect 372988 998242 373040 998248
rect 372344 997756 372396 997762
rect 372344 997698 372396 997704
rect 372356 996441 372384 997698
rect 372528 997620 372580 997626
rect 372528 997562 372580 997568
rect 372540 996985 372568 997562
rect 372526 996976 372582 996985
rect 372526 996911 372582 996920
rect 372342 996432 372398 996441
rect 372342 996367 372398 996376
rect 372342 996024 372398 996033
rect 372172 995982 372342 996010
rect 372342 995959 372398 995968
rect 373000 994634 373028 998242
rect 374656 997801 374684 1006402
rect 377404 1006188 377456 1006194
rect 377404 1006130 377456 1006136
rect 376024 1005304 376076 1005310
rect 376024 1005246 376076 1005252
rect 374642 997792 374698 997801
rect 374642 997727 374698 997736
rect 376036 994770 376064 1005246
rect 377416 997830 377444 1006130
rect 378784 1005440 378836 1005446
rect 378784 1005382 378836 1005388
rect 378796 998782 378824 1005382
rect 378784 998776 378836 998782
rect 378784 998718 378836 998724
rect 378600 998708 378652 998714
rect 378600 998650 378652 998656
rect 378612 998306 378640 998650
rect 378600 998300 378652 998306
rect 378600 998242 378652 998248
rect 377404 997824 377456 997830
rect 377404 997766 377456 997772
rect 380176 995450 380204 1006810
rect 429200 1006800 429252 1006806
rect 429198 1006768 429200 1006777
rect 429252 1006768 429254 1006777
rect 429198 1006703 429254 1006712
rect 431684 1006664 431736 1006670
rect 431682 1006632 431684 1006641
rect 431736 1006632 431738 1006641
rect 431682 1006567 431738 1006576
rect 428372 1006528 428424 1006534
rect 428370 1006496 428372 1006505
rect 428424 1006496 428426 1006505
rect 428370 1006431 428426 1006440
rect 427542 1006360 427598 1006369
rect 402244 1006324 402296 1006330
rect 427542 1006295 427544 1006304
rect 402244 1006266 402296 1006272
rect 427596 1006295 427598 1006304
rect 427544 1006266 427596 1006272
rect 382832 1006052 382884 1006058
rect 382832 1005994 382884 1006000
rect 400864 1006052 400916 1006058
rect 400864 1005994 400916 1006000
rect 380900 1001224 380952 1001230
rect 380900 1001166 380952 1001172
rect 380912 995897 380940 1001166
rect 382648 998912 382700 998918
rect 382648 998854 382700 998860
rect 382464 998300 382516 998306
rect 382464 998242 382516 998248
rect 380898 995888 380954 995897
rect 380898 995823 380954 995832
rect 382186 995888 382242 995897
rect 382186 995823 382242 995832
rect 380164 995444 380216 995450
rect 380164 995386 380216 995392
rect 382200 995314 382228 995823
rect 382476 995353 382504 998242
rect 382660 995761 382688 998854
rect 382646 995752 382702 995761
rect 382646 995687 382702 995696
rect 382462 995344 382518 995353
rect 382188 995308 382240 995314
rect 382462 995279 382518 995288
rect 382188 995250 382240 995256
rect 382844 995081 382872 1005994
rect 383568 998776 383620 998782
rect 383620 998724 383700 998730
rect 383568 998718 383700 998724
rect 383580 998702 383700 998718
rect 383292 998572 383344 998578
rect 383292 998514 383344 998520
rect 383108 997824 383160 997830
rect 383108 997766 383160 997772
rect 383120 995586 383148 997766
rect 383108 995580 383160 995586
rect 383108 995522 383160 995528
rect 383304 995450 383332 998514
rect 383476 998436 383528 998442
rect 383476 998378 383528 998384
rect 383108 995444 383160 995450
rect 383108 995386 383160 995392
rect 383292 995444 383344 995450
rect 383292 995386 383344 995392
rect 382830 995072 382886 995081
rect 382830 995007 382886 995016
rect 383120 994809 383148 995386
rect 383106 994800 383162 994809
rect 376024 994764 376076 994770
rect 383106 994735 383162 994744
rect 376024 994706 376076 994712
rect 372988 994628 373040 994634
rect 372988 994570 373040 994576
rect 383488 994537 383516 998378
rect 383672 995330 383700 998702
rect 399944 997144 399996 997150
rect 399944 997086 399996 997092
rect 399956 996985 399984 997086
rect 399942 996976 399998 996985
rect 399942 996911 399998 996920
rect 400494 996704 400550 996713
rect 400494 996639 400550 996648
rect 400034 996432 400090 996441
rect 400034 996367 400090 996376
rect 399852 995852 399904 995858
rect 399852 995794 399904 995800
rect 385038 995752 385094 995761
rect 389362 995752 389418 995761
rect 385094 995710 385342 995738
rect 385038 995687 385094 995696
rect 389730 995752 389786 995761
rect 389418 995710 389666 995738
rect 389362 995687 389418 995696
rect 392214 995752 392270 995761
rect 392150 995710 392214 995738
rect 389730 995687 389786 995696
rect 396630 995752 396686 995761
rect 396382 995710 396630 995738
rect 392214 995687 392270 995696
rect 396630 995687 396686 995696
rect 386326 995616 386382 995625
rect 385696 995586 385986 995602
rect 385684 995580 385986 995586
rect 385736 995574 385986 995580
rect 386326 995551 386382 995560
rect 385684 995522 385736 995528
rect 384316 995438 384698 995466
rect 384316 995330 384344 995438
rect 383672 995302 384344 995330
rect 386340 995314 386368 995551
rect 386328 995308 386380 995314
rect 386328 995250 386380 995256
rect 386512 995308 386564 995314
rect 386512 995250 386564 995256
rect 386524 994809 386552 995250
rect 387812 994809 387840 995452
rect 388364 995178 388392 995452
rect 388640 995450 389022 995466
rect 389744 995450 389772 995687
rect 388628 995444 389022 995450
rect 388680 995438 389022 995444
rect 389088 995444 389140 995450
rect 388628 995386 388680 995392
rect 389088 995386 389140 995392
rect 389732 995444 389784 995450
rect 389732 995386 389784 995392
rect 388902 995344 388958 995353
rect 389100 995330 389128 995386
rect 388958 995302 389128 995330
rect 388902 995279 388958 995288
rect 388352 995172 388404 995178
rect 388352 995114 388404 995120
rect 386510 994800 386566 994809
rect 386510 994735 386566 994744
rect 387798 994800 387854 994809
rect 387798 994735 387854 994744
rect 392688 994537 392716 995452
rect 393332 995042 393360 995452
rect 393320 995036 393372 995042
rect 393320 994978 393372 994984
rect 393976 994770 394004 995452
rect 395186 995438 395292 995466
rect 395264 995382 395292 995438
rect 395252 995376 395304 995382
rect 395252 995318 395304 995324
rect 393964 994764 394016 994770
rect 393964 994706 394016 994712
rect 397012 994634 397040 995452
rect 397656 994906 397684 995452
rect 398852 995246 398880 995452
rect 399864 995382 399892 995794
rect 400048 995761 400076 996367
rect 400034 995752 400090 995761
rect 400034 995687 400090 995696
rect 400508 995489 400536 996639
rect 400876 995994 400904 1005994
rect 402256 996130 402284 1006266
rect 429198 1006224 429254 1006233
rect 429198 1006159 429200 1006168
rect 429252 1006159 429254 1006168
rect 429200 1006130 429252 1006136
rect 421838 1006088 421894 1006097
rect 421838 1006023 421894 1006032
rect 425150 1006088 425206 1006097
rect 431682 1006088 431738 1006097
rect 425150 1006023 425152 1006032
rect 421852 1005582 421880 1006023
rect 425204 1006023 425206 1006032
rect 429752 1006052 429804 1006058
rect 425152 1005994 425204 1006000
rect 431682 1006023 431684 1006032
rect 429752 1005994 429804 1006000
rect 431736 1006023 431738 1006032
rect 431684 1005994 431736 1006000
rect 428372 1005848 428424 1005854
rect 428370 1005816 428372 1005825
rect 428424 1005816 428426 1005825
rect 428370 1005751 428426 1005760
rect 423496 1005712 423548 1005718
rect 423494 1005680 423496 1005689
rect 423548 1005680 423550 1005689
rect 423494 1005615 423550 1005624
rect 421840 1005576 421892 1005582
rect 421840 1005518 421892 1005524
rect 425704 1005576 425756 1005582
rect 425704 1005518 425756 1005524
rect 423496 1005440 423548 1005446
rect 423494 1005408 423496 1005417
rect 423548 1005408 423550 1005417
rect 423494 1005343 423550 1005352
rect 425518 1005136 425574 1005145
rect 425518 1005071 425520 1005080
rect 425572 1005071 425574 1005080
rect 425520 1005042 425572 1005048
rect 422666 1004864 422722 1004873
rect 420460 1004828 420512 1004834
rect 422666 1004799 422668 1004808
rect 420460 1004770 420512 1004776
rect 422720 1004799 422722 1004808
rect 422668 1004770 422720 1004776
rect 419448 1001972 419500 1001978
rect 419448 1001914 419500 1001920
rect 414478 996432 414534 996441
rect 414478 996367 414534 996376
rect 402244 996124 402296 996130
rect 402244 996066 402296 996072
rect 400864 995988 400916 995994
rect 400864 995930 400916 995936
rect 400494 995480 400550 995489
rect 400494 995415 400550 995424
rect 399852 995376 399904 995382
rect 399852 995318 399904 995324
rect 398840 995240 398892 995246
rect 398840 995182 398892 995188
rect 397644 994900 397696 994906
rect 397644 994842 397696 994848
rect 397000 994628 397052 994634
rect 397000 994570 397052 994576
rect 383474 994528 383530 994537
rect 383474 994463 383530 994472
rect 392674 994528 392730 994537
rect 392674 994463 392730 994472
rect 414492 994294 414520 996367
rect 416134 995752 416190 995761
rect 416134 995687 416190 995696
rect 415398 995480 415454 995489
rect 415398 995415 415400 995424
rect 415452 995415 415454 995424
rect 415400 995386 415452 995392
rect 416148 995293 416176 995687
rect 416136 995287 416188 995293
rect 416136 995229 416188 995235
rect 419460 994702 419488 1001914
rect 420472 994974 420500 1004770
rect 424324 1003944 424376 1003950
rect 424322 1003912 424324 1003921
rect 424376 1003912 424378 1003921
rect 424322 1003847 424378 1003856
rect 424692 1002720 424744 1002726
rect 424690 1002688 424692 1002697
rect 424744 1002688 424746 1002697
rect 424690 1002623 424746 1002632
rect 423588 1002108 423640 1002114
rect 423588 1002050 423640 1002056
rect 421470 1002008 421526 1002017
rect 421470 1001943 421472 1001952
rect 421524 1001943 421526 1001952
rect 421472 1001914 421524 1001920
rect 423600 1001230 423628 1002050
rect 425518 1002008 425574 1002017
rect 425518 1001943 425520 1001952
rect 425572 1001943 425574 1001952
rect 425520 1001914 425572 1001920
rect 425716 1001366 425744 1005518
rect 427174 1005408 427230 1005417
rect 427174 1005343 427176 1005352
rect 427228 1005343 427230 1005352
rect 427176 1005314 427228 1005320
rect 428002 1005000 428058 1005009
rect 428002 1004935 428004 1004944
rect 428056 1004935 428058 1004944
rect 428004 1004906 428056 1004912
rect 429764 1002590 429792 1005994
rect 432420 1005712 432472 1005718
rect 432420 1005654 432472 1005660
rect 432432 1005446 432460 1005654
rect 437492 1005582 437520 1007082
rect 553950 1007040 554006 1007049
rect 553950 1006975 553952 1006984
rect 554004 1006975 554006 1006984
rect 562324 1007004 562376 1007010
rect 553952 1006946 554004 1006952
rect 562324 1006946 562376 1006952
rect 505008 1006936 505060 1006942
rect 505006 1006904 505008 1006913
rect 513380 1006936 513432 1006942
rect 505060 1006904 505062 1006913
rect 513380 1006878 513432 1006884
rect 555974 1006904 556030 1006913
rect 505006 1006839 505062 1006848
rect 507858 1006768 507914 1006777
rect 507858 1006703 507860 1006712
rect 507912 1006703 507914 1006712
rect 507860 1006674 507912 1006680
rect 505374 1006632 505430 1006641
rect 469864 1006596 469916 1006602
rect 505374 1006567 505376 1006576
rect 469864 1006538 469916 1006544
rect 505428 1006567 505430 1006576
rect 505376 1006538 505428 1006544
rect 440884 1006528 440936 1006534
rect 440884 1006470 440936 1006476
rect 437480 1005576 437532 1005582
rect 437480 1005518 437532 1005524
rect 432420 1005440 432472 1005446
rect 432420 1005382 432472 1005388
rect 431224 1005100 431276 1005106
rect 431224 1005042 431276 1005048
rect 439504 1005100 439556 1005106
rect 439504 1005042 439556 1005048
rect 429752 1002584 429804 1002590
rect 429752 1002526 429804 1002532
rect 426346 1002144 426402 1002153
rect 426346 1002079 426348 1002088
rect 426400 1002079 426402 1002088
rect 426348 1002050 426400 1002056
rect 428188 1001904 428240 1001910
rect 428188 1001846 428240 1001852
rect 425704 1001360 425756 1001366
rect 425704 1001302 425756 1001308
rect 423588 1001224 423640 1001230
rect 423588 1001166 423640 1001172
rect 428200 998442 428228 1001846
rect 428188 998436 428240 998442
rect 428188 998378 428240 998384
rect 430854 998336 430910 998345
rect 430854 998271 430856 998280
rect 430908 998271 430910 998280
rect 430856 998242 430908 998248
rect 430026 998200 430082 998209
rect 430026 998135 430028 998144
rect 430080 998135 430082 998144
rect 430028 998106 430080 998112
rect 430026 997928 430082 997937
rect 430026 997863 430028 997872
rect 430080 997863 430082 997872
rect 430028 997834 430080 997840
rect 431236 997762 431264 1005042
rect 432878 1004728 432934 1004737
rect 432878 1004663 432880 1004672
rect 432932 1004663 432934 1004672
rect 438124 1004692 438176 1004698
rect 432880 1004634 432932 1004640
rect 438124 1004634 438176 1004640
rect 433984 998300 434036 998306
rect 433984 998242 434036 998248
rect 432604 998164 432656 998170
rect 432604 998106 432656 998112
rect 432050 998064 432106 998073
rect 432050 997999 432052 998008
rect 432104 997999 432106 998008
rect 432052 997970 432104 997976
rect 432052 997892 432104 997898
rect 432052 997834 432104 997840
rect 431224 997756 431276 997762
rect 431224 997698 431276 997704
rect 432064 997150 432092 997834
rect 432616 997490 432644 998106
rect 433996 997626 434024 998242
rect 436744 998028 436796 998034
rect 436744 997970 436796 997976
rect 435362 997792 435418 997801
rect 435362 997727 435418 997736
rect 433984 997620 434036 997626
rect 433984 997562 434036 997568
rect 432604 997484 432656 997490
rect 432604 997426 432656 997432
rect 432052 997144 432104 997150
rect 432052 997086 432104 997092
rect 420460 994968 420512 994974
rect 420460 994910 420512 994916
rect 419448 994696 419500 994702
rect 419448 994638 419500 994644
rect 381176 994288 381228 994294
rect 381176 994230 381228 994236
rect 414480 994288 414532 994294
rect 414480 994230 414532 994236
rect 370504 985992 370556 985998
rect 370504 985934 370556 985940
rect 381188 983634 381216 994230
rect 414112 991636 414164 991642
rect 414112 991578 414164 991584
rect 397828 985992 397880 985998
rect 397828 985934 397880 985940
rect 364996 983606 365470 983634
rect 381188 983606 381662 983634
rect 397840 983620 397868 985934
rect 414124 983620 414152 991578
rect 435376 991506 435404 997727
rect 430304 991500 430356 991506
rect 430304 991442 430356 991448
rect 435364 991500 435416 991506
rect 435364 991442 435416 991448
rect 430316 983620 430344 991442
rect 436756 985998 436784 997970
rect 438136 986134 438164 1004634
rect 439516 1001502 439544 1005042
rect 439504 1001496 439556 1001502
rect 439504 1001438 439556 1001444
rect 440896 998850 440924 1006470
rect 451924 1006188 451976 1006194
rect 451924 1006130 451976 1006136
rect 445024 1005712 445076 1005718
rect 445024 1005654 445076 1005660
rect 443644 1003944 443696 1003950
rect 443644 1003886 443696 1003892
rect 440884 998844 440936 998850
rect 440884 998786 440936 998792
rect 439688 997756 439740 997762
rect 439688 997698 439740 997704
rect 439700 996441 439728 997698
rect 439872 997620 439924 997626
rect 439872 997562 439924 997568
rect 439884 996985 439912 997562
rect 440056 997484 440108 997490
rect 440056 997426 440108 997432
rect 440068 997257 440096 997426
rect 440054 997248 440110 997257
rect 440054 997183 440110 997192
rect 439870 996976 439926 996985
rect 439870 996911 439926 996920
rect 439686 996432 439742 996441
rect 439686 996367 439742 996376
rect 443656 994265 443684 1003886
rect 445036 998578 445064 1005654
rect 448980 1002720 449032 1002726
rect 448980 1002662 449032 1002668
rect 446404 1001360 446456 1001366
rect 446404 1001302 446456 1001308
rect 446416 998714 446444 1001302
rect 448520 998844 448572 998850
rect 448520 998786 448572 998792
rect 446404 998708 446456 998714
rect 446404 998650 446456 998656
rect 445024 998572 445076 998578
rect 445024 998514 445076 998520
rect 448532 995625 448560 998786
rect 448992 997082 449020 1002662
rect 448980 997076 449032 997082
rect 448980 997018 449032 997024
rect 451936 996169 451964 1006130
rect 454684 1005848 454736 1005854
rect 454684 1005790 454736 1005796
rect 451922 996160 451978 996169
rect 451922 996095 451978 996104
rect 448518 995616 448574 995625
rect 448518 995551 448574 995560
rect 454696 995110 454724 1005790
rect 467104 1005576 467156 1005582
rect 467104 1005518 467156 1005524
rect 457444 1005440 457496 1005446
rect 457444 1005382 457496 1005388
rect 454684 995104 454736 995110
rect 454684 995046 454736 995052
rect 457456 994537 457484 1005382
rect 463700 1005304 463752 1005310
rect 463700 1005246 463752 1005252
rect 458180 1001496 458232 1001502
rect 458180 1001438 458232 1001444
rect 458192 998714 458220 1001438
rect 462228 1001224 462280 1001230
rect 462228 1001166 462280 1001172
rect 462240 998850 462268 1001166
rect 458364 998844 458416 998850
rect 458364 998786 458416 998792
rect 462228 998844 462280 998850
rect 462228 998786 462280 998792
rect 458180 998708 458232 998714
rect 458180 998650 458232 998656
rect 458376 995353 458404 998786
rect 463712 998578 463740 1005246
rect 464988 1002584 465040 1002590
rect 464988 1002526 465040 1002532
rect 461584 998572 461636 998578
rect 461584 998514 461636 998520
rect 463700 998572 463752 998578
rect 463700 998514 463752 998520
rect 458362 995344 458418 995353
rect 458362 995279 458418 995288
rect 461596 994838 461624 998514
rect 465000 995081 465028 1002526
rect 464986 995072 465042 995081
rect 464986 995007 465042 995016
rect 461584 994832 461636 994838
rect 461584 994774 461636 994780
rect 457442 994528 457498 994537
rect 457442 994463 457498 994472
rect 446128 994288 446180 994294
rect 443642 994256 443698 994265
rect 446128 994230 446180 994236
rect 443642 994191 443698 994200
rect 438124 986128 438176 986134
rect 438124 986070 438176 986076
rect 436744 985992 436796 985998
rect 436744 985934 436796 985940
rect 446140 983634 446168 994230
rect 467116 993993 467144 1005518
rect 469876 995897 469904 1006538
rect 506202 1006496 506258 1006505
rect 506202 1006431 506204 1006440
rect 506256 1006431 506258 1006440
rect 506204 1006402 506256 1006408
rect 498842 1006088 498898 1006097
rect 471244 1006052 471296 1006058
rect 471244 1005994 471296 1006000
rect 496728 1006052 496780 1006058
rect 498842 1006023 498844 1006032
rect 496728 1005994 496780 1006000
rect 498896 1006023 498898 1006032
rect 498844 1005994 498896 1006000
rect 471256 997754 471284 1005994
rect 472256 998844 472308 998850
rect 472256 998786 472308 998792
rect 472072 998436 472124 998442
rect 472072 998378 472124 998384
rect 471256 997726 471468 997754
rect 470508 997076 470560 997082
rect 470508 997018 470560 997024
rect 469862 995888 469918 995897
rect 469862 995823 469918 995832
rect 470520 994566 470548 997018
rect 471058 996160 471114 996169
rect 471058 996095 471114 996104
rect 471242 996160 471298 996169
rect 471242 996095 471298 996104
rect 471072 994809 471100 996095
rect 471256 995081 471284 996095
rect 471242 995072 471298 995081
rect 471242 995007 471298 995016
rect 471058 994800 471114 994809
rect 471058 994735 471114 994744
rect 470508 994560 470560 994566
rect 470508 994502 470560 994508
rect 471440 994430 471468 997726
rect 471428 994424 471480 994430
rect 471428 994366 471480 994372
rect 472084 994294 472112 998378
rect 472268 995081 472296 998786
rect 472440 998708 472492 998714
rect 472440 998650 472492 998656
rect 472452 995586 472480 998650
rect 472624 998572 472676 998578
rect 472624 998514 472676 998520
rect 472636 996713 472664 998514
rect 488908 997756 488960 997762
rect 488908 997698 488960 997704
rect 488920 997257 488948 997698
rect 489092 997620 489144 997626
rect 489092 997562 489144 997568
rect 488906 997248 488962 997257
rect 488906 997183 488962 997192
rect 489104 996985 489132 997562
rect 489090 996976 489146 996985
rect 489090 996911 489146 996920
rect 472622 996704 472678 996713
rect 472622 996639 472678 996648
rect 489826 996704 489882 996713
rect 489826 996639 489882 996648
rect 490010 996704 490066 996713
rect 490010 996639 490066 996648
rect 474738 995616 474794 995625
rect 473372 995586 473662 995602
rect 472440 995580 472492 995586
rect 472440 995522 472492 995528
rect 473360 995580 473662 995586
rect 473412 995574 473662 995580
rect 474794 995574 474950 995602
rect 474738 995551 474794 995560
rect 473360 995522 473412 995528
rect 474016 995438 474306 995466
rect 476408 995438 476790 995466
rect 477052 995438 477342 995466
rect 474016 995081 474044 995438
rect 476408 995081 476436 995438
rect 477052 995081 477080 995438
rect 472254 995072 472310 995081
rect 472254 995007 472310 995016
rect 474002 995072 474058 995081
rect 474002 995007 474058 995016
rect 476394 995072 476450 995081
rect 476394 995007 476450 995016
rect 477038 995072 477094 995081
rect 477038 995007 477094 995016
rect 474462 994800 474518 994809
rect 474462 994735 474518 994744
rect 472072 994288 472124 994294
rect 472072 994230 472124 994236
rect 474476 993993 474504 994735
rect 477972 994294 478000 995452
rect 477960 994288 478012 994294
rect 478616 994265 478644 995452
rect 480824 995438 481114 995466
rect 480824 995081 480852 995438
rect 480810 995072 480866 995081
rect 480810 995007 480866 995016
rect 481652 994537 481680 995452
rect 482296 994566 482324 995452
rect 482940 994566 482968 995452
rect 484136 995081 484164 995452
rect 484122 995072 484178 995081
rect 484122 995007 484178 995016
rect 484582 995072 484638 995081
rect 484582 995007 484638 995016
rect 482284 994560 482336 994566
rect 481638 994528 481694 994537
rect 482284 994502 482336 994508
rect 482928 994560 482980 994566
rect 482928 994502 482980 994508
rect 481638 994463 481694 994472
rect 484596 994430 484624 995007
rect 484584 994424 484636 994430
rect 484584 994366 484636 994372
rect 485332 994265 485360 995452
rect 485976 995110 486004 995452
rect 486344 995438 486634 995466
rect 486344 995353 486372 995438
rect 486330 995344 486386 995353
rect 486330 995279 486386 995288
rect 485964 995104 486016 995110
rect 485964 995046 486016 995052
rect 487816 994809 487844 995452
rect 487802 994800 487858 994809
rect 487802 994735 487858 994744
rect 489840 994566 489868 996639
rect 490024 994838 490052 996639
rect 496740 994838 496768 1005994
rect 499488 1005440 499540 1005446
rect 500500 1005440 500552 1005446
rect 499488 1005382 499540 1005388
rect 500498 1005408 500500 1005417
rect 500552 1005408 500554 1005417
rect 498844 1005304 498896 1005310
rect 498842 1005272 498844 1005281
rect 498896 1005272 498898 1005281
rect 498842 1005207 498898 1005216
rect 498108 1004964 498160 1004970
rect 498108 1004906 498160 1004912
rect 497924 1004828 497976 1004834
rect 497924 1004770 497976 1004776
rect 497936 1001230 497964 1004770
rect 497924 1001224 497976 1001230
rect 497924 1001166 497976 1001172
rect 498120 1000498 498148 1004906
rect 499500 1000550 499528 1005382
rect 500498 1005343 500554 1005352
rect 500498 1005000 500554 1005009
rect 500498 1004935 500500 1004944
rect 500552 1004935 500554 1004944
rect 500500 1004906 500552 1004912
rect 499670 1004864 499726 1004873
rect 499670 1004799 499672 1004808
rect 499724 1004799 499726 1004808
rect 499672 1004770 499724 1004776
rect 513392 1004086 513420 1006878
rect 555974 1006839 555976 1006848
rect 556028 1006839 556030 1006848
rect 555976 1006810 556028 1006816
rect 556802 1006768 556858 1006777
rect 520924 1006732 520976 1006738
rect 556802 1006703 556804 1006712
rect 520924 1006674 520976 1006680
rect 556856 1006703 556858 1006712
rect 556804 1006674 556856 1006680
rect 518164 1006596 518216 1006602
rect 518164 1006538 518216 1006544
rect 516784 1005304 516836 1005310
rect 516784 1005246 516836 1005252
rect 513380 1004080 513432 1004086
rect 513380 1004022 513432 1004028
rect 509882 1002552 509938 1002561
rect 509882 1002487 509884 1002496
rect 509936 1002487 509938 1002496
rect 515404 1002516 515456 1002522
rect 509884 1002458 509936 1002464
rect 515404 1002458 515456 1002464
rect 501694 1002416 501750 1002425
rect 501694 1002351 501696 1002360
rect 501748 1002351 501750 1002360
rect 503720 1002380 503772 1002386
rect 501696 1002322 501748 1002328
rect 503720 1002322 503772 1002328
rect 503350 1002280 503406 1002289
rect 500592 1002244 500644 1002250
rect 503350 1002215 503352 1002224
rect 500592 1002186 500644 1002192
rect 503404 1002215 503406 1002224
rect 503352 1002186 503404 1002192
rect 499488 1000544 499540 1000550
rect 498120 1000470 498240 1000498
rect 499488 1000486 499540 1000492
rect 500316 1000544 500368 1000550
rect 500316 1000486 500368 1000492
rect 498212 997082 498240 1000470
rect 498200 997076 498252 997082
rect 498200 997018 498252 997024
rect 490012 994832 490064 994838
rect 490012 994774 490064 994780
rect 496728 994832 496780 994838
rect 496728 994774 496780 994780
rect 489828 994560 489880 994566
rect 489828 994502 489880 994508
rect 500328 994430 500356 1000486
rect 500604 997490 500632 1002186
rect 501694 1002144 501750 1002153
rect 500972 1002102 501694 1002130
rect 500776 1001972 500828 1001978
rect 500776 1001914 500828 1001920
rect 500788 998442 500816 1001914
rect 500972 998850 501000 1002102
rect 501694 1002079 501750 1002088
rect 502522 1002144 502578 1002153
rect 502522 1002079 502524 1002088
rect 502576 1002079 502578 1002088
rect 502524 1002050 502576 1002056
rect 501326 1002008 501382 1002017
rect 501326 1001943 501328 1001952
rect 501380 1001943 501382 1001952
rect 502154 1002008 502210 1002017
rect 503350 1002008 503406 1002017
rect 502154 1001943 502210 1001952
rect 502352 1001966 503350 1001994
rect 501328 1001914 501380 1001920
rect 500960 998844 501012 998850
rect 500960 998786 501012 998792
rect 502168 998578 502196 1001943
rect 502156 998572 502208 998578
rect 502156 998514 502208 998520
rect 500776 998436 500828 998442
rect 500776 998378 500828 998384
rect 500592 997484 500644 997490
rect 500592 997426 500644 997432
rect 502352 994566 502380 1001966
rect 503350 1001943 503406 1001952
rect 503732 1000550 503760 1002322
rect 504178 1002280 504234 1002289
rect 504178 1002215 504180 1002224
rect 504232 1002215 504234 1002224
rect 510068 1002244 510120 1002250
rect 504180 1002186 504232 1002192
rect 510068 1002186 510120 1002192
rect 505744 1002108 505796 1002114
rect 505744 1002050 505796 1002056
rect 504546 1002008 504602 1002017
rect 504546 1001943 504548 1001952
rect 504600 1001943 504602 1001952
rect 504548 1001914 504600 1001920
rect 503720 1000544 503772 1000550
rect 503720 1000486 503772 1000492
rect 505374 999016 505430 999025
rect 505374 998951 505376 998960
rect 505428 998951 505430 998960
rect 505376 998922 505428 998928
rect 505756 995110 505784 1002050
rect 506848 1001972 506900 1001978
rect 506848 1001914 506900 1001920
rect 506860 997754 506888 1001914
rect 507398 999152 507454 999161
rect 507398 999087 507400 999096
rect 507452 999087 507454 999096
rect 509240 999116 509292 999122
rect 507400 999058 507452 999064
rect 509240 999058 509292 999064
rect 507030 998744 507086 998753
rect 507030 998679 507032 998688
rect 507084 998679 507086 998688
rect 507032 998650 507084 998656
rect 509054 998336 509110 998345
rect 509054 998271 509056 998280
rect 509108 998271 509110 998280
rect 509056 998242 509108 998248
rect 508226 998200 508282 998209
rect 508226 998135 508228 998144
rect 508280 998135 508282 998144
rect 508228 998106 508280 998112
rect 508228 997960 508280 997966
rect 508226 997928 508228 997937
rect 508280 997928 508282 997937
rect 508226 997863 508282 997872
rect 509252 997762 509280 999058
rect 510080 998714 510108 1002186
rect 511448 998980 511500 998986
rect 511448 998922 511500 998928
rect 509884 998708 509936 998714
rect 509884 998650 509936 998656
rect 510068 998708 510120 998714
rect 510068 998650 510120 998656
rect 509896 997762 509924 998650
rect 511264 998164 511316 998170
rect 511264 998106 511316 998112
rect 510712 997960 510764 997966
rect 510712 997902 510764 997908
rect 509240 997756 509292 997762
rect 506860 997726 507072 997754
rect 507044 995518 507072 997726
rect 509240 997698 509292 997704
rect 509884 997756 509936 997762
rect 509884 997698 509936 997704
rect 510724 997626 510752 997902
rect 510712 997620 510764 997626
rect 510712 997562 510764 997568
rect 511276 996130 511304 998106
rect 511460 997257 511488 998922
rect 514024 998300 514076 998306
rect 514024 998242 514076 998248
rect 512642 997792 512698 997801
rect 512642 997727 512698 997736
rect 511446 997248 511502 997257
rect 511446 997183 511502 997192
rect 511264 996124 511316 996130
rect 511264 996066 511316 996072
rect 507032 995512 507084 995518
rect 507032 995454 507084 995460
rect 505744 995104 505796 995110
rect 505744 995046 505796 995052
rect 502340 994560 502392 994566
rect 502340 994502 502392 994508
rect 500316 994424 500368 994430
rect 500316 994366 500368 994372
rect 477960 994230 478012 994236
rect 478602 994256 478658 994265
rect 478602 994191 478658 994200
rect 485318 994256 485374 994265
rect 485318 994191 485374 994200
rect 511078 994256 511134 994265
rect 511078 994191 511134 994200
rect 467102 993984 467158 993993
rect 467102 993919 467158 993928
rect 474462 993984 474518 993993
rect 474462 993919 474518 993928
rect 478972 991500 479024 991506
rect 478972 991442 479024 991448
rect 462780 986128 462832 986134
rect 462780 986070 462832 986076
rect 446140 983606 446522 983634
rect 462792 983620 462820 986070
rect 478984 983620 479012 991442
rect 495164 985992 495216 985998
rect 495164 985934 495216 985940
rect 495176 983620 495204 985934
rect 511092 983634 511120 994191
rect 512656 990146 512684 997727
rect 513656 994832 513708 994838
rect 513656 994774 513708 994780
rect 513840 994832 513892 994838
rect 513840 994774 513892 994780
rect 513668 994294 513696 994774
rect 513852 994566 513880 994774
rect 513840 994560 513892 994566
rect 513840 994502 513892 994508
rect 513656 994288 513708 994294
rect 513656 994230 513708 994236
rect 512644 990140 512696 990146
rect 512644 990082 512696 990088
rect 514036 985998 514064 998242
rect 514208 994560 514260 994566
rect 514208 994502 514260 994508
rect 514220 994294 514248 994502
rect 514208 994288 514260 994294
rect 514208 994230 514260 994236
rect 515416 986134 515444 1002458
rect 516796 1001894 516824 1005246
rect 516796 1001866 517100 1001894
rect 516876 1000544 516928 1000550
rect 516876 1000486 516928 1000492
rect 516690 998608 516746 998617
rect 516888 998578 516916 1000486
rect 516690 998543 516692 998552
rect 516744 998543 516746 998552
rect 516876 998572 516928 998578
rect 516692 998514 516744 998520
rect 516876 998514 516928 998520
rect 516876 997756 516928 997762
rect 516876 997698 516928 997704
rect 516692 997484 516744 997490
rect 516692 997426 516744 997432
rect 516704 996713 516732 997426
rect 516888 996985 516916 997698
rect 516874 996976 516930 996985
rect 516874 996911 516930 996920
rect 516690 996704 516746 996713
rect 516690 996639 516746 996648
rect 517072 993682 517100 1001866
rect 517520 998844 517572 998850
rect 517520 998786 517572 998792
rect 517532 995858 517560 998786
rect 517704 997076 517756 997082
rect 517704 997018 517756 997024
rect 517520 995852 517572 995858
rect 517520 995794 517572 995800
rect 517716 994294 517744 997018
rect 518176 995353 518204 1006538
rect 518900 1004080 518952 1004086
rect 518900 1004022 518952 1004028
rect 518912 1001894 518940 1004022
rect 518912 1001866 519124 1001894
rect 518898 998608 518954 998617
rect 518898 998543 518954 998552
rect 518912 995625 518940 998543
rect 519096 996441 519124 1001866
rect 519082 996432 519138 996441
rect 519082 996367 519138 996376
rect 518898 995616 518954 995625
rect 518898 995551 518954 995560
rect 518162 995344 518218 995353
rect 518162 995279 518218 995288
rect 520936 995081 520964 1006674
rect 555146 1006496 555202 1006505
rect 555146 1006431 555148 1006440
rect 555200 1006431 555202 1006440
rect 555148 1006402 555200 1006408
rect 551466 1006360 551522 1006369
rect 551466 1006295 551468 1006304
rect 551520 1006295 551522 1006304
rect 556804 1006324 556856 1006330
rect 551468 1006266 551520 1006272
rect 556804 1006266 556856 1006272
rect 555424 1006188 555476 1006194
rect 555424 1006130 555476 1006136
rect 550270 1006088 550326 1006097
rect 522304 1006052 522356 1006058
rect 522304 1005994 522356 1006000
rect 549168 1006052 549220 1006058
rect 550270 1006023 550272 1006032
rect 549168 1005994 549220 1006000
rect 550324 1006023 550326 1006032
rect 554778 1006088 554834 1006097
rect 554778 1006023 554780 1006032
rect 550272 1005994 550324 1006000
rect 554832 1006023 554834 1006032
rect 554780 1005994 554832 1006000
rect 521292 1001224 521344 1001230
rect 521292 1001166 521344 1001172
rect 520922 995072 520978 995081
rect 520922 995007 520978 995016
rect 517704 994288 517756 994294
rect 517704 994230 517756 994236
rect 521304 993818 521332 1001166
rect 522316 995994 522344 1005994
rect 523868 998912 523920 998918
rect 523868 998854 523920 998860
rect 523684 998436 523736 998442
rect 523684 998378 523736 998384
rect 523498 996704 523554 996713
rect 523498 996639 523554 996648
rect 522304 995988 522356 995994
rect 522304 995930 522356 995936
rect 523316 995852 523368 995858
rect 523316 995794 523368 995800
rect 523328 994265 523356 995794
rect 523512 994994 523540 996639
rect 523696 996169 523724 998378
rect 523880 997665 523908 998854
rect 524052 998572 524104 998578
rect 524052 998514 524104 998520
rect 523866 997656 523922 997665
rect 523866 997591 523922 997600
rect 524064 997257 524092 998514
rect 549180 998442 549208 1005994
rect 551468 1005304 551520 1005310
rect 551466 1005272 551468 1005281
rect 551520 1005272 551522 1005281
rect 551466 1005207 551522 1005216
rect 554778 1003368 554834 1003377
rect 554608 1003338 554778 1003354
rect 553400 1003332 553452 1003338
rect 553400 1003274 553452 1003280
rect 554596 1003332 554778 1003338
rect 554648 1003326 554778 1003332
rect 554778 1003303 554834 1003312
rect 554596 1003274 554648 1003280
rect 553122 1002688 553178 1002697
rect 553122 1002623 553124 1002632
rect 553176 1002623 553178 1002632
rect 553124 1002594 553176 1002600
rect 553216 1002176 553268 1002182
rect 553216 1002118 553268 1002124
rect 550272 1001224 550324 1001230
rect 550270 1001192 550272 1001201
rect 550324 1001192 550326 1001201
rect 550270 1001127 550326 1001136
rect 549168 998436 549220 998442
rect 549168 998378 549220 998384
rect 550548 998300 550600 998306
rect 550548 998242 550600 998248
rect 552940 998300 552992 998306
rect 552940 998242 552992 998248
rect 550560 997558 550588 998242
rect 552294 997792 552350 997801
rect 551940 997750 552294 997778
rect 550548 997552 550600 997558
rect 550548 997494 550600 997500
rect 540336 997416 540388 997422
rect 540336 997358 540388 997364
rect 524050 997248 524106 997257
rect 524050 997183 524106 997192
rect 540348 996985 540376 997358
rect 540334 996976 540390 996985
rect 540334 996911 540390 996920
rect 524050 996432 524106 996441
rect 524050 996367 524106 996376
rect 523682 996160 523738 996169
rect 523682 996095 523738 996104
rect 524064 995330 524092 996367
rect 529754 995752 529810 995761
rect 532146 995752 532202 995761
rect 529810 995710 530058 995738
rect 529754 995687 529810 995696
rect 532882 995752 532938 995761
rect 532202 995710 532542 995738
rect 532146 995687 532202 995696
rect 532882 995687 532938 995696
rect 535274 995752 535330 995761
rect 536562 995752 536618 995761
rect 535330 995710 535578 995738
rect 535274 995687 535330 995696
rect 536618 995710 536774 995738
rect 536562 995687 536618 995696
rect 529018 995616 529074 995625
rect 529074 995574 529414 995602
rect 529018 995551 529074 995560
rect 527916 995512 527968 995518
rect 524616 995438 525090 995466
rect 525260 995438 525734 995466
rect 526088 995438 526378 995466
rect 527968 995460 528218 995466
rect 527916 995454 528218 995460
rect 527928 995438 528218 995454
rect 524616 995330 524644 995438
rect 524064 995302 524644 995330
rect 525260 994994 525288 995438
rect 523512 994966 525288 994994
rect 523500 994560 523552 994566
rect 523500 994502 523552 994508
rect 523684 994560 523736 994566
rect 526088 994537 526116 995438
rect 528756 995110 528784 995452
rect 532896 995178 532924 995687
rect 533526 995616 533582 995625
rect 533582 995574 533738 995602
rect 533526 995551 533582 995560
rect 533094 995438 533384 995466
rect 533356 995178 533384 995438
rect 528928 995172 528980 995178
rect 528928 995114 528980 995120
rect 532884 995172 532936 995178
rect 532884 995114 532936 995120
rect 533344 995172 533396 995178
rect 533344 995114 533396 995120
rect 534080 995172 534132 995178
rect 534080 995114 534132 995120
rect 528744 995104 528796 995110
rect 528744 995046 528796 995052
rect 523684 994502 523736 994508
rect 526074 994528 526130 994537
rect 523314 994256 523370 994265
rect 523314 994191 523370 994200
rect 523512 994158 523540 994502
rect 523696 994294 523724 994502
rect 526074 994463 526130 994472
rect 523684 994288 523736 994294
rect 528940 994265 528968 995114
rect 534092 994430 534120 995114
rect 534368 994566 534396 995452
rect 537128 995438 537418 995466
rect 537128 995353 537156 995438
rect 537114 995344 537170 995353
rect 537114 995279 537170 995288
rect 534356 994560 534408 994566
rect 534356 994502 534408 994508
rect 534080 994424 534132 994430
rect 534080 994366 534132 994372
rect 538048 994294 538076 995452
rect 539244 994838 539272 995452
rect 551940 994838 551968 997750
rect 552294 997727 552350 997736
rect 552296 997280 552348 997286
rect 552294 997248 552296 997257
rect 552348 997248 552350 997257
rect 552294 997183 552350 997192
rect 552952 996554 552980 998242
rect 553228 996810 553256 1002118
rect 553412 999122 553440 1003274
rect 553768 1002652 553820 1002658
rect 553768 1002594 553820 1002600
rect 553400 999116 553452 999122
rect 553400 999058 553452 999064
rect 553780 998578 553808 1002594
rect 553952 1002176 554004 1002182
rect 553950 1002144 553952 1002153
rect 554004 1002144 554006 1002153
rect 553950 1002079 554006 1002088
rect 553768 998572 553820 998578
rect 553768 998514 553820 998520
rect 555436 997422 555464 1006130
rect 555974 1004864 556030 1004873
rect 555974 1004799 555976 1004808
rect 556028 1004799 556030 1004808
rect 555976 1004770 556028 1004776
rect 556344 999116 556396 999122
rect 556344 999058 556396 999064
rect 555424 997416 555476 997422
rect 555424 997358 555476 997364
rect 553216 996804 553268 996810
rect 553216 996746 553268 996752
rect 553122 996568 553178 996577
rect 552952 996526 553122 996554
rect 553122 996503 553178 996512
rect 556356 996334 556384 999058
rect 556816 998714 556844 1006266
rect 558826 1006224 558882 1006233
rect 562336 1006194 562364 1006946
rect 569408 1006868 569460 1006874
rect 569408 1006810 569460 1006816
rect 564440 1006732 564492 1006738
rect 564440 1006674 564492 1006680
rect 558826 1006159 558828 1006168
rect 558880 1006159 558882 1006168
rect 562324 1006188 562376 1006194
rect 558828 1006130 558880 1006136
rect 562324 1006130 562376 1006136
rect 564452 1005446 564480 1006674
rect 567844 1006188 567896 1006194
rect 567844 1006130 567896 1006136
rect 564440 1005440 564492 1005446
rect 564440 1005382 564492 1005388
rect 557170 1005000 557226 1005009
rect 557170 1004935 557172 1004944
rect 557224 1004935 557226 1004944
rect 558920 1004964 558972 1004970
rect 557172 1004906 557224 1004912
rect 558920 1004906 558972 1004912
rect 558184 1004828 558236 1004834
rect 558184 1004770 558236 1004776
rect 557630 1004728 557686 1004737
rect 557630 1004663 557632 1004672
rect 557684 1004663 557686 1004672
rect 557632 1004634 557684 1004640
rect 557998 1002280 558054 1002289
rect 557998 1002215 558000 1002224
rect 558052 1002215 558054 1002224
rect 558000 1002186 558052 1002192
rect 557998 1002008 558054 1002017
rect 557998 1001943 558000 1001952
rect 558052 1001943 558054 1001952
rect 558000 1001914 558052 1001920
rect 558196 1000006 558224 1004770
rect 558932 1003950 558960 1004906
rect 560850 1004728 560906 1004737
rect 559564 1004692 559616 1004698
rect 560850 1004663 560852 1004672
rect 559564 1004634 559616 1004640
rect 560904 1004663 560906 1004672
rect 566464 1004692 566516 1004698
rect 560852 1004634 560904 1004640
rect 566464 1004634 566516 1004640
rect 558920 1003944 558972 1003950
rect 558920 1003886 558972 1003892
rect 558826 1002688 558882 1002697
rect 558826 1002623 558828 1002632
rect 558880 1002623 558882 1002632
rect 558828 1002594 558880 1002600
rect 558184 1000000 558236 1000006
rect 558184 999942 558236 999948
rect 556804 998708 556856 998714
rect 556804 998650 556856 998656
rect 556344 996328 556396 996334
rect 556344 996270 556396 996276
rect 539232 994832 539284 994838
rect 539232 994774 539284 994780
rect 551928 994832 551980 994838
rect 551928 994774 551980 994780
rect 538036 994288 538088 994294
rect 523684 994230 523736 994236
rect 528926 994256 528982 994265
rect 538036 994230 538088 994236
rect 528926 994191 528982 994200
rect 523500 994152 523552 994158
rect 523500 994094 523552 994100
rect 521292 993812 521344 993818
rect 521292 993754 521344 993760
rect 517060 993676 517112 993682
rect 517060 993618 517112 993624
rect 559576 991506 559604 1004634
rect 562508 1002652 562560 1002658
rect 562508 1002594 562560 1002600
rect 560850 1002552 560906 1002561
rect 560850 1002487 560852 1002496
rect 560904 1002487 560906 1002496
rect 560852 1002458 560904 1002464
rect 560482 1002416 560538 1002425
rect 560482 1002351 560484 1002360
rect 560536 1002351 560538 1002360
rect 560484 1002322 560536 1002328
rect 560944 1002244 560996 1002250
rect 560944 1002186 560996 1002192
rect 560022 1002144 560078 1002153
rect 560022 1002079 560024 1002088
rect 560076 1002079 560078 1002088
rect 560024 1002050 560076 1002056
rect 560300 1001972 560352 1001978
rect 560300 1001914 560352 1001920
rect 560312 995994 560340 1001914
rect 560300 995988 560352 995994
rect 560300 995930 560352 995936
rect 560956 992934 560984 1002186
rect 562324 1002108 562376 1002114
rect 562324 1002050 562376 1002056
rect 561678 1002008 561734 1002017
rect 561678 1001943 561680 1001952
rect 561732 1001943 561734 1001952
rect 561680 1001914 561732 1001920
rect 560944 992928 560996 992934
rect 560944 992870 560996 992876
rect 559564 991500 559616 991506
rect 559564 991442 559616 991448
rect 562336 990146 562364 1002050
rect 562520 993070 562548 1002594
rect 565084 1002516 565136 1002522
rect 565084 1002458 565136 1002464
rect 563060 1002380 563112 1002386
rect 563060 1002322 563112 1002328
rect 563072 996130 563100 1002322
rect 563704 1001972 563756 1001978
rect 563704 1001914 563756 1001920
rect 563060 996124 563112 996130
rect 563060 996066 563112 996072
rect 562508 993064 562560 993070
rect 562508 993006 562560 993012
rect 543832 990140 543884 990146
rect 543832 990082 543884 990088
rect 562324 990140 562376 990146
rect 562324 990082 562376 990088
rect 515404 986128 515456 986134
rect 515404 986070 515456 986076
rect 527640 986128 527692 986134
rect 527640 986070 527692 986076
rect 514024 985992 514076 985998
rect 514024 985934 514076 985940
rect 511092 983606 511474 983634
rect 527652 983620 527680 986070
rect 543844 983620 543872 990082
rect 563716 987426 563744 1001914
rect 564440 998436 564492 998442
rect 564440 998378 564492 998384
rect 564452 996674 564480 998378
rect 564440 996668 564492 996674
rect 564440 996610 564492 996616
rect 563704 987420 563756 987426
rect 563704 987362 563756 987368
rect 565096 985998 565124 1002458
rect 565820 1000000 565872 1000006
rect 565820 999942 565872 999948
rect 565832 996946 565860 999942
rect 565820 996940 565872 996946
rect 565820 996882 565872 996888
rect 566476 986134 566504 1004634
rect 567856 1000142 567884 1006130
rect 569224 1005304 569276 1005310
rect 569224 1005246 569276 1005252
rect 569236 1001894 569264 1005246
rect 569420 1001894 569448 1006810
rect 570328 1006460 570380 1006466
rect 570328 1006402 570380 1006408
rect 570340 1004154 570368 1006402
rect 573548 1006052 573600 1006058
rect 573548 1005994 573600 1006000
rect 570604 1005440 570656 1005446
rect 570604 1005382 570656 1005388
rect 570328 1004148 570380 1004154
rect 570328 1004090 570380 1004096
rect 569236 1001866 569356 1001894
rect 569420 1001866 569540 1001894
rect 567844 1000136 567896 1000142
rect 567844 1000078 567896 1000084
rect 567476 998708 567528 998714
rect 567476 998650 567528 998656
rect 567488 996198 567516 998650
rect 569132 998572 569184 998578
rect 569132 998514 569184 998520
rect 568856 996668 568908 996674
rect 568856 996610 568908 996616
rect 567476 996192 567528 996198
rect 567476 996134 567528 996140
rect 568868 994430 568896 996610
rect 569144 995110 569172 998514
rect 569132 995104 569184 995110
rect 569132 995046 569184 995052
rect 568856 994424 568908 994430
rect 568856 994366 568908 994372
rect 569328 993954 569356 1001866
rect 569512 997694 569540 1001866
rect 569500 997688 569552 997694
rect 569500 997630 569552 997636
rect 570616 994294 570644 1005382
rect 573364 1004148 573416 1004154
rect 573364 1004090 573416 1004096
rect 570788 1003944 570840 1003950
rect 570788 1003886 570840 1003892
rect 570800 994673 570828 1003886
rect 571340 1000136 571392 1000142
rect 571340 1000078 571392 1000084
rect 571352 997150 571380 1000078
rect 571340 997144 571392 997150
rect 571340 997086 571392 997092
rect 572810 994936 572866 994945
rect 572810 994871 572866 994880
rect 570786 994664 570842 994673
rect 570786 994599 570842 994608
rect 570604 994288 570656 994294
rect 570604 994230 570656 994236
rect 569316 993948 569368 993954
rect 569316 993890 569368 993896
rect 572824 990894 572852 994871
rect 573376 994566 573404 1004090
rect 573560 997286 573588 1005994
rect 574100 1001224 574152 1001230
rect 574100 1001166 574152 1001172
rect 573548 997280 573600 997286
rect 573548 997222 573600 997228
rect 573364 994560 573416 994566
rect 573364 994502 573416 994508
rect 574112 994090 574140 1001166
rect 617340 1000544 617392 1000550
rect 617340 1000486 617392 1000492
rect 625436 1000544 625488 1000550
rect 625436 1000486 625488 1000492
rect 590936 999320 590988 999326
rect 590936 999262 590988 999268
rect 590384 997416 590436 997422
rect 590384 997358 590436 997364
rect 590396 996418 590424 997358
rect 590566 996976 590622 996985
rect 590566 996911 590568 996920
rect 590620 996911 590622 996920
rect 590568 996882 590620 996888
rect 590568 996736 590620 996742
rect 590566 996704 590568 996713
rect 590620 996704 590622 996713
rect 590566 996639 590622 996648
rect 590566 996432 590622 996441
rect 590396 996390 590566 996418
rect 590566 996367 590622 996376
rect 590384 996328 590436 996334
rect 590384 996270 590436 996276
rect 590396 995058 590424 996270
rect 590568 996192 590620 996198
rect 590568 996134 590620 996140
rect 590580 995353 590608 996134
rect 590566 995344 590622 995353
rect 590566 995279 590622 995288
rect 590566 995072 590622 995081
rect 590396 995030 590566 995058
rect 590566 995007 590622 995016
rect 590948 994566 590976 999262
rect 617352 998442 617380 1000486
rect 625068 999320 625120 999326
rect 625068 999262 625120 999268
rect 618168 999184 618220 999190
rect 618168 999126 618220 999132
rect 591120 998436 591172 998442
rect 591120 998378 591172 998384
rect 617340 998436 617392 998442
rect 617340 998378 617392 998384
rect 591132 997150 591160 998378
rect 591304 997824 591356 997830
rect 591304 997766 591356 997772
rect 591316 997286 591344 997766
rect 618180 997558 618208 999126
rect 623688 997688 623740 997694
rect 623688 997630 623740 997636
rect 618168 997552 618220 997558
rect 618168 997494 618220 997500
rect 591304 997280 591356 997286
rect 591304 997222 591356 997228
rect 591120 997144 591172 997150
rect 591120 997086 591172 997092
rect 623700 995586 623728 997630
rect 625080 997257 625108 999262
rect 625066 997248 625122 997257
rect 625066 997183 625122 997192
rect 625250 997248 625306 997257
rect 625250 997183 625306 997192
rect 623688 995580 623740 995586
rect 623688 995522 623740 995528
rect 625264 995178 625292 997183
rect 625252 995172 625304 995178
rect 625252 995114 625304 995120
rect 625114 995104 625166 995110
rect 625166 995052 625200 995058
rect 625114 995046 625200 995052
rect 625126 995030 625200 995046
rect 590936 994560 590988 994566
rect 590936 994502 590988 994508
rect 591304 994560 591356 994566
rect 625172 994537 625200 995030
rect 591304 994502 591356 994508
rect 625158 994528 625214 994537
rect 591316 994294 591344 994502
rect 625158 994463 625214 994472
rect 625448 994294 625476 1000486
rect 625620 999184 625672 999190
rect 625620 999126 625672 999132
rect 625632 996033 625660 999126
rect 625804 997824 625856 997830
rect 625804 997766 625856 997772
rect 625618 996024 625674 996033
rect 625618 995959 625674 995968
rect 625816 995761 625844 997766
rect 630310 995786 630366 995795
rect 625802 995752 625858 995761
rect 625802 995687 625858 995696
rect 627182 995752 627238 995761
rect 629206 995752 629262 995761
rect 627238 995710 627532 995738
rect 627182 995687 627238 995696
rect 629206 995687 629262 995696
rect 629850 995752 629906 995761
rect 629906 995710 630016 995738
rect 635646 995752 635702 995761
rect 630366 995730 630568 995738
rect 630310 995721 630568 995730
rect 630324 995710 630568 995721
rect 629850 995687 629906 995696
rect 635646 995687 635702 995696
rect 637026 995752 637082 995761
rect 637082 995710 637376 995738
rect 637026 995687 637082 995696
rect 626552 995586 626888 995602
rect 626540 995580 626888 995586
rect 626592 995574 626888 995580
rect 626540 995522 626592 995528
rect 629220 995518 629248 995687
rect 635186 995616 635242 995625
rect 635242 995574 635536 995602
rect 635186 995551 635242 995560
rect 629208 995512 629260 995518
rect 627932 995438 628176 995466
rect 631508 995512 631560 995518
rect 629208 995454 629260 995460
rect 630876 995438 631212 995466
rect 631560 995460 631856 995466
rect 631508 995454 631856 995460
rect 631520 995438 631856 995454
rect 634004 995438 634340 995466
rect 634832 995438 634892 995466
rect 627932 994809 627960 995438
rect 627918 994800 627974 994809
rect 627918 994735 627974 994744
rect 630876 994294 630904 995438
rect 634004 995178 634032 995438
rect 633992 995172 634044 995178
rect 633992 995114 634044 995120
rect 634832 994838 634860 995438
rect 634820 994832 634872 994838
rect 635660 994809 635688 995687
rect 635844 995438 636180 995466
rect 638572 995438 638908 995466
rect 635844 995353 635872 995438
rect 635830 995344 635886 995353
rect 635830 995279 635886 995288
rect 638880 995110 638908 995438
rect 639064 995438 639216 995466
rect 639524 995438 639860 995466
rect 640996 995438 641056 995466
rect 638868 995104 638920 995110
rect 638868 995046 638920 995052
rect 634820 994774 634872 994780
rect 635646 994800 635702 994809
rect 635646 994735 635702 994744
rect 639064 994566 639092 995438
rect 639052 994560 639104 994566
rect 639052 994502 639104 994508
rect 639524 994430 639552 995438
rect 640800 995104 640852 995110
rect 640996 995081 641024 995438
rect 660304 995147 660356 995153
rect 660304 995089 660356 995095
rect 640800 995046 640852 995052
rect 640982 995072 641038 995081
rect 639512 994424 639564 994430
rect 639512 994366 639564 994372
rect 591304 994288 591356 994294
rect 591304 994230 591356 994236
rect 625436 994288 625488 994294
rect 625436 994230 625488 994236
rect 630864 994288 630916 994294
rect 630864 994230 630916 994236
rect 574100 994084 574152 994090
rect 574100 994026 574152 994032
rect 572812 990888 572864 990894
rect 572812 990830 572864 990836
rect 576308 990888 576360 990894
rect 576308 990830 576360 990836
rect 566464 986128 566516 986134
rect 566464 986070 566516 986076
rect 560116 985992 560168 985998
rect 560116 985934 560168 985940
rect 565084 985992 565136 985998
rect 565084 985934 565136 985940
rect 560128 983620 560156 985934
rect 576320 983620 576348 990830
rect 608784 987420 608836 987426
rect 608784 987362 608836 987368
rect 592500 986128 592552 986134
rect 592500 986070 592552 986076
rect 592512 983620 592540 986070
rect 608796 983620 608824 987362
rect 624976 985992 625028 985998
rect 624976 985934 625028 985940
rect 624988 983620 625016 985934
rect 640812 983634 640840 995046
rect 640982 995007 641038 995016
rect 660316 994702 660344 995089
rect 660304 994696 660356 994702
rect 660304 994638 660356 994644
rect 660764 994628 660816 994634
rect 660764 994570 660816 994576
rect 660776 993682 660804 994570
rect 660948 994560 661000 994566
rect 660948 994502 661000 994508
rect 660960 993818 660988 994502
rect 660948 993812 661000 993818
rect 660948 993754 661000 993760
rect 660764 993676 660816 993682
rect 660764 993618 660816 993624
rect 660304 993064 660356 993070
rect 660304 993006 660356 993012
rect 658924 991500 658976 991506
rect 658924 991442 658976 991448
rect 640812 983606 641194 983634
rect 62118 976032 62174 976041
rect 62118 975967 62174 975976
rect 62132 975730 62160 975967
rect 651654 975896 651710 975905
rect 651654 975831 651710 975840
rect 651668 975730 651696 975831
rect 62120 975724 62172 975730
rect 62120 975666 62172 975672
rect 651656 975724 651708 975730
rect 651656 975666 651708 975672
rect 62118 962976 62174 962985
rect 62118 962911 62174 962920
rect 62132 961926 62160 962911
rect 651470 962568 651526 962577
rect 651470 962503 651526 962512
rect 651484 961926 651512 962503
rect 62120 961920 62172 961926
rect 62120 961862 62172 961868
rect 651472 961920 651524 961926
rect 651472 961862 651524 961868
rect 62118 949920 62174 949929
rect 62118 949855 62174 949864
rect 62132 946014 62160 949855
rect 652206 949376 652262 949385
rect 652206 949311 652262 949320
rect 652220 948122 652248 949311
rect 652208 948116 652260 948122
rect 652208 948058 652260 948064
rect 62120 946008 62172 946014
rect 62120 945950 62172 945956
rect 651472 937032 651524 937038
rect 651472 936974 651524 936980
rect 651484 936193 651512 936974
rect 651470 936184 651526 936193
rect 651470 936119 651526 936128
rect 658936 936057 658964 991442
rect 660316 937281 660344 993006
rect 667204 992928 667256 992934
rect 667204 992870 667256 992876
rect 664444 975724 664496 975730
rect 664444 975666 664496 975672
rect 661682 957808 661738 957817
rect 661682 957743 661738 957752
rect 660302 937272 660358 937281
rect 660302 937207 660358 937216
rect 661696 937038 661724 957743
rect 663064 948116 663116 948122
rect 663064 948058 663116 948064
rect 663076 941769 663104 948058
rect 664456 947345 664484 975666
rect 665824 961920 665876 961926
rect 665824 961862 665876 961868
rect 664442 947336 664498 947345
rect 664442 947271 664498 947280
rect 663062 941760 663118 941769
rect 663062 941695 663118 941704
rect 665836 939865 665864 961862
rect 665822 939856 665878 939865
rect 665822 939791 665878 939800
rect 667216 937825 667244 992870
rect 668584 990140 668636 990146
rect 668584 990082 668636 990088
rect 668596 938505 668624 990082
rect 675036 966709 675418 966737
rect 674378 966104 674434 966113
rect 674378 966039 674434 966048
rect 673366 962840 673422 962849
rect 673366 962775 673422 962784
rect 673090 962568 673146 962577
rect 673090 962503 673146 962512
rect 672906 958760 672962 958769
rect 672906 958695 672962 958704
rect 672920 939794 672948 958695
rect 672920 939766 673040 939794
rect 668582 938496 668638 938505
rect 668582 938431 668638 938440
rect 672170 938088 672226 938097
rect 672170 938023 672226 938032
rect 667202 937816 667258 937825
rect 667202 937751 667258 937760
rect 672184 937281 672212 938023
rect 672814 937816 672870 937825
rect 672814 937751 672870 937760
rect 672630 937544 672686 937553
rect 672630 937479 672686 937488
rect 672170 937272 672226 937281
rect 672170 937207 672226 937216
rect 661684 937032 661736 937038
rect 661684 936974 661736 936980
rect 671802 936728 671858 936737
rect 671802 936663 671858 936672
rect 658922 936048 658978 936057
rect 658922 935983 658978 935992
rect 671618 935776 671674 935785
rect 671618 935711 671674 935720
rect 62118 923808 62174 923817
rect 62118 923743 62174 923752
rect 62132 923302 62160 923743
rect 62120 923296 62172 923302
rect 62120 923238 62172 923244
rect 651470 922720 651526 922729
rect 651470 922655 651526 922664
rect 651484 921874 651512 922655
rect 651472 921868 651524 921874
rect 651472 921810 651524 921816
rect 661684 921868 661736 921874
rect 661684 921810 661736 921816
rect 62118 910752 62174 910761
rect 62118 910687 62174 910696
rect 62132 909498 62160 910687
rect 652390 909528 652446 909537
rect 62120 909492 62172 909498
rect 652390 909463 652392 909472
rect 62120 909434 62172 909440
rect 652444 909463 652446 909472
rect 652392 909434 652444 909440
rect 62118 897832 62174 897841
rect 62118 897767 62174 897776
rect 62132 897054 62160 897767
rect 62120 897048 62172 897054
rect 62120 896990 62172 896996
rect 651470 896200 651526 896209
rect 651470 896135 651526 896144
rect 651484 895694 651512 896135
rect 651472 895688 651524 895694
rect 651472 895630 651524 895636
rect 54482 892256 54538 892265
rect 54482 892191 54538 892200
rect 55862 892256 55918 892265
rect 55862 892191 55918 892200
rect 651654 882872 651710 882881
rect 651654 882807 651710 882816
rect 651668 881890 651696 882807
rect 651656 881884 651708 881890
rect 651656 881826 651708 881832
rect 62118 871720 62174 871729
rect 62118 871655 62174 871664
rect 62132 870874 62160 871655
rect 62120 870868 62172 870874
rect 62120 870810 62172 870816
rect 651470 869680 651526 869689
rect 651470 869615 651526 869624
rect 651484 869446 651512 869615
rect 651472 869440 651524 869446
rect 651472 869382 651524 869388
rect 658924 869440 658976 869446
rect 658924 869382 658976 869388
rect 62762 858664 62818 858673
rect 62762 858599 62818 858608
rect 62118 845608 62174 845617
rect 62118 845543 62174 845552
rect 62132 844626 62160 845543
rect 54484 844620 54536 844626
rect 54484 844562 54536 844568
rect 62120 844620 62172 844626
rect 62120 844562 62172 844568
rect 53102 799232 53158 799241
rect 53102 799167 53158 799176
rect 54496 774353 54524 844562
rect 62118 832552 62174 832561
rect 62118 832487 62174 832496
rect 62132 832182 62160 832487
rect 55864 832176 55916 832182
rect 55864 832118 55916 832124
rect 62120 832176 62172 832182
rect 62120 832118 62172 832124
rect 54482 774344 54538 774353
rect 54482 774279 54538 774288
rect 55876 772857 55904 832118
rect 62118 819496 62174 819505
rect 62118 819431 62174 819440
rect 62132 818378 62160 819431
rect 62120 818372 62172 818378
rect 62120 818314 62172 818320
rect 62118 806576 62174 806585
rect 62118 806511 62174 806520
rect 62132 806002 62160 806511
rect 62120 805996 62172 806002
rect 62120 805938 62172 805944
rect 62776 788633 62804 858599
rect 652390 856352 652446 856361
rect 652390 856287 652446 856296
rect 652404 855642 652432 856287
rect 652392 855636 652444 855642
rect 652392 855578 652444 855584
rect 652022 843024 652078 843033
rect 652022 842959 652078 842968
rect 651470 829832 651526 829841
rect 651470 829767 651526 829776
rect 651484 829462 651512 829767
rect 651472 829456 651524 829462
rect 651472 829398 651524 829404
rect 651470 816504 651526 816513
rect 651470 816439 651526 816448
rect 651484 815658 651512 816439
rect 651472 815652 651524 815658
rect 651472 815594 651524 815600
rect 651470 803312 651526 803321
rect 651470 803247 651472 803256
rect 651524 803247 651526 803256
rect 651472 803218 651524 803224
rect 62946 793656 63002 793665
rect 62946 793591 63002 793600
rect 62762 788624 62818 788633
rect 62762 788559 62818 788568
rect 62762 780464 62818 780473
rect 62762 780399 62818 780408
rect 55862 772848 55918 772857
rect 55862 772783 55918 772792
rect 62118 767408 62174 767417
rect 62118 767343 62120 767352
rect 62172 767343 62174 767352
rect 62120 767314 62172 767320
rect 62118 754352 62174 754361
rect 62118 754287 62174 754296
rect 62132 753574 62160 754287
rect 51724 753568 51776 753574
rect 51724 753510 51776 753516
rect 62120 753568 62172 753574
rect 62120 753510 62172 753516
rect 50342 730552 50398 730561
rect 50342 730487 50398 730496
rect 50344 714876 50396 714882
rect 50344 714818 50396 714824
rect 48962 669352 49018 669361
rect 48962 669287 49018 669296
rect 47584 662448 47636 662454
rect 47584 662390 47636 662396
rect 47398 638072 47454 638081
rect 47398 638007 47454 638016
rect 47412 620401 47440 638007
rect 47398 620392 47454 620401
rect 47398 620327 47454 620336
rect 47216 611108 47268 611114
rect 47216 611050 47268 611056
rect 45376 610904 45428 610910
rect 45376 610846 45428 610852
rect 45190 598904 45246 598913
rect 45190 598839 45246 598848
rect 45190 598496 45246 598505
rect 45190 598431 45246 598440
rect 45006 598088 45062 598097
rect 45006 598023 45062 598032
rect 45204 582374 45232 598431
rect 47596 582457 47624 662390
rect 50356 627337 50384 714818
rect 51736 691393 51764 753510
rect 62776 743073 62804 780399
rect 62762 743064 62818 743073
rect 62762 742999 62818 743008
rect 62960 741713 62988 793591
rect 651470 789984 651526 789993
rect 651470 789919 651526 789928
rect 651484 789410 651512 789919
rect 651472 789404 651524 789410
rect 651472 789346 651524 789352
rect 651470 776656 651526 776665
rect 651470 776591 651526 776600
rect 651484 775606 651512 776591
rect 651472 775600 651524 775606
rect 651472 775542 651524 775548
rect 651470 763328 651526 763337
rect 651470 763263 651472 763272
rect 651524 763263 651526 763272
rect 651472 763234 651524 763240
rect 651470 750136 651526 750145
rect 651470 750071 651526 750080
rect 651484 749426 651512 750071
rect 651472 749420 651524 749426
rect 651472 749362 651524 749368
rect 62946 741704 63002 741713
rect 62946 741639 63002 741648
rect 62118 741296 62174 741305
rect 62118 741231 62174 741240
rect 62132 741130 62160 741231
rect 54484 741124 54536 741130
rect 54484 741066 54536 741072
rect 62120 741124 62172 741130
rect 62120 741066 62172 741072
rect 51722 691384 51778 691393
rect 51722 691319 51778 691328
rect 53104 688696 53156 688702
rect 53104 688638 53156 688644
rect 51724 674892 51776 674898
rect 51724 674834 51776 674840
rect 51736 646649 51764 674834
rect 51722 646640 51778 646649
rect 51722 646575 51778 646584
rect 53116 644745 53144 688638
rect 54496 688129 54524 741066
rect 62762 728240 62818 728249
rect 62762 728175 62818 728184
rect 62118 715320 62174 715329
rect 62118 715255 62174 715264
rect 62132 714882 62160 715255
rect 62120 714876 62172 714882
rect 62120 714818 62172 714824
rect 62118 702264 62174 702273
rect 62118 702199 62174 702208
rect 62132 701078 62160 702199
rect 55864 701072 55916 701078
rect 55864 701014 55916 701020
rect 62120 701072 62172 701078
rect 62120 701014 62172 701020
rect 54482 688120 54538 688129
rect 54482 688055 54538 688064
rect 54484 647896 54536 647902
rect 54484 647838 54536 647844
rect 53102 644736 53158 644745
rect 53102 644671 53158 644680
rect 51724 636268 51776 636274
rect 51724 636210 51776 636216
rect 50342 627328 50398 627337
rect 50342 627263 50398 627272
rect 48964 623824 49016 623830
rect 48964 623766 49016 623772
rect 48976 601361 49004 623766
rect 51736 601769 51764 636210
rect 51722 601760 51778 601769
rect 51722 601695 51778 601704
rect 48962 601352 49018 601361
rect 48962 601287 49018 601296
rect 54496 600953 54524 647838
rect 55876 643249 55904 701014
rect 62776 697921 62804 728175
rect 651470 723480 651526 723489
rect 651470 723415 651526 723424
rect 651484 723178 651512 723415
rect 651472 723172 651524 723178
rect 651472 723114 651524 723120
rect 652036 718321 652064 842959
rect 652574 736808 652630 736817
rect 652574 736743 652630 736752
rect 652588 735622 652616 736743
rect 652576 735616 652628 735622
rect 652576 735558 652628 735564
rect 652022 718312 652078 718321
rect 652022 718247 652078 718256
rect 658936 716009 658964 869382
rect 660304 829456 660356 829462
rect 660304 829398 660356 829404
rect 660316 778977 660344 829398
rect 660302 778968 660358 778977
rect 660302 778903 660358 778912
rect 660304 763224 660356 763230
rect 660304 763166 660356 763172
rect 658922 716000 658978 716009
rect 658922 715935 658978 715944
rect 652574 710288 652630 710297
rect 652574 710223 652630 710232
rect 652588 709374 652616 710223
rect 652576 709368 652628 709374
rect 652576 709310 652628 709316
rect 62762 697912 62818 697921
rect 62762 697847 62818 697856
rect 652392 696992 652444 696998
rect 652390 696960 652392 696969
rect 652444 696960 652446 696969
rect 652390 696895 652446 696904
rect 62118 689208 62174 689217
rect 62118 689143 62174 689152
rect 62132 688702 62160 689143
rect 62120 688696 62172 688702
rect 62120 688638 62172 688644
rect 652022 683632 652078 683641
rect 652022 683567 652078 683576
rect 62118 676152 62174 676161
rect 62118 676087 62174 676096
rect 62132 674898 62160 676087
rect 62120 674892 62172 674898
rect 62120 674834 62172 674840
rect 651470 670440 651526 670449
rect 651470 670375 651526 670384
rect 651484 669390 651512 670375
rect 651472 669384 651524 669390
rect 651472 669326 651524 669332
rect 62118 663096 62174 663105
rect 62118 663031 62174 663040
rect 62132 662454 62160 663031
rect 62120 662448 62172 662454
rect 62120 662390 62172 662396
rect 651470 657112 651526 657121
rect 651470 657047 651526 657056
rect 651484 656946 651512 657047
rect 651472 656940 651524 656946
rect 651472 656882 651524 656888
rect 62118 650040 62174 650049
rect 62118 649975 62174 649984
rect 62132 647902 62160 649975
rect 62120 647896 62172 647902
rect 62120 647838 62172 647844
rect 651470 643784 651526 643793
rect 651470 643719 651526 643728
rect 55862 643240 55918 643249
rect 55862 643175 55918 643184
rect 651484 643142 651512 643719
rect 651472 643136 651524 643142
rect 651472 643078 651524 643084
rect 62118 637120 62174 637129
rect 62118 637055 62174 637064
rect 62132 636274 62160 637055
rect 62120 636268 62172 636274
rect 62120 636210 62172 636216
rect 651470 630592 651526 630601
rect 651470 630527 651526 630536
rect 651484 629338 651512 630527
rect 651472 629332 651524 629338
rect 651472 629274 651524 629280
rect 62118 624064 62174 624073
rect 62118 623999 62174 624008
rect 62132 623830 62160 623999
rect 62120 623824 62172 623830
rect 62120 623766 62172 623772
rect 651470 617264 651526 617273
rect 651470 617199 651526 617208
rect 651484 616894 651512 617199
rect 651472 616888 651524 616894
rect 651472 616830 651524 616836
rect 62118 611008 62174 611017
rect 62118 610943 62174 610952
rect 62132 608666 62160 610943
rect 56048 608660 56100 608666
rect 56048 608602 56100 608608
rect 62120 608660 62172 608666
rect 62120 608602 62172 608608
rect 54482 600944 54538 600953
rect 54482 600879 54538 600888
rect 48964 597576 49016 597582
rect 48964 597518 49016 597524
rect 47582 582448 47638 582457
rect 47582 582383 47638 582392
rect 45020 582346 45232 582374
rect 44822 556472 44878 556481
rect 44822 556407 44878 556416
rect 44362 556064 44418 556073
rect 44362 555999 44418 556008
rect 44178 548720 44234 548729
rect 44178 548655 44234 548664
rect 43626 547768 43682 547777
rect 43626 547703 43682 547712
rect 43640 379514 43668 547703
rect 43810 547088 43866 547097
rect 43810 547023 43866 547032
rect 43456 379486 43576 379514
rect 43640 379486 43760 379514
rect 43350 375456 43406 375465
rect 43350 375391 43406 375400
rect 42798 365800 42854 365809
rect 42798 365735 42854 365744
rect 42536 364398 42656 364426
rect 42430 364304 42486 364313
rect 42430 364239 42486 364248
rect 42444 363950 42472 364239
rect 42182 363922 42472 363950
rect 41786 363624 41842 363633
rect 41786 363559 41842 363568
rect 41800 363256 41828 363559
rect 42628 362794 42656 364398
rect 42168 362766 42288 362794
rect 42168 362712 42196 362766
rect 42260 362726 42288 362766
rect 42536 362766 42656 362794
rect 42536 362726 42564 362766
rect 42260 362698 42564 362726
rect 41800 360097 41828 360264
rect 41786 360088 41842 360097
rect 41786 360023 41842 360032
rect 42154 359952 42210 359961
rect 42154 359887 42210 359896
rect 42168 359584 42196 359887
rect 41786 359408 41842 359417
rect 41786 359343 41842 359352
rect 41800 358972 41828 359343
rect 41786 358728 41842 358737
rect 41786 358663 41842 358672
rect 41800 358428 41828 358663
rect 42430 356960 42486 356969
rect 42430 356895 42486 356904
rect 42168 356425 42196 356592
rect 42154 356416 42210 356425
rect 42154 356351 42210 356360
rect 42444 355926 42472 356895
rect 42182 355898 42472 355926
rect 43364 355881 43392 375391
rect 43350 355872 43406 355881
rect 43350 355807 43406 355816
rect 41878 355736 41934 355745
rect 41878 355671 41934 355680
rect 41892 355300 41920 355671
rect 43548 355314 43576 379486
rect 43732 355586 43760 379486
rect 43824 355722 43852 547023
rect 44192 536897 44220 548655
rect 44178 536888 44234 536897
rect 44178 536823 44234 536832
rect 44376 428913 44404 555999
rect 45020 555665 45048 582346
rect 48976 557841 49004 597518
rect 51724 583772 51776 583778
rect 51724 583714 51776 583720
rect 48962 557832 49018 557841
rect 48962 557767 49018 557776
rect 51736 557569 51764 583714
rect 55864 558136 55916 558142
rect 55864 558078 55916 558084
rect 51722 557560 51778 557569
rect 51722 557495 51778 557504
rect 45558 556880 45614 556889
rect 45558 556815 45614 556824
rect 45006 555656 45062 555665
rect 45006 555591 45062 555600
rect 44822 555248 44878 555257
rect 44822 555183 44878 555192
rect 44638 554432 44694 554441
rect 44638 554367 44694 554376
rect 44362 428904 44418 428913
rect 44362 428839 44418 428848
rect 44178 428496 44234 428505
rect 44178 428431 44234 428440
rect 43994 419520 44050 419529
rect 43994 419455 44050 419464
rect 44008 355858 44036 419455
rect 44192 385665 44220 428431
rect 44454 427680 44510 427689
rect 44454 427615 44510 427624
rect 44178 385656 44234 385665
rect 44178 385591 44234 385600
rect 44468 384849 44496 427615
rect 44652 427281 44680 554367
rect 44836 428097 44864 555183
rect 45006 551576 45062 551585
rect 45006 551511 45062 551520
rect 45020 529689 45048 551511
rect 45190 550760 45246 550769
rect 45190 550695 45246 550704
rect 45204 532817 45232 550695
rect 45374 549128 45430 549137
rect 45374 549063 45430 549072
rect 45388 537169 45416 549063
rect 45374 537160 45430 537169
rect 45374 537095 45430 537104
rect 45190 532808 45246 532817
rect 45190 532743 45246 532752
rect 45006 529680 45062 529689
rect 45006 529615 45062 529624
rect 45572 429729 45600 556815
rect 47584 545148 47636 545154
rect 47584 545090 47636 545096
rect 46204 506524 46256 506530
rect 46204 506466 46256 506472
rect 45558 429720 45614 429729
rect 45558 429655 45614 429664
rect 45006 429312 45062 429321
rect 45006 429247 45062 429256
rect 44822 428088 44878 428097
rect 44822 428023 44878 428032
rect 44638 427272 44694 427281
rect 44638 427207 44694 427216
rect 44638 421560 44694 421569
rect 44638 421495 44694 421504
rect 44652 407017 44680 421495
rect 44822 420744 44878 420753
rect 44822 420679 44878 420688
rect 44638 407008 44694 407017
rect 44638 406943 44694 406952
rect 44638 385248 44694 385257
rect 44638 385183 44694 385192
rect 44454 384840 44510 384849
rect 44454 384775 44510 384784
rect 44652 379514 44680 385183
rect 44836 379514 44864 420679
rect 45020 386753 45048 429247
rect 45190 426864 45246 426873
rect 45190 426799 45246 426808
rect 45006 386744 45062 386753
rect 45006 386679 45062 386688
rect 45006 384432 45062 384441
rect 45006 384367 45062 384376
rect 44652 379486 44772 379514
rect 44836 379486 44956 379514
rect 44454 377904 44510 377913
rect 44454 377839 44510 377848
rect 44270 377496 44326 377505
rect 44270 377431 44326 377440
rect 44284 356697 44312 377431
rect 44468 364993 44496 377839
rect 44454 364984 44510 364993
rect 44454 364919 44510 364928
rect 44744 360194 44772 379486
rect 44744 360166 44864 360194
rect 44270 356688 44326 356697
rect 44270 356623 44326 356632
rect 44008 355830 44312 355858
rect 44284 355722 44312 355830
rect 43824 355694 44220 355722
rect 44284 355706 44680 355722
rect 44284 355700 44692 355706
rect 44284 355694 44640 355700
rect 44192 355586 44220 355694
rect 44640 355642 44692 355648
rect 43732 355558 43944 355586
rect 44192 355558 44772 355586
rect 43916 355450 43944 355558
rect 43916 355422 44128 355450
rect 43548 355286 44036 355314
rect 44008 354634 44036 355286
rect 44100 354906 44128 355422
rect 44100 354890 44615 354906
rect 44100 354884 44627 354890
rect 44100 354878 44575 354884
rect 44575 354826 44627 354832
rect 44575 354680 44627 354686
rect 44008 354628 44575 354634
rect 44008 354622 44627 354628
rect 44008 354606 44615 354622
rect 44744 354498 44772 355558
rect 44836 354634 44864 360166
rect 44928 357434 44956 379486
rect 45020 360194 45048 384367
rect 45204 384033 45232 426799
rect 45558 426456 45614 426465
rect 45558 426391 45614 426400
rect 45374 422376 45430 422385
rect 45374 422311 45430 422320
rect 45388 405657 45416 422311
rect 45374 405648 45430 405657
rect 45374 405583 45430 405592
rect 45572 399809 45600 426391
rect 45558 399800 45614 399809
rect 45558 399735 45614 399744
rect 45374 386064 45430 386073
rect 45374 385999 45430 386008
rect 45190 384024 45246 384033
rect 45190 383959 45246 383968
rect 45190 383616 45246 383625
rect 45190 383551 45246 383560
rect 45204 379514 45232 383551
rect 45204 379486 45324 379514
rect 45020 360166 45232 360194
rect 44928 357406 45048 357434
rect 45020 355842 45048 357406
rect 45008 355836 45060 355842
rect 45008 355778 45060 355784
rect 44836 354606 44956 354634
rect 44744 354482 44839 354498
rect 44744 354476 44851 354482
rect 44744 354470 44799 354476
rect 44799 354418 44851 354424
rect 44686 354340 44738 354346
rect 44686 354282 44738 354288
rect 43902 354240 43958 354249
rect 44698 354226 44726 354282
rect 43958 354198 44726 354226
rect 43902 354175 43958 354184
rect 44730 353832 44786 353841
rect 44928 353818 44956 354606
rect 45204 354090 45232 360166
rect 44786 353790 44956 353818
rect 45020 354062 45232 354090
rect 44730 353767 44786 353776
rect 28538 351248 28594 351257
rect 28538 351183 28594 351192
rect 8588 345100 8616 345236
rect 9048 345100 9076 345236
rect 9508 345100 9536 345236
rect 9968 345100 9996 345236
rect 10428 345100 10456 345236
rect 10888 345100 10916 345236
rect 11348 345100 11376 345236
rect 11808 345100 11836 345236
rect 12268 345100 12296 345236
rect 12728 345100 12756 345236
rect 13188 345100 13216 345236
rect 13648 345100 13676 345236
rect 14108 345100 14136 345236
rect 28552 343913 28580 351183
rect 40222 345400 40278 345409
rect 40222 345335 40278 345344
rect 40236 345098 40264 345335
rect 28908 345092 28960 345098
rect 28908 345034 28960 345040
rect 40224 345092 40276 345098
rect 40224 345034 40276 345040
rect 28920 344321 28948 345034
rect 28906 344312 28962 344321
rect 28906 344247 28962 344256
rect 28538 343904 28594 343913
rect 28538 343839 28594 343848
rect 45020 341737 45048 354062
rect 45296 345014 45324 379486
rect 45204 344986 45324 345014
rect 45006 341728 45062 341737
rect 45006 341663 45062 341672
rect 45204 340921 45232 344986
rect 45388 343369 45416 385999
rect 45558 380760 45614 380769
rect 45558 380695 45614 380704
rect 45572 356969 45600 380695
rect 45742 379944 45798 379953
rect 45742 379879 45798 379888
rect 45756 359961 45784 379879
rect 46216 367033 46244 506466
rect 47596 430137 47624 545090
rect 50344 532772 50396 532778
rect 50344 532714 50396 532720
rect 48964 491972 49016 491978
rect 48964 491914 49016 491920
rect 47582 430128 47638 430137
rect 47582 430063 47638 430072
rect 46938 423600 46994 423609
rect 46938 423535 46994 423544
rect 46952 400217 46980 423535
rect 47584 415472 47636 415478
rect 47584 415414 47636 415420
rect 46938 400208 46994 400217
rect 46938 400143 46994 400152
rect 46938 383208 46994 383217
rect 46938 383143 46994 383152
rect 46202 367024 46258 367033
rect 46202 366959 46258 366968
rect 46388 362976 46440 362982
rect 46388 362918 46440 362924
rect 45742 359952 45798 359961
rect 45742 359887 45798 359896
rect 45558 356960 45614 356969
rect 45558 356895 45614 356904
rect 45650 356688 45706 356697
rect 45480 356646 45650 356674
rect 45480 353274 45508 356646
rect 45650 356623 45706 356632
rect 45926 355872 45982 355881
rect 45652 355836 45704 355842
rect 45926 355807 45982 355816
rect 45652 355778 45704 355784
rect 45664 354074 45692 355778
rect 45652 354068 45704 354074
rect 45652 354010 45704 354016
rect 45940 353802 45968 355807
rect 45928 353796 45980 353802
rect 45928 353738 45980 353744
rect 45480 353258 45600 353274
rect 45480 353252 45612 353258
rect 45480 353246 45560 353252
rect 45560 353194 45612 353200
rect 45374 343360 45430 343369
rect 45374 343295 45430 343304
rect 45190 340912 45246 340921
rect 45190 340847 45246 340856
rect 45558 340096 45614 340105
rect 45558 340031 45614 340040
rect 35806 339824 35862 339833
rect 35806 339759 35862 339768
rect 35820 339522 35848 339759
rect 35808 339516 35860 339522
rect 35808 339458 35860 339464
rect 37924 339516 37976 339522
rect 37924 339458 37976 339464
rect 35806 339008 35862 339017
rect 35806 338943 35862 338952
rect 31022 338600 31078 338609
rect 31022 338535 31078 338544
rect 31036 329089 31064 338535
rect 35820 338162 35848 338943
rect 35808 338156 35860 338162
rect 35808 338098 35860 338104
rect 36544 338156 36596 338162
rect 36544 338098 36596 338104
rect 31022 329080 31078 329089
rect 31022 329015 31078 329024
rect 36556 328409 36584 338098
rect 37936 334529 37964 339458
rect 45374 337240 45430 337249
rect 45374 337175 45430 337184
rect 45388 337090 45416 337175
rect 45388 337062 45508 337090
rect 42890 334656 42946 334665
rect 42890 334591 42946 334600
rect 43258 334656 43314 334665
rect 43258 334591 43314 334600
rect 44178 334656 44234 334665
rect 44178 334591 44234 334600
rect 37922 334520 37978 334529
rect 37922 334455 37978 334464
rect 42614 334384 42670 334393
rect 42670 334342 42840 334370
rect 42614 334319 42670 334328
rect 36542 328400 36598 328409
rect 36542 328335 36598 328344
rect 41786 326768 41842 326777
rect 41786 326703 41842 326712
rect 41800 326264 41828 326703
rect 42614 326496 42670 326505
rect 42614 326431 42670 326440
rect 41786 325408 41842 325417
rect 41786 325343 41842 325352
rect 41800 325040 41828 325343
rect 41878 324728 41934 324737
rect 41878 324663 41934 324672
rect 41892 324428 41920 324663
rect 42182 323734 42472 323762
rect 42062 322824 42118 322833
rect 42062 322759 42118 322768
rect 42076 322592 42104 322759
rect 42444 321473 42472 323734
rect 42430 321464 42486 321473
rect 42430 321399 42486 321408
rect 42182 321354 42288 321382
rect 42260 321314 42288 321354
rect 42628 321314 42656 326431
rect 42260 321286 42656 321314
rect 41786 321056 41842 321065
rect 41786 320991 41842 321000
rect 41800 320725 41828 320991
rect 42812 320226 42840 334342
rect 42904 328454 42932 334591
rect 42904 328426 43024 328454
rect 42996 326505 43024 328426
rect 42982 326496 43038 326505
rect 42982 326431 43038 326440
rect 43272 322833 43300 334591
rect 43258 322824 43314 322833
rect 43258 322759 43314 322768
rect 42536 320198 42840 320226
rect 42536 320090 42564 320198
rect 42182 320062 42564 320090
rect 42182 319518 42472 319546
rect 42444 319025 42472 319518
rect 42430 319016 42486 319025
rect 42430 318951 42486 318960
rect 44192 317393 44220 334591
rect 42430 317384 42486 317393
rect 42430 317319 42486 317328
rect 44178 317384 44234 317393
rect 44178 317319 44234 317328
rect 42444 317059 42472 317319
rect 42182 317031 42472 317059
rect 42430 316432 42486 316441
rect 42182 316390 42430 316418
rect 42430 316367 42486 316376
rect 45480 316033 45508 337062
rect 45572 331214 45600 340031
rect 46204 336796 46256 336802
rect 46204 336738 46256 336744
rect 45572 331186 45692 331214
rect 42154 316024 42210 316033
rect 42154 315959 42210 315968
rect 45466 316024 45522 316033
rect 45466 315959 45522 315968
rect 42168 315757 42196 315959
rect 41786 315616 41842 315625
rect 41786 315551 41842 315560
rect 41800 315180 41828 315551
rect 45664 313721 45692 331186
rect 42154 313712 42210 313721
rect 42154 313647 42210 313656
rect 45650 313712 45706 313721
rect 45650 313647 45706 313656
rect 42168 313344 42196 313647
rect 42430 312760 42486 312769
rect 42182 312718 42430 312746
rect 42430 312695 42486 312704
rect 41786 312624 41842 312633
rect 41786 312559 41842 312568
rect 41800 312052 41828 312559
rect 44730 311808 44786 311817
rect 44730 311743 44786 311752
rect 44178 311536 44234 311545
rect 44178 311471 44234 311480
rect 41786 303104 41842 303113
rect 41786 303039 41842 303048
rect 8588 301988 8616 302124
rect 9048 301988 9076 302124
rect 9508 301988 9536 302124
rect 9968 301988 9996 302124
rect 10428 301988 10456 302124
rect 10888 301988 10916 302124
rect 11348 301988 11376 302124
rect 11808 301988 11836 302124
rect 12268 301988 12296 302124
rect 12728 301988 12756 302124
rect 13188 301988 13216 302124
rect 13648 301988 13676 302124
rect 14108 301988 14136 302124
rect 41800 300937 41828 303039
rect 41786 300928 41842 300937
rect 41786 300863 41842 300872
rect 44192 299305 44220 311471
rect 44546 311264 44602 311273
rect 44546 311199 44602 311208
rect 44178 299296 44234 299305
rect 44178 299231 44234 299240
rect 44270 298888 44326 298897
rect 44270 298823 44326 298832
rect 43258 298072 43314 298081
rect 43258 298007 43314 298016
rect 42890 297256 42946 297265
rect 42890 297191 42946 297200
rect 41786 296848 41842 296857
rect 41786 296783 41842 296792
rect 32402 294808 32458 294817
rect 32402 294743 32458 294752
rect 32416 284986 32444 294743
rect 41800 292777 41828 296783
rect 42062 296032 42118 296041
rect 42062 295967 42118 295976
rect 41786 292768 41842 292777
rect 41786 292703 41842 292712
rect 42076 292369 42104 295967
rect 42062 292360 42118 292369
rect 42062 292295 42118 292304
rect 42246 291136 42302 291145
rect 42246 291071 42302 291080
rect 42062 290456 42118 290465
rect 42062 290391 42118 290400
rect 41326 290320 41382 290329
rect 41326 290255 41382 290264
rect 41340 285122 41368 290255
rect 42076 289921 42104 290391
rect 42260 289921 42288 291071
rect 42062 289912 42118 289921
rect 42062 289847 42118 289856
rect 42246 289912 42302 289921
rect 42246 289847 42302 289856
rect 41708 285122 42380 285138
rect 41328 285116 41380 285122
rect 41328 285058 41380 285064
rect 41696 285116 42380 285122
rect 41748 285110 42380 285116
rect 41696 285058 41748 285064
rect 32404 284980 32456 284986
rect 32404 284922 32456 284928
rect 41696 284980 41748 284986
rect 41696 284922 41748 284928
rect 41708 284866 41736 284922
rect 41708 284838 42288 284866
rect 42260 283059 42288 284838
rect 42182 283031 42288 283059
rect 42352 281874 42380 285110
rect 42182 281846 42380 281874
rect 41970 281480 42026 281489
rect 41970 281415 42026 281424
rect 41984 281180 42012 281415
rect 42182 280554 42472 280582
rect 42154 279848 42210 279857
rect 42154 279783 42210 279792
rect 42168 279344 42196 279783
rect 42444 278769 42472 280554
rect 42430 278760 42486 278769
rect 42430 278695 42486 278704
rect 42430 278216 42486 278225
rect 42168 278066 42196 278188
rect 42260 278174 42430 278202
rect 42260 278066 42288 278174
rect 42430 278151 42486 278160
rect 42168 278038 42288 278066
rect 41786 277944 41842 277953
rect 41786 277879 41842 277888
rect 41800 277508 41828 277879
rect 42338 277672 42394 277681
rect 42338 277607 42394 277616
rect 42062 277128 42118 277137
rect 42062 277063 42118 277072
rect 42076 276896 42104 277063
rect 42062 276584 42118 276593
rect 42062 276519 42118 276528
rect 42076 276352 42104 276519
rect 41786 274272 41842 274281
rect 41786 274207 41842 274216
rect 41800 273836 41828 274207
rect 42062 273456 42118 273465
rect 42062 273391 42118 273400
rect 42076 273224 42104 273391
rect 42062 272912 42118 272921
rect 42062 272847 42118 272856
rect 42076 272544 42104 272847
rect 42352 272014 42380 277607
rect 42182 271986 42380 272014
rect 41786 270464 41842 270473
rect 41786 270399 41842 270408
rect 42430 270464 42486 270473
rect 42430 270399 42486 270408
rect 41800 270164 41828 270399
rect 42444 269535 42472 270399
rect 42182 269507 42472 269535
rect 41786 269104 41842 269113
rect 41786 269039 41842 269048
rect 41800 268872 41828 269039
rect 42904 267734 42932 297191
rect 43074 293584 43130 293593
rect 43074 293519 43130 293528
rect 43088 273465 43116 293519
rect 43074 273456 43130 273465
rect 43074 273391 43130 273400
rect 42904 267706 43116 267734
rect 40682 267064 40738 267073
rect 40682 266999 40738 267008
rect 8588 258740 8616 258876
rect 9048 258740 9076 258876
rect 9508 258740 9536 258876
rect 9968 258740 9996 258876
rect 10428 258740 10456 258876
rect 10888 258740 10916 258876
rect 11348 258740 11376 258876
rect 11808 258740 11836 258876
rect 12268 258740 12296 258876
rect 12728 258740 12756 258876
rect 13188 258740 13216 258876
rect 13648 258740 13676 258876
rect 14108 258740 14136 258876
rect 35806 257136 35862 257145
rect 35806 257071 35862 257080
rect 35820 256766 35848 257071
rect 40696 256766 40724 266999
rect 35808 256760 35860 256766
rect 35808 256702 35860 256708
rect 40684 256760 40736 256766
rect 40684 256702 40736 256708
rect 42890 254824 42946 254833
rect 42890 254759 42946 254768
rect 35622 253464 35678 253473
rect 35622 253399 35678 253408
rect 35438 253056 35494 253065
rect 35438 252991 35494 253000
rect 35452 252618 35480 252991
rect 35636 252890 35664 253399
rect 35806 253056 35862 253065
rect 35806 252991 35862 253000
rect 35624 252884 35676 252890
rect 35624 252826 35676 252832
rect 35820 252754 35848 252991
rect 41696 252884 41748 252890
rect 41696 252826 41748 252832
rect 41708 252770 41736 252826
rect 35808 252748 35860 252754
rect 35808 252690 35860 252696
rect 40684 252748 40736 252754
rect 41708 252742 41920 252770
rect 40684 252690 40736 252696
rect 35440 252612 35492 252618
rect 35440 252554 35492 252560
rect 35806 252240 35862 252249
rect 35806 252175 35862 252184
rect 35820 251258 35848 252175
rect 35808 251252 35860 251258
rect 35808 251194 35860 251200
rect 36544 251252 36596 251258
rect 36544 251194 36596 251200
rect 36556 242894 36584 251194
rect 36544 242888 36596 242894
rect 36544 242830 36596 242836
rect 40696 242593 40724 252690
rect 41696 252612 41748 252618
rect 41696 252554 41748 252560
rect 41708 248414 41736 252554
rect 41892 252498 41920 252742
rect 41892 252470 42472 252498
rect 42444 248414 42472 252470
rect 41708 248386 42288 248414
rect 42444 248386 42564 248414
rect 41696 242888 41748 242894
rect 41694 242856 41696 242865
rect 41748 242856 41750 242865
rect 41694 242791 41750 242800
rect 40682 242584 40738 242593
rect 40682 242519 40738 242528
rect 41786 240136 41842 240145
rect 41786 240071 41842 240080
rect 41800 239836 41828 240071
rect 42076 238513 42104 238649
rect 42062 238504 42118 238513
rect 42062 238439 42118 238448
rect 42260 238014 42288 248386
rect 42536 238762 42564 248386
rect 42706 242856 42762 242865
rect 42706 242791 42762 242800
rect 42536 238734 42656 238762
rect 42182 237986 42288 238014
rect 42628 237538 42656 238734
rect 42536 237510 42656 237538
rect 42536 237425 42564 237510
rect 42522 237416 42578 237425
rect 42522 237351 42578 237360
rect 41800 235929 41828 236164
rect 41786 235920 41842 235929
rect 41786 235855 41842 235864
rect 42430 235920 42486 235929
rect 42430 235855 42486 235864
rect 42444 234983 42472 235855
rect 42182 234955 42472 234983
rect 42720 234614 42748 242791
rect 42536 234586 42748 234614
rect 42246 234560 42302 234569
rect 42246 234495 42302 234504
rect 42260 234342 42288 234495
rect 42182 234314 42288 234342
rect 42338 234152 42394 234161
rect 42338 234087 42394 234096
rect 42352 233695 42380 234087
rect 42182 233667 42380 233695
rect 42338 233200 42394 233209
rect 42168 233158 42338 233186
rect 42168 233104 42196 233158
rect 42338 233135 42394 233144
rect 42338 231840 42394 231849
rect 42338 231775 42394 231784
rect 42352 230670 42380 231775
rect 42182 230642 42380 230670
rect 42154 230344 42210 230353
rect 42154 230279 42210 230288
rect 42168 229976 42196 230279
rect 42338 229392 42394 229401
rect 42182 229350 42338 229378
rect 42338 229327 42394 229336
rect 42536 228834 42564 234586
rect 42182 228806 42564 228834
rect 42430 227624 42486 227633
rect 42430 227559 42486 227568
rect 41970 227352 42026 227361
rect 41970 227287 42026 227296
rect 41984 226984 42012 227287
rect 42168 226358 42288 226386
rect 42168 226304 42196 226358
rect 42260 226318 42288 226358
rect 42444 226318 42472 227559
rect 42904 226522 42932 254759
rect 43088 254425 43116 267706
rect 43272 255241 43300 298007
rect 43442 294400 43498 294409
rect 43442 294335 43498 294344
rect 43456 270473 43484 294335
rect 43626 293176 43682 293185
rect 43626 293111 43682 293120
rect 43640 279857 43668 293111
rect 43810 291952 43866 291961
rect 43810 291887 43866 291896
rect 43626 279848 43682 279857
rect 43626 279783 43682 279792
rect 43824 277137 43852 291887
rect 43810 277128 43866 277137
rect 43810 277063 43866 277072
rect 43442 270464 43498 270473
rect 43442 270399 43498 270408
rect 43718 256456 43774 256465
rect 43718 256391 43774 256400
rect 43442 255640 43498 255649
rect 43442 255575 43498 255584
rect 43258 255232 43314 255241
rect 43258 255167 43314 255176
rect 43456 255082 43484 255575
rect 43364 255054 43484 255082
rect 43074 254416 43130 254425
rect 43074 254351 43130 254360
rect 43074 249112 43130 249121
rect 43074 249047 43130 249056
rect 43088 231849 43116 249047
rect 43364 248414 43392 255054
rect 43534 251152 43590 251161
rect 43534 251087 43590 251096
rect 43364 248386 43484 248414
rect 43258 242584 43314 242593
rect 43258 242519 43314 242528
rect 43074 231840 43130 231849
rect 43074 231775 43130 231784
rect 43272 226522 43300 242519
rect 43456 234614 43484 248386
rect 42904 226494 43024 226522
rect 42260 226290 42472 226318
rect 42430 225720 42486 225729
rect 42182 225678 42430 225706
rect 42430 225655 42486 225664
rect 42996 224954 43024 226494
rect 43180 226494 43300 226522
rect 43364 234586 43484 234614
rect 43180 225729 43208 226494
rect 43166 225720 43222 225729
rect 43166 225655 43222 225664
rect 42904 224926 43024 224954
rect 43364 224954 43392 234586
rect 43548 227633 43576 251087
rect 43534 227624 43590 227633
rect 43534 227559 43590 227568
rect 43364 224926 43484 224954
rect 40682 222864 40738 222873
rect 40682 222799 40738 222808
rect 35530 217968 35586 217977
rect 35530 217903 35586 217912
rect 8588 215492 8616 215628
rect 9048 215492 9076 215628
rect 9508 215492 9536 215628
rect 9968 215492 9996 215628
rect 10428 215492 10456 215628
rect 10888 215492 10916 215628
rect 11348 215492 11376 215628
rect 11808 215492 11836 215628
rect 12268 215492 12296 215628
rect 12728 215492 12756 215628
rect 13188 215492 13216 215628
rect 13648 215492 13676 215628
rect 14108 215492 14136 215628
rect 35544 214305 35572 217903
rect 35530 214296 35586 214305
rect 35530 214231 35586 214240
rect 35806 214296 35862 214305
rect 35806 214231 35862 214240
rect 35820 213994 35848 214231
rect 40696 213994 40724 222799
rect 35808 213988 35860 213994
rect 35808 213930 35860 213936
rect 40684 213988 40736 213994
rect 40684 213930 40736 213936
rect 42904 212129 42932 224926
rect 43456 212945 43484 224926
rect 43732 213761 43760 256391
rect 44284 256057 44312 298823
rect 44560 298489 44588 311199
rect 44744 300121 44772 311743
rect 44730 300112 44786 300121
rect 44730 300047 44786 300056
rect 44730 299704 44786 299713
rect 44730 299639 44786 299648
rect 44546 298480 44602 298489
rect 44546 298415 44602 298424
rect 44744 296714 44772 299639
rect 45468 298172 45520 298178
rect 45468 298114 45520 298120
rect 45480 296714 45508 298114
rect 44652 296686 44772 296714
rect 44836 296686 45508 296714
rect 44454 291544 44510 291553
rect 44454 291479 44510 291488
rect 44468 278225 44496 291479
rect 44454 278216 44510 278225
rect 44454 278151 44510 278160
rect 44652 256873 44680 296686
rect 44638 256864 44694 256873
rect 44638 256799 44694 256808
rect 44270 256048 44326 256057
rect 44270 255983 44326 255992
rect 44178 254008 44234 254017
rect 44178 253943 44234 253952
rect 43718 213752 43774 213761
rect 43718 213687 43774 213696
rect 43442 212936 43498 212945
rect 43442 212871 43498 212880
rect 43442 212528 43498 212537
rect 43442 212463 43498 212472
rect 42890 212120 42946 212129
rect 42890 212055 42946 212064
rect 35806 211440 35862 211449
rect 35806 211375 35862 211384
rect 35820 211206 35848 211375
rect 35808 211200 35860 211206
rect 35808 211142 35860 211148
rect 41696 211200 41748 211206
rect 41696 211142 41748 211148
rect 41708 209001 41736 211142
rect 42798 209400 42854 209409
rect 42798 209335 42854 209344
rect 35806 208992 35862 209001
rect 35806 208927 35862 208936
rect 41694 208992 41750 209001
rect 41694 208927 41750 208936
rect 35820 208418 35848 208927
rect 35808 208412 35860 208418
rect 35808 208354 35860 208360
rect 40040 208412 40092 208418
rect 40040 208354 40092 208360
rect 40052 207777 40080 208354
rect 40038 207768 40094 207777
rect 40038 207703 40094 207712
rect 35622 204096 35678 204105
rect 35622 204031 35678 204040
rect 35636 202201 35664 204031
rect 35806 203688 35862 203697
rect 35806 203623 35862 203632
rect 35820 202910 35848 203623
rect 35808 202904 35860 202910
rect 35808 202846 35860 202852
rect 37924 202904 37976 202910
rect 37924 202846 37976 202852
rect 35622 202192 35678 202201
rect 35622 202127 35678 202136
rect 37936 197849 37964 202846
rect 37922 197840 37978 197849
rect 37922 197775 37978 197784
rect 41786 197160 41842 197169
rect 41786 197095 41842 197104
rect 41800 196656 41828 197095
rect 41878 195800 41934 195809
rect 41878 195735 41934 195744
rect 41892 195432 41920 195735
rect 41786 195256 41842 195265
rect 41786 195191 41842 195200
rect 41800 194820 41828 195191
rect 42246 194984 42302 194993
rect 42246 194919 42302 194928
rect 42260 193225 42288 194919
rect 42246 193216 42302 193225
rect 42246 193151 42302 193160
rect 42168 192930 42196 192984
rect 42338 192944 42394 192953
rect 42168 192902 42338 192930
rect 42338 192879 42394 192888
rect 42168 191706 42196 191760
rect 42338 191720 42394 191729
rect 42168 191678 42338 191706
rect 42338 191655 42394 191664
rect 42430 191176 42486 191185
rect 42168 191026 42196 191148
rect 42260 191134 42430 191162
rect 42260 191026 42288 191134
rect 42430 191111 42486 191120
rect 42168 190998 42288 191026
rect 42430 190496 42486 190505
rect 42182 190454 42430 190482
rect 42430 190431 42486 190440
rect 42430 189952 42486 189961
rect 42182 189910 42430 189938
rect 42430 189887 42486 189896
rect 42430 187640 42486 187649
rect 42430 187575 42486 187584
rect 42444 187459 42472 187575
rect 42182 187431 42472 187459
rect 41786 187232 41842 187241
rect 41786 187167 41842 187176
rect 41800 186796 41828 187167
rect 42338 186280 42394 186289
rect 42338 186215 42394 186224
rect 42168 186017 42196 186184
rect 42154 186008 42210 186017
rect 42154 185943 42210 185952
rect 42352 185619 42380 186215
rect 42182 185591 42380 185619
rect 42430 184920 42486 184929
rect 42430 184855 42486 184864
rect 42444 183779 42472 184855
rect 42182 183751 42472 183779
rect 42430 183152 42486 183161
rect 42182 183110 42430 183138
rect 42430 183087 42486 183096
rect 42812 182491 42840 209335
rect 43258 208040 43314 208049
rect 43258 207975 43314 207984
rect 42982 206408 43038 206417
rect 42982 206343 43038 206352
rect 42996 191185 43024 206343
rect 42982 191176 43038 191185
rect 42982 191111 43038 191120
rect 43272 183161 43300 207975
rect 43456 206281 43484 212463
rect 44192 211313 44220 253943
rect 44638 251968 44694 251977
rect 44638 251903 44694 251912
rect 44652 251818 44680 251903
rect 44652 251790 44772 251818
rect 44546 248704 44602 248713
rect 44546 248639 44602 248648
rect 44362 248296 44418 248305
rect 44362 248231 44418 248240
rect 44376 235929 44404 248231
rect 44362 235920 44418 235929
rect 44362 235855 44418 235864
rect 44560 234161 44588 248639
rect 44744 238754 44772 251790
rect 44652 238726 44772 238754
rect 44652 234614 44680 238726
rect 44652 234586 44772 234614
rect 44546 234152 44602 234161
rect 44546 234087 44602 234096
rect 44546 233200 44602 233209
rect 44744 233186 44772 234586
rect 44602 233158 44772 233186
rect 44546 233135 44602 233144
rect 44836 214985 44864 296686
rect 45006 295216 45062 295225
rect 45006 295151 45062 295160
rect 45020 276593 45048 295151
rect 45190 293992 45246 294001
rect 45190 293927 45246 293936
rect 45006 276584 45062 276593
rect 45006 276519 45062 276528
rect 45204 272921 45232 293927
rect 45190 272912 45246 272921
rect 45190 272847 45246 272856
rect 46216 257961 46244 336738
rect 46400 303113 46428 362918
rect 46952 356425 46980 383143
rect 47122 379128 47178 379137
rect 47122 379063 47178 379072
rect 47136 364313 47164 379063
rect 47122 364304 47178 364313
rect 47122 364239 47178 364248
rect 46938 356416 46994 356425
rect 46938 356351 46994 356360
rect 47596 345409 47624 415414
rect 47768 389292 47820 389298
rect 47768 389234 47820 389240
rect 47582 345400 47638 345409
rect 47582 345335 47638 345344
rect 46938 338464 46994 338473
rect 46938 338399 46994 338408
rect 46952 319025 46980 338399
rect 47582 333160 47638 333169
rect 47582 333095 47638 333104
rect 46938 319016 46994 319025
rect 46938 318951 46994 318960
rect 46386 303104 46442 303113
rect 46386 303039 46442 303048
rect 46202 257952 46258 257961
rect 46202 257887 46258 257896
rect 45834 250744 45890 250753
rect 45834 250679 45890 250688
rect 45558 250336 45614 250345
rect 45558 250271 45614 250280
rect 45572 230353 45600 250271
rect 45558 230344 45614 230353
rect 45558 230279 45614 230288
rect 45848 229401 45876 250679
rect 46018 249520 46074 249529
rect 46018 249455 46074 249464
rect 46032 234569 46060 249455
rect 46202 247888 46258 247897
rect 46202 247823 46258 247832
rect 46018 234560 46074 234569
rect 46018 234495 46074 234504
rect 45834 229392 45890 229401
rect 45834 229327 45890 229336
rect 44822 214976 44878 214985
rect 44822 214911 44878 214920
rect 44178 211304 44234 211313
rect 44178 211239 44234 211248
rect 44178 210488 44234 210497
rect 44178 210423 44234 210432
rect 43810 206816 43866 206825
rect 43810 206751 43866 206760
rect 43442 206272 43498 206281
rect 43442 206207 43498 206216
rect 43626 205592 43682 205601
rect 43626 205527 43682 205536
rect 43442 202192 43498 202201
rect 43442 202127 43498 202136
rect 43258 183152 43314 183161
rect 43258 183087 43314 183096
rect 42182 182463 42840 182491
rect 43456 42838 43484 202127
rect 43640 190505 43668 205527
rect 43824 192953 43852 206751
rect 43994 205184 44050 205193
rect 43994 205119 44050 205128
rect 43810 192944 43866 192953
rect 43810 192879 43866 192888
rect 44008 191729 44036 205119
rect 43994 191720 44050 191729
rect 43994 191655 44050 191664
rect 43626 190496 43682 190505
rect 43626 190431 43682 190440
rect 44192 184929 44220 210423
rect 44546 208584 44602 208593
rect 44546 208519 44602 208528
rect 44362 206000 44418 206009
rect 44362 205935 44418 205944
rect 44376 187649 44404 205935
rect 44560 189961 44588 208519
rect 44822 204776 44878 204785
rect 44822 204711 44878 204720
rect 44546 189952 44602 189961
rect 44546 189887 44602 189896
rect 44362 187640 44418 187649
rect 44362 187575 44418 187584
rect 44178 184920 44234 184929
rect 44178 184855 44234 184864
rect 44836 74534 44864 204711
rect 44836 74506 45508 74534
rect 45480 50386 45508 74506
rect 46216 53106 46244 247823
rect 46938 247072 46994 247081
rect 46938 247007 46994 247016
rect 46952 238513 46980 247007
rect 46938 238504 46994 238513
rect 46938 238439 46994 238448
rect 46386 203552 46442 203561
rect 46386 203487 46442 203496
rect 46204 53100 46256 53106
rect 46204 53042 46256 53048
rect 46400 51746 46428 203487
rect 46388 51740 46440 51746
rect 46388 51682 46440 51688
rect 45468 50380 45520 50386
rect 45468 50322 45520 50328
rect 47596 49026 47624 333095
rect 47780 300529 47808 389234
rect 48976 387025 49004 491914
rect 50356 430953 50384 532714
rect 54484 518968 54536 518974
rect 54484 518910 54536 518916
rect 51724 480276 51776 480282
rect 51724 480218 51776 480224
rect 50528 440292 50580 440298
rect 50528 440234 50580 440240
rect 50342 430944 50398 430953
rect 50342 430879 50398 430888
rect 48962 387016 49018 387025
rect 48962 386951 49018 386960
rect 50540 351257 50568 440234
rect 51736 386753 51764 480218
rect 51908 466472 51960 466478
rect 51908 466414 51960 466420
rect 51722 386744 51778 386753
rect 51722 386679 51778 386688
rect 51920 386481 51948 466414
rect 53104 454096 53156 454102
rect 53104 454038 53156 454044
rect 51906 386472 51962 386481
rect 51906 386407 51962 386416
rect 51724 375420 51776 375426
rect 51724 375362 51776 375368
rect 50526 351248 50582 351257
rect 50526 351183 50582 351192
rect 48962 334112 49018 334121
rect 48962 334047 49018 334056
rect 47766 300520 47822 300529
rect 47766 300455 47822 300464
rect 47766 247480 47822 247489
rect 47766 247415 47822 247424
rect 47780 53242 47808 247415
rect 47950 213344 48006 213353
rect 47950 213279 48006 213288
rect 47964 190505 47992 213279
rect 48134 210896 48190 210905
rect 48134 210831 48190 210840
rect 48148 194449 48176 210831
rect 48778 206272 48834 206281
rect 48778 206207 48834 206216
rect 48134 194440 48190 194449
rect 48134 194375 48190 194384
rect 48792 192409 48820 206207
rect 48778 192400 48834 192409
rect 48778 192335 48834 192344
rect 47950 190496 48006 190505
rect 47950 190431 48006 190440
rect 47768 53236 47820 53242
rect 47768 53178 47820 53184
rect 48976 51882 49004 334047
rect 51736 301345 51764 375362
rect 53116 321473 53144 454038
rect 54496 430545 54524 518910
rect 54482 430536 54538 430545
rect 54482 430471 54538 430480
rect 54484 427848 54536 427854
rect 54484 427790 54536 427796
rect 54496 344321 54524 427790
rect 55876 408513 55904 558078
rect 56060 540297 56088 608602
rect 651470 603936 651526 603945
rect 651470 603871 651526 603880
rect 651484 603158 651512 603871
rect 651472 603152 651524 603158
rect 651472 603094 651524 603100
rect 62118 597952 62174 597961
rect 62118 597887 62174 597896
rect 62132 597582 62160 597887
rect 62120 597576 62172 597582
rect 62120 597518 62172 597524
rect 651470 590744 651526 590753
rect 651470 590679 651472 590688
rect 651524 590679 651526 590688
rect 651472 590650 651524 590656
rect 62118 584896 62174 584905
rect 62118 584831 62174 584840
rect 62132 583778 62160 584831
rect 62120 583772 62172 583778
rect 62120 583714 62172 583720
rect 652036 583001 652064 683567
rect 660316 625297 660344 763166
rect 661696 760481 661724 921810
rect 663064 909492 663116 909498
rect 663064 909434 663116 909440
rect 663076 760889 663104 909434
rect 671344 895688 671396 895694
rect 671344 895630 671396 895636
rect 664444 881884 664496 881890
rect 664444 881826 664496 881832
rect 664456 868737 664484 881826
rect 669226 879200 669282 879209
rect 669226 879135 669282 879144
rect 664442 868728 664498 868737
rect 664442 868663 664498 868672
rect 668214 868184 668270 868193
rect 668214 868119 668270 868128
rect 664444 855636 664496 855642
rect 664444 855578 664496 855584
rect 663062 760880 663118 760889
rect 663062 760815 663118 760824
rect 661682 760472 661738 760481
rect 661682 760407 661738 760416
rect 663064 723172 663116 723178
rect 663064 723114 663116 723120
rect 661684 696992 661736 696998
rect 661684 696934 661736 696940
rect 660302 625288 660358 625297
rect 660302 625223 660358 625232
rect 660304 616888 660356 616894
rect 660304 616830 660356 616836
rect 660316 599593 660344 616830
rect 660302 599584 660358 599593
rect 660302 599519 660358 599528
rect 652022 582992 652078 583001
rect 652022 582927 652078 582936
rect 661696 581097 661724 696934
rect 663076 689353 663104 723114
rect 664456 716553 664484 855578
rect 667204 803208 667256 803214
rect 667204 803150 667256 803156
rect 666282 777064 666338 777073
rect 666282 776999 666338 777008
rect 665824 749420 665876 749426
rect 665824 749362 665876 749368
rect 664442 716544 664498 716553
rect 664442 716479 664498 716488
rect 664444 709368 664496 709374
rect 664444 709310 664496 709316
rect 663062 689344 663118 689353
rect 663062 689279 663118 689288
rect 661868 669384 661920 669390
rect 661868 669326 661920 669332
rect 661880 643793 661908 669326
rect 661866 643784 661922 643793
rect 661866 643719 661922 643728
rect 662052 590708 662104 590714
rect 662052 590650 662104 590656
rect 661682 581088 661738 581097
rect 661682 581023 661738 581032
rect 651470 577416 651526 577425
rect 651470 577351 651526 577360
rect 651484 576910 651512 577351
rect 651472 576904 651524 576910
rect 651472 576846 651524 576852
rect 62118 571840 62174 571849
rect 62118 571775 62174 571784
rect 62132 569265 62160 571775
rect 62118 569256 62174 569265
rect 62118 569191 62174 569200
rect 651654 564088 651710 564097
rect 651654 564023 651710 564032
rect 651668 563106 651696 564023
rect 651656 563100 651708 563106
rect 651656 563042 651708 563048
rect 658924 563100 658976 563106
rect 658924 563042 658976 563048
rect 62118 558784 62174 558793
rect 62118 558719 62174 558728
rect 62132 558142 62160 558719
rect 62120 558136 62172 558142
rect 62120 558078 62172 558084
rect 658936 554033 658964 563042
rect 658922 554024 658978 554033
rect 658922 553959 658978 553968
rect 651470 550896 651526 550905
rect 651470 550831 651526 550840
rect 651484 550662 651512 550831
rect 651472 550656 651524 550662
rect 651472 550598 651524 550604
rect 660304 550656 660356 550662
rect 660304 550598 660356 550604
rect 62118 545864 62174 545873
rect 62118 545799 62174 545808
rect 62132 545154 62160 545799
rect 62120 545148 62172 545154
rect 62120 545090 62172 545096
rect 56046 540288 56102 540297
rect 56046 540223 56102 540232
rect 651470 537568 651526 537577
rect 651470 537503 651526 537512
rect 651484 536858 651512 537503
rect 651472 536852 651524 536858
rect 651472 536794 651524 536800
rect 62118 532808 62174 532817
rect 62118 532743 62120 532752
rect 62172 532743 62174 532752
rect 62120 532714 62172 532720
rect 651838 524240 651894 524249
rect 651838 524175 651894 524184
rect 651852 523054 651880 524175
rect 651840 523048 651892 523054
rect 651840 522990 651892 522996
rect 62118 519752 62174 519761
rect 62118 519687 62174 519696
rect 62132 518974 62160 519687
rect 62120 518968 62172 518974
rect 62120 518910 62172 518916
rect 651470 511048 651526 511057
rect 651470 510983 651526 510992
rect 651484 510678 651512 510983
rect 651472 510672 651524 510678
rect 651472 510614 651524 510620
rect 659108 510672 659160 510678
rect 659108 510614 659160 510620
rect 62118 506696 62174 506705
rect 62118 506631 62174 506640
rect 62132 506530 62160 506631
rect 62120 506524 62172 506530
rect 62120 506466 62172 506472
rect 651470 497720 651526 497729
rect 651470 497655 651526 497664
rect 651484 496874 651512 497655
rect 651472 496868 651524 496874
rect 651472 496810 651524 496816
rect 62118 493640 62174 493649
rect 62118 493575 62174 493584
rect 62132 491978 62160 493575
rect 62120 491972 62172 491978
rect 62120 491914 62172 491920
rect 651470 484528 651526 484537
rect 651470 484463 651472 484472
rect 651524 484463 651526 484472
rect 651472 484434 651524 484440
rect 62118 480584 62174 480593
rect 62118 480519 62174 480528
rect 62132 480282 62160 480519
rect 62120 480276 62172 480282
rect 62120 480218 62172 480224
rect 651470 471200 651526 471209
rect 651470 471135 651526 471144
rect 651484 470626 651512 471135
rect 651472 470620 651524 470626
rect 651472 470562 651524 470568
rect 62118 467528 62174 467537
rect 62118 467463 62174 467472
rect 62132 466478 62160 467463
rect 62120 466472 62172 466478
rect 62120 466414 62172 466420
rect 652390 457872 652446 457881
rect 652390 457807 652446 457816
rect 652404 456822 652432 457807
rect 652392 456816 652444 456822
rect 652392 456758 652444 456764
rect 62118 454608 62174 454617
rect 62118 454543 62174 454552
rect 62132 454102 62160 454543
rect 62120 454096 62172 454102
rect 62120 454038 62172 454044
rect 651470 444544 651526 444553
rect 651470 444479 651472 444488
rect 651524 444479 651526 444488
rect 651472 444450 651524 444456
rect 62118 441552 62174 441561
rect 62118 441487 62174 441496
rect 62132 440298 62160 441487
rect 62120 440292 62172 440298
rect 62120 440234 62172 440240
rect 651470 431352 651526 431361
rect 651470 431287 651526 431296
rect 651484 430642 651512 431287
rect 651472 430636 651524 430642
rect 651472 430578 651524 430584
rect 62118 428496 62174 428505
rect 62118 428431 62174 428440
rect 62132 427854 62160 428431
rect 62120 427848 62172 427854
rect 62120 427790 62172 427796
rect 651838 418024 651894 418033
rect 651838 417959 651894 417968
rect 651852 416838 651880 417959
rect 651840 416832 651892 416838
rect 651840 416774 651892 416780
rect 62120 415472 62172 415478
rect 62118 415440 62120 415449
rect 62172 415440 62174 415449
rect 62118 415375 62174 415384
rect 55862 408504 55918 408513
rect 55862 408439 55918 408448
rect 651470 404696 651526 404705
rect 651470 404631 651526 404640
rect 651484 404394 651512 404631
rect 651472 404388 651524 404394
rect 651472 404330 651524 404336
rect 62118 402384 62174 402393
rect 62118 402319 62174 402328
rect 62132 401674 62160 402319
rect 55864 401668 55916 401674
rect 55864 401610 55916 401616
rect 62120 401668 62172 401674
rect 62120 401610 62172 401616
rect 54482 344312 54538 344321
rect 54482 344247 54538 344256
rect 53288 322992 53340 322998
rect 53288 322934 53340 322940
rect 53102 321464 53158 321473
rect 53102 321399 53158 321408
rect 51722 301336 51778 301345
rect 51722 301271 51778 301280
rect 49146 290456 49202 290465
rect 49146 290391 49202 290400
rect 49160 52018 49188 290391
rect 50342 290184 50398 290193
rect 50342 290119 50398 290128
rect 49514 208992 49570 209001
rect 49514 208927 49570 208936
rect 49528 196489 49556 208927
rect 49514 196480 49570 196489
rect 49514 196415 49570 196424
rect 50356 53378 50384 290119
rect 51722 289912 51778 289921
rect 51722 289847 51778 289856
rect 50526 246528 50582 246537
rect 50526 246463 50582 246472
rect 50344 53372 50396 53378
rect 50344 53314 50396 53320
rect 49148 52012 49200 52018
rect 49148 51954 49200 51960
rect 48964 51876 49016 51882
rect 48964 51818 49016 51824
rect 50540 50522 50568 246463
rect 50528 50516 50580 50522
rect 50528 50458 50580 50464
rect 51736 49162 51764 289847
rect 53300 257553 53328 322934
rect 54484 310548 54536 310554
rect 54484 310490 54536 310496
rect 53286 257544 53342 257553
rect 53286 257479 53342 257488
rect 54496 217977 54524 310490
rect 55876 278769 55904 401610
rect 652574 391504 652630 391513
rect 652574 391439 652630 391448
rect 652588 390590 652616 391439
rect 652576 390584 652628 390590
rect 652576 390526 652628 390532
rect 658924 390584 658976 390590
rect 658924 390526 658976 390532
rect 62118 389328 62174 389337
rect 62118 389263 62120 389272
rect 62172 389263 62174 389272
rect 62120 389234 62172 389240
rect 652022 378176 652078 378185
rect 652022 378111 652078 378120
rect 62118 376272 62174 376281
rect 62118 376207 62174 376216
rect 62132 375426 62160 376207
rect 62120 375420 62172 375426
rect 62120 375362 62172 375368
rect 651654 364848 651710 364857
rect 651654 364783 651710 364792
rect 651668 364410 651696 364783
rect 651656 364404 651708 364410
rect 651656 364346 651708 364352
rect 62118 363352 62174 363361
rect 62118 363287 62174 363296
rect 62132 362982 62160 363287
rect 62120 362976 62172 362982
rect 62120 362918 62172 362924
rect 651470 351656 651526 351665
rect 651470 351591 651526 351600
rect 651484 350606 651512 351591
rect 651472 350600 651524 350606
rect 651472 350542 651524 350548
rect 62762 350296 62818 350305
rect 62762 350231 62818 350240
rect 62118 337240 62174 337249
rect 62118 337175 62174 337184
rect 62132 336802 62160 337175
rect 62120 336796 62172 336802
rect 62120 336738 62172 336744
rect 62118 324184 62174 324193
rect 62118 324119 62174 324128
rect 62132 322998 62160 324119
rect 62120 322992 62172 322998
rect 62120 322934 62172 322940
rect 62118 311128 62174 311137
rect 62118 311063 62174 311072
rect 62132 310554 62160 311063
rect 62120 310548 62172 310554
rect 62120 310490 62172 310496
rect 62118 298208 62174 298217
rect 62118 298143 62120 298152
rect 62172 298143 62174 298152
rect 62120 298114 62172 298120
rect 55862 278760 55918 278769
rect 55862 278695 55918 278704
rect 62776 267073 62804 350231
rect 651470 338328 651526 338337
rect 651470 338263 651526 338272
rect 651484 338162 651512 338263
rect 651472 338156 651524 338162
rect 651472 338098 651524 338104
rect 651470 325000 651526 325009
rect 651470 324935 651526 324944
rect 651484 324358 651512 324935
rect 651472 324352 651524 324358
rect 651472 324294 651524 324300
rect 651470 311808 651526 311817
rect 651470 311743 651526 311752
rect 651484 310554 651512 311743
rect 651472 310548 651524 310554
rect 651472 310490 651524 310496
rect 651470 285288 651526 285297
rect 651470 285223 651526 285232
rect 62946 285152 63002 285161
rect 62946 285087 63002 285096
rect 62762 267064 62818 267073
rect 62762 266999 62818 267008
rect 62764 228540 62816 228546
rect 62764 228482 62816 228488
rect 57888 227044 57940 227050
rect 57888 226986 57940 226992
rect 56508 222488 56560 222494
rect 56508 222430 56560 222436
rect 56324 218204 56376 218210
rect 56324 218146 56376 218152
rect 55680 218068 55732 218074
rect 55680 218010 55732 218016
rect 54482 217968 54538 217977
rect 54482 217903 54538 217912
rect 55692 217138 55720 218010
rect 56336 217274 56364 218146
rect 56520 218074 56548 222430
rect 57900 218074 57928 226986
rect 61292 225616 61344 225622
rect 61292 225558 61344 225564
rect 60648 224528 60700 224534
rect 60648 224470 60700 224476
rect 58992 224256 59044 224262
rect 58992 224198 59044 224204
rect 56508 218068 56560 218074
rect 56508 218010 56560 218016
rect 57336 218068 57388 218074
rect 57336 218010 57388 218016
rect 57888 218068 57940 218074
rect 57888 218010 57940 218016
rect 58164 218068 58216 218074
rect 58164 218010 58216 218016
rect 56336 217246 56502 217274
rect 55646 217110 55720 217138
rect 55646 216988 55674 217110
rect 56474 216988 56502 217246
rect 57348 217138 57376 218010
rect 58176 217138 58204 218010
rect 59004 217274 59032 224198
rect 59820 218612 59872 218618
rect 59820 218554 59872 218560
rect 57302 217110 57376 217138
rect 58130 217110 58204 217138
rect 58958 217246 59032 217274
rect 57302 216988 57330 217110
rect 58130 216988 58158 217110
rect 58958 216988 58986 217246
rect 59832 217138 59860 218554
rect 60660 217274 60688 224470
rect 61304 218074 61332 225558
rect 61476 221604 61528 221610
rect 61476 221546 61528 221552
rect 61292 218068 61344 218074
rect 61292 218010 61344 218016
rect 61488 217274 61516 221546
rect 62304 218884 62356 218890
rect 62304 218826 62356 218832
rect 59786 217110 59860 217138
rect 60614 217246 60688 217274
rect 61442 217246 61516 217274
rect 59786 216988 59814 217110
rect 60614 216988 60642 217246
rect 61442 216988 61470 217246
rect 62316 217138 62344 218826
rect 62776 218210 62804 228482
rect 62960 222873 62988 285087
rect 651484 284374 651512 285223
rect 651472 284368 651524 284374
rect 651472 284310 651524 284316
rect 65904 274666 65932 277780
rect 67008 274718 67036 277780
rect 66996 274712 67048 274718
rect 65904 274638 66300 274666
rect 66996 274654 67048 274660
rect 66272 268394 66300 274638
rect 68204 271318 68232 277780
rect 68192 271312 68244 271318
rect 68192 271254 68244 271260
rect 69400 269822 69428 277780
rect 70596 275330 70624 277780
rect 70584 275324 70636 275330
rect 70584 275266 70636 275272
rect 71792 274990 71820 277780
rect 71780 274984 71832 274990
rect 71780 274926 71832 274932
rect 71044 274712 71096 274718
rect 71044 274654 71096 274660
rect 69388 269816 69440 269822
rect 69388 269758 69440 269764
rect 66260 268388 66312 268394
rect 66260 268330 66312 268336
rect 71056 267034 71084 274654
rect 72988 271182 73016 277780
rect 74092 275194 74120 277780
rect 75302 277766 75868 277794
rect 74080 275188 74132 275194
rect 74080 275130 74132 275136
rect 73804 274984 73856 274990
rect 73804 274926 73856 274932
rect 72976 271176 73028 271182
rect 72976 271118 73028 271124
rect 73816 267170 73844 274926
rect 75840 269958 75868 277766
rect 76484 275602 76512 277780
rect 76472 275596 76524 275602
rect 76472 275538 76524 275544
rect 77208 275188 77260 275194
rect 77208 275130 77260 275136
rect 77220 273970 77248 275130
rect 77208 273964 77260 273970
rect 77208 273906 77260 273912
rect 77680 272542 77708 277780
rect 78876 272950 78904 277780
rect 78864 272944 78916 272950
rect 78864 272886 78916 272892
rect 77668 272536 77720 272542
rect 77668 272478 77720 272484
rect 80072 270094 80100 277780
rect 81268 275738 81296 277780
rect 81256 275732 81308 275738
rect 81256 275674 81308 275680
rect 82372 274242 82400 277780
rect 83582 277766 84148 277794
rect 82360 274236 82412 274242
rect 82360 274178 82412 274184
rect 80060 270088 80112 270094
rect 80060 270030 80112 270036
rect 75828 269952 75880 269958
rect 75828 269894 75880 269900
rect 84120 269686 84148 277766
rect 84764 274106 84792 277780
rect 85960 275466 85988 277780
rect 86868 275596 86920 275602
rect 86868 275538 86920 275544
rect 85948 275460 86000 275466
rect 85948 275402 86000 275408
rect 84752 274100 84804 274106
rect 84752 274042 84804 274048
rect 84108 269680 84160 269686
rect 84108 269622 84160 269628
rect 86880 268938 86908 275538
rect 87156 272678 87184 277780
rect 88352 276010 88380 277780
rect 89548 277394 89576 277780
rect 89548 277366 89668 277394
rect 88340 276004 88392 276010
rect 88340 275946 88392 275952
rect 89640 275890 89668 277366
rect 89640 275862 89760 275890
rect 88984 275732 89036 275738
rect 88984 275674 89036 275680
rect 87144 272672 87196 272678
rect 87144 272614 87196 272620
rect 86868 268932 86920 268938
rect 86868 268874 86920 268880
rect 88996 267714 89024 275674
rect 89732 271454 89760 275862
rect 90652 274718 90680 277780
rect 91862 277766 92428 277794
rect 90640 274712 90692 274718
rect 90640 274654 90692 274660
rect 89720 271448 89772 271454
rect 89720 271390 89772 271396
rect 92400 268530 92428 277766
rect 93044 271726 93072 277780
rect 94240 272814 94268 277780
rect 95436 275874 95464 277780
rect 95424 275868 95476 275874
rect 95424 275810 95476 275816
rect 96632 275602 96660 277780
rect 97750 277766 97948 277794
rect 98946 277766 99328 277794
rect 100142 277766 100708 277794
rect 96620 275596 96672 275602
rect 96620 275538 96672 275544
rect 95884 274712 95936 274718
rect 95884 274654 95936 274660
rect 94228 272808 94280 272814
rect 94228 272750 94280 272756
rect 93032 271720 93084 271726
rect 93032 271662 93084 271668
rect 92388 268524 92440 268530
rect 92388 268466 92440 268472
rect 88984 267708 89036 267714
rect 88984 267650 89036 267656
rect 95896 267578 95924 274654
rect 97920 270230 97948 277766
rect 97908 270224 97960 270230
rect 97908 270166 97960 270172
rect 99300 268666 99328 277766
rect 99288 268660 99340 268666
rect 99288 268602 99340 268608
rect 95884 267572 95936 267578
rect 95884 267514 95936 267520
rect 100680 267306 100708 277766
rect 101324 274378 101352 277780
rect 101312 274372 101364 274378
rect 101312 274314 101364 274320
rect 102520 268802 102548 277780
rect 103716 275738 103744 277780
rect 104912 277394 104940 277780
rect 104912 277366 105032 277394
rect 104808 275868 104860 275874
rect 104808 275810 104860 275816
rect 103704 275732 103756 275738
rect 103704 275674 103756 275680
rect 104820 274650 104848 275810
rect 104808 274644 104860 274650
rect 104808 274586 104860 274592
rect 105004 273086 105032 277366
rect 106016 274786 106044 277780
rect 107226 277766 107608 277794
rect 108422 277766 108988 277794
rect 109618 277766 110276 277794
rect 106004 274780 106056 274786
rect 106004 274722 106056 274728
rect 104992 273080 105044 273086
rect 104992 273022 105044 273028
rect 102508 268796 102560 268802
rect 102508 268738 102560 268744
rect 107580 267442 107608 277766
rect 108960 269074 108988 277766
rect 110248 270366 110276 277766
rect 110800 275194 110828 277780
rect 110788 275188 110840 275194
rect 110788 275130 110840 275136
rect 110420 274780 110472 274786
rect 110420 274722 110472 274728
rect 110432 271862 110460 274722
rect 110420 271856 110472 271862
rect 110420 271798 110472 271804
rect 111996 271590 112024 277780
rect 113192 275874 113220 277780
rect 113180 275868 113232 275874
rect 113180 275810 113232 275816
rect 114296 273222 114324 277780
rect 115506 277766 115888 277794
rect 114284 273216 114336 273222
rect 114284 273158 114336 273164
rect 111984 271584 112036 271590
rect 111984 271526 112036 271532
rect 115860 270502 115888 277766
rect 116688 270638 116716 277780
rect 117898 277766 118648 277794
rect 116676 270632 116728 270638
rect 116676 270574 116728 270580
rect 115848 270496 115900 270502
rect 115848 270438 115900 270444
rect 110236 270360 110288 270366
rect 110236 270302 110288 270308
rect 118620 269414 118648 277766
rect 119080 269550 119108 277780
rect 120290 277766 120948 277794
rect 120920 271726 120948 277766
rect 121380 274514 121408 277780
rect 122590 277766 122788 277794
rect 121368 274508 121420 274514
rect 121368 274450 121420 274456
rect 120724 271720 120776 271726
rect 120724 271662 120776 271668
rect 120908 271720 120960 271726
rect 120908 271662 120960 271668
rect 119804 269680 119856 269686
rect 119804 269622 119856 269628
rect 119068 269544 119120 269550
rect 119068 269486 119120 269492
rect 118608 269408 118660 269414
rect 118608 269350 118660 269356
rect 108948 269068 109000 269074
rect 108948 269010 109000 269016
rect 107568 267436 107620 267442
rect 107568 267378 107620 267384
rect 100668 267300 100720 267306
rect 100668 267242 100720 267248
rect 73804 267164 73856 267170
rect 73804 267106 73856 267112
rect 71044 267028 71096 267034
rect 71044 266970 71096 266976
rect 119816 266490 119844 269622
rect 120736 266762 120764 271662
rect 122760 268258 122788 277766
rect 123772 273834 123800 277780
rect 124982 277766 125548 277794
rect 126178 277766 126928 277794
rect 123760 273828 123812 273834
rect 123760 273770 123812 273776
rect 122748 268252 122800 268258
rect 122748 268194 122800 268200
rect 125520 267986 125548 277766
rect 126900 269550 126928 277766
rect 127360 272406 127388 277780
rect 127348 272400 127400 272406
rect 127348 272342 127400 272348
rect 128556 271046 128584 277780
rect 129660 274922 129688 277780
rect 129648 274916 129700 274922
rect 129648 274858 129700 274864
rect 128544 271040 128596 271046
rect 128544 270982 128596 270988
rect 130856 270910 130884 277780
rect 132066 277766 132448 277794
rect 133262 277766 133828 277794
rect 130844 270904 130896 270910
rect 130844 270846 130896 270852
rect 126888 269544 126940 269550
rect 126888 269486 126940 269492
rect 125508 267980 125560 267986
rect 125508 267922 125560 267928
rect 132420 266898 132448 277766
rect 133800 268122 133828 277766
rect 134444 273698 134472 277780
rect 135640 275058 135668 277780
rect 135628 275052 135680 275058
rect 135628 274994 135680 275000
rect 136548 274916 136600 274922
rect 136548 274858 136600 274864
rect 134432 273692 134484 273698
rect 134432 273634 134484 273640
rect 136560 269793 136588 274858
rect 136546 269784 136602 269793
rect 136546 269719 136602 269728
rect 136836 269278 136864 277780
rect 137940 270774 137968 277780
rect 138664 272944 138716 272950
rect 138664 272886 138716 272892
rect 138480 271312 138532 271318
rect 138480 271254 138532 271260
rect 137928 270768 137980 270774
rect 137928 270710 137980 270716
rect 136824 269272 136876 269278
rect 136824 269214 136876 269220
rect 137284 268388 137336 268394
rect 137284 268330 137336 268336
rect 133788 268116 133840 268122
rect 133788 268058 133840 268064
rect 132408 266892 132460 266898
rect 132408 266834 132460 266840
rect 120724 266756 120776 266762
rect 120724 266698 120776 266704
rect 119804 266484 119856 266490
rect 119804 266426 119856 266432
rect 137296 264316 137324 268330
rect 138112 267028 138164 267034
rect 138112 266970 138164 266976
rect 138124 264316 138152 266970
rect 138492 264330 138520 271254
rect 138676 266626 138704 272886
rect 139136 272270 139164 277780
rect 140136 275324 140188 275330
rect 140136 275266 140188 275272
rect 139124 272264 139176 272270
rect 139124 272206 139176 272212
rect 139768 269816 139820 269822
rect 139952 269816 140004 269822
rect 139768 269758 139820 269764
rect 139950 269784 139952 269793
rect 140004 269784 140006 269793
rect 138664 266620 138716 266626
rect 138664 266562 138716 266568
rect 138492 264302 138966 264330
rect 139780 264316 139808 269758
rect 139950 269719 140006 269728
rect 140148 264330 140176 275266
rect 140332 274786 140360 277780
rect 141542 277766 141832 277794
rect 140320 274780 140372 274786
rect 140320 274722 140372 274728
rect 141804 272950 141832 277766
rect 142724 275330 142752 277780
rect 143356 276004 143408 276010
rect 143356 275946 143408 275952
rect 142712 275324 142764 275330
rect 142712 275266 142764 275272
rect 141792 272944 141844 272950
rect 141792 272886 141844 272892
rect 141608 272264 141660 272270
rect 141608 272206 141660 272212
rect 141424 267164 141476 267170
rect 141424 267106 141476 267112
rect 140148 264302 140622 264330
rect 141436 264316 141464 267106
rect 141620 267034 141648 272206
rect 142160 271176 142212 271182
rect 142160 271118 142212 271124
rect 141608 267028 141660 267034
rect 141608 266970 141660 266976
rect 142172 264330 142200 271118
rect 143368 269958 143396 275946
rect 143540 273964 143592 273970
rect 143540 273906 143592 273912
rect 142620 269952 142672 269958
rect 142620 269894 142672 269900
rect 143356 269952 143408 269958
rect 143356 269894 143408 269900
rect 142632 267734 142660 269894
rect 142632 267706 142752 267734
rect 142724 264330 142752 267706
rect 143552 264330 143580 273906
rect 143920 272270 143948 277780
rect 144644 274780 144696 274786
rect 144644 274722 144696 274728
rect 144656 273562 144684 274722
rect 145024 273970 145052 277780
rect 146220 274786 146248 277780
rect 147430 277766 147628 277794
rect 146760 275460 146812 275466
rect 146760 275402 146812 275408
rect 146208 274780 146260 274786
rect 146208 274722 146260 274728
rect 145564 274236 145616 274242
rect 145564 274178 145616 274184
rect 145012 273964 145064 273970
rect 145012 273906 145064 273912
rect 144644 273556 144696 273562
rect 144644 273498 144696 273504
rect 145104 272536 145156 272542
rect 145104 272478 145156 272484
rect 143908 272264 143960 272270
rect 143908 272206 143960 272212
rect 144736 268932 144788 268938
rect 144736 268874 144788 268880
rect 144552 267708 144604 267714
rect 144552 267650 144604 267656
rect 144564 267170 144592 267650
rect 144552 267164 144604 267170
rect 144552 267106 144604 267112
rect 142172 264302 142278 264330
rect 142724 264302 143106 264330
rect 143552 264302 143934 264330
rect 144748 264316 144776 268874
rect 144920 267708 144972 267714
rect 144920 267650 144972 267656
rect 144932 266490 144960 267650
rect 144920 266484 144972 266490
rect 144920 266426 144972 266432
rect 145116 264330 145144 272478
rect 145576 266558 145604 274178
rect 146772 270094 146800 275402
rect 146392 270088 146444 270094
rect 146392 270030 146444 270036
rect 146760 270088 146812 270094
rect 146760 270030 146812 270036
rect 145564 266552 145616 266558
rect 145564 266494 145616 266500
rect 145116 264302 145590 264330
rect 146404 264316 146432 270030
rect 147600 268394 147628 277766
rect 148324 274100 148376 274106
rect 148324 274042 148376 274048
rect 147588 268388 147640 268394
rect 147588 268330 147640 268336
rect 147588 267980 147640 267986
rect 147588 267922 147640 267928
rect 147600 267170 147628 267922
rect 147404 267164 147456 267170
rect 147404 267106 147456 267112
rect 147588 267164 147640 267170
rect 147588 267106 147640 267112
rect 147416 267050 147444 267106
rect 147416 267022 147720 267050
rect 147220 266416 147272 266422
rect 147220 266358 147272 266364
rect 147232 264316 147260 266358
rect 147692 264330 147720 267022
rect 148336 266422 148364 274042
rect 148612 271182 148640 277780
rect 149808 274922 149836 277780
rect 149796 274916 149848 274922
rect 149796 274858 149848 274864
rect 149888 274780 149940 274786
rect 149888 274722 149940 274728
rect 148600 271176 148652 271182
rect 148600 271118 148652 271124
rect 149900 267170 149928 274722
rect 151004 271318 151032 277780
rect 152004 272672 152056 272678
rect 152004 272614 152056 272620
rect 150992 271312 151044 271318
rect 150992 271254 151044 271260
rect 151084 270632 151136 270638
rect 151084 270574 151136 270580
rect 150532 267708 150584 267714
rect 150532 267650 150584 267656
rect 149060 267164 149112 267170
rect 149060 267106 149112 267112
rect 149888 267164 149940 267170
rect 149888 267106 149940 267112
rect 149072 266626 149100 267106
rect 149060 266620 149112 266626
rect 149060 266562 149112 266568
rect 148876 266552 148928 266558
rect 148876 266494 148928 266500
rect 148324 266416 148376 266422
rect 148324 266358 148376 266364
rect 147692 264302 148074 264330
rect 148888 264316 148916 266494
rect 149704 266416 149756 266422
rect 149704 266358 149756 266364
rect 149716 264316 149744 266358
rect 150544 264316 150572 267650
rect 151096 266490 151124 270574
rect 151360 270088 151412 270094
rect 151360 270030 151412 270036
rect 151084 266484 151136 266490
rect 151084 266426 151136 266432
rect 151372 264316 151400 270030
rect 152016 264330 152044 272614
rect 152200 272542 152228 277780
rect 152188 272536 152240 272542
rect 152188 272478 152240 272484
rect 153304 272134 153332 277780
rect 153292 272128 153344 272134
rect 153292 272070 153344 272076
rect 152648 271448 152700 271454
rect 152648 271390 152700 271396
rect 152660 264330 152688 271390
rect 153844 270088 153896 270094
rect 153844 270030 153896 270036
rect 152016 264302 152214 264330
rect 152660 264302 153042 264330
rect 153856 264316 153884 270030
rect 154500 269958 154528 277780
rect 155710 277766 155908 277794
rect 154488 269952 154540 269958
rect 154488 269894 154540 269900
rect 155880 268530 155908 277766
rect 156892 276010 156920 277780
rect 156880 276004 156932 276010
rect 156880 275946 156932 275952
rect 156604 275596 156656 275602
rect 156604 275538 156656 275544
rect 156052 272808 156104 272814
rect 156052 272750 156104 272756
rect 155500 268524 155552 268530
rect 155500 268466 155552 268472
rect 155868 268524 155920 268530
rect 155868 268466 155920 268472
rect 154672 267572 154724 267578
rect 154672 267514 154724 267520
rect 154684 264316 154712 267514
rect 155512 264316 155540 268466
rect 156064 264330 156092 272750
rect 156616 266762 156644 275538
rect 157616 274644 157668 274650
rect 157616 274586 157668 274592
rect 156420 266756 156472 266762
rect 156420 266698 156472 266704
rect 156604 266756 156656 266762
rect 156604 266698 156656 266704
rect 156432 264602 156460 266698
rect 156432 264574 156736 264602
rect 156708 264330 156736 264574
rect 157628 264330 157656 274586
rect 158088 274106 158116 277780
rect 159298 277766 159956 277794
rect 158076 274100 158128 274106
rect 158076 274042 158128 274048
rect 158812 270224 158864 270230
rect 158812 270166 158864 270172
rect 156064 264302 156354 264330
rect 156708 264302 157182 264330
rect 157628 264302 158010 264330
rect 158824 264316 158852 270166
rect 159928 270094 159956 277766
rect 160100 275732 160152 275738
rect 160100 275674 160152 275680
rect 160112 274242 160140 275674
rect 160480 275466 160508 277780
rect 160468 275460 160520 275466
rect 160468 275402 160520 275408
rect 161584 274718 161612 277780
rect 162124 275188 162176 275194
rect 162124 275130 162176 275136
rect 161572 274712 161624 274718
rect 161572 274654 161624 274660
rect 160928 274372 160980 274378
rect 160928 274314 160980 274320
rect 160100 274236 160152 274242
rect 160100 274178 160152 274184
rect 159916 270088 159968 270094
rect 159916 270030 159968 270036
rect 160468 268660 160520 268666
rect 160468 268602 160520 268608
rect 159640 266756 159692 266762
rect 159640 266698 159692 266704
rect 159652 264316 159680 266698
rect 160480 264316 160508 268602
rect 160940 264330 160968 274314
rect 162136 267578 162164 275130
rect 162780 268666 162808 277780
rect 163976 275602 164004 277780
rect 163964 275596 164016 275602
rect 163964 275538 164016 275544
rect 163136 274712 163188 274718
rect 163136 274654 163188 274660
rect 163148 268802 163176 274654
rect 164240 274236 164292 274242
rect 164240 274178 164292 274184
rect 163320 273080 163372 273086
rect 163320 273022 163372 273028
rect 162952 268796 163004 268802
rect 162952 268738 163004 268744
rect 163136 268796 163188 268802
rect 163136 268738 163188 268744
rect 162768 268660 162820 268666
rect 162768 268602 162820 268608
rect 162124 267572 162176 267578
rect 162124 267514 162176 267520
rect 162124 267300 162176 267306
rect 162124 267242 162176 267248
rect 160940 264302 161322 264330
rect 162136 264316 162164 267242
rect 162964 264316 162992 268738
rect 163332 264330 163360 273022
rect 164252 264330 164280 274178
rect 164976 271856 165028 271862
rect 164976 271798 165028 271804
rect 164988 264330 165016 271798
rect 165172 271454 165200 277780
rect 166382 277766 166948 277794
rect 165160 271448 165212 271454
rect 165160 271390 165212 271396
rect 166920 270230 166948 277766
rect 167564 273086 167592 277780
rect 167736 275460 167788 275466
rect 167736 275402 167788 275408
rect 167552 273080 167604 273086
rect 167552 273022 167604 273028
rect 166908 270224 166960 270230
rect 166908 270166 166960 270172
rect 166908 269408 166960 269414
rect 166908 269350 166960 269356
rect 166264 269068 166316 269074
rect 166264 269010 166316 269016
rect 163332 264302 163806 264330
rect 164252 264302 164634 264330
rect 164988 264302 165462 264330
rect 166276 264316 166304 269010
rect 166920 267306 166948 269350
rect 167748 267442 167776 275402
rect 168668 272678 168696 277780
rect 169878 277766 170168 277794
rect 169944 275868 169996 275874
rect 169944 275810 169996 275816
rect 169024 273216 169076 273222
rect 169024 273158 169076 273164
rect 168656 272672 168708 272678
rect 168656 272614 168708 272620
rect 168380 271584 168432 271590
rect 168380 271526 168432 271532
rect 167920 270360 167972 270366
rect 167920 270302 167972 270308
rect 167092 267436 167144 267442
rect 167092 267378 167144 267384
rect 167736 267436 167788 267442
rect 167736 267378 167788 267384
rect 166908 267300 166960 267306
rect 166908 267242 166960 267248
rect 167104 264316 167132 267378
rect 167932 264316 167960 270302
rect 168392 264330 168420 271526
rect 169036 266762 169064 273158
rect 169576 267572 169628 267578
rect 169576 267514 169628 267520
rect 169024 266756 169076 266762
rect 169024 266698 169076 266704
rect 168392 264302 168774 264330
rect 169588 264316 169616 267514
rect 169956 264330 169984 275810
rect 170140 274718 170168 277766
rect 171060 275466 171088 277780
rect 172270 277766 172468 277794
rect 171048 275460 171100 275466
rect 171048 275402 171100 275408
rect 170128 274712 170180 274718
rect 170128 274654 170180 274660
rect 171784 272128 171836 272134
rect 171784 272070 171836 272076
rect 171232 270496 171284 270502
rect 171232 270438 171284 270444
rect 169956 264302 170430 264330
rect 171244 264316 171272 270438
rect 171796 267714 171824 272070
rect 172440 270502 172468 277766
rect 173072 274712 173124 274718
rect 173072 274654 173124 274660
rect 172428 270496 172480 270502
rect 172428 270438 172480 270444
rect 173084 270366 173112 274654
rect 173452 271590 173480 277780
rect 174662 277766 175136 277794
rect 173440 271584 173492 271590
rect 173440 271526 173492 271532
rect 173072 270360 173124 270366
rect 173072 270302 173124 270308
rect 173716 269680 173768 269686
rect 173716 269622 173768 269628
rect 171784 267708 171836 267714
rect 171784 267650 171836 267656
rect 172060 266756 172112 266762
rect 172060 266698 172112 266704
rect 172072 264316 172100 266698
rect 172888 266484 172940 266490
rect 172888 266426 172940 266432
rect 172900 264316 172928 266426
rect 173728 264316 173756 269622
rect 175108 267306 175136 277766
rect 175844 271862 175872 277780
rect 176752 274508 176804 274514
rect 176752 274450 176804 274456
rect 175832 271856 175884 271862
rect 175832 271798 175884 271804
rect 175280 271720 175332 271726
rect 175280 271662 175332 271668
rect 174544 267300 174596 267306
rect 174544 267242 174596 267248
rect 175096 267300 175148 267306
rect 175096 267242 175148 267248
rect 174556 264316 174584 267242
rect 175292 264330 175320 271662
rect 176200 268252 176252 268258
rect 176200 268194 176252 268200
rect 175292 264302 175398 264330
rect 176212 264316 176240 268194
rect 176764 264330 176792 274450
rect 176948 274242 176976 277780
rect 178144 275738 178172 277780
rect 178132 275732 178184 275738
rect 178132 275674 178184 275680
rect 176936 274236 176988 274242
rect 176936 274178 176988 274184
rect 177488 273828 177540 273834
rect 177488 273770 177540 273776
rect 177500 264330 177528 273770
rect 178684 269544 178736 269550
rect 178684 269486 178736 269492
rect 176764 264302 177054 264330
rect 177500 264302 177882 264330
rect 178696 264316 178724 269486
rect 179340 268938 179368 277780
rect 180536 272814 180564 277780
rect 181732 275874 181760 277780
rect 181720 275868 181772 275874
rect 181720 275810 181772 275816
rect 182088 275052 182140 275058
rect 182088 274994 182140 275000
rect 180524 272808 180576 272814
rect 180524 272750 180576 272756
rect 179880 272400 179932 272406
rect 179880 272342 179932 272348
rect 179328 268932 179380 268938
rect 179328 268874 179380 268880
rect 179512 266620 179564 266626
rect 179512 266562 179564 266568
rect 179524 264316 179552 266562
rect 179892 264330 179920 272342
rect 181352 271040 181404 271046
rect 181352 270982 181404 270988
rect 181168 269816 181220 269822
rect 181168 269758 181220 269764
rect 179892 264302 180366 264330
rect 181180 264316 181208 269758
rect 181364 267734 181392 270982
rect 182100 269822 182128 274994
rect 182928 274514 182956 277780
rect 184138 277766 184796 277794
rect 183468 275324 183520 275330
rect 183468 275266 183520 275272
rect 182916 274508 182968 274514
rect 182916 274450 182968 274456
rect 182456 270904 182508 270910
rect 182456 270846 182508 270852
rect 182088 269816 182140 269822
rect 182088 269758 182140 269764
rect 182180 269272 182232 269278
rect 182180 269214 182232 269220
rect 181364 267706 181576 267734
rect 181548 264330 181576 267706
rect 182192 266422 182220 269214
rect 182180 266416 182232 266422
rect 182180 266358 182232 266364
rect 182468 264330 182496 270846
rect 183480 269550 183508 275266
rect 184204 273080 184256 273086
rect 184204 273022 184256 273028
rect 183468 269544 183520 269550
rect 183468 269486 183520 269492
rect 183652 268116 183704 268122
rect 183652 268058 183704 268064
rect 181548 264302 182022 264330
rect 182468 264302 182850 264330
rect 183664 264316 183692 268058
rect 184216 267034 184244 273022
rect 184768 269686 184796 277766
rect 185228 274718 185256 277780
rect 186424 275330 186452 277780
rect 186412 275324 186464 275330
rect 186412 275266 186464 275272
rect 185584 274916 185636 274922
rect 185584 274858 185636 274864
rect 185216 274712 185268 274718
rect 185216 274654 185268 274660
rect 185032 273692 185084 273698
rect 185032 273634 185084 273640
rect 184756 269680 184808 269686
rect 184756 269622 184808 269628
rect 184020 267028 184072 267034
rect 184020 266970 184072 266976
rect 184204 267028 184256 267034
rect 184204 266970 184256 266976
rect 184032 266762 184060 266970
rect 184480 266892 184532 266898
rect 184480 266834 184532 266840
rect 184020 266756 184072 266762
rect 184020 266698 184072 266704
rect 184492 264316 184520 266834
rect 185044 264330 185072 273634
rect 185596 269074 185624 274858
rect 187148 274712 187200 274718
rect 187148 274654 187200 274660
rect 186964 269816 187016 269822
rect 186964 269758 187016 269764
rect 185584 269068 185636 269074
rect 185584 269010 185636 269016
rect 186136 266416 186188 266422
rect 186136 266358 186188 266364
rect 185044 264302 185334 264330
rect 186148 264316 186176 266358
rect 186976 264316 187004 269758
rect 187160 267578 187188 274654
rect 187620 273086 187648 277780
rect 188816 275330 188844 277780
rect 187792 275324 187844 275330
rect 187792 275266 187844 275272
rect 188804 275324 188856 275330
rect 188804 275266 188856 275272
rect 187804 274378 187832 275266
rect 187792 274372 187844 274378
rect 187792 274314 187844 274320
rect 187792 273556 187844 273562
rect 187792 273498 187844 273504
rect 187608 273080 187660 273086
rect 187608 273022 187660 273028
rect 187804 272898 187832 273498
rect 187712 272870 187832 272898
rect 189816 272944 189868 272950
rect 189816 272886 189868 272892
rect 187332 269816 187384 269822
rect 187332 269758 187384 269764
rect 187344 269550 187372 269758
rect 187332 269544 187384 269550
rect 187332 269486 187384 269492
rect 187148 267572 187200 267578
rect 187148 267514 187200 267520
rect 187712 265674 187740 272870
rect 187884 270768 187936 270774
rect 187884 270710 187936 270716
rect 187700 265668 187752 265674
rect 187700 265610 187752 265616
rect 187896 265554 187924 270710
rect 189448 266756 189500 266762
rect 189448 266698 189500 266704
rect 188252 265668 188304 265674
rect 188252 265610 188304 265616
rect 187804 265526 187924 265554
rect 187804 264316 187832 265526
rect 188264 264330 188292 265610
rect 188264 264302 188646 264330
rect 189460 264316 189488 266698
rect 189828 264330 189856 272886
rect 190012 271046 190040 277780
rect 191208 272950 191236 277780
rect 191196 272944 191248 272950
rect 191196 272886 191248 272892
rect 190736 272264 190788 272270
rect 190736 272206 190788 272212
rect 190000 271040 190052 271046
rect 190000 270982 190052 270988
rect 190748 264330 190776 272206
rect 192312 271726 192340 277780
rect 193508 273970 193536 277780
rect 194704 277394 194732 277780
rect 194612 277366 194732 277394
rect 193864 276004 193916 276010
rect 193864 275946 193916 275952
rect 192484 273964 192536 273970
rect 192484 273906 192536 273912
rect 193496 273964 193548 273970
rect 193496 273906 193548 273912
rect 192300 271720 192352 271726
rect 192300 271662 192352 271668
rect 191932 269816 191984 269822
rect 191932 269758 191984 269764
rect 189828 264302 190302 264330
rect 190748 264302 191130 264330
rect 191944 264316 191972 269758
rect 192496 264330 192524 273906
rect 193588 268388 193640 268394
rect 193588 268330 193640 268336
rect 192496 264302 192786 264330
rect 193600 264316 193628 268330
rect 193876 267034 193904 275946
rect 194612 269822 194640 277366
rect 195900 274650 195928 277780
rect 197110 277766 197308 277794
rect 198306 277766 198688 277794
rect 195888 274644 195940 274650
rect 195888 274586 195940 274592
rect 195980 271312 196032 271318
rect 195980 271254 196032 271260
rect 194784 271176 194836 271182
rect 194784 271118 194836 271124
rect 194600 269816 194652 269822
rect 194600 269758 194652 269764
rect 194416 267164 194468 267170
rect 194416 267106 194468 267112
rect 193864 267028 193916 267034
rect 193864 266970 193916 266976
rect 194428 264316 194456 267106
rect 194796 264330 194824 271118
rect 195992 264330 196020 271254
rect 196900 269068 196952 269074
rect 196900 269010 196952 269016
rect 194796 264302 195270 264330
rect 195992 264302 196098 264330
rect 196912 264316 196940 269010
rect 197280 268394 197308 277766
rect 197544 272536 197596 272542
rect 197544 272478 197596 272484
rect 197268 268388 197320 268394
rect 197268 268330 197320 268336
rect 197556 264330 197584 272478
rect 198660 269958 198688 277766
rect 199488 272542 199516 277780
rect 200592 277394 200620 277780
rect 200500 277366 200620 277394
rect 199660 274508 199712 274514
rect 199660 274450 199712 274456
rect 199476 272536 199528 272542
rect 199476 272478 199528 272484
rect 198188 269952 198240 269958
rect 198188 269894 198240 269900
rect 198648 269952 198700 269958
rect 198648 269894 198700 269900
rect 198200 264330 198228 269894
rect 199384 267708 199436 267714
rect 199384 267650 199436 267656
rect 197556 264302 197754 264330
rect 198200 264302 198582 264330
rect 199396 264316 199424 267650
rect 199672 267170 199700 274450
rect 200500 270910 200528 277366
rect 201788 276010 201816 277780
rect 201776 276004 201828 276010
rect 201776 275946 201828 275952
rect 202144 275596 202196 275602
rect 202144 275538 202196 275544
rect 200672 274100 200724 274106
rect 200672 274042 200724 274048
rect 200488 270904 200540 270910
rect 200488 270846 200540 270852
rect 200212 268524 200264 268530
rect 200212 268466 200264 268472
rect 199660 267164 199712 267170
rect 199660 267106 199712 267112
rect 200224 264316 200252 268466
rect 200684 264330 200712 274042
rect 201868 267028 201920 267034
rect 201868 266970 201920 266976
rect 200684 264302 201066 264330
rect 201880 264316 201908 266970
rect 202156 266422 202184 275538
rect 202696 270088 202748 270094
rect 202696 270030 202748 270036
rect 202144 266416 202196 266422
rect 202144 266358 202196 266364
rect 202708 264316 202736 270030
rect 202984 268530 203012 277780
rect 203904 277766 204194 277794
rect 205390 277766 205588 277794
rect 203904 268802 203932 277766
rect 205560 270094 205588 277766
rect 206284 274644 206336 274650
rect 206284 274586 206336 274592
rect 205732 271448 205784 271454
rect 205732 271390 205784 271396
rect 205548 270088 205600 270094
rect 205548 270030 205600 270036
rect 203524 268796 203576 268802
rect 203524 268738 203576 268744
rect 203892 268796 203944 268802
rect 203892 268738 203944 268744
rect 202972 268524 203024 268530
rect 202972 268466 203024 268472
rect 203536 264316 203564 268738
rect 205180 268660 205232 268666
rect 205180 268602 205232 268608
rect 204352 267436 204404 267442
rect 204352 267378 204404 267384
rect 204364 264316 204392 267378
rect 205192 264316 205220 268602
rect 205744 264330 205772 271390
rect 206296 267034 206324 274586
rect 206572 274106 206600 277780
rect 207782 277766 208348 277794
rect 206560 274100 206612 274106
rect 206560 274042 206612 274048
rect 207664 271856 207716 271862
rect 207664 271798 207716 271804
rect 207388 270224 207440 270230
rect 207388 270166 207440 270172
rect 206284 267028 206336 267034
rect 206284 266970 206336 266976
rect 206836 266416 206888 266422
rect 206836 266358 206888 266364
rect 205744 264302 206034 264330
rect 206848 264316 206876 266358
rect 207400 264330 207428 270166
rect 207676 267714 207704 271798
rect 208320 269550 208348 277766
rect 208492 272672 208544 272678
rect 208492 272614 208544 272620
rect 208308 269544 208360 269550
rect 208308 269486 208360 269492
rect 207664 267708 207716 267714
rect 207664 267650 207716 267656
rect 207400 264302 207690 264330
rect 208504 264316 208532 272614
rect 208872 271182 208900 277780
rect 210068 274514 210096 277780
rect 210792 275460 210844 275466
rect 210792 275402 210844 275408
rect 210056 274508 210108 274514
rect 210056 274450 210108 274456
rect 208860 271176 208912 271182
rect 208860 271118 208912 271124
rect 210804 270502 210832 275402
rect 211264 273086 211292 277780
rect 211988 273216 212040 273222
rect 211988 273158 212040 273164
rect 211252 273080 211304 273086
rect 211252 273022 211304 273028
rect 208676 270496 208728 270502
rect 208676 270438 208728 270444
rect 210792 270496 210844 270502
rect 210792 270438 210844 270444
rect 211804 270496 211856 270502
rect 211804 270438 211856 270444
rect 208688 266626 208716 270438
rect 210148 270360 210200 270366
rect 210148 270302 210200 270308
rect 209320 266892 209372 266898
rect 209320 266834 209372 266840
rect 208676 266620 208728 266626
rect 208676 266562 208728 266568
rect 209332 264316 209360 266834
rect 210160 264316 210188 270302
rect 210976 266620 211028 266626
rect 210976 266562 211028 266568
rect 210988 264316 211016 266562
rect 211816 264316 211844 270438
rect 212000 267442 212028 273158
rect 212460 270366 212488 277780
rect 213670 277766 213868 277794
rect 212632 271584 212684 271590
rect 212632 271526 212684 271532
rect 212448 270360 212500 270366
rect 212448 270302 212500 270308
rect 211988 267436 212040 267442
rect 211988 267378 212040 267384
rect 212644 264316 212672 271526
rect 213840 270230 213868 277766
rect 214656 274236 214708 274242
rect 214656 274178 214708 274184
rect 213828 270224 213880 270230
rect 213828 270166 213880 270172
rect 213828 269680 213880 269686
rect 213828 269622 213880 269628
rect 213460 267708 213512 267714
rect 213460 267650 213512 267656
rect 213472 264316 213500 267650
rect 213840 266626 213868 269622
rect 214288 267300 214340 267306
rect 214288 267242 214340 267248
rect 213828 266620 213880 266626
rect 213828 266562 213880 266568
rect 214300 264316 214328 267242
rect 214668 264330 214696 274178
rect 214852 271862 214880 277780
rect 214840 271856 214892 271862
rect 214840 271798 214892 271804
rect 215956 271318 215984 277780
rect 217166 277766 217456 277794
rect 216864 275732 216916 275738
rect 216864 275674 216916 275680
rect 215944 271312 215996 271318
rect 215944 271254 215996 271260
rect 216128 271040 216180 271046
rect 216128 270982 216180 270988
rect 215944 268932 215996 268938
rect 215944 268874 215996 268880
rect 214668 264302 215142 264330
rect 215956 264316 215984 268874
rect 216140 266898 216168 270982
rect 216876 267734 216904 275674
rect 217232 272808 217284 272814
rect 217232 272750 217284 272756
rect 216784 267706 216904 267734
rect 216128 266892 216180 266898
rect 216128 266834 216180 266840
rect 216784 264316 216812 267706
rect 217244 264330 217272 272750
rect 217428 272678 217456 277766
rect 218348 275466 218376 277780
rect 218888 275868 218940 275874
rect 218888 275810 218940 275816
rect 218336 275460 218388 275466
rect 218336 275402 218388 275408
rect 217416 272672 217468 272678
rect 217416 272614 217468 272620
rect 218428 267164 218480 267170
rect 218428 267106 218480 267112
rect 217244 264302 217626 264330
rect 218440 264316 218468 267106
rect 218900 264330 218928 275810
rect 219544 268666 219572 277780
rect 220556 277766 220754 277794
rect 220556 274242 220584 277766
rect 221936 275602 221964 277780
rect 223146 277766 223528 277794
rect 223500 276026 223528 277766
rect 222108 276004 222160 276010
rect 223500 275998 223620 276026
rect 222108 275946 222160 275952
rect 221924 275596 221976 275602
rect 221924 275538 221976 275544
rect 220912 274372 220964 274378
rect 220912 274314 220964 274320
rect 220544 274236 220596 274242
rect 220544 274178 220596 274184
rect 220084 273080 220136 273086
rect 220084 273022 220136 273028
rect 219532 268660 219584 268666
rect 219532 268602 219584 268608
rect 220096 267306 220124 273022
rect 220084 267300 220136 267306
rect 220084 267242 220136 267248
rect 220084 266620 220136 266626
rect 220084 266562 220136 266568
rect 218900 264302 219282 264330
rect 220096 264316 220124 266562
rect 220924 264316 220952 274314
rect 222120 271862 222148 275946
rect 222844 275324 222896 275330
rect 222844 275266 222896 275272
rect 221464 271856 221516 271862
rect 221464 271798 221516 271804
rect 222108 271856 222160 271862
rect 222108 271798 222160 271804
rect 221476 267170 221504 271798
rect 221740 267572 221792 267578
rect 221740 267514 221792 267520
rect 221464 267164 221516 267170
rect 221464 267106 221516 267112
rect 221752 264316 221780 267514
rect 222568 267436 222620 267442
rect 222568 267378 222620 267384
rect 222580 264316 222608 267378
rect 222856 266422 222884 275266
rect 223592 271454 223620 275998
rect 224236 275126 224264 277780
rect 225432 275330 225460 277780
rect 225420 275324 225472 275330
rect 225420 275266 225472 275272
rect 224224 275120 224276 275126
rect 224224 275062 224276 275068
rect 226156 275120 226208 275126
rect 226156 275062 226208 275068
rect 224868 272944 224920 272950
rect 224920 272892 225000 272898
rect 224868 272886 225000 272892
rect 224880 272870 225000 272886
rect 223580 271448 223632 271454
rect 223580 271390 223632 271396
rect 224224 270904 224276 270910
rect 224224 270846 224276 270852
rect 224236 267442 224264 270846
rect 224224 267436 224276 267442
rect 224224 267378 224276 267384
rect 223396 266892 223448 266898
rect 223396 266834 223448 266840
rect 222844 266416 222896 266422
rect 222844 266358 222896 266364
rect 223408 264316 223436 266834
rect 224224 266416 224276 266422
rect 224224 266358 224276 266364
rect 224236 264316 224264 266358
rect 224972 264330 225000 272870
rect 225512 271720 225564 271726
rect 225512 271662 225564 271668
rect 225524 264330 225552 271662
rect 226168 271590 226196 275062
rect 226340 273964 226392 273970
rect 226340 273906 226392 273912
rect 226156 271584 226208 271590
rect 226156 271526 226208 271532
rect 226352 264330 226380 273906
rect 226628 269686 226656 277780
rect 227824 277394 227852 277780
rect 228836 277766 229034 277794
rect 230230 277766 230428 277794
rect 227824 277366 227944 277394
rect 227260 269816 227312 269822
rect 227260 269758 227312 269764
rect 226616 269680 226668 269686
rect 226616 269622 226668 269628
rect 227272 264330 227300 269758
rect 227916 268802 227944 277366
rect 228836 272814 228864 277766
rect 228824 272808 228876 272814
rect 228824 272750 228876 272756
rect 230400 269958 230428 277766
rect 231412 272542 231440 277780
rect 232530 277766 233188 277794
rect 230572 272536 230624 272542
rect 230572 272478 230624 272484
rect 231400 272536 231452 272542
rect 231400 272478 231452 272484
rect 230020 269952 230072 269958
rect 230020 269894 230072 269900
rect 230388 269952 230440 269958
rect 230388 269894 230440 269900
rect 227720 268796 227772 268802
rect 227720 268738 227772 268744
rect 227904 268796 227956 268802
rect 227904 268738 227956 268744
rect 227732 267578 227760 268738
rect 229192 268388 229244 268394
rect 229192 268330 229244 268336
rect 227720 267572 227772 267578
rect 227720 267514 227772 267520
rect 228364 267028 228416 267034
rect 228364 266970 228416 266976
rect 224972 264302 225078 264330
rect 225524 264302 225906 264330
rect 226352 264302 226734 264330
rect 227272 264302 227562 264330
rect 228376 264316 228404 266970
rect 229204 264316 229232 268330
rect 230032 264316 230060 269894
rect 230584 264330 230612 272478
rect 232136 271856 232188 271862
rect 232136 271798 232188 271804
rect 230756 269544 230808 269550
rect 230756 269486 230808 269492
rect 230768 266422 230796 269486
rect 231676 267436 231728 267442
rect 231676 267378 231728 267384
rect 230756 266416 230808 266422
rect 230756 266358 230808 266364
rect 230584 264302 230874 264330
rect 231688 264316 231716 267378
rect 232148 264330 232176 271798
rect 233160 270502 233188 277766
rect 233148 270496 233200 270502
rect 233148 270438 233200 270444
rect 233332 268524 233384 268530
rect 233332 268466 233384 268472
rect 232148 264302 232530 264330
rect 233344 264316 233372 268466
rect 233712 268394 233740 277780
rect 233884 275596 233936 275602
rect 233884 275538 233936 275544
rect 233700 268388 233752 268394
rect 233700 268330 233752 268336
rect 233896 267442 233924 275538
rect 234908 273970 234936 277780
rect 236104 275602 236132 277780
rect 236092 275596 236144 275602
rect 236092 275538 236144 275544
rect 235448 274100 235500 274106
rect 235448 274042 235500 274048
rect 234896 273964 234948 273970
rect 234896 273906 234948 273912
rect 234988 270088 235040 270094
rect 234988 270030 235040 270036
rect 234160 267572 234212 267578
rect 234160 267514 234212 267520
rect 233884 267436 233936 267442
rect 233884 267378 233936 267384
rect 234172 264316 234200 267514
rect 235000 264316 235028 270030
rect 235460 264330 235488 274042
rect 237300 270638 237328 277780
rect 237472 275460 237524 275466
rect 237472 275402 237524 275408
rect 237484 271726 237512 275402
rect 238496 274718 238524 277780
rect 238484 274712 238536 274718
rect 238484 274654 238536 274660
rect 237840 274508 237892 274514
rect 237840 274450 237892 274456
rect 237472 271720 237524 271726
rect 237472 271662 237524 271668
rect 237472 271176 237524 271182
rect 237472 271118 237524 271124
rect 237288 270632 237340 270638
rect 237288 270574 237340 270580
rect 237288 270496 237340 270502
rect 237288 270438 237340 270444
rect 237300 267034 237328 270438
rect 237288 267028 237340 267034
rect 237288 266970 237340 266976
rect 236644 266416 236696 266422
rect 236644 266358 236696 266364
rect 235460 264302 235842 264330
rect 236656 264316 236684 266358
rect 237484 264316 237512 271118
rect 237852 264330 237880 274450
rect 239600 274106 239628 277780
rect 239772 274712 239824 274718
rect 239772 274654 239824 274660
rect 239588 274100 239640 274106
rect 239588 274042 239640 274048
rect 239784 270094 239812 274654
rect 240600 274236 240652 274242
rect 240600 274178 240652 274184
rect 240612 270994 240640 274178
rect 240796 271182 240824 277780
rect 242006 277766 242388 277794
rect 242360 272678 242388 277766
rect 242164 272672 242216 272678
rect 242164 272614 242216 272620
rect 242348 272672 242400 272678
rect 242348 272614 242400 272620
rect 242176 271402 242204 272614
rect 242176 271374 242296 271402
rect 242072 271312 242124 271318
rect 242072 271254 242124 271260
rect 240784 271176 240836 271182
rect 240784 271118 240836 271124
rect 240612 270966 240732 270994
rect 239956 270360 240008 270366
rect 239956 270302 240008 270308
rect 239772 270088 239824 270094
rect 239772 270030 239824 270036
rect 239128 267300 239180 267306
rect 239128 267242 239180 267248
rect 237852 264302 238326 264330
rect 239140 264316 239168 267242
rect 239968 264316 239996 270302
rect 240508 270224 240560 270230
rect 240508 270166 240560 270172
rect 240520 264330 240548 270166
rect 240704 266558 240732 270966
rect 241612 267164 241664 267170
rect 241612 267106 241664 267112
rect 240692 266552 240744 266558
rect 240692 266494 240744 266500
rect 240520 264302 240810 264330
rect 241624 264316 241652 267106
rect 242084 264330 242112 271254
rect 242268 266422 242296 271374
rect 243188 271318 243216 277780
rect 244384 275466 244412 277780
rect 244372 275460 244424 275466
rect 244372 275402 244424 275408
rect 245108 275324 245160 275330
rect 245108 275266 245160 275272
rect 243728 271720 243780 271726
rect 243728 271662 243780 271668
rect 243176 271312 243228 271318
rect 243176 271254 243228 271260
rect 242256 266416 242308 266422
rect 242256 266358 242308 266364
rect 243268 266416 243320 266422
rect 243268 266358 243320 266364
rect 242084 264302 242466 264330
rect 243280 264316 243308 266358
rect 243740 264330 243768 271662
rect 244924 268660 244976 268666
rect 244924 268602 244976 268608
rect 243740 264302 244122 264330
rect 244936 264316 244964 268602
rect 245120 266762 245148 275266
rect 245580 268530 245608 277780
rect 246776 277394 246804 277780
rect 246776 277366 246896 277394
rect 245568 268524 245620 268530
rect 245568 268466 245620 268472
rect 246580 267436 246632 267442
rect 246580 267378 246632 267384
rect 245108 266756 245160 266762
rect 245108 266698 245160 266704
rect 245752 266552 245804 266558
rect 245752 266494 245804 266500
rect 245764 264316 245792 266494
rect 246592 264316 246620 267378
rect 246868 267170 246896 277366
rect 247132 271584 247184 271590
rect 247132 271526 247184 271532
rect 246856 267164 246908 267170
rect 246856 267106 246908 267112
rect 247144 265674 247172 271526
rect 247880 271454 247908 277780
rect 249090 277766 249656 277794
rect 249064 272808 249116 272814
rect 249064 272750 249116 272756
rect 247316 271448 247368 271454
rect 247316 271390 247368 271396
rect 247868 271448 247920 271454
rect 247868 271390 247920 271396
rect 247132 265668 247184 265674
rect 247132 265610 247184 265616
rect 247328 264330 247356 271390
rect 249076 266898 249104 272750
rect 249628 270230 249656 277766
rect 250272 275330 250300 277780
rect 251088 275596 251140 275602
rect 251088 275538 251140 275544
rect 250260 275324 250312 275330
rect 250260 275266 250312 275272
rect 249616 270224 249668 270230
rect 249616 270166 249668 270172
rect 249892 269816 249944 269822
rect 249892 269758 249944 269764
rect 249064 266892 249116 266898
rect 249064 266834 249116 266840
rect 249064 266756 249116 266762
rect 249064 266698 249116 266704
rect 247868 265668 247920 265674
rect 247868 265610 247920 265616
rect 247880 264330 247908 265610
rect 247328 264302 247434 264330
rect 247880 264302 248262 264330
rect 249076 264316 249104 266698
rect 249904 264316 249932 269758
rect 251100 269074 251128 275538
rect 251468 269822 251496 277780
rect 252678 277766 252968 277794
rect 252940 272542 252968 277766
rect 252744 272536 252796 272542
rect 252744 272478 252796 272484
rect 252928 272536 252980 272542
rect 252928 272478 252980 272484
rect 252008 270496 252060 270502
rect 252008 270438 252060 270444
rect 251456 269816 251508 269822
rect 251456 269758 251508 269764
rect 251088 269068 251140 269074
rect 251088 269010 251140 269016
rect 250720 268796 250772 268802
rect 250720 268738 250772 268744
rect 250732 264316 250760 268738
rect 251548 266892 251600 266898
rect 251548 266834 251600 266840
rect 251560 264316 251588 266834
rect 252020 266422 252048 270438
rect 252376 269952 252428 269958
rect 252376 269894 252428 269900
rect 252008 266416 252060 266422
rect 252008 266358 252060 266364
rect 252388 264316 252416 269894
rect 252756 264330 252784 272478
rect 253860 270366 253888 277780
rect 254584 275460 254636 275466
rect 254584 275402 254636 275408
rect 253848 270360 253900 270366
rect 253848 270302 253900 270308
rect 253204 270088 253256 270094
rect 253204 270030 253256 270036
rect 253216 269686 253244 270030
rect 253204 269680 253256 269686
rect 253204 269622 253256 269628
rect 254596 267306 254624 275402
rect 255056 274666 255084 277780
rect 255056 274638 255360 274666
rect 255332 268394 255360 274638
rect 256160 273970 256188 277780
rect 257370 277766 258028 277794
rect 255504 273964 255556 273970
rect 255504 273906 255556 273912
rect 256148 273964 256200 273970
rect 256148 273906 256200 273912
rect 254860 268388 254912 268394
rect 254860 268330 254912 268336
rect 255320 268388 255372 268394
rect 255320 268330 255372 268336
rect 254584 267300 254636 267306
rect 254584 267242 254636 267248
rect 254032 267028 254084 267034
rect 254032 266970 254084 266976
rect 252756 264302 253230 264330
rect 254044 264316 254072 266970
rect 254872 264316 254900 268330
rect 255516 264330 255544 273906
rect 256516 269068 256568 269074
rect 256516 269010 256568 269016
rect 255516 264302 255714 264330
rect 256528 264316 256556 269010
rect 258000 266898 258028 277766
rect 258552 277394 258580 277780
rect 258460 277366 258580 277394
rect 258460 269958 258488 277366
rect 258632 274100 258684 274106
rect 258632 274042 258684 274048
rect 258448 269952 258500 269958
rect 258448 269894 258500 269900
rect 258172 269680 258224 269686
rect 258172 269622 258224 269628
rect 257988 266892 258040 266898
rect 257988 266834 258040 266840
rect 257344 266416 257396 266422
rect 257344 266358 257396 266364
rect 257356 264316 257384 266358
rect 258184 264316 258212 269622
rect 258644 264330 258672 274042
rect 259552 272672 259604 272678
rect 259552 272614 259604 272620
rect 259564 265674 259592 272614
rect 259748 271590 259776 277780
rect 260944 275466 260972 277780
rect 260932 275460 260984 275466
rect 260932 275402 260984 275408
rect 259736 271584 259788 271590
rect 259736 271526 259788 271532
rect 261024 271312 261076 271318
rect 261024 271254 261076 271260
rect 259828 271176 259880 271182
rect 259828 271118 259880 271124
rect 259552 265668 259604 265674
rect 259552 265610 259604 265616
rect 258644 264302 259026 264330
rect 259840 264316 259868 271118
rect 260380 265668 260432 265674
rect 260380 265610 260432 265616
rect 260392 264330 260420 265610
rect 261036 264330 261064 271254
rect 262140 271182 262168 277780
rect 263258 277766 263548 277794
rect 264454 277766 264928 277794
rect 265650 277766 266216 277794
rect 262128 271176 262180 271182
rect 262128 271118 262180 271124
rect 263324 270224 263376 270230
rect 263324 270166 263376 270172
rect 263140 268524 263192 268530
rect 263140 268466 263192 268472
rect 262312 267300 262364 267306
rect 262312 267242 262364 267248
rect 260392 264302 260682 264330
rect 261036 264302 261510 264330
rect 262324 264316 262352 267242
rect 263152 264316 263180 268466
rect 263336 266422 263364 270166
rect 263520 268530 263548 277766
rect 264336 271448 264388 271454
rect 264336 271390 264388 271396
rect 263508 268524 263560 268530
rect 263508 268466 263560 268472
rect 263968 267164 264020 267170
rect 263968 267106 264020 267112
rect 263324 266416 263376 266422
rect 263324 266358 263376 266364
rect 263980 264316 264008 267106
rect 264348 264330 264376 271390
rect 264900 269278 264928 277766
rect 265072 270360 265124 270366
rect 265072 270302 265124 270308
rect 264888 269272 264940 269278
rect 264888 269214 264940 269220
rect 265084 266830 265112 270302
rect 266188 270094 266216 277766
rect 266832 275330 266860 277780
rect 266360 275324 266412 275330
rect 266360 275266 266412 275272
rect 266820 275324 266872 275330
rect 266820 275266 266872 275272
rect 266176 270088 266228 270094
rect 266176 270030 266228 270036
rect 265072 266824 265124 266830
rect 265072 266766 265124 266772
rect 265624 266416 265676 266422
rect 265624 266358 265676 266364
rect 264348 264302 264822 264330
rect 265636 264316 265664 266358
rect 266372 264330 266400 275266
rect 268028 272542 268056 277780
rect 267740 272536 267792 272542
rect 267740 272478 267792 272484
rect 268016 272536 268068 272542
rect 268016 272478 268068 272484
rect 267280 269816 267332 269822
rect 267280 269758 267332 269764
rect 266372 264302 266478 264330
rect 267292 264316 267320 269758
rect 267752 264330 267780 272478
rect 269224 270230 269252 277780
rect 270420 277394 270448 277780
rect 270328 277366 270448 277394
rect 269212 270224 269264 270230
rect 269212 270166 269264 270172
rect 270328 269822 270356 277366
rect 271524 273970 271552 277780
rect 272734 277766 273116 277794
rect 270592 273964 270644 273970
rect 270592 273906 270644 273912
rect 271512 273964 271564 273970
rect 271512 273906 271564 273912
rect 270316 269816 270368 269822
rect 270316 269758 270368 269764
rect 269120 269272 269172 269278
rect 269120 269214 269172 269220
rect 268936 266824 268988 266830
rect 268936 266766 268988 266772
rect 267752 264302 268134 264330
rect 268948 264316 268976 266766
rect 269132 266422 269160 269214
rect 269764 268388 269816 268394
rect 269764 268330 269816 268336
rect 269120 266416 269172 266422
rect 269120 266358 269172 266364
rect 269776 264316 269804 268330
rect 270604 264316 270632 273906
rect 272616 271584 272668 271590
rect 272616 271526 272668 271532
rect 272248 269952 272300 269958
rect 272248 269894 272300 269900
rect 271420 267028 271472 267034
rect 271420 266970 271472 266976
rect 271432 264316 271460 266970
rect 272260 264316 272288 269894
rect 272628 264330 272656 271526
rect 273088 269958 273116 277766
rect 273916 275466 273944 277780
rect 273536 275460 273588 275466
rect 273536 275402 273588 275408
rect 273904 275460 273956 275466
rect 273904 275402 273956 275408
rect 273076 269952 273128 269958
rect 273076 269894 273128 269900
rect 273548 264330 273576 275402
rect 275112 271318 275140 277780
rect 275100 271312 275152 271318
rect 275100 271254 275152 271260
rect 276308 271182 276336 277780
rect 276664 275324 276716 275330
rect 276664 275266 276716 275272
rect 274640 271176 274692 271182
rect 274640 271118 274692 271124
rect 276296 271176 276348 271182
rect 276296 271118 276348 271124
rect 274652 264330 274680 271118
rect 275560 268524 275612 268530
rect 275560 268466 275612 268472
rect 272628 264302 273102 264330
rect 273548 264302 273930 264330
rect 274652 264302 274758 264330
rect 275572 264316 275600 268466
rect 276676 267034 276704 275266
rect 277504 274990 277532 277780
rect 278700 277394 278728 277780
rect 278608 277366 278728 277394
rect 277492 274984 277544 274990
rect 277492 274926 277544 274932
rect 277216 270088 277268 270094
rect 277216 270030 277268 270036
rect 276664 267028 276716 267034
rect 276664 266970 276716 266976
rect 276388 266416 276440 266422
rect 276388 266358 276440 266364
rect 276400 264316 276428 266358
rect 277228 264316 277256 270030
rect 278044 267028 278096 267034
rect 278044 266970 278096 266976
rect 278056 264316 278084 266970
rect 278608 266422 278636 277366
rect 279804 272542 279832 277780
rect 280804 273964 280856 273970
rect 280804 273906 280856 273912
rect 278780 272536 278832 272542
rect 278780 272478 278832 272484
rect 279792 272536 279844 272542
rect 279792 272478 279844 272484
rect 278596 266416 278648 266422
rect 278596 266358 278648 266364
rect 278792 264330 278820 272478
rect 279700 270224 279752 270230
rect 279700 270166 279752 270172
rect 278792 264302 278898 264330
rect 279712 264316 279740 270166
rect 280528 269816 280580 269822
rect 280528 269758 280580 269764
rect 280540 264316 280568 269758
rect 280816 267734 280844 273906
rect 281000 273766 281028 277780
rect 282210 277766 282776 277794
rect 280988 273760 281040 273766
rect 280988 273702 281040 273708
rect 282184 269952 282236 269958
rect 282184 269894 282236 269900
rect 280816 267706 280936 267734
rect 280908 264330 280936 267706
rect 280908 264302 281382 264330
rect 282196 264316 282224 269894
rect 282748 269142 282776 277766
rect 282920 275460 282972 275466
rect 282920 275402 282972 275408
rect 282736 269136 282788 269142
rect 282736 269078 282788 269084
rect 282932 264330 282960 275402
rect 283392 274854 283420 277780
rect 284588 275330 284616 277780
rect 284576 275324 284628 275330
rect 284576 275266 284628 275272
rect 284300 274984 284352 274990
rect 284300 274926 284352 274932
rect 283380 274848 283432 274854
rect 283380 274790 283432 274796
rect 283472 271312 283524 271318
rect 283472 271254 283524 271260
rect 283484 264330 283512 271254
rect 284312 265674 284340 274926
rect 285784 274718 285812 277780
rect 286888 277394 286916 277780
rect 286796 277366 286916 277394
rect 285772 274712 285824 274718
rect 285772 274654 285824 274660
rect 284484 271176 284536 271182
rect 284484 271118 284536 271124
rect 284300 265668 284352 265674
rect 284300 265610 284352 265616
rect 284496 264330 284524 271118
rect 286796 269958 286824 277366
rect 286968 274712 287020 274718
rect 286968 274654 287020 274660
rect 286784 269952 286836 269958
rect 286784 269894 286836 269900
rect 286980 267034 287008 274654
rect 287520 273760 287572 273766
rect 287520 273702 287572 273708
rect 287152 272536 287204 272542
rect 287152 272478 287204 272484
rect 286968 267028 287020 267034
rect 286968 266970 287020 266976
rect 286324 266416 286376 266422
rect 286324 266358 286376 266364
rect 285220 265668 285272 265674
rect 285220 265610 285272 265616
rect 285232 264330 285260 265610
rect 282932 264302 283038 264330
rect 283484 264302 283866 264330
rect 284496 264302 284694 264330
rect 285232 264302 285522 264330
rect 286336 264316 286364 266358
rect 287164 264316 287192 272478
rect 287532 264330 287560 273702
rect 288084 272950 288112 277780
rect 289280 274922 289308 277780
rect 290096 275324 290148 275330
rect 290096 275266 290148 275272
rect 289268 274916 289320 274922
rect 289268 274858 289320 274864
rect 289084 274848 289136 274854
rect 289084 274790 289136 274796
rect 288072 272944 288124 272950
rect 288072 272886 288124 272892
rect 288808 269136 288860 269142
rect 288808 269078 288860 269084
rect 287532 264302 288006 264330
rect 288820 264316 288848 269078
rect 289096 267734 289124 274790
rect 289096 267706 289216 267734
rect 289188 264330 289216 267706
rect 290108 264330 290136 275266
rect 290476 274718 290504 277780
rect 290464 274712 290516 274718
rect 290464 274654 290516 274660
rect 290464 272944 290516 272950
rect 290464 272886 290516 272892
rect 290476 266422 290504 272886
rect 291672 270366 291700 277780
rect 292868 270502 292896 277780
rect 294064 275126 294092 277780
rect 295168 275210 295196 277780
rect 295168 275182 295380 275210
rect 294052 275120 294104 275126
rect 294052 275062 294104 275068
rect 295156 275120 295208 275126
rect 295156 275062 295208 275068
rect 293408 274916 293460 274922
rect 293408 274858 293460 274864
rect 292856 270496 292908 270502
rect 292856 270438 292908 270444
rect 291660 270360 291712 270366
rect 291660 270302 291712 270308
rect 292120 269952 292172 269958
rect 292120 269894 292172 269900
rect 291292 267028 291344 267034
rect 291292 266970 291344 266976
rect 290464 266416 290516 266422
rect 290464 266358 290516 266364
rect 289188 264302 289662 264330
rect 290108 264302 290490 264330
rect 291304 264316 291332 266970
rect 292132 264316 292160 269894
rect 292948 266416 293000 266422
rect 292948 266358 293000 266364
rect 292960 264316 292988 266358
rect 293420 264330 293448 274858
rect 294144 274712 294196 274718
rect 294144 274654 294196 274660
rect 294156 264330 294184 274654
rect 295168 267034 295196 275062
rect 295352 269142 295380 275182
rect 296364 274718 296392 277780
rect 297574 277766 297956 277794
rect 296352 274712 296404 274718
rect 296352 274654 296404 274660
rect 296260 270496 296312 270502
rect 296260 270438 296312 270444
rect 295524 270360 295576 270366
rect 295524 270302 295576 270308
rect 295340 269136 295392 269142
rect 295340 269078 295392 269084
rect 295536 267734 295564 270302
rect 295444 267706 295564 267734
rect 295156 267028 295208 267034
rect 295156 266970 295208 266976
rect 293420 264302 293802 264330
rect 294156 264302 294630 264330
rect 295444 264316 295472 267706
rect 296272 264316 296300 270438
rect 297548 269136 297600 269142
rect 297548 269078 297600 269084
rect 297088 267028 297140 267034
rect 297088 266970 297140 266976
rect 297100 264316 297128 266970
rect 297560 264330 297588 269078
rect 297928 266422 297956 277766
rect 298756 275398 298784 277780
rect 299952 275738 299980 277780
rect 300964 277766 301162 277794
rect 299940 275732 299992 275738
rect 299940 275674 299992 275680
rect 300768 275732 300820 275738
rect 300768 275674 300820 275680
rect 298744 275392 298796 275398
rect 298744 275334 298796 275340
rect 300032 275392 300084 275398
rect 300032 275334 300084 275340
rect 298376 274712 298428 274718
rect 298376 274654 298428 274660
rect 297916 266416 297968 266422
rect 297916 266358 297968 266364
rect 298388 264330 298416 274654
rect 299572 266416 299624 266422
rect 299572 266358 299624 266364
rect 297560 264302 297942 264330
rect 298388 264302 298770 264330
rect 299584 264316 299612 266358
rect 300044 264330 300072 275334
rect 300780 267734 300808 275674
rect 300964 267734 300992 277766
rect 302344 277394 302372 277780
rect 303448 277394 303476 277780
rect 303724 277766 304658 277794
rect 305012 277766 305854 277794
rect 306392 277766 307050 277794
rect 307772 277766 308246 277794
rect 302344 277366 302464 277394
rect 303448 277366 303568 277394
rect 300780 267706 300900 267734
rect 300964 267706 301084 267734
rect 300872 264330 300900 267706
rect 301056 266422 301084 267706
rect 301044 266416 301096 266422
rect 301044 266358 301096 266364
rect 302056 266416 302108 266422
rect 302056 266358 302108 266364
rect 300044 264302 300426 264330
rect 300872 264302 301254 264330
rect 302068 264316 302096 266358
rect 302436 264330 302464 277366
rect 303540 267734 303568 277366
rect 303724 267734 303752 277766
rect 303540 267706 303660 267734
rect 303724 267706 304120 267734
rect 303632 264330 303660 267706
rect 304092 264330 304120 267706
rect 305012 264330 305040 277766
rect 306392 266370 306420 277766
rect 307772 267734 307800 277766
rect 309428 277394 309456 277780
rect 310546 277766 310928 277794
rect 309428 277366 309548 277394
rect 306208 266342 306420 266370
rect 307496 267706 307800 267734
rect 302436 264302 302910 264330
rect 303632 264302 303738 264330
rect 304092 264302 304566 264330
rect 305012 264302 305394 264330
rect 306208 264316 306236 266342
rect 307496 264330 307524 267706
rect 308680 266552 308732 266558
rect 308680 266494 308732 266500
rect 307852 266416 307904 266422
rect 307852 266358 307904 266364
rect 307050 264302 307524 264330
rect 307864 264316 307892 266358
rect 308692 264316 308720 266494
rect 309520 266422 309548 277366
rect 309784 270156 309836 270162
rect 309784 270098 309836 270104
rect 309508 266416 309560 266422
rect 309508 266358 309560 266364
rect 309796 264330 309824 270098
rect 310900 266558 310928 277766
rect 311360 277766 311742 277794
rect 311912 277766 312938 277794
rect 313292 277766 314134 277794
rect 314672 277766 315330 277794
rect 316052 277766 316526 277794
rect 311360 270162 311388 277766
rect 311348 270156 311400 270162
rect 311348 270098 311400 270104
rect 310888 266552 310940 266558
rect 310888 266494 310940 266500
rect 311164 266552 311216 266558
rect 311164 266494 311216 266500
rect 310336 266416 310388 266422
rect 310336 266358 310388 266364
rect 309534 264302 309824 264330
rect 310348 264316 310376 266358
rect 311176 264316 311204 266494
rect 311912 266422 311940 277766
rect 312820 267300 312872 267306
rect 312820 267242 312872 267248
rect 311900 266416 311952 266422
rect 311900 266358 311952 266364
rect 312360 266416 312412 266422
rect 312360 266358 312412 266364
rect 312372 264330 312400 266358
rect 312018 264302 312400 264330
rect 312832 264316 312860 267242
rect 313292 266558 313320 277766
rect 314476 269816 314528 269822
rect 314476 269758 314528 269764
rect 313648 267436 313700 267442
rect 313648 267378 313700 267384
rect 313280 266552 313332 266558
rect 313280 266494 313332 266500
rect 313660 264316 313688 267378
rect 314488 264316 314516 269758
rect 314672 266422 314700 277766
rect 315764 271312 315816 271318
rect 315764 271254 315816 271260
rect 314660 266416 314712 266422
rect 314660 266358 314712 266364
rect 315776 264330 315804 271254
rect 316052 267306 316080 277766
rect 317708 277394 317736 277780
rect 318826 277766 319024 277794
rect 317708 277366 317828 277394
rect 316960 270292 317012 270298
rect 316960 270234 317012 270240
rect 316040 267300 316092 267306
rect 316040 267242 316092 267248
rect 316132 266892 316184 266898
rect 316132 266834 316184 266840
rect 315330 264302 315804 264330
rect 316144 264316 316172 266834
rect 316972 264316 317000 270234
rect 317800 267442 317828 277366
rect 318616 271788 318668 271794
rect 318616 271730 318668 271736
rect 317788 267436 317840 267442
rect 317788 267378 317840 267384
rect 317788 266416 317840 266422
rect 317788 266358 317840 266364
rect 317800 264316 317828 266358
rect 318628 264316 318656 271730
rect 318996 269822 319024 277766
rect 320008 271318 320036 277780
rect 320192 277766 321218 277794
rect 321572 277766 322414 277794
rect 323136 277766 323610 277794
rect 319996 271312 320048 271318
rect 319996 271254 320048 271260
rect 318984 269816 319036 269822
rect 318984 269758 319036 269764
rect 319444 269136 319496 269142
rect 319444 269078 319496 269084
rect 319456 264316 319484 269078
rect 320192 266898 320220 277766
rect 321572 270298 321600 277766
rect 321560 270292 321612 270298
rect 321560 270234 321612 270240
rect 321928 270224 321980 270230
rect 321928 270166 321980 270172
rect 321100 269272 321152 269278
rect 321100 269214 321152 269220
rect 320180 266892 320232 266898
rect 320180 266834 320232 266840
rect 320272 266756 320324 266762
rect 320272 266698 320324 266704
rect 320284 264316 320312 266698
rect 321112 264316 321140 269214
rect 321940 264316 321968 270166
rect 322756 268388 322808 268394
rect 322756 268330 322808 268336
rect 322768 264316 322796 268330
rect 323136 266422 323164 277766
rect 324792 271794 324820 277780
rect 325712 277766 326002 277794
rect 327106 277766 327488 277794
rect 324780 271788 324832 271794
rect 324780 271730 324832 271736
rect 325516 271312 325568 271318
rect 325516 271254 325568 271260
rect 323584 270088 323636 270094
rect 323584 270030 323636 270036
rect 323124 266416 323176 266422
rect 323124 266358 323176 266364
rect 323596 264316 323624 270030
rect 324412 267028 324464 267034
rect 324412 266970 324464 266976
rect 324424 264316 324452 266970
rect 325528 264330 325556 271254
rect 325712 269142 325740 277766
rect 326436 275460 326488 275466
rect 326436 275402 326488 275408
rect 325700 269136 325752 269142
rect 325700 269078 325752 269084
rect 326448 264330 326476 275402
rect 326896 269952 326948 269958
rect 326896 269894 326948 269900
rect 325266 264302 325556 264330
rect 326094 264302 326476 264330
rect 326908 264316 326936 269894
rect 327460 266762 327488 277766
rect 327920 277766 328302 277794
rect 328472 277766 329498 277794
rect 329852 277766 330694 277794
rect 331232 277766 331890 277794
rect 332612 277766 333086 277794
rect 327920 269278 327948 277766
rect 328472 270230 328500 277766
rect 329472 275324 329524 275330
rect 329472 275266 329524 275272
rect 328460 270224 328512 270230
rect 328460 270166 328512 270172
rect 327908 269272 327960 269278
rect 327908 269214 327960 269220
rect 327448 266756 327500 266762
rect 327448 266698 327500 266704
rect 327724 266552 327776 266558
rect 327724 266494 327776 266500
rect 327736 264316 327764 266494
rect 329484 266422 329512 275266
rect 329656 269816 329708 269822
rect 329656 269758 329708 269764
rect 328552 266416 328604 266422
rect 328552 266358 328604 266364
rect 329472 266416 329524 266422
rect 329472 266358 329524 266364
rect 328564 264316 328592 266358
rect 329668 264330 329696 269758
rect 329852 268394 329880 277766
rect 331036 272672 331088 272678
rect 331036 272614 331088 272620
rect 329840 268388 329892 268394
rect 329840 268330 329892 268336
rect 330208 266688 330260 266694
rect 330208 266630 330260 266636
rect 329406 264302 329696 264330
rect 330220 264316 330248 266630
rect 331048 264316 331076 272614
rect 331232 270094 331260 277766
rect 332612 270494 332640 277766
rect 334176 271318 334204 277780
rect 335372 275466 335400 277780
rect 335924 277766 336582 277794
rect 336752 277766 337778 277794
rect 335360 275460 335412 275466
rect 335360 275402 335412 275408
rect 334624 271448 334676 271454
rect 334624 271390 334676 271396
rect 334164 271312 334216 271318
rect 334164 271254 334216 271260
rect 333888 271176 333940 271182
rect 333888 271118 333940 271124
rect 332520 270466 332640 270494
rect 331220 270088 331272 270094
rect 331220 270030 331272 270036
rect 332324 270088 332376 270094
rect 332324 270030 332376 270036
rect 331864 266892 331916 266898
rect 331864 266834 331916 266840
rect 331876 264316 331904 266834
rect 332336 266558 332364 270030
rect 332520 267034 332548 270466
rect 333520 268524 333572 268530
rect 333520 268466 333572 268472
rect 332508 267028 332560 267034
rect 332508 266970 332560 266976
rect 332324 266552 332376 266558
rect 332324 266494 332376 266500
rect 332692 266416 332744 266422
rect 332692 266358 332744 266364
rect 332704 264316 332732 266358
rect 333532 264316 333560 268466
rect 333900 266422 333928 271118
rect 334348 267436 334400 267442
rect 334348 267378 334400 267384
rect 333888 266416 333940 266422
rect 333888 266358 333940 266364
rect 334360 264316 334388 267378
rect 334636 266694 334664 271390
rect 335924 269958 335952 277766
rect 336752 270094 336780 277766
rect 338960 275330 338988 277780
rect 339512 277766 340170 277794
rect 338948 275324 339000 275330
rect 338948 275266 339000 275272
rect 338948 275188 339000 275194
rect 338948 275130 339000 275136
rect 338028 272536 338080 272542
rect 338028 272478 338080 272484
rect 336740 270088 336792 270094
rect 336740 270030 336792 270036
rect 335912 269952 335964 269958
rect 335912 269894 335964 269900
rect 336832 269952 336884 269958
rect 336832 269894 336884 269900
rect 335636 269476 335688 269482
rect 335636 269418 335688 269424
rect 335176 268388 335228 268394
rect 335176 268330 335228 268336
rect 334624 266688 334676 266694
rect 334624 266630 334676 266636
rect 335188 264316 335216 268330
rect 335648 266898 335676 269418
rect 335636 266892 335688 266898
rect 335636 266834 335688 266840
rect 336004 266892 336056 266898
rect 336004 266834 336056 266840
rect 336016 264316 336044 266834
rect 336844 264316 336872 269894
rect 338040 264330 338068 272478
rect 338960 264330 338988 275130
rect 339316 270156 339368 270162
rect 339316 270098 339368 270104
rect 337686 264302 338068 264330
rect 338514 264302 338988 264330
rect 339328 264316 339356 270098
rect 339512 269822 339540 277766
rect 341352 271454 341380 277780
rect 341524 275460 341576 275466
rect 341524 275402 341576 275408
rect 341340 271448 341392 271454
rect 341340 271390 341392 271396
rect 340604 271312 340656 271318
rect 340604 271254 340656 271260
rect 339500 269816 339552 269822
rect 339500 269758 339552 269764
rect 340616 264330 340644 271254
rect 341536 270162 341564 275402
rect 342456 272678 342484 277780
rect 343666 277766 343864 277794
rect 342904 274236 342956 274242
rect 342904 274178 342956 274184
rect 342444 272672 342496 272678
rect 342444 272614 342496 272620
rect 342168 271448 342220 271454
rect 342168 271390 342220 271396
rect 341524 270156 341576 270162
rect 341524 270098 341576 270104
rect 341800 270088 341852 270094
rect 341800 270030 341852 270036
rect 340972 266416 341024 266422
rect 340972 266358 341024 266364
rect 340170 264302 340644 264330
rect 340984 264316 341012 266358
rect 341812 264316 341840 270030
rect 342180 266422 342208 271390
rect 342916 267442 342944 274178
rect 343836 269482 343864 277766
rect 344480 277766 344862 277794
rect 345124 277766 346058 277794
rect 344480 271182 344508 277766
rect 344468 271176 344520 271182
rect 344468 271118 344520 271124
rect 344652 271176 344704 271182
rect 344652 271118 344704 271124
rect 343824 269476 343876 269482
rect 343824 269418 343876 269424
rect 342904 267436 342956 267442
rect 342904 267378 342956 267384
rect 343456 267300 343508 267306
rect 343456 267242 343508 267248
rect 342628 267164 342680 267170
rect 342628 267106 342680 267112
rect 342168 266416 342220 266422
rect 342168 266358 342220 266364
rect 342640 264316 342668 267106
rect 343468 264316 343496 267242
rect 344664 264330 344692 271118
rect 345124 268530 345152 277766
rect 347240 274242 347268 277780
rect 347792 277766 348450 277794
rect 347228 274236 347280 274242
rect 347228 274178 347280 274184
rect 346308 273964 346360 273970
rect 346308 273906 346360 273912
rect 345112 268524 345164 268530
rect 345112 268466 345164 268472
rect 345940 268524 345992 268530
rect 345940 268466 345992 268472
rect 345112 266416 345164 266422
rect 345112 266358 345164 266364
rect 344310 264302 344692 264330
rect 345124 264316 345152 266358
rect 345952 264316 345980 268466
rect 346320 266422 346348 273906
rect 347044 273284 347096 273290
rect 347044 273226 347096 273232
rect 347056 266898 347084 273226
rect 347596 269816 347648 269822
rect 347596 269758 347648 269764
rect 347044 266892 347096 266898
rect 347044 266834 347096 266840
rect 346768 266552 346820 266558
rect 346768 266494 346820 266500
rect 346308 266416 346360 266422
rect 346308 266358 346360 266364
rect 346780 264316 346808 266494
rect 347608 264316 347636 269758
rect 347792 268394 347820 277766
rect 349632 273290 349660 277780
rect 350552 277766 350750 277794
rect 349620 273284 349672 273290
rect 349620 273226 349672 273232
rect 350264 273284 350316 273290
rect 350264 273226 350316 273232
rect 348424 270224 348476 270230
rect 348424 270166 348476 270172
rect 347780 268388 347832 268394
rect 347780 268330 347832 268336
rect 348436 264316 348464 270166
rect 350080 268388 350132 268394
rect 350080 268330 350132 268336
rect 349252 266416 349304 266422
rect 349252 266358 349304 266364
rect 349264 264316 349292 266358
rect 350092 264316 350120 268330
rect 350276 266422 350304 273226
rect 350552 269958 350580 277766
rect 350724 275596 350776 275602
rect 350724 275538 350776 275544
rect 350736 271182 350764 275538
rect 351932 272542 351960 277780
rect 353128 275330 353156 277780
rect 354324 275466 354352 277780
rect 354312 275460 354364 275466
rect 354312 275402 354364 275408
rect 353116 275324 353168 275330
rect 353116 275266 353168 275272
rect 353944 275324 353996 275330
rect 353944 275266 353996 275272
rect 352932 272808 352984 272814
rect 352932 272750 352984 272756
rect 351920 272536 351972 272542
rect 351920 272478 351972 272484
rect 350724 271176 350776 271182
rect 350724 271118 350776 271124
rect 351828 271176 351880 271182
rect 351828 271118 351880 271124
rect 350540 269952 350592 269958
rect 350540 269894 350592 269900
rect 351644 269680 351696 269686
rect 351644 269622 351696 269628
rect 350908 267436 350960 267442
rect 350908 267378 350960 267384
rect 350264 266416 350316 266422
rect 350264 266358 350316 266364
rect 350920 264316 350948 267378
rect 351656 266558 351684 269622
rect 351644 266552 351696 266558
rect 351644 266494 351696 266500
rect 351840 265690 351868 271118
rect 351748 265662 351868 265690
rect 351748 264316 351776 265662
rect 352944 264330 352972 272750
rect 353956 267306 353984 275266
rect 355324 271720 355376 271726
rect 355324 271662 355376 271668
rect 354220 269952 354272 269958
rect 354220 269894 354272 269900
rect 353944 267300 353996 267306
rect 353944 267242 353996 267248
rect 353392 267028 353444 267034
rect 353392 266970 353444 266976
rect 352590 264302 352972 264330
rect 353404 264316 353432 266970
rect 354232 264316 354260 269894
rect 355336 267034 355364 271662
rect 355520 271318 355548 277780
rect 356336 275324 356388 275330
rect 356336 275266 356388 275272
rect 356348 273290 356376 275266
rect 356336 273284 356388 273290
rect 356336 273226 356388 273232
rect 356520 271856 356572 271862
rect 356520 271798 356572 271804
rect 355508 271312 355560 271318
rect 355508 271254 355560 271260
rect 356532 267170 356560 271798
rect 356716 271454 356744 277780
rect 357452 277766 357926 277794
rect 356704 271448 356756 271454
rect 356704 271390 356756 271396
rect 356704 270360 356756 270366
rect 356704 270302 356756 270308
rect 356520 267164 356572 267170
rect 356520 267106 356572 267112
rect 355324 267028 355376 267034
rect 355324 266970 355376 266976
rect 355876 267028 355928 267034
rect 355876 266970 355928 266976
rect 355048 266552 355100 266558
rect 355048 266494 355100 266500
rect 355060 264316 355088 266494
rect 355888 264316 355916 266970
rect 356716 264316 356744 270302
rect 357452 270094 357480 277766
rect 358636 272536 358688 272542
rect 358636 272478 358688 272484
rect 357440 270088 357492 270094
rect 357440 270030 357492 270036
rect 358360 266756 358412 266762
rect 358360 266698 358412 266704
rect 357532 266416 357584 266422
rect 357532 266358 357584 266364
rect 357544 264316 357572 266358
rect 358372 264316 358400 266698
rect 358648 266422 358676 272478
rect 359016 271862 359044 277780
rect 360212 275466 360240 277780
rect 361408 275602 361436 277780
rect 361396 275596 361448 275602
rect 361396 275538 361448 275544
rect 362224 275596 362276 275602
rect 362224 275538 362276 275544
rect 360200 275460 360252 275466
rect 360200 275402 360252 275408
rect 360292 274712 360344 274718
rect 360292 274654 360344 274660
rect 360108 274100 360160 274106
rect 360108 274042 360160 274048
rect 359004 271856 359056 271862
rect 359004 271798 359056 271804
rect 359004 270496 359056 270502
rect 359004 270438 359056 270444
rect 359016 266558 359044 270438
rect 360120 267734 360148 274042
rect 360304 268530 360332 274654
rect 360844 271448 360896 271454
rect 360844 271390 360896 271396
rect 360292 268524 360344 268530
rect 360292 268466 360344 268472
rect 360028 267706 360148 267734
rect 359188 267300 359240 267306
rect 359188 267242 359240 267248
rect 359004 266552 359056 266558
rect 359004 266494 359056 266500
rect 358636 266416 358688 266422
rect 358636 266358 358688 266364
rect 359200 264316 359228 267242
rect 360028 264316 360056 267706
rect 360856 266762 360884 271390
rect 361028 268524 361080 268530
rect 361028 268466 361080 268472
rect 361040 267442 361068 268466
rect 361028 267436 361080 267442
rect 361028 267378 361080 267384
rect 360844 266756 360896 266762
rect 360844 266698 360896 266704
rect 362236 266626 362264 275538
rect 362604 273970 362632 277780
rect 363052 275460 363104 275466
rect 363052 275402 363104 275408
rect 362868 274372 362920 274378
rect 362868 274314 362920 274320
rect 362592 273964 362644 273970
rect 362592 273906 362644 273912
rect 362880 267734 362908 274314
rect 363064 270230 363092 275402
rect 363800 274718 363828 277780
rect 364352 277766 365010 277794
rect 365732 277766 366114 277794
rect 363788 274712 363840 274718
rect 363788 274654 363840 274660
rect 364156 271312 364208 271318
rect 364156 271254 364208 271260
rect 363052 270224 363104 270230
rect 363052 270166 363104 270172
rect 363052 268660 363104 268666
rect 363052 268602 363104 268608
rect 363064 267734 363092 268602
rect 362788 267706 362908 267734
rect 362972 267706 363092 267734
rect 360844 266620 360896 266626
rect 360844 266562 360896 266568
rect 362224 266620 362276 266626
rect 362224 266562 362276 266568
rect 360856 264316 360884 266562
rect 362788 266490 362816 267706
rect 361672 266484 361724 266490
rect 361672 266426 361724 266432
rect 362776 266484 362828 266490
rect 362776 266426 362828 266432
rect 361684 264316 361712 266426
rect 362972 266370 363000 267706
rect 363328 267164 363380 267170
rect 363328 267106 363380 267112
rect 362880 266342 363000 266370
rect 362880 264330 362908 266342
rect 362526 264302 362908 264330
rect 363340 264316 363368 267106
rect 364168 264316 364196 271254
rect 364352 269686 364380 277766
rect 364984 270224 365036 270230
rect 364984 270166 365036 270172
rect 364340 269680 364392 269686
rect 364340 269622 364392 269628
rect 364996 264316 365024 270166
rect 365732 269822 365760 277766
rect 367296 275466 367324 277780
rect 367284 275460 367336 275466
rect 367284 275402 367336 275408
rect 368492 275330 368520 277780
rect 369124 275460 369176 275466
rect 369124 275402 369176 275408
rect 368480 275324 368532 275330
rect 368480 275266 368532 275272
rect 367100 274712 367152 274718
rect 367100 274654 367152 274660
rect 366916 274236 366968 274242
rect 366916 274178 366968 274184
rect 365720 269816 365772 269822
rect 365720 269758 365772 269764
rect 365812 267436 365864 267442
rect 365812 267378 365864 267384
rect 365824 264316 365852 267378
rect 366928 264330 366956 274178
rect 367112 268394 367140 274654
rect 368388 272672 368440 272678
rect 368388 272614 368440 272620
rect 367100 268388 367152 268394
rect 367100 268330 367152 268336
rect 368204 267708 368256 267714
rect 368204 267650 368256 267656
rect 367468 266416 367520 266422
rect 367468 266358 367520 266364
rect 366666 264302 366956 264330
rect 367480 264316 367508 266358
rect 368216 264330 368244 267650
rect 368400 266422 368428 272614
rect 369136 267034 369164 275402
rect 369688 274718 369716 277780
rect 369872 277766 370898 277794
rect 369676 274712 369728 274718
rect 369676 274654 369728 274660
rect 369400 270088 369452 270094
rect 369400 270030 369452 270036
rect 369124 267028 369176 267034
rect 369124 266970 369176 266976
rect 368388 266416 368440 266422
rect 368388 266358 368440 266364
rect 369412 264330 369440 270030
rect 369872 268530 369900 277766
rect 370504 275732 370556 275738
rect 370504 275674 370556 275680
rect 369860 268524 369912 268530
rect 369860 268466 369912 268472
rect 370320 268524 370372 268530
rect 370320 268466 370372 268472
rect 370332 264330 370360 268466
rect 370516 267170 370544 275674
rect 372080 271182 372108 277780
rect 373000 277766 373290 277794
rect 373000 272814 373028 277766
rect 373264 272944 373316 272950
rect 373264 272886 373316 272892
rect 372988 272808 373040 272814
rect 372988 272750 373040 272756
rect 372528 271584 372580 271590
rect 372528 271526 372580 271532
rect 372068 271176 372120 271182
rect 372068 271118 372120 271124
rect 372344 269816 372396 269822
rect 372344 269758 372396 269764
rect 370780 267572 370832 267578
rect 370780 267514 370832 267520
rect 370504 267164 370556 267170
rect 370504 267106 370556 267112
rect 368216 264302 368322 264330
rect 369150 264302 369440 264330
rect 369978 264302 370360 264330
rect 370792 264316 370820 267514
rect 371608 266416 371660 266422
rect 371608 266358 371660 266364
rect 371620 264316 371648 266358
rect 372356 264330 372384 269758
rect 372540 266422 372568 271526
rect 373276 267306 373304 272886
rect 374380 271726 374408 277780
rect 375392 277766 375590 277794
rect 375104 275324 375156 275330
rect 375104 275266 375156 275272
rect 374368 271720 374420 271726
rect 374368 271662 374420 271668
rect 374920 268388 374972 268394
rect 374920 268330 374972 268336
rect 373264 267300 373316 267306
rect 373264 267242 373316 267248
rect 373264 267164 373316 267170
rect 373264 267106 373316 267112
rect 372528 266416 372580 266422
rect 372528 266358 372580 266364
rect 372356 264302 372462 264330
rect 373276 264316 373304 267106
rect 374092 266416 374144 266422
rect 374092 266358 374144 266364
rect 374104 264316 374132 266358
rect 374932 264316 374960 268330
rect 375116 266422 375144 275266
rect 375392 269958 375420 277766
rect 376772 270502 376800 277780
rect 377968 275466 377996 277780
rect 378152 277766 379178 277794
rect 377956 275460 378008 275466
rect 377956 275402 378008 275408
rect 377772 273964 377824 273970
rect 377772 273906 377824 273912
rect 376760 270496 376812 270502
rect 376760 270438 376812 270444
rect 377588 270496 377640 270502
rect 377588 270438 377640 270444
rect 375380 269952 375432 269958
rect 375380 269894 375432 269900
rect 376576 269952 376628 269958
rect 376576 269894 376628 269900
rect 375748 267300 375800 267306
rect 375748 267242 375800 267248
rect 375104 266416 375156 266422
rect 375104 266358 375156 266364
rect 375760 264316 375788 267242
rect 376588 264316 376616 269894
rect 377600 267714 377628 270438
rect 377588 267708 377640 267714
rect 377588 267650 377640 267656
rect 377784 264330 377812 273906
rect 378152 270366 378180 277766
rect 380360 272542 380388 277780
rect 380716 272808 380768 272814
rect 380716 272750 380768 272756
rect 380348 272536 380400 272542
rect 380348 272478 380400 272484
rect 380532 272536 380584 272542
rect 380532 272478 380584 272484
rect 379428 271176 379480 271182
rect 379428 271118 379480 271124
rect 378140 270360 378192 270366
rect 378140 270302 378192 270308
rect 378232 267028 378284 267034
rect 378232 266970 378284 266976
rect 377430 264302 377812 264330
rect 378244 264316 378272 266970
rect 379440 264330 379468 271118
rect 379888 266416 379940 266422
rect 379888 266358 379940 266364
rect 379086 264302 379468 264330
rect 379900 264316 379928 266358
rect 380544 264330 380572 272478
rect 380728 266422 380756 272750
rect 381556 271454 381584 277780
rect 382004 275460 382056 275466
rect 382004 275402 382056 275408
rect 381544 271448 381596 271454
rect 381544 271390 381596 271396
rect 381544 271040 381596 271046
rect 381544 270982 381596 270988
rect 381556 267578 381584 270982
rect 381544 267572 381596 267578
rect 381544 267514 381596 267520
rect 380716 266416 380768 266422
rect 380716 266358 380768 266364
rect 382016 264330 382044 275402
rect 382660 272950 382688 277780
rect 383856 274106 383884 277780
rect 385052 275602 385080 277780
rect 385040 275596 385092 275602
rect 385040 275538 385092 275544
rect 386052 274712 386104 274718
rect 386052 274654 386104 274660
rect 383844 274100 383896 274106
rect 383844 274042 383896 274048
rect 384948 274100 385000 274106
rect 384948 274042 385000 274048
rect 382924 273080 382976 273086
rect 382924 273022 382976 273028
rect 382648 272944 382700 272950
rect 382648 272886 382700 272892
rect 382372 268932 382424 268938
rect 382372 268874 382424 268880
rect 380544 264302 380742 264330
rect 381570 264302 382044 264330
rect 382384 264316 382412 268874
rect 382936 267442 382964 273022
rect 384028 269680 384080 269686
rect 384028 269622 384080 269628
rect 383200 267708 383252 267714
rect 383200 267650 383252 267656
rect 382924 267436 382976 267442
rect 382924 267378 382976 267384
rect 383212 264316 383240 267650
rect 384040 264316 384068 269622
rect 384960 267734 384988 274042
rect 386064 271318 386092 274654
rect 386248 274378 386276 277780
rect 386432 277766 387458 277794
rect 386236 274372 386288 274378
rect 386236 274314 386288 274320
rect 386052 271312 386104 271318
rect 386052 271254 386104 271260
rect 385684 270360 385736 270366
rect 385684 270302 385736 270308
rect 384868 267706 384988 267734
rect 384868 264316 384896 267706
rect 385696 264316 385724 270302
rect 386432 268666 386460 277766
rect 388640 275738 388668 277780
rect 389180 276004 389232 276010
rect 389180 275946 389232 275952
rect 388628 275732 388680 275738
rect 388628 275674 388680 275680
rect 388168 275596 388220 275602
rect 388168 275538 388220 275544
rect 387708 271720 387760 271726
rect 387708 271662 387760 271668
rect 387340 268796 387392 268802
rect 387340 268738 387392 268744
rect 386420 268660 386472 268666
rect 386420 268602 386472 268608
rect 386512 266416 386564 266422
rect 386512 266358 386564 266364
rect 386524 264316 386552 266358
rect 387352 264316 387380 268738
rect 387720 266422 387748 271662
rect 388180 269686 388208 275538
rect 389192 274242 389220 275946
rect 389744 274718 389772 277780
rect 390572 277766 390954 277794
rect 389732 274712 389784 274718
rect 389732 274654 389784 274660
rect 389180 274236 389232 274242
rect 389180 274178 389232 274184
rect 390284 274236 390336 274242
rect 390284 274178 390336 274184
rect 388628 272944 388680 272950
rect 388628 272886 388680 272892
rect 388640 272678 388668 272886
rect 388628 272672 388680 272678
rect 388628 272614 388680 272620
rect 389088 270904 389140 270910
rect 389088 270846 389140 270852
rect 388168 269680 388220 269686
rect 388168 269622 388220 269628
rect 389100 267734 389128 270846
rect 389008 267706 389128 267734
rect 388168 266756 388220 266762
rect 388168 266698 388220 266704
rect 387708 266416 387760 266422
rect 387708 266358 387760 266364
rect 388180 264316 388208 266698
rect 389008 264316 389036 267706
rect 390296 264330 390324 274178
rect 390572 270230 390600 277766
rect 392136 273086 392164 277780
rect 393332 276010 393360 277780
rect 393320 276004 393372 276010
rect 393320 275946 393372 275952
rect 393596 275868 393648 275874
rect 393596 275810 393648 275816
rect 392584 274508 392636 274514
rect 392584 274450 392636 274456
rect 392124 273080 392176 273086
rect 392124 273022 392176 273028
rect 391848 272944 391900 272950
rect 391848 272886 391900 272892
rect 390560 270224 390612 270230
rect 390560 270166 390612 270172
rect 390652 267572 390704 267578
rect 390652 267514 390704 267520
rect 389850 264302 390324 264330
rect 390664 264316 390692 267514
rect 391860 264330 391888 272886
rect 392308 270224 392360 270230
rect 392308 270166 392360 270172
rect 391506 264302 391888 264330
rect 392320 264316 392348 270166
rect 392596 267170 392624 274450
rect 393608 272678 393636 275810
rect 394528 272814 394556 277780
rect 394712 277766 395738 277794
rect 396092 277766 396934 277794
rect 397472 277766 398038 277794
rect 394516 272808 394568 272814
rect 394516 272750 394568 272756
rect 393596 272672 393648 272678
rect 393596 272614 393648 272620
rect 393964 272672 394016 272678
rect 393964 272614 394016 272620
rect 393976 267306 394004 272614
rect 394332 271856 394384 271862
rect 394332 271798 394384 271804
rect 393964 267300 394016 267306
rect 393964 267242 394016 267248
rect 392584 267164 392636 267170
rect 392584 267106 392636 267112
rect 393136 266892 393188 266898
rect 393136 266834 393188 266840
rect 393148 264316 393176 266834
rect 394344 264330 394372 271798
rect 394712 270502 394740 277766
rect 395896 274372 395948 274378
rect 395896 274314 395948 274320
rect 394700 270496 394752 270502
rect 394700 270438 394752 270444
rect 394700 269544 394752 269550
rect 394700 269486 394752 269492
rect 394712 267714 394740 269486
rect 394700 267708 394752 267714
rect 394700 267650 394752 267656
rect 394792 266552 394844 266558
rect 394792 266494 394844 266500
rect 393990 264302 394372 264330
rect 394804 264316 394832 266494
rect 395908 264330 395936 274314
rect 396092 270094 396120 277766
rect 397276 272808 397328 272814
rect 397276 272750 397328 272756
rect 396264 270496 396316 270502
rect 396264 270438 396316 270444
rect 396080 270088 396132 270094
rect 396080 270030 396132 270036
rect 396276 266762 396304 270438
rect 397092 267436 397144 267442
rect 397092 267378 397144 267384
rect 396264 266756 396316 266762
rect 396264 266698 396316 266704
rect 396448 266416 396500 266422
rect 396448 266358 396500 266364
rect 395646 264302 395936 264330
rect 396460 264316 396488 266358
rect 397104 264330 397132 267378
rect 397288 266422 397316 272750
rect 397472 268530 397500 277766
rect 398104 271448 398156 271454
rect 398104 271390 398156 271396
rect 397460 268524 397512 268530
rect 397460 268466 397512 268472
rect 398116 266558 398144 271390
rect 399220 271046 399248 277780
rect 400416 271590 400444 277780
rect 401626 277766 401824 277794
rect 400588 276004 400640 276010
rect 400588 275946 400640 275952
rect 400404 271584 400456 271590
rect 400404 271526 400456 271532
rect 400128 271312 400180 271318
rect 400128 271254 400180 271260
rect 399208 271040 399260 271046
rect 399208 270982 399260 270988
rect 398472 267708 398524 267714
rect 398472 267650 398524 267656
rect 398104 266552 398156 266558
rect 398104 266494 398156 266500
rect 397276 266416 397328 266422
rect 397276 266358 397328 266364
rect 398484 264330 398512 267650
rect 399760 267300 399812 267306
rect 399760 267242 399812 267248
rect 398932 266416 398984 266422
rect 398932 266358 398984 266364
rect 397104 264302 397302 264330
rect 398130 264302 398512 264330
rect 398944 264316 398972 266358
rect 399772 264316 399800 267242
rect 400140 266422 400168 271254
rect 400600 268938 400628 275946
rect 401324 271040 401376 271046
rect 401324 270982 401376 270988
rect 400588 268932 400640 268938
rect 400588 268874 400640 268880
rect 400588 268524 400640 268530
rect 400588 268466 400640 268472
rect 400128 266416 400180 266422
rect 400128 266358 400180 266364
rect 400600 264316 400628 268466
rect 401336 264330 401364 270982
rect 401796 269822 401824 277766
rect 402808 274514 402836 277780
rect 404004 275330 404032 277780
rect 404556 277766 405214 277794
rect 403992 275324 404044 275330
rect 403992 275266 404044 275272
rect 403992 274848 404044 274854
rect 403992 274790 404044 274796
rect 402796 274508 402848 274514
rect 402796 274450 402848 274456
rect 403072 270088 403124 270094
rect 403072 270030 403124 270036
rect 401784 269816 401836 269822
rect 401784 269758 401836 269764
rect 401600 269408 401652 269414
rect 401600 269350 401652 269356
rect 401612 266898 401640 269350
rect 402244 268660 402296 268666
rect 402244 268602 402296 268608
rect 401600 266892 401652 266898
rect 401600 266834 401652 266840
rect 401336 264302 401442 264330
rect 402256 264316 402284 268602
rect 403084 264316 403112 270030
rect 404004 269958 404032 274790
rect 404176 273080 404228 273086
rect 404176 273022 404228 273028
rect 403992 269952 404044 269958
rect 403992 269894 404044 269900
rect 404188 264330 404216 273022
rect 404360 269680 404412 269686
rect 404360 269622 404412 269628
rect 404372 267578 404400 269622
rect 404556 268394 404584 277766
rect 406304 272678 406332 277780
rect 407500 274854 407528 277780
rect 407488 274848 407540 274854
rect 407488 274790 407540 274796
rect 407120 274712 407172 274718
rect 407120 274654 407172 274660
rect 406844 274508 406896 274514
rect 406844 274450 406896 274456
rect 406292 272672 406344 272678
rect 406292 272614 406344 272620
rect 404544 268388 404596 268394
rect 404544 268330 404596 268336
rect 404360 267572 404412 267578
rect 404360 267514 404412 267520
rect 404728 267164 404780 267170
rect 404728 267106 404780 267112
rect 403926 264302 404216 264330
rect 404740 264316 404768 267106
rect 405556 266892 405608 266898
rect 405556 266834 405608 266840
rect 405568 264316 405596 266834
rect 406856 264330 406884 274450
rect 407132 271182 407160 274654
rect 408696 273970 408724 277780
rect 408684 273964 408736 273970
rect 408684 273906 408736 273912
rect 409892 273290 409920 277780
rect 410064 275732 410116 275738
rect 410064 275674 410116 275680
rect 409144 273284 409196 273290
rect 409144 273226 409196 273232
rect 409880 273284 409932 273290
rect 409880 273226 409932 273232
rect 408408 272672 408460 272678
rect 408408 272614 408460 272620
rect 407120 271176 407172 271182
rect 407120 271118 407172 271124
rect 407212 268388 407264 268394
rect 407212 268330 407264 268336
rect 406410 264302 406884 264330
rect 407224 264316 407252 268330
rect 408420 264330 408448 272614
rect 409156 267034 409184 273226
rect 410076 272950 410104 275674
rect 411088 274718 411116 277780
rect 412284 275874 412312 277780
rect 412272 275868 412324 275874
rect 412272 275810 412324 275816
rect 411260 275324 411312 275330
rect 411260 275266 411312 275272
rect 411076 274712 411128 274718
rect 411076 274654 411128 274660
rect 410064 272944 410116 272950
rect 410064 272886 410116 272892
rect 411272 271946 411300 275266
rect 412456 272944 412508 272950
rect 412456 272886 412508 272892
rect 410904 271918 411300 271946
rect 409788 271584 409840 271590
rect 409788 271526 409840 271532
rect 409604 267572 409656 267578
rect 409604 267514 409656 267520
rect 409144 267028 409196 267034
rect 409144 266970 409196 266976
rect 408868 266416 408920 266422
rect 408868 266358 408920 266364
rect 408066 264302 408448 264330
rect 408880 264316 408908 266358
rect 409616 264330 409644 267514
rect 409800 266422 409828 271526
rect 409788 266416 409840 266422
rect 409788 266358 409840 266364
rect 410904 264330 410932 271918
rect 412180 266756 412232 266762
rect 412180 266698 412232 266704
rect 411352 266416 411404 266422
rect 411352 266358 411404 266364
rect 409616 264302 409722 264330
rect 410550 264302 410932 264330
rect 411364 264316 411392 266358
rect 412192 264316 412220 266698
rect 412468 266422 412496 272886
rect 413388 272542 413416 277780
rect 414584 275466 414612 277780
rect 415780 276010 415808 277780
rect 416792 277766 416990 277794
rect 415768 276004 415820 276010
rect 415768 275946 415820 275952
rect 415308 275868 415360 275874
rect 415308 275810 415360 275816
rect 414572 275460 414624 275466
rect 414572 275402 414624 275408
rect 413928 273964 413980 273970
rect 413928 273906 413980 273912
rect 413376 272536 413428 272542
rect 413376 272478 413428 272484
rect 413008 269952 413060 269958
rect 413008 269894 413060 269900
rect 412456 266416 412508 266422
rect 412456 266358 412508 266364
rect 413020 264316 413048 269894
rect 413940 267734 413968 273906
rect 415124 272536 415176 272542
rect 415124 272478 415176 272484
rect 413848 267706 413968 267734
rect 413848 264316 413876 267706
rect 415136 264330 415164 272478
rect 415320 270910 415348 275810
rect 416412 275460 416464 275466
rect 416412 275402 416464 275408
rect 415308 270904 415360 270910
rect 415308 270846 415360 270852
rect 416424 266422 416452 275402
rect 416596 271176 416648 271182
rect 416596 271118 416648 271124
rect 415492 266416 415544 266422
rect 415492 266358 415544 266364
rect 416412 266416 416464 266422
rect 416412 266358 416464 266364
rect 414690 264302 415164 264330
rect 415504 264316 415532 266358
rect 416608 264330 416636 271118
rect 416792 269550 416820 277766
rect 418172 275602 418200 277780
rect 418160 275596 418212 275602
rect 418160 275538 418212 275544
rect 418344 275596 418396 275602
rect 418344 275538 418396 275544
rect 418356 272814 418384 275538
rect 419368 274106 419396 277780
rect 419552 277766 420578 277794
rect 421392 277766 421682 277794
rect 422312 277766 422878 277794
rect 423692 277766 424074 277794
rect 419356 274100 419408 274106
rect 419356 274042 419408 274048
rect 419172 273216 419224 273222
rect 419172 273158 419224 273164
rect 418344 272808 418396 272814
rect 418344 272750 418396 272756
rect 416780 269544 416832 269550
rect 416780 269486 416832 269492
rect 417148 269272 417200 269278
rect 417148 269214 417200 269220
rect 416346 264302 416636 264330
rect 417160 264316 417188 269214
rect 418988 268932 419040 268938
rect 418988 268874 419040 268880
rect 419000 267306 419028 268874
rect 418988 267300 419040 267306
rect 418988 267242 419040 267248
rect 417976 266756 418028 266762
rect 417976 266698 418028 266704
rect 417988 264316 418016 266698
rect 419184 264330 419212 273158
rect 419552 270366 419580 277766
rect 420920 275188 420972 275194
rect 420920 275130 420972 275136
rect 420932 274378 420960 275130
rect 420920 274372 420972 274378
rect 420920 274314 420972 274320
rect 421392 271726 421420 277766
rect 421564 274100 421616 274106
rect 421564 274042 421616 274048
rect 421380 271720 421432 271726
rect 421380 271662 421432 271668
rect 419540 270360 419592 270366
rect 419540 270302 419592 270308
rect 419632 269544 419684 269550
rect 419632 269486 419684 269492
rect 418830 264302 419212 264330
rect 419644 264316 419672 269486
rect 420460 268116 420512 268122
rect 420460 268058 420512 268064
rect 420472 264316 420500 268058
rect 421288 267300 421340 267306
rect 421288 267242 421340 267248
rect 421300 264316 421328 267242
rect 421576 266626 421604 274042
rect 421748 271720 421800 271726
rect 421748 271662 421800 271668
rect 421760 267714 421788 271662
rect 422312 269074 422340 277766
rect 423692 270502 423720 277766
rect 425256 275874 425284 277780
rect 425244 275868 425296 275874
rect 425244 275810 425296 275816
rect 426256 274848 426308 274854
rect 426256 274790 426308 274796
rect 424968 274644 425020 274650
rect 424968 274586 425020 274592
rect 423680 270496 423732 270502
rect 423680 270438 423732 270444
rect 424600 270496 424652 270502
rect 424600 270438 424652 270444
rect 422300 269068 422352 269074
rect 422300 269010 422352 269016
rect 422300 268796 422352 268802
rect 422300 268738 422352 268744
rect 421748 267708 421800 267714
rect 421748 267650 421800 267656
rect 422312 267442 422340 268738
rect 422300 267436 422352 267442
rect 422300 267378 422352 267384
rect 422116 267028 422168 267034
rect 422116 266970 422168 266976
rect 421564 266620 421616 266626
rect 421564 266562 421616 266568
rect 422128 264316 422156 266970
rect 422944 266620 422996 266626
rect 422944 266562 422996 266568
rect 422956 264316 422984 266562
rect 423772 266416 423824 266422
rect 423772 266358 423824 266364
rect 423784 264316 423812 266358
rect 424612 264316 424640 270438
rect 424980 266422 425008 274586
rect 426072 272808 426124 272814
rect 426072 272750 426124 272756
rect 425704 271040 425756 271046
rect 425704 270982 425756 270988
rect 425716 266898 425744 270982
rect 425704 266892 425756 266898
rect 425704 266834 425756 266840
rect 424968 266416 425020 266422
rect 424968 266358 425020 266364
rect 425428 266416 425480 266422
rect 425428 266358 425480 266364
rect 425440 264316 425468 266358
rect 426084 264330 426112 272750
rect 426268 271862 426296 274790
rect 426452 274242 426480 277780
rect 426636 277766 427662 277794
rect 426440 274236 426492 274242
rect 426440 274178 426492 274184
rect 426256 271856 426308 271862
rect 426256 271798 426308 271804
rect 426636 269686 426664 277766
rect 427820 276004 427872 276010
rect 427820 275946 427872 275952
rect 426900 273828 426952 273834
rect 426900 273770 426952 273776
rect 426624 269680 426676 269686
rect 426624 269622 426676 269628
rect 426912 266422 426940 273770
rect 427084 271856 427136 271862
rect 427084 271798 427136 271804
rect 427096 271454 427124 271798
rect 427084 271448 427136 271454
rect 427084 271390 427136 271396
rect 427268 271448 427320 271454
rect 427268 271390 427320 271396
rect 427280 271046 427308 271390
rect 427268 271040 427320 271046
rect 427268 270982 427320 270988
rect 427832 270910 427860 275946
rect 428844 275738 428872 277780
rect 429396 277766 429962 277794
rect 430592 277766 431158 277794
rect 428832 275732 428884 275738
rect 428832 275674 428884 275680
rect 429200 275732 429252 275738
rect 429200 275674 429252 275680
rect 429016 273556 429068 273562
rect 429016 273498 429068 273504
rect 427820 270904 427872 270910
rect 427820 270846 427872 270852
rect 428464 270632 428516 270638
rect 428464 270574 428516 270580
rect 427360 269680 427412 269686
rect 427360 269622 427412 269628
rect 426900 266416 426952 266422
rect 426900 266358 426952 266364
rect 427372 264330 427400 269622
rect 428476 266762 428504 270574
rect 428464 266756 428516 266762
rect 428464 266698 428516 266704
rect 427912 266484 427964 266490
rect 427912 266426 427964 266432
rect 426084 264302 426282 264330
rect 427110 264302 427400 264330
rect 427924 264316 427952 266426
rect 429028 264330 429056 273498
rect 429212 273086 429240 275674
rect 429200 273080 429252 273086
rect 429200 273022 429252 273028
rect 429396 270230 429424 277766
rect 429568 270360 429620 270366
rect 429568 270302 429620 270308
rect 429384 270224 429436 270230
rect 429384 270166 429436 270172
rect 428766 264302 429056 264330
rect 429580 264316 429608 270302
rect 430592 269414 430620 277766
rect 432340 274854 432368 277780
rect 432972 275868 433024 275874
rect 432972 275810 433024 275816
rect 432328 274848 432380 274854
rect 432328 274790 432380 274796
rect 431684 271040 431736 271046
rect 431684 270982 431736 270988
rect 430580 269408 430632 269414
rect 430580 269350 430632 269356
rect 430396 266756 430448 266762
rect 430396 266698 430448 266704
rect 430408 264316 430436 266698
rect 431696 264330 431724 270982
rect 431960 267844 432012 267850
rect 431960 267786 432012 267792
rect 431972 267170 432000 267786
rect 432984 267734 433012 275810
rect 433536 271862 433564 277780
rect 434732 275194 434760 277780
rect 435928 275602 435956 277780
rect 436112 277766 437046 277794
rect 435916 275596 435968 275602
rect 435916 275538 435968 275544
rect 434720 275188 434772 275194
rect 434720 275130 434772 275136
rect 435640 274780 435692 274786
rect 435640 274722 435692 274728
rect 434628 273080 434680 273086
rect 434628 273022 434680 273028
rect 433524 271856 433576 271862
rect 433524 271798 433576 271804
rect 433156 270768 433208 270774
rect 433156 270710 433208 270716
rect 432892 267706 433012 267734
rect 431960 267164 432012 267170
rect 431960 267106 432012 267112
rect 432052 266756 432104 266762
rect 432052 266698 432104 266704
rect 432064 266422 432092 266698
rect 432052 266416 432104 266422
rect 432052 266358 432104 266364
rect 432328 266416 432380 266422
rect 432328 266358 432380 266364
rect 432340 264330 432368 266358
rect 431250 264302 431724 264330
rect 432078 264302 432368 264330
rect 432892 264316 432920 267706
rect 433168 266422 433196 270710
rect 434444 269136 434496 269142
rect 434444 269078 434496 269084
rect 433156 266416 433208 266422
rect 433156 266358 433208 266364
rect 433708 266416 433760 266422
rect 433708 266358 433760 266364
rect 433720 264316 433748 266358
rect 434456 264330 434484 269078
rect 434640 266422 434668 273022
rect 435652 271318 435680 274722
rect 435640 271312 435692 271318
rect 435640 271254 435692 271260
rect 435364 270904 435416 270910
rect 435364 270846 435416 270852
rect 435376 267578 435404 270846
rect 436112 268802 436140 277766
rect 437480 275188 437532 275194
rect 437480 275130 437532 275136
rect 437492 274514 437520 275130
rect 437480 274508 437532 274514
rect 437480 274450 437532 274456
rect 438228 271726 438256 277780
rect 439424 274786 439452 277780
rect 440252 277766 440634 277794
rect 441632 277766 441830 277794
rect 439412 274780 439464 274786
rect 439412 274722 439464 274728
rect 438768 274236 438820 274242
rect 438768 274178 438820 274184
rect 438216 271720 438268 271726
rect 438216 271662 438268 271668
rect 436928 271448 436980 271454
rect 436928 271390 436980 271396
rect 436940 270910 436968 271390
rect 436928 270904 436980 270910
rect 436928 270846 436980 270852
rect 436100 268796 436152 268802
rect 436100 268738 436152 268744
rect 436192 268252 436244 268258
rect 436192 268194 436244 268200
rect 435640 267708 435692 267714
rect 435640 267650 435692 267656
rect 435364 267572 435416 267578
rect 435364 267514 435416 267520
rect 434628 266416 434680 266422
rect 434628 266358 434680 266364
rect 435652 264330 435680 267650
rect 434456 264302 434562 264330
rect 435390 264302 435680 264330
rect 436204 264316 436232 268194
rect 437848 267980 437900 267986
rect 437848 267922 437900 267928
rect 437020 266416 437072 266422
rect 437020 266358 437072 266364
rect 437032 264316 437060 266358
rect 437860 264316 437888 267922
rect 438780 267734 438808 274178
rect 439320 272400 439372 272406
rect 439320 272342 439372 272348
rect 438688 267706 438808 267734
rect 438688 264316 438716 267706
rect 439332 266626 439360 272342
rect 440252 268938 440280 277766
rect 440884 274508 440936 274514
rect 440884 274450 440936 274456
rect 440240 268932 440292 268938
rect 440240 268874 440292 268880
rect 440332 267436 440384 267442
rect 440332 267378 440384 267384
rect 439320 266620 439372 266626
rect 439320 266562 439372 266568
rect 439504 266620 439556 266626
rect 439504 266562 439556 266568
rect 439516 264316 439544 266562
rect 440344 264316 440372 267378
rect 440896 266422 440924 274450
rect 441160 268796 441212 268802
rect 441160 268738 441212 268744
rect 440884 266416 440936 266422
rect 440884 266358 440936 266364
rect 441172 264316 441200 268738
rect 441632 268530 441660 277766
rect 443012 276010 443040 277780
rect 443288 277766 444222 277794
rect 444392 277766 445326 277794
rect 443000 276004 443052 276010
rect 443000 275946 443052 275952
rect 442908 271720 442960 271726
rect 442908 271662 442960 271668
rect 441620 268524 441672 268530
rect 441620 268466 441672 268472
rect 442724 268524 442776 268530
rect 442724 268466 442776 268472
rect 441988 266416 442040 266422
rect 441988 266358 442040 266364
rect 442000 264316 442028 266358
rect 442736 264330 442764 268466
rect 442920 266422 442948 271662
rect 443288 268666 443316 277766
rect 443736 276004 443788 276010
rect 443736 275946 443788 275952
rect 443748 271590 443776 275946
rect 443736 271584 443788 271590
rect 443736 271526 443788 271532
rect 444392 270094 444420 277766
rect 446508 275738 446536 277780
rect 447152 277766 447718 277794
rect 446496 275732 446548 275738
rect 446496 275674 446548 275680
rect 446772 275732 446824 275738
rect 446772 275674 446824 275680
rect 445024 270904 445076 270910
rect 445024 270846 445076 270852
rect 444380 270088 444432 270094
rect 444380 270030 444432 270036
rect 443644 268932 443696 268938
rect 443644 268874 443696 268880
rect 443276 268660 443328 268666
rect 443276 268602 443328 268608
rect 442908 266416 442960 266422
rect 442908 266358 442960 266364
rect 442736 264302 442842 264330
rect 443656 264316 443684 268874
rect 444472 266552 444524 266558
rect 444472 266494 444524 266500
rect 444484 264316 444512 266494
rect 445036 266422 445064 270846
rect 446128 268660 446180 268666
rect 446128 268602 446180 268608
rect 445300 267572 445352 267578
rect 445300 267514 445352 267520
rect 445024 266416 445076 266422
rect 445024 266358 445076 266364
rect 445312 264316 445340 267514
rect 446140 264316 446168 268602
rect 446784 268530 446812 275674
rect 446956 270224 447008 270230
rect 446956 270166 447008 270172
rect 446772 268524 446824 268530
rect 446772 268466 446824 268472
rect 446404 267028 446456 267034
rect 446404 266970 446456 266976
rect 446416 266762 446444 266970
rect 446404 266756 446456 266762
rect 446404 266698 446456 266704
rect 446968 264316 446996 270166
rect 447152 267850 447180 277766
rect 447784 271856 447836 271862
rect 447784 271798 447836 271804
rect 447140 267844 447192 267850
rect 447140 267786 447192 267792
rect 447796 266558 447824 271798
rect 448900 271318 448928 277780
rect 449164 275596 449216 275602
rect 449164 275538 449216 275544
rect 448888 271312 448940 271318
rect 448888 271254 448940 271260
rect 448612 268524 448664 268530
rect 448612 268466 448664 268472
rect 447784 266552 447836 266558
rect 447784 266494 447836 266500
rect 447784 266416 447836 266422
rect 447784 266358 447836 266364
rect 447796 264316 447824 266358
rect 448624 264316 448652 268466
rect 449176 266422 449204 275538
rect 450096 275194 450124 277780
rect 451306 277766 451504 277794
rect 450084 275188 450136 275194
rect 450084 275130 450136 275136
rect 449900 275052 449952 275058
rect 449900 274994 449952 275000
rect 449912 273970 449940 274994
rect 449900 273964 449952 273970
rect 449900 273906 449952 273912
rect 451096 273964 451148 273970
rect 451096 273906 451148 273912
rect 449900 269408 449952 269414
rect 449900 269350 449952 269356
rect 449912 267170 449940 269350
rect 449900 267164 449952 267170
rect 449900 267106 449952 267112
rect 450268 267164 450320 267170
rect 450268 267106 450320 267112
rect 449440 266756 449492 266762
rect 449440 266698 449492 266704
rect 449164 266416 449216 266422
rect 449164 266358 449216 266364
rect 449452 264316 449480 266698
rect 450280 264316 450308 267106
rect 451108 264316 451136 273906
rect 451476 268394 451504 277766
rect 452488 272678 452516 277780
rect 453592 276010 453620 277780
rect 453580 276004 453632 276010
rect 453580 275946 453632 275952
rect 453948 274780 454000 274786
rect 453948 274722 454000 274728
rect 453960 272950 453988 274722
rect 453948 272944 454000 272950
rect 453948 272886 454000 272892
rect 452476 272672 452528 272678
rect 452476 272614 452528 272620
rect 453856 272672 453908 272678
rect 453856 272614 453908 272620
rect 451740 272264 451792 272270
rect 451740 272206 451792 272212
rect 451464 268388 451516 268394
rect 451464 268330 451516 268336
rect 451752 267034 451780 272206
rect 453304 271584 453356 271590
rect 453304 271526 453356 271532
rect 451740 267028 451792 267034
rect 451740 266970 451792 266976
rect 451924 267028 451976 267034
rect 451924 266970 451976 266976
rect 451936 266914 451964 266970
rect 451246 266898 451964 266914
rect 451234 266892 451964 266898
rect 451286 266886 451964 266892
rect 451234 266834 451286 266840
rect 453316 266830 453344 271526
rect 453304 266824 453356 266830
rect 453304 266766 453356 266772
rect 452752 266688 452804 266694
rect 452752 266630 452804 266636
rect 451924 266416 451976 266422
rect 451924 266358 451976 266364
rect 451936 264316 451964 266358
rect 452764 264316 452792 266630
rect 453868 264330 453896 272614
rect 454788 271454 454816 277780
rect 455984 275330 456012 277780
rect 456984 276004 457036 276010
rect 456984 275946 457036 275952
rect 455972 275324 456024 275330
rect 455972 275266 456024 275272
rect 455880 275188 455932 275194
rect 455880 275130 455932 275136
rect 456800 275188 456852 275194
rect 456800 275130 456852 275136
rect 454776 271448 454828 271454
rect 454776 271390 454828 271396
rect 454684 271312 454736 271318
rect 454684 271254 454736 271260
rect 454408 266552 454460 266558
rect 454408 266494 454460 266500
rect 453606 264302 453896 264330
rect 454420 264316 454448 266494
rect 454696 266422 454724 271254
rect 455892 267734 455920 275130
rect 456812 273222 456840 275130
rect 456800 273216 456852 273222
rect 456800 273158 456852 273164
rect 456996 270774 457024 275946
rect 457180 274786 457208 277780
rect 457168 274780 457220 274786
rect 457168 274722 457220 274728
rect 458376 274106 458404 277780
rect 458364 274100 458416 274106
rect 458364 274042 458416 274048
rect 459376 274100 459428 274106
rect 459376 274042 459428 274048
rect 458088 272944 458140 272950
rect 458088 272886 458140 272892
rect 457444 271448 457496 271454
rect 457444 271390 457496 271396
rect 456984 270768 457036 270774
rect 456984 270710 457036 270716
rect 455800 267706 455920 267734
rect 455236 266824 455288 266830
rect 455236 266766 455288 266772
rect 454684 266416 454736 266422
rect 454684 266358 454736 266364
rect 455248 264316 455276 266766
rect 455800 266694 455828 267706
rect 456432 266892 456484 266898
rect 456432 266834 456484 266840
rect 455788 266688 455840 266694
rect 455788 266630 455840 266636
rect 456444 264330 456472 266834
rect 457456 266558 457484 271390
rect 457720 269816 457772 269822
rect 457720 269758 457772 269764
rect 457444 266552 457496 266558
rect 457444 266494 457496 266500
rect 456892 266416 456944 266422
rect 456892 266358 456944 266364
rect 456090 264302 456472 264330
rect 456904 264316 456932 266358
rect 457732 264316 457760 269758
rect 458100 266422 458128 272886
rect 459192 266620 459244 266626
rect 459192 266562 459244 266568
rect 458088 266416 458140 266422
rect 458088 266358 458140 266364
rect 458548 266416 458600 266422
rect 458548 266358 458600 266364
rect 458560 264316 458588 266358
rect 459204 264330 459232 266562
rect 459388 266422 459416 274042
rect 459572 269958 459600 277780
rect 460676 275058 460704 277780
rect 460664 275052 460716 275058
rect 460664 274994 460716 275000
rect 460020 273692 460072 273698
rect 460020 273634 460072 273640
rect 459560 269952 459612 269958
rect 459560 269894 459612 269900
rect 460032 267034 460060 273634
rect 461872 272542 461900 277780
rect 463068 275466 463096 277780
rect 463988 277766 464278 277794
rect 465092 277766 465474 277794
rect 463056 275460 463108 275466
rect 463056 275402 463108 275408
rect 463148 273216 463200 273222
rect 463148 273158 463200 273164
rect 461860 272536 461912 272542
rect 461860 272478 461912 272484
rect 461860 269952 461912 269958
rect 461860 269894 461912 269900
rect 461032 268388 461084 268394
rect 461032 268330 461084 268336
rect 460020 267028 460072 267034
rect 460020 266970 460072 266976
rect 460204 266484 460256 266490
rect 460204 266426 460256 266432
rect 459376 266416 459428 266422
rect 459376 266358 459428 266364
rect 459204 264302 459402 264330
rect 460216 264316 460244 266426
rect 461044 264316 461072 268330
rect 461872 264316 461900 269894
rect 463160 264330 463188 273158
rect 463516 272536 463568 272542
rect 463516 272478 463568 272484
rect 462714 264302 463188 264330
rect 463528 264316 463556 272478
rect 463988 271182 464016 277766
rect 464160 274780 464212 274786
rect 464160 274722 464212 274728
rect 463976 271176 464028 271182
rect 463976 271118 464028 271124
rect 464172 267306 464200 274722
rect 464528 271176 464580 271182
rect 464528 271118 464580 271124
rect 464540 267734 464568 271118
rect 465092 269278 465120 277766
rect 465724 270768 465776 270774
rect 465724 270710 465776 270716
rect 465080 269272 465132 269278
rect 465080 269214 465132 269220
rect 464356 267706 464568 267734
rect 465540 267708 465592 267714
rect 464160 267300 464212 267306
rect 464160 267242 464212 267248
rect 464356 266778 464384 267706
rect 465540 267650 465592 267656
rect 465552 267306 465580 267650
rect 465540 267300 465592 267306
rect 465540 267242 465592 267248
rect 465172 267028 465224 267034
rect 465172 266970 465224 266976
rect 464172 266750 464384 266778
rect 464172 266626 464200 266750
rect 464160 266620 464212 266626
rect 464160 266562 464212 266568
rect 464344 266620 464396 266626
rect 464344 266562 464396 266568
rect 464356 264316 464384 266562
rect 465184 264316 465212 266970
rect 465736 266626 465764 270710
rect 466656 270638 466684 277780
rect 467656 275460 467708 275466
rect 467656 275402 467708 275408
rect 466644 270632 466696 270638
rect 466644 270574 466696 270580
rect 466000 270088 466052 270094
rect 466000 270030 466052 270036
rect 465724 266620 465776 266626
rect 465724 266562 465776 266568
rect 466012 264316 466040 270030
rect 466828 267708 466880 267714
rect 466828 267650 466880 267656
rect 466840 264316 466868 267650
rect 467668 264316 467696 275402
rect 467852 275194 467880 277780
rect 468036 277766 468970 277794
rect 469232 277766 470166 277794
rect 467840 275188 467892 275194
rect 467840 275130 467892 275136
rect 468036 269550 468064 277766
rect 468208 275188 468260 275194
rect 468208 275130 468260 275136
rect 468024 269544 468076 269550
rect 468024 269486 468076 269492
rect 468220 267986 468248 275130
rect 468760 269272 468812 269278
rect 468760 269214 468812 269220
rect 468208 267980 468260 267986
rect 468208 267922 468260 267928
rect 468772 264330 468800 269214
rect 469232 268274 469260 277766
rect 470968 274916 471020 274922
rect 470968 274858 471020 274864
rect 470980 269822 471008 274858
rect 471348 274786 471376 277780
rect 471992 277766 472558 277794
rect 471336 274780 471388 274786
rect 471336 274722 471388 274728
rect 471244 274372 471296 274378
rect 471244 274314 471296 274320
rect 470968 269816 471020 269822
rect 470968 269758 471020 269764
rect 469048 268246 469260 268274
rect 469048 268122 469076 268246
rect 469036 268116 469088 268122
rect 469036 268058 469088 268064
rect 469220 268116 469272 268122
rect 469220 268058 469272 268064
rect 469232 266898 469260 268058
rect 471256 267306 471284 274314
rect 471612 269816 471664 269822
rect 471612 269758 471664 269764
rect 471624 267734 471652 269758
rect 471992 269414 472020 277766
rect 473740 272406 473768 277780
rect 474936 274650 474964 277780
rect 476146 277766 476344 277794
rect 474924 274644 474976 274650
rect 474924 274586 474976 274592
rect 475384 274644 475436 274650
rect 475384 274586 475436 274592
rect 473728 272400 473780 272406
rect 473728 272342 473780 272348
rect 474648 272400 474700 272406
rect 474648 272342 474700 272348
rect 473084 272128 473136 272134
rect 473084 272070 473136 272076
rect 471980 269408 472032 269414
rect 471980 269350 472032 269356
rect 471440 267706 471652 267734
rect 471244 267300 471296 267306
rect 471244 267242 471296 267248
rect 469220 266892 469272 266898
rect 469220 266834 469272 266840
rect 470140 266892 470192 266898
rect 470140 266834 470192 266840
rect 469312 266620 469364 266626
rect 469312 266562 469364 266568
rect 468510 264302 468800 264330
rect 469324 264316 469352 266562
rect 470152 264316 470180 266834
rect 471440 264330 471468 267706
rect 471796 267300 471848 267306
rect 471796 267242 471848 267248
rect 470994 264302 471468 264330
rect 471808 264316 471836 267242
rect 473096 264330 473124 272070
rect 474280 269544 474332 269550
rect 474280 269486 474332 269492
rect 473266 266656 473322 266665
rect 473266 266591 473268 266600
rect 473320 266591 473322 266600
rect 473452 266620 473504 266626
rect 473268 266562 473320 266568
rect 473452 266562 473504 266568
rect 472650 264302 473124 264330
rect 473464 264316 473492 266562
rect 474292 264316 474320 269486
rect 474660 266626 474688 272342
rect 475396 267306 475424 274586
rect 476316 270502 476344 277766
rect 477236 273834 477264 277780
rect 477224 273828 477276 273834
rect 477224 273770 477276 273776
rect 478432 272814 478460 277780
rect 478892 277766 479642 277794
rect 478420 272808 478472 272814
rect 478420 272750 478472 272756
rect 478696 271992 478748 271998
rect 478696 271934 478748 271940
rect 478144 270632 478196 270638
rect 478144 270574 478196 270580
rect 476304 270496 476356 270502
rect 476304 270438 476356 270444
rect 476764 269408 476816 269414
rect 476764 269350 476816 269356
rect 475384 267300 475436 267306
rect 475384 267242 475436 267248
rect 475936 267300 475988 267306
rect 475936 267242 475988 267248
rect 474830 266656 474886 266665
rect 474648 266620 474700 266626
rect 474830 266591 474832 266600
rect 474648 266562 474700 266568
rect 474884 266591 474886 266600
rect 474832 266562 474884 266568
rect 475108 266076 475160 266082
rect 475108 266018 475160 266024
rect 475120 264316 475148 266018
rect 475948 264316 475976 267242
rect 476776 264316 476804 269350
rect 477592 267708 477644 267714
rect 477592 267650 477644 267656
rect 477604 264316 477632 267650
rect 478156 266626 478184 270574
rect 478144 266620 478196 266626
rect 478144 266562 478196 266568
rect 478708 264330 478736 271934
rect 478892 269686 478920 277766
rect 480824 272270 480852 277780
rect 482020 273562 482048 277780
rect 483216 277394 483244 277780
rect 483124 277366 483244 277394
rect 482928 274780 482980 274786
rect 482928 274722 482980 274728
rect 482008 273556 482060 273562
rect 482008 273498 482060 273504
rect 481364 273420 481416 273426
rect 481364 273362 481416 273368
rect 480812 272264 480864 272270
rect 480812 272206 480864 272212
rect 479248 270496 479300 270502
rect 479248 270438 479300 270444
rect 478880 269680 478932 269686
rect 478880 269622 478932 269628
rect 478446 264302 478736 264330
rect 479260 264316 479288 270438
rect 480076 265668 480128 265674
rect 480076 265610 480128 265616
rect 480088 264316 480116 265610
rect 481376 264330 481404 273362
rect 482744 272808 482796 272814
rect 482744 272750 482796 272756
rect 481732 266620 481784 266626
rect 481732 266562 481784 266568
rect 480930 264302 481404 264330
rect 481744 264316 481772 266562
rect 482756 264330 482784 272750
rect 482940 272134 482968 274722
rect 482928 272128 482980 272134
rect 482928 272070 482980 272076
rect 483124 270366 483152 277366
rect 484320 273698 484348 277780
rect 484308 273692 484360 273698
rect 484308 273634 484360 273640
rect 483756 272128 483808 272134
rect 483756 272070 483808 272076
rect 483112 270360 483164 270366
rect 483112 270302 483164 270308
rect 483768 264330 483796 272070
rect 485516 271046 485544 277780
rect 486712 276010 486740 277780
rect 486700 276004 486752 276010
rect 486700 275946 486752 275952
rect 486884 276004 486936 276010
rect 486884 275946 486936 275952
rect 486896 273222 486924 275946
rect 487908 275874 487936 277780
rect 488736 277766 489118 277794
rect 487896 275868 487948 275874
rect 487896 275810 487948 275816
rect 488448 274508 488500 274514
rect 488448 274450 488500 274456
rect 488460 273834 488488 274450
rect 488448 273828 488500 273834
rect 488448 273770 488500 273776
rect 487988 273692 488040 273698
rect 487988 273634 488040 273640
rect 487068 273556 487120 273562
rect 487068 273498 487120 273504
rect 486884 273216 486936 273222
rect 486884 273158 486936 273164
rect 485504 271040 485556 271046
rect 485504 270982 485556 270988
rect 486700 270360 486752 270366
rect 486700 270302 486752 270308
rect 484216 269680 484268 269686
rect 484216 269622 484268 269628
rect 482586 264302 482784 264330
rect 483414 264302 483796 264330
rect 484228 264316 484256 269622
rect 485228 267572 485280 267578
rect 485228 267514 485280 267520
rect 485240 266626 485268 267514
rect 485228 266620 485280 266626
rect 485228 266562 485280 266568
rect 485872 266620 485924 266626
rect 485872 266562 485924 266568
rect 485044 265940 485096 265946
rect 485044 265882 485096 265888
rect 485056 264316 485084 265882
rect 485884 264316 485912 266562
rect 486712 264316 486740 270302
rect 487080 266626 487108 273498
rect 487068 266620 487120 266626
rect 487068 266562 487120 266568
rect 488000 264330 488028 273634
rect 488736 273086 488764 277766
rect 488908 275868 488960 275874
rect 488908 275810 488960 275816
rect 488724 273080 488776 273086
rect 488724 273022 488776 273028
rect 488356 272264 488408 272270
rect 488356 272206 488408 272212
rect 487554 264302 488028 264330
rect 488368 264316 488396 272206
rect 488540 271040 488592 271046
rect 488540 270982 488592 270988
rect 488552 267850 488580 270982
rect 488920 268258 488948 275810
rect 490300 273254 490328 277780
rect 491312 277766 491510 277794
rect 491312 274666 491340 277766
rect 492600 275874 492628 277780
rect 492588 275868 492640 275874
rect 492588 275810 492640 275816
rect 490564 274644 490616 274650
rect 490564 274586 490616 274592
rect 490748 274644 490800 274650
rect 490748 274586 490800 274592
rect 491036 274638 491340 274666
rect 490576 274378 490604 274586
rect 490564 274372 490616 274378
rect 490564 274314 490616 274320
rect 490760 274242 490788 274586
rect 491036 274514 491064 274638
rect 491024 274508 491076 274514
rect 491024 274450 491076 274456
rect 491208 274508 491260 274514
rect 491208 274450 491260 274456
rect 490748 274236 490800 274242
rect 490748 274178 490800 274184
rect 490932 274236 490984 274242
rect 490932 274178 490984 274184
rect 490944 273834 490972 274178
rect 490932 273828 490984 273834
rect 490932 273770 490984 273776
rect 490208 273226 490328 273254
rect 490208 269142 490236 273226
rect 490196 269136 490248 269142
rect 490196 269078 490248 269084
rect 488908 268252 488960 268258
rect 488908 268194 488960 268200
rect 488540 267844 488592 267850
rect 488540 267786 488592 267792
rect 489184 267844 489236 267850
rect 489184 267786 489236 267792
rect 489196 264316 489224 267786
rect 490012 266620 490064 266626
rect 490012 266562 490064 266568
rect 490024 264316 490052 266562
rect 491220 264330 491248 274450
rect 493796 274242 493824 277780
rect 494992 275194 495020 277780
rect 495164 276004 495216 276010
rect 495164 275946 495216 275952
rect 495440 276004 495492 276010
rect 495440 275946 495492 275952
rect 495176 275194 495204 275946
rect 494980 275188 495032 275194
rect 494980 275130 495032 275136
rect 495164 275188 495216 275194
rect 495164 275130 495216 275136
rect 494704 275052 494756 275058
rect 494704 274994 494756 275000
rect 493784 274236 493836 274242
rect 493784 274178 493836 274184
rect 492036 273828 492088 273834
rect 492036 273770 492088 273776
rect 492048 264330 492076 273770
rect 493692 273216 493744 273222
rect 493692 273158 493744 273164
rect 492772 268116 492824 268122
rect 492772 268058 492824 268064
rect 492784 267714 492812 268058
rect 492772 267708 492824 267714
rect 492772 267650 492824 267656
rect 492956 267708 493008 267714
rect 492956 267650 493008 267656
rect 492968 267594 492996 267650
rect 490866 264302 491248 264330
rect 491694 264302 492076 264330
rect 492508 267566 492996 267594
rect 492508 264316 492536 267566
rect 493704 264330 493732 273158
rect 494336 270360 494388 270366
rect 494334 270328 494336 270337
rect 494520 270360 494572 270366
rect 494388 270328 494390 270337
rect 494520 270302 494572 270308
rect 494334 270263 494390 270272
rect 494150 270056 494206 270065
rect 494150 269991 494206 270000
rect 493350 264302 493732 264330
rect 494164 264316 494192 269991
rect 494532 269686 494560 270302
rect 494520 269680 494572 269686
rect 494520 269622 494572 269628
rect 494716 267442 494744 274994
rect 495452 272406 495480 275946
rect 496188 274650 496216 277780
rect 496176 274644 496228 274650
rect 496176 274586 496228 274592
rect 496268 274236 496320 274242
rect 496268 274178 496320 274184
rect 495440 272400 495492 272406
rect 495440 272342 495492 272348
rect 494886 270328 494942 270337
rect 494886 270263 494942 270272
rect 494900 269686 494928 270263
rect 494888 269680 494940 269686
rect 494888 269622 494940 269628
rect 494704 267436 494756 267442
rect 494704 267378 494756 267384
rect 494980 265804 495032 265810
rect 494980 265746 495032 265752
rect 494992 264316 495020 265746
rect 496280 264330 496308 274178
rect 496636 273080 496688 273086
rect 496636 273022 496688 273028
rect 495834 264302 496308 264330
rect 496648 264316 496676 273022
rect 497384 270910 497412 277780
rect 498200 275868 498252 275874
rect 498200 275810 498252 275816
rect 497372 270904 497424 270910
rect 497372 270846 497424 270852
rect 498212 268122 498240 275810
rect 498580 275058 498608 277780
rect 499592 277766 499790 277794
rect 500512 277766 500894 277794
rect 498568 275052 498620 275058
rect 498568 274994 498620 275000
rect 499120 269068 499172 269074
rect 499120 269010 499172 269016
rect 498200 268116 498252 268122
rect 498200 268058 498252 268064
rect 497464 267436 497516 267442
rect 497464 267378 497516 267384
rect 497476 264316 497504 267378
rect 498568 266348 498620 266354
rect 498568 266290 498620 266296
rect 498580 264330 498608 266290
rect 498318 264302 498608 264330
rect 499132 264316 499160 269010
rect 499592 268802 499620 277766
rect 500512 271726 500540 277766
rect 502076 275738 502104 277780
rect 502536 277766 503286 277794
rect 504008 277766 504482 277794
rect 502064 275732 502116 275738
rect 502064 275674 502116 275680
rect 501972 274508 502024 274514
rect 501972 274450 502024 274456
rect 501604 272400 501656 272406
rect 501604 272342 501656 272348
rect 500500 271720 500552 271726
rect 500500 271662 500552 271668
rect 500868 271720 500920 271726
rect 500868 271662 500920 271668
rect 499580 268796 499632 268802
rect 499580 268738 499632 268744
rect 500684 268116 500736 268122
rect 500684 268058 500736 268064
rect 499762 267200 499818 267209
rect 499762 267135 499764 267144
rect 499816 267135 499818 267144
rect 499948 267164 500000 267170
rect 499764 267106 499816 267112
rect 499948 267106 500000 267112
rect 499960 264316 499988 267106
rect 500696 264330 500724 268058
rect 500880 267170 500908 271662
rect 501050 267200 501106 267209
rect 500868 267164 500920 267170
rect 501050 267135 501052 267144
rect 500868 267106 500920 267112
rect 501104 267135 501106 267144
rect 501052 267106 501104 267112
rect 501616 266354 501644 272342
rect 501604 266348 501656 266354
rect 501604 266290 501656 266296
rect 501984 264330 502012 274450
rect 502338 269648 502394 269657
rect 502338 269583 502394 269592
rect 502352 267578 502380 269583
rect 502536 268938 502564 277766
rect 504008 271862 504036 277766
rect 504548 276004 504600 276010
rect 504548 275946 504600 275952
rect 504916 276004 504968 276010
rect 504916 275946 504968 275952
rect 504560 275466 504588 275946
rect 504548 275460 504600 275466
rect 504548 275402 504600 275408
rect 504732 274508 504784 274514
rect 504732 274450 504784 274456
rect 504744 274394 504772 274450
rect 504192 274366 504772 274394
rect 504192 274242 504220 274366
rect 504180 274236 504232 274242
rect 504180 274178 504232 274184
rect 503996 271856 504048 271862
rect 503996 271798 504048 271804
rect 504732 271856 504784 271862
rect 504732 271798 504784 271804
rect 504178 270600 504234 270609
rect 504178 270535 504234 270544
rect 504192 270230 504220 270535
rect 504180 270224 504232 270230
rect 504180 270166 504232 270172
rect 504364 270224 504416 270230
rect 504364 270166 504416 270172
rect 504376 269686 504404 270166
rect 504364 269680 504416 269686
rect 504548 269680 504600 269686
rect 504364 269622 504416 269628
rect 504546 269648 504548 269657
rect 504600 269648 504602 269657
rect 504546 269583 504602 269592
rect 502524 268932 502576 268938
rect 502524 268874 502576 268880
rect 503076 268932 503128 268938
rect 503076 268874 503128 268880
rect 503088 268666 503116 268874
rect 504088 268796 504140 268802
rect 504088 268738 504140 268744
rect 503076 268660 503128 268666
rect 503076 268602 503128 268608
rect 503260 268660 503312 268666
rect 503260 268602 503312 268608
rect 502340 267572 502392 267578
rect 502340 267514 502392 267520
rect 502800 267572 502852 267578
rect 502800 267514 502852 267520
rect 502812 264330 502840 267514
rect 500696 264302 500802 264330
rect 501630 264302 502012 264330
rect 502458 264302 502840 264330
rect 503272 264316 503300 268602
rect 504100 268530 504128 268738
rect 504088 268524 504140 268530
rect 504088 268466 504140 268472
rect 504272 268524 504324 268530
rect 504272 268466 504324 268472
rect 504284 268258 504312 268466
rect 504272 268252 504324 268258
rect 504272 268194 504324 268200
rect 504744 267734 504772 271798
rect 504560 267706 504772 267734
rect 504560 264330 504588 267706
rect 504114 264302 504588 264330
rect 504928 264316 504956 275946
rect 505664 275874 505692 277780
rect 505652 275868 505704 275874
rect 505652 275810 505704 275816
rect 506860 275058 506888 277780
rect 507964 277394 507992 277780
rect 507872 277366 507992 277394
rect 507032 276004 507084 276010
rect 507032 275946 507084 275952
rect 507044 275058 507072 275946
rect 507216 275868 507268 275874
rect 507216 275810 507268 275816
rect 505100 275052 505152 275058
rect 505100 274994 505152 275000
rect 506848 275052 506900 275058
rect 506848 274994 506900 275000
rect 507032 275052 507084 275058
rect 507032 274994 507084 275000
rect 505112 268938 505140 274994
rect 505100 268932 505152 268938
rect 505100 268874 505152 268880
rect 505744 268252 505796 268258
rect 505744 268194 505796 268200
rect 505756 264316 505784 268194
rect 507228 267578 507256 275810
rect 507676 270904 507728 270910
rect 507676 270846 507728 270852
rect 506204 267572 506256 267578
rect 506204 267514 506256 267520
rect 506480 267572 506532 267578
rect 506480 267514 506532 267520
rect 507216 267572 507268 267578
rect 507216 267514 507268 267520
rect 507400 267572 507452 267578
rect 507400 267514 507452 267520
rect 506216 267209 506244 267514
rect 506492 267322 506520 267514
rect 506400 267294 506520 267322
rect 506202 267200 506258 267209
rect 506400 267170 506428 267294
rect 506202 267135 506258 267144
rect 506388 267164 506440 267170
rect 506388 267106 506440 267112
rect 506572 267164 506624 267170
rect 506572 267106 506624 267112
rect 506584 264316 506612 267106
rect 507412 264316 507440 267514
rect 507688 267170 507716 270846
rect 507872 270609 507900 277366
rect 508044 276004 508096 276010
rect 508044 275946 508096 275952
rect 508056 271726 508084 275946
rect 509160 275738 509188 277780
rect 509344 277766 510370 277794
rect 509148 275732 509200 275738
rect 509148 275674 509200 275680
rect 508044 271720 508096 271726
rect 508044 271662 508096 271668
rect 508964 271720 509016 271726
rect 508964 271662 509016 271668
rect 507858 270600 507914 270609
rect 507858 270535 507914 270544
rect 508228 268932 508280 268938
rect 508228 268874 508280 268880
rect 507858 267200 507914 267209
rect 507676 267164 507728 267170
rect 507858 267135 507860 267144
rect 507676 267106 507728 267112
rect 507912 267135 507914 267144
rect 507860 267106 507912 267112
rect 508240 264316 508268 268874
rect 508976 264330 509004 271662
rect 509344 268802 509372 277766
rect 511552 271590 511580 277780
rect 512748 275874 512776 277780
rect 513944 277394 513972 277780
rect 513852 277366 513972 277394
rect 512736 275868 512788 275874
rect 512736 275810 512788 275816
rect 512920 275868 512972 275874
rect 512920 275810 512972 275816
rect 512184 275732 512236 275738
rect 512184 275674 512236 275680
rect 512196 275330 512224 275674
rect 512184 275324 512236 275330
rect 512184 275266 512236 275272
rect 511540 271584 511592 271590
rect 511540 271526 511592 271532
rect 511908 271584 511960 271590
rect 511908 271526 511960 271532
rect 511724 271448 511776 271454
rect 511722 271416 511724 271425
rect 511776 271416 511778 271425
rect 511722 271351 511778 271360
rect 509882 269784 509938 269793
rect 509882 269719 509938 269728
rect 509332 268796 509384 268802
rect 509332 268738 509384 268744
rect 508976 264302 509082 264330
rect 509896 264316 509924 269719
rect 510712 268796 510764 268802
rect 510712 268738 510764 268744
rect 510724 264316 510752 268738
rect 511920 264330 511948 271526
rect 512932 266762 512960 275810
rect 513852 273970 513880 277366
rect 514024 276004 514076 276010
rect 514024 275946 514076 275952
rect 514036 275058 514064 275946
rect 514024 275052 514076 275058
rect 514024 274994 514076 275000
rect 513840 273964 513892 273970
rect 513840 273906 513892 273912
rect 513194 272368 513250 272377
rect 513194 272303 513250 272312
rect 512920 266756 512972 266762
rect 512920 266698 512972 266704
rect 512368 266416 512420 266422
rect 512368 266358 512420 266364
rect 511566 264302 511948 264330
rect 512380 264316 512408 266358
rect 513208 264316 513236 272303
rect 515140 271454 515168 277780
rect 515496 275868 515548 275874
rect 515496 275810 515548 275816
rect 515128 271448 515180 271454
rect 515312 271448 515364 271454
rect 515128 271390 515180 271396
rect 515310 271416 515312 271425
rect 515364 271416 515366 271425
rect 515310 271351 515366 271360
rect 514484 271312 514536 271318
rect 514484 271254 514536 271260
rect 514300 268796 514352 268802
rect 514300 268738 514352 268744
rect 514312 268682 514340 268738
rect 513760 268666 514340 268682
rect 513748 268660 514340 268666
rect 513800 268654 514340 268660
rect 513748 268602 513800 268608
rect 513380 266756 513432 266762
rect 513380 266698 513432 266704
rect 513392 266286 513420 266698
rect 513380 266280 513432 266286
rect 513380 266222 513432 266228
rect 514496 264330 514524 271254
rect 515508 266762 515536 275810
rect 516244 275738 516272 277780
rect 516428 277766 517454 277794
rect 516232 275732 516284 275738
rect 516232 275674 516284 275680
rect 516428 272678 516456 277766
rect 516784 275868 516836 275874
rect 516784 275810 516836 275816
rect 516598 274136 516654 274145
rect 516598 274071 516600 274080
rect 516652 274071 516654 274080
rect 516600 274042 516652 274048
rect 516416 272672 516468 272678
rect 516416 272614 516468 272620
rect 516600 272672 516652 272678
rect 516600 272614 516652 272620
rect 516612 272490 516640 272614
rect 516060 272462 516640 272490
rect 515496 266756 515548 266762
rect 515496 266698 515548 266704
rect 514852 266416 514904 266422
rect 514852 266358 514904 266364
rect 514050 264302 514524 264330
rect 514864 264316 514892 266358
rect 516060 264330 516088 272462
rect 516508 266756 516560 266762
rect 516508 266698 516560 266704
rect 515706 264302 516088 264330
rect 516520 264316 516548 266698
rect 516796 266422 516824 275810
rect 518440 274236 518492 274242
rect 518440 274178 518492 274184
rect 518452 272377 518480 274178
rect 518438 272368 518494 272377
rect 518438 272303 518494 272312
rect 518636 271454 518664 277780
rect 519832 276010 519860 277780
rect 520292 277766 521042 277794
rect 521856 277766 522238 277794
rect 523144 277766 523434 277794
rect 524538 277766 524736 277794
rect 519820 276004 519872 276010
rect 519820 275946 519872 275952
rect 520004 276004 520056 276010
rect 520004 275946 520056 275952
rect 519188 275862 519584 275890
rect 519188 275738 519216 275862
rect 519556 275754 519584 275862
rect 519176 275732 519228 275738
rect 519176 275674 519228 275680
rect 519360 275732 519412 275738
rect 519556 275726 519768 275754
rect 519360 275674 519412 275680
rect 519372 275330 519400 275674
rect 519740 275602 519768 275726
rect 519544 275596 519596 275602
rect 519544 275538 519596 275544
rect 519728 275596 519780 275602
rect 519728 275538 519780 275544
rect 519556 275330 519584 275538
rect 519360 275324 519412 275330
rect 519360 275266 519412 275272
rect 519544 275324 519596 275330
rect 519544 275266 519596 275272
rect 519726 274136 519782 274145
rect 519726 274071 519782 274080
rect 519740 273970 519768 274071
rect 519728 273964 519780 273970
rect 519728 273906 519780 273912
rect 520016 271674 520044 275946
rect 519924 271646 520044 271674
rect 518624 271448 518676 271454
rect 518624 271390 518676 271396
rect 518438 268560 518494 268569
rect 518438 268495 518494 268504
rect 518990 268560 519046 268569
rect 519046 268530 519400 268546
rect 519046 268524 519412 268530
rect 519046 268518 519360 268524
rect 518990 268495 519046 268504
rect 517336 266484 517388 266490
rect 517336 266426 517388 266432
rect 516784 266416 516836 266422
rect 516784 266358 516836 266364
rect 517348 264316 517376 266426
rect 518452 264330 518480 268495
rect 519360 268466 519412 268472
rect 519174 268424 519230 268433
rect 518820 268394 519174 268410
rect 518808 268388 519174 268394
rect 518860 268382 519174 268388
rect 519174 268359 519230 268368
rect 518808 268330 518860 268336
rect 519924 267734 519952 271646
rect 520096 271448 520148 271454
rect 520096 271390 520148 271396
rect 519832 267706 519952 267734
rect 518898 267336 518954 267345
rect 518898 267271 518900 267280
rect 518952 267271 518954 267280
rect 519176 267300 519228 267306
rect 518900 267242 518952 267248
rect 519176 267242 519228 267248
rect 519188 267034 519216 267242
rect 519176 267028 519228 267034
rect 519176 266970 519228 266976
rect 519360 267028 519412 267034
rect 519360 266970 519412 266976
rect 519176 266892 519228 266898
rect 519176 266834 519228 266840
rect 518714 266792 518770 266801
rect 518714 266727 518716 266736
rect 518768 266727 518770 266736
rect 518898 266792 518954 266801
rect 519188 266778 519216 266834
rect 518954 266750 519216 266778
rect 518898 266727 518954 266736
rect 518716 266698 518768 266704
rect 519372 264330 519400 266970
rect 518190 264302 518480 264330
rect 519018 264302 519400 264330
rect 519832 264316 519860 267706
rect 520108 267034 520136 271390
rect 520292 268394 520320 277766
rect 521106 273728 521162 273737
rect 521106 273663 521162 273672
rect 520462 268424 520518 268433
rect 520280 268388 520332 268394
rect 520462 268359 520464 268368
rect 520280 268330 520332 268336
rect 520516 268359 520518 268368
rect 520464 268330 520516 268336
rect 520096 267028 520148 267034
rect 520096 266970 520148 266976
rect 520280 267028 520332 267034
rect 520280 266970 520332 266976
rect 520292 266354 520320 266970
rect 520280 266348 520332 266354
rect 520280 266290 520332 266296
rect 521120 264330 521148 273663
rect 521856 272950 521884 277766
rect 522396 276412 522448 276418
rect 522396 276354 522448 276360
rect 522212 276276 522264 276282
rect 522212 276218 522264 276224
rect 522224 275738 522252 276218
rect 522212 275732 522264 275738
rect 522212 275674 522264 275680
rect 522408 275602 522436 276354
rect 522396 275596 522448 275602
rect 522396 275538 522448 275544
rect 523144 274922 523172 277766
rect 523132 274916 523184 274922
rect 523132 274858 523184 274864
rect 523316 274916 523368 274922
rect 523316 274858 523368 274864
rect 521844 272944 521896 272950
rect 521844 272886 521896 272892
rect 521474 272504 521530 272513
rect 521474 272439 521530 272448
rect 520674 264302 521148 264330
rect 521488 264316 521516 272439
rect 523328 269793 523356 274858
rect 524708 274530 524736 277766
rect 525260 277766 525734 277794
rect 524880 276140 524932 276146
rect 524880 276082 524932 276088
rect 524892 275874 524920 276082
rect 524880 275868 524932 275874
rect 524880 275810 524932 275816
rect 524432 274502 524736 274530
rect 524432 274394 524460 274502
rect 524248 274366 524460 274394
rect 524248 273970 524276 274366
rect 524236 273964 524288 273970
rect 524236 273906 524288 273912
rect 524420 273964 524472 273970
rect 524420 273906 524472 273912
rect 524432 273850 524460 273906
rect 524248 273822 524460 273850
rect 524248 273737 524276 273822
rect 524234 273728 524290 273737
rect 524234 273663 524290 273672
rect 524386 273006 524736 273034
rect 524386 272950 524414 273006
rect 524374 272944 524426 272950
rect 524374 272886 524426 272892
rect 524512 272944 524564 272950
rect 524512 272886 524564 272892
rect 524524 272678 524552 272886
rect 524708 272762 524736 273006
rect 524708 272734 525104 272762
rect 524328 272672 524380 272678
rect 524328 272614 524380 272620
rect 524512 272672 524564 272678
rect 524512 272614 524564 272620
rect 524880 272672 524932 272678
rect 524880 272614 524932 272620
rect 523958 271688 524014 271697
rect 523958 271623 524014 271632
rect 523972 271454 524000 271623
rect 523960 271448 524012 271454
rect 523960 271390 524012 271396
rect 524144 271448 524196 271454
rect 524144 271390 524196 271396
rect 523960 270904 524012 270910
rect 523958 270872 523960 270881
rect 524012 270872 524014 270881
rect 523958 270807 524014 270816
rect 523314 269784 523370 269793
rect 523314 269719 523370 269728
rect 521658 269512 521714 269521
rect 521658 269447 521714 269456
rect 521672 267306 521700 269447
rect 521660 267300 521712 267306
rect 521660 267242 521712 267248
rect 522948 267300 523000 267306
rect 522948 267242 523000 267248
rect 523960 267300 524012 267306
rect 523960 267242 524012 267248
rect 522960 267034 522988 267242
rect 523972 267186 524000 267242
rect 523604 267170 524000 267186
rect 523592 267164 524000 267170
rect 523644 267158 524000 267164
rect 523592 267106 523644 267112
rect 522948 267028 523000 267034
rect 522948 266970 523000 266976
rect 523132 267028 523184 267034
rect 523132 266970 523184 266976
rect 522672 266348 522724 266354
rect 522672 266290 522724 266296
rect 522684 264330 522712 266290
rect 522330 264302 522712 264330
rect 523144 264316 523172 266970
rect 524156 264330 524184 271390
rect 524340 267034 524368 272614
rect 524604 272536 524656 272542
rect 524892 272513 524920 272614
rect 525076 272542 525104 272734
rect 525064 272536 525116 272542
rect 524604 272478 524656 272484
rect 524878 272504 524934 272513
rect 524616 272241 524644 272478
rect 525064 272478 525116 272484
rect 524878 272439 524934 272448
rect 524602 272232 524658 272241
rect 524602 272167 524658 272176
rect 525260 271810 525288 277766
rect 526916 276418 526944 277780
rect 527192 277766 528126 277794
rect 526904 276412 526956 276418
rect 526904 276354 526956 276360
rect 525798 275768 525854 275777
rect 525798 275703 525854 275712
rect 524616 271782 525288 271810
rect 524616 271182 524644 271782
rect 524786 271688 524842 271697
rect 524786 271623 524842 271632
rect 524800 271182 524828 271623
rect 524604 271176 524656 271182
rect 524604 271118 524656 271124
rect 524788 271176 524840 271182
rect 524788 271118 524840 271124
rect 524880 270904 524932 270910
rect 524878 270872 524880 270881
rect 524932 270872 524934 270881
rect 524878 270807 524934 270816
rect 525812 269226 525840 275703
rect 526258 271144 526314 271153
rect 526258 271079 526314 271088
rect 526272 270774 526300 271079
rect 526260 270768 526312 270774
rect 526260 270710 526312 270716
rect 526444 270768 526496 270774
rect 526444 270710 526496 270716
rect 525720 269198 525840 269226
rect 525522 268696 525578 268705
rect 525522 268631 525578 268640
rect 524510 267064 524566 267073
rect 524328 267028 524380 267034
rect 524510 266999 524566 267008
rect 524788 267028 524840 267034
rect 524328 266970 524380 266976
rect 524524 266880 524552 266999
rect 524788 266970 524840 266976
rect 524386 266852 524552 266880
rect 524386 266762 524414 266852
rect 524374 266756 524426 266762
rect 524374 266698 524426 266704
rect 524512 266756 524564 266762
rect 524512 266698 524564 266704
rect 524524 266354 524552 266698
rect 524512 266348 524564 266354
rect 524512 266290 524564 266296
rect 523986 264302 524184 264330
rect 524800 264316 524828 266970
rect 525536 264330 525564 268631
rect 525720 267034 525748 269198
rect 525890 267064 525946 267073
rect 525708 267028 525760 267034
rect 525890 266999 525892 267008
rect 525708 266970 525760 266976
rect 525944 266999 525946 267008
rect 525892 266970 525944 266976
rect 525536 264302 525642 264330
rect 526456 264316 526484 270710
rect 527192 268546 527220 277766
rect 527822 274680 527878 274689
rect 527822 274615 527878 274624
rect 527836 274106 527864 274615
rect 527824 274100 527876 274106
rect 527824 274042 527876 274048
rect 528008 274100 528060 274106
rect 528008 274042 528060 274048
rect 527008 268518 527220 268546
rect 527008 268394 527036 268518
rect 526996 268388 527048 268394
rect 526996 268330 527048 268336
rect 527180 268388 527232 268394
rect 527180 268330 527232 268336
rect 527192 267345 527220 268330
rect 527178 267336 527234 267345
rect 527178 267271 527234 267280
rect 527638 267336 527694 267345
rect 527638 267271 527694 267280
rect 527652 264330 527680 267271
rect 527298 264302 527680 264330
rect 528020 264330 528048 274042
rect 529308 273254 529336 277780
rect 530504 276282 530532 277780
rect 530492 276276 530544 276282
rect 530492 276218 530544 276224
rect 530858 275768 530914 275777
rect 530308 275732 530360 275738
rect 530858 275703 530860 275712
rect 530308 275674 530360 275680
rect 530912 275703 530914 275712
rect 530860 275674 530912 275680
rect 529216 273226 529336 273254
rect 529020 271312 529072 271318
rect 529020 271254 529072 271260
rect 529032 270774 529060 271254
rect 528652 270768 528704 270774
rect 528650 270736 528652 270745
rect 529020 270768 529072 270774
rect 528704 270736 528706 270745
rect 529020 270710 529072 270716
rect 528650 270671 528706 270680
rect 528468 270224 528520 270230
rect 528520 270172 529060 270178
rect 528468 270166 529060 270172
rect 528480 270150 529060 270166
rect 529032 270094 529060 270150
rect 529020 270088 529072 270094
rect 529020 270030 529072 270036
rect 529216 269958 529244 273226
rect 529388 271448 529440 271454
rect 529388 271390 529440 271396
rect 529400 271182 529428 271390
rect 529388 271176 529440 271182
rect 529572 271176 529624 271182
rect 529388 271118 529440 271124
rect 529570 271144 529572 271153
rect 529624 271144 529626 271153
rect 529570 271079 529626 271088
rect 529754 271144 529810 271153
rect 529754 271079 529810 271088
rect 529768 270042 529796 271079
rect 529400 270014 529796 270042
rect 529204 269952 529256 269958
rect 529204 269894 529256 269900
rect 529400 264330 529428 270014
rect 530320 269958 530348 275674
rect 531608 273254 531636 277780
rect 531516 273226 531636 273254
rect 531516 272241 531544 273226
rect 531502 272232 531558 272241
rect 531502 272167 531558 272176
rect 532804 271182 532832 277780
rect 532988 277766 534014 277794
rect 534184 277766 535210 277794
rect 535472 277766 536406 277794
rect 532792 271176 532844 271182
rect 532792 271118 532844 271124
rect 532988 270178 533016 277766
rect 534184 273254 534212 277766
rect 535090 275360 535146 275369
rect 535090 275295 535146 275304
rect 534184 273226 534396 273254
rect 534078 272776 534134 272785
rect 534078 272711 534134 272720
rect 534092 272626 534120 272711
rect 534000 272598 534120 272626
rect 534000 272542 534028 272598
rect 533988 272536 534040 272542
rect 533526 272504 533582 272513
rect 534172 272536 534224 272542
rect 533988 272478 534040 272484
rect 534170 272504 534172 272513
rect 534224 272504 534226 272513
rect 533526 272439 533582 272448
rect 534170 272439 534226 272448
rect 533160 271176 533212 271182
rect 533160 271118 533212 271124
rect 533172 270745 533200 271118
rect 533158 270736 533214 270745
rect 533158 270671 533214 270680
rect 532712 270150 533016 270178
rect 531410 270056 531466 270065
rect 531410 269991 531466 270000
rect 529756 269952 529808 269958
rect 529756 269894 529808 269900
rect 530308 269952 530360 269958
rect 530308 269894 530360 269900
rect 530584 269952 530636 269958
rect 530584 269894 530636 269900
rect 528020 264302 528126 264330
rect 528954 264302 529428 264330
rect 529768 264316 529796 269894
rect 530596 264316 530624 269894
rect 531424 264316 531452 269991
rect 532712 269521 532740 270150
rect 532884 269952 532936 269958
rect 532884 269894 532936 269900
rect 533068 269952 533120 269958
rect 533068 269894 533120 269900
rect 532896 269793 532924 269894
rect 532882 269784 532938 269793
rect 532882 269719 532938 269728
rect 532698 269512 532754 269521
rect 532698 269447 532754 269456
rect 532238 266928 532294 266937
rect 532238 266863 532294 266872
rect 532252 264316 532280 266863
rect 533080 264316 533108 269894
rect 533540 264330 533568 272439
rect 534368 270881 534396 273226
rect 533894 270872 533950 270881
rect 533894 270807 533950 270816
rect 534354 270872 534410 270881
rect 534354 270807 534410 270816
rect 533908 270230 533936 270807
rect 533896 270224 533948 270230
rect 533896 270166 533948 270172
rect 534034 270224 534086 270230
rect 534034 270166 534086 270172
rect 534046 270042 534074 270166
rect 533908 270014 534074 270042
rect 533908 269793 533936 270014
rect 533894 269784 533950 269793
rect 533894 269719 533950 269728
rect 533894 268696 533950 268705
rect 533950 268654 534074 268682
rect 533894 268631 533950 268640
rect 534046 268530 534074 268654
rect 533896 268524 533948 268530
rect 533896 268466 533948 268472
rect 534034 268524 534086 268530
rect 534034 268466 534086 268472
rect 533908 268138 533936 268466
rect 533908 268110 534074 268138
rect 534046 267986 534074 268110
rect 533896 267980 533948 267986
rect 533896 267922 533948 267928
rect 534034 267980 534086 267986
rect 534034 267922 534086 267928
rect 533908 267753 533936 267922
rect 533894 267744 533950 267753
rect 533894 267679 533950 267688
rect 533710 267336 533766 267345
rect 533766 267294 534074 267322
rect 533710 267271 533766 267280
rect 533894 267200 533950 267209
rect 533894 267135 533950 267144
rect 533908 267034 533936 267135
rect 534046 267034 534074 267294
rect 534170 267200 534226 267209
rect 534170 267135 534226 267144
rect 533896 267028 533948 267034
rect 533896 266970 533948 266976
rect 534034 267028 534086 267034
rect 534034 266970 534086 266976
rect 534184 266898 534212 267135
rect 533988 266892 534040 266898
rect 533988 266834 534040 266840
rect 534172 266892 534224 266898
rect 534172 266834 534224 266840
rect 534000 266778 534028 266834
rect 534000 266750 534120 266778
rect 534092 266665 534120 266750
rect 534078 266656 534134 266665
rect 534078 266591 534134 266600
rect 535104 264330 535132 275295
rect 535472 267753 535500 277766
rect 536838 275632 536894 275641
rect 536838 275567 536840 275576
rect 536892 275567 536894 275576
rect 537024 275596 537076 275602
rect 536840 275538 536892 275544
rect 537024 275538 537076 275544
rect 536746 273864 536802 273873
rect 536746 273799 536802 273808
rect 535918 269512 535974 269521
rect 535918 269447 535974 269456
rect 535458 267744 535514 267753
rect 535458 267679 535514 267688
rect 535932 264330 535960 269447
rect 536760 264330 536788 273799
rect 537036 273254 537064 275538
rect 537588 275330 537616 277780
rect 538784 277394 538812 277780
rect 539612 277766 539902 277794
rect 538784 277366 538904 277394
rect 537942 275632 537998 275641
rect 537760 275596 537812 275602
rect 537942 275567 537944 275576
rect 537760 275538 537812 275544
rect 537996 275567 537998 275576
rect 537944 275538 537996 275544
rect 537772 275330 537800 275538
rect 538232 275466 538536 275482
rect 538220 275460 538536 275466
rect 538272 275454 538536 275460
rect 538220 275402 538272 275408
rect 537576 275324 537628 275330
rect 537576 275266 537628 275272
rect 537760 275324 537812 275330
rect 537760 275266 537812 275272
rect 538508 274786 538536 275454
rect 538678 275360 538734 275369
rect 538678 275295 538680 275304
rect 538732 275295 538734 275304
rect 538680 275266 538732 275272
rect 538678 274952 538734 274961
rect 538678 274887 538734 274896
rect 538312 274780 538364 274786
rect 538312 274722 538364 274728
rect 538496 274780 538548 274786
rect 538496 274722 538548 274728
rect 538324 274666 538352 274722
rect 538692 274666 538720 274887
rect 538324 274638 538720 274666
rect 538876 273254 538904 277366
rect 537036 273226 537248 273254
rect 537024 269272 537076 269278
rect 537022 269240 537024 269249
rect 537076 269240 537078 269249
rect 537022 269175 537078 269184
rect 537220 266898 537248 273226
rect 538692 273226 538904 273254
rect 537944 269816 537996 269822
rect 537944 269758 537996 269764
rect 538126 269784 538182 269793
rect 537956 269550 537984 269758
rect 538126 269719 538182 269728
rect 537944 269544 537996 269550
rect 537944 269486 537996 269492
rect 537574 267608 537630 267617
rect 537574 267543 537630 267552
rect 537208 266892 537260 266898
rect 537208 266834 537260 266840
rect 537392 266892 537444 266898
rect 537392 266834 537444 266840
rect 537404 266665 537432 266834
rect 537390 266656 537446 266665
rect 537390 266591 537446 266600
rect 537588 264330 537616 267543
rect 538140 264602 538168 269719
rect 538692 269249 538720 273226
rect 539612 270722 539640 277766
rect 541084 277394 541112 277780
rect 540992 277366 541112 277394
rect 541820 277766 542294 277794
rect 543200 277766 543490 277794
rect 540992 275466 541020 277366
rect 540980 275460 541032 275466
rect 540980 275402 541032 275408
rect 541164 275460 541216 275466
rect 541164 275402 541216 275408
rect 541176 274961 541204 275402
rect 541162 274952 541218 274961
rect 541162 274887 541218 274896
rect 538876 270694 539640 270722
rect 540520 270768 540572 270774
rect 540520 270710 540572 270716
rect 538876 270638 538904 270694
rect 538864 270632 538916 270638
rect 538864 270574 538916 270580
rect 539506 270600 539562 270609
rect 539506 270535 539562 270544
rect 538864 270088 538916 270094
rect 538864 270030 538916 270036
rect 538876 269822 538904 270030
rect 538864 269816 538916 269822
rect 538864 269758 538916 269764
rect 538678 269240 538734 269249
rect 538678 269175 538734 269184
rect 539230 268152 539286 268161
rect 539230 268087 539286 268096
rect 533540 264302 533922 264330
rect 534750 264302 535132 264330
rect 535578 264302 535960 264330
rect 536406 264302 536788 264330
rect 537234 264302 537616 264330
rect 538048 264574 538168 264602
rect 538048 264316 538076 264574
rect 539244 264330 539272 268087
rect 539520 266898 539548 270535
rect 539508 266892 539560 266898
rect 539508 266834 539560 266840
rect 539692 266892 539744 266898
rect 539692 266834 539744 266840
rect 538890 264302 539272 264330
rect 539704 264316 539732 266834
rect 540532 264316 540560 270710
rect 541820 270094 541848 277766
rect 543200 274689 543228 277766
rect 544672 275466 544700 277780
rect 544660 275460 544712 275466
rect 544660 275402 544712 275408
rect 544844 275460 544896 275466
rect 544844 275402 544896 275408
rect 543186 274680 543242 274689
rect 543186 274615 543242 274624
rect 544856 272785 544884 275402
rect 545868 274786 545896 277780
rect 546512 277766 547078 277794
rect 547892 277766 548182 277794
rect 546040 275460 546092 275466
rect 546040 275402 546092 275408
rect 546224 275460 546276 275466
rect 546224 275402 546276 275408
rect 546052 274786 546080 275402
rect 545856 274780 545908 274786
rect 545856 274722 545908 274728
rect 546040 274780 546092 274786
rect 546040 274722 546092 274728
rect 544842 272776 544898 272785
rect 544842 272711 544898 272720
rect 543002 272504 543058 272513
rect 543002 272439 543058 272448
rect 540980 270088 541032 270094
rect 540980 270030 541032 270036
rect 541808 270088 541860 270094
rect 541808 270030 541860 270036
rect 541992 270088 542044 270094
rect 541992 270030 542044 270036
rect 540992 269550 541020 270030
rect 540980 269544 541032 269550
rect 540980 269486 541032 269492
rect 541348 269544 541400 269550
rect 542004 269521 542032 270030
rect 541348 269486 541400 269492
rect 541990 269512 542046 269521
rect 541360 264316 541388 269486
rect 541990 269447 542046 269456
rect 542174 267336 542230 267345
rect 542174 267271 542230 267280
rect 542188 264316 542216 267271
rect 543016 264316 543044 272439
rect 546236 271561 546264 275402
rect 543554 271552 543610 271561
rect 543554 271487 543610 271496
rect 546222 271552 546278 271561
rect 546222 271487 546278 271496
rect 543568 270774 543596 271487
rect 543556 270768 543608 270774
rect 543556 270710 543608 270716
rect 543694 270768 543746 270774
rect 543694 270710 543746 270716
rect 543554 270600 543610 270609
rect 543706 270586 543734 270710
rect 543610 270558 543734 270586
rect 543554 270535 543610 270544
rect 546512 269498 546540 277766
rect 546236 269470 546540 269498
rect 546236 269414 546264 269470
rect 546224 269408 546276 269414
rect 546224 269350 546276 269356
rect 546408 269408 546460 269414
rect 546408 269350 546460 269356
rect 543554 267608 543610 267617
rect 543554 267543 543610 267552
rect 543568 267458 543596 267543
rect 543568 267430 543734 267458
rect 543706 267306 543734 267430
rect 543556 267300 543608 267306
rect 543556 267242 543608 267248
rect 543694 267300 543746 267306
rect 543694 267242 543746 267248
rect 543568 266642 543596 267242
rect 543568 266626 543734 266642
rect 543568 266620 543746 266626
rect 543568 266614 543694 266620
rect 543694 266562 543746 266568
rect 546420 266354 546448 269350
rect 547510 268424 547566 268433
rect 547510 268359 547512 268368
rect 547564 268359 547566 268368
rect 547696 268388 547748 268394
rect 547512 268330 547564 268336
rect 547696 268330 547748 268336
rect 547708 268161 547736 268330
rect 547694 268152 547750 268161
rect 547694 268087 547750 268096
rect 546408 266348 546460 266354
rect 546408 266290 546460 266296
rect 547892 266082 547920 277766
rect 549364 277394 549392 277780
rect 549640 277766 550574 277794
rect 549640 277394 549668 277766
rect 549272 277366 549392 277394
rect 549456 277366 549668 277394
rect 549272 268433 549300 277366
rect 549456 269278 549484 277366
rect 551756 271046 551784 277780
rect 552492 277766 552966 277794
rect 553412 277766 554162 277794
rect 554792 277766 555266 277794
rect 552492 271998 552520 277766
rect 552480 271992 552532 271998
rect 552480 271934 552532 271940
rect 552848 271992 552900 271998
rect 552848 271934 552900 271940
rect 551744 271040 551796 271046
rect 551744 270982 551796 270988
rect 552664 271040 552716 271046
rect 552664 270982 552716 270988
rect 552202 270736 552258 270745
rect 552202 270671 552258 270680
rect 552216 270502 552244 270671
rect 552676 270638 552704 270982
rect 552664 270632 552716 270638
rect 552664 270574 552716 270580
rect 552204 270496 552256 270502
rect 552204 270438 552256 270444
rect 552388 270496 552440 270502
rect 552388 270438 552440 270444
rect 552400 269906 552428 270438
rect 552308 269878 552428 269906
rect 552308 269822 552336 269878
rect 552296 269816 552348 269822
rect 552296 269758 552348 269764
rect 552480 269816 552532 269822
rect 552480 269758 552532 269764
rect 552492 269634 552520 269758
rect 552400 269606 552520 269634
rect 552400 269550 552428 269606
rect 552388 269544 552440 269550
rect 552388 269486 552440 269492
rect 551928 269408 551980 269414
rect 551980 269356 552336 269362
rect 551928 269350 552336 269356
rect 551940 269334 552336 269350
rect 552308 269278 552336 269334
rect 549444 269272 549496 269278
rect 549444 269214 549496 269220
rect 549628 269272 549680 269278
rect 549628 269214 549680 269220
rect 552296 269272 552348 269278
rect 552296 269214 552348 269220
rect 549258 268424 549314 268433
rect 549258 268359 549314 268368
rect 549640 266490 549668 269214
rect 552860 267442 552888 271934
rect 553412 270745 553440 277766
rect 553398 270736 553454 270745
rect 553398 270671 553454 270680
rect 553032 269680 553084 269686
rect 553032 269622 553084 269628
rect 553044 269414 553072 269622
rect 553032 269408 553084 269414
rect 553032 269350 553084 269356
rect 552848 267436 552900 267442
rect 552848 267378 552900 267384
rect 553032 267436 553084 267442
rect 553032 267378 553084 267384
rect 553044 266626 553072 267378
rect 553032 266620 553084 266626
rect 553032 266562 553084 266568
rect 549628 266484 549680 266490
rect 549628 266426 549680 266432
rect 547880 266076 547932 266082
rect 547880 266018 547932 266024
rect 554792 265674 554820 277766
rect 556448 273426 556476 277780
rect 557644 277394 557672 277780
rect 557552 277366 557672 277394
rect 556436 273420 556488 273426
rect 556436 273362 556488 273368
rect 557552 269414 557580 277366
rect 558840 274786 558868 277780
rect 558828 274780 558880 274786
rect 558828 274722 558880 274728
rect 560036 272134 560064 277780
rect 560312 277766 561246 277794
rect 561692 277766 562442 277794
rect 560024 272128 560076 272134
rect 560024 272070 560076 272076
rect 560312 270366 560340 277766
rect 560300 270360 560352 270366
rect 560300 270302 560352 270308
rect 558920 269680 558972 269686
rect 558920 269622 558972 269628
rect 557540 269408 557592 269414
rect 557540 269350 557592 269356
rect 558932 267714 558960 269622
rect 558920 267708 558972 267714
rect 558920 267650 558972 267656
rect 561692 265946 561720 277766
rect 563532 273562 563560 277780
rect 564452 277766 564742 277794
rect 563520 273556 563572 273562
rect 563520 273498 563572 273504
rect 564452 270502 564480 277766
rect 565924 273698 565952 277780
rect 565912 273692 565964 273698
rect 565912 273634 565964 273640
rect 567120 272270 567148 277780
rect 567304 277766 568330 277794
rect 568592 277766 569526 277794
rect 567108 272264 567160 272270
rect 567108 272206 567160 272212
rect 564440 270496 564492 270502
rect 564440 270438 564492 270444
rect 567304 267850 567332 277766
rect 568592 269550 568620 277766
rect 570708 274650 570736 277780
rect 570696 274644 570748 274650
rect 570696 274586 570748 274592
rect 570880 274644 570932 274650
rect 570880 274586 570932 274592
rect 568580 269544 568632 269550
rect 568580 269486 568632 269492
rect 567292 267844 567344 267850
rect 567292 267786 567344 267792
rect 570892 267442 570920 274586
rect 571812 273834 571840 277780
rect 572732 277766 573022 277794
rect 571800 273828 571852 273834
rect 571800 273770 571852 273776
rect 572732 269686 572760 277766
rect 574204 273222 574232 277780
rect 574480 277766 575414 277794
rect 575584 277766 576610 277794
rect 574192 273216 574244 273222
rect 574192 273158 574244 273164
rect 574480 270337 574508 277766
rect 574466 270328 574522 270337
rect 574466 270263 574522 270272
rect 572720 269680 572772 269686
rect 572720 269622 572772 269628
rect 570880 267436 570932 267442
rect 570880 267378 570932 267384
rect 561680 265940 561732 265946
rect 561680 265882 561732 265888
rect 575584 265810 575612 277766
rect 577792 274514 577820 277780
rect 578528 277766 578910 277794
rect 577780 274508 577832 274514
rect 577780 274450 577832 274456
rect 578528 273086 578556 277766
rect 578884 273216 578936 273222
rect 578884 273158 578936 273164
rect 578516 273080 578568 273086
rect 578516 273022 578568 273028
rect 578896 267578 578924 273158
rect 580092 271998 580120 277780
rect 580264 273080 580316 273086
rect 580264 273022 580316 273028
rect 580080 271992 580132 271998
rect 580080 271934 580132 271940
rect 578884 267572 578936 267578
rect 578884 267514 578936 267520
rect 580276 266898 580304 273022
rect 581288 272406 581316 277780
rect 582484 277394 582512 277780
rect 582392 277366 582512 277394
rect 581276 272400 581328 272406
rect 581276 272342 581328 272348
rect 582392 269074 582420 277366
rect 583680 275058 583708 277780
rect 584048 277766 584890 277794
rect 583668 275052 583720 275058
rect 583668 274994 583720 275000
rect 582380 269068 582432 269074
rect 582380 269010 582432 269016
rect 581644 268796 581696 268802
rect 581644 268738 581696 268744
rect 581828 268796 581880 268802
rect 581828 268738 581880 268744
rect 581656 268122 581684 268738
rect 580448 268116 580500 268122
rect 580448 268058 580500 268064
rect 581644 268116 581696 268122
rect 581644 268058 581696 268064
rect 580460 267850 580488 268058
rect 581840 267986 581868 268738
rect 581828 267980 581880 267986
rect 581828 267922 581880 267928
rect 584048 267850 584076 277766
rect 585784 274508 585836 274514
rect 585784 274450 585836 274456
rect 580448 267844 580500 267850
rect 580448 267786 580500 267792
rect 584036 267844 584088 267850
rect 584036 267786 584088 267792
rect 585796 267170 585824 274450
rect 586072 274378 586100 277780
rect 587176 274650 587204 277780
rect 587912 277766 588386 277794
rect 587164 274644 587216 274650
rect 587164 274586 587216 274592
rect 586060 274372 586112 274378
rect 586060 274314 586112 274320
rect 587912 268122 587940 277766
rect 589568 271862 589596 277780
rect 590764 275194 590792 277780
rect 591040 277766 591974 277794
rect 590752 275188 590804 275194
rect 590752 275130 590804 275136
rect 589556 271856 589608 271862
rect 589556 271798 589608 271804
rect 590660 269068 590712 269074
rect 590660 269010 590712 269016
rect 590672 268666 590700 269010
rect 590660 268660 590712 268666
rect 590660 268602 590712 268608
rect 591040 268258 591068 277766
rect 591488 271720 591540 271726
rect 591488 271662 591540 271668
rect 591500 271046 591528 271662
rect 591488 271040 591540 271046
rect 591488 270982 591540 270988
rect 593156 270910 593184 277780
rect 594352 273222 594380 277780
rect 594812 277766 595470 277794
rect 594340 273216 594392 273222
rect 594340 273158 594392 273164
rect 593144 270904 593196 270910
rect 593144 270846 593196 270852
rect 594812 268938 594840 277766
rect 596652 271862 596680 277780
rect 597848 274922 597876 277780
rect 599044 277394 599072 277780
rect 598952 277366 599072 277394
rect 597836 274916 597888 274922
rect 597836 274858 597888 274864
rect 598952 274666 598980 277366
rect 598860 274638 598980 274666
rect 596640 271856 596692 271862
rect 596640 271798 596692 271804
rect 594800 268932 594852 268938
rect 594800 268874 594852 268880
rect 598860 268802 598888 274638
rect 600240 271590 600268 277780
rect 601436 274378 601464 277780
rect 601424 274372 601476 274378
rect 601424 274314 601476 274320
rect 602540 274242 602568 277780
rect 602528 274236 602580 274242
rect 602528 274178 602580 274184
rect 603736 271726 603764 277780
rect 604932 276010 604960 277780
rect 604920 276004 604972 276010
rect 604920 275946 604972 275952
rect 606128 272814 606156 277780
rect 606116 272808 606168 272814
rect 606116 272750 606168 272756
rect 603724 271720 603776 271726
rect 603724 271662 603776 271668
rect 600228 271584 600280 271590
rect 600228 271526 600280 271532
rect 607324 270774 607352 277780
rect 607600 277766 608534 277794
rect 608704 277766 609730 277794
rect 607312 270768 607364 270774
rect 607312 270710 607364 270716
rect 607600 269278 607628 277766
rect 607864 271584 607916 271590
rect 607864 271526 607916 271532
rect 607588 269272 607640 269278
rect 607588 269214 607640 269220
rect 598848 268796 598900 268802
rect 598848 268738 598900 268744
rect 591028 268252 591080 268258
rect 591028 268194 591080 268200
rect 587900 268116 587952 268122
rect 587900 268058 587952 268064
rect 607876 267345 607904 271526
rect 608704 268666 608732 277766
rect 610820 271454 610848 277780
rect 612016 275874 612044 277780
rect 612004 275868 612056 275874
rect 612004 275810 612056 275816
rect 611360 275188 611412 275194
rect 611360 275130 611412 275136
rect 611372 272950 611400 275130
rect 613212 273970 613240 277780
rect 613384 274236 613436 274242
rect 613384 274178 613436 274184
rect 613200 273964 613252 273970
rect 613200 273906 613252 273912
rect 611360 272944 611412 272950
rect 611360 272886 611412 272892
rect 610808 271448 610860 271454
rect 610808 271390 610860 271396
rect 608692 268660 608744 268666
rect 608692 268602 608744 268608
rect 607862 267336 607918 267345
rect 607862 267271 607918 267280
rect 585784 267164 585836 267170
rect 585784 267106 585836 267112
rect 580264 266892 580316 266898
rect 580264 266834 580316 266840
rect 613396 266762 613424 274178
rect 614408 272678 614436 277780
rect 615604 274242 615632 277780
rect 616800 275194 616828 277780
rect 616788 275188 616840 275194
rect 616788 275130 616840 275136
rect 615592 274236 615644 274242
rect 615592 274178 615644 274184
rect 614396 272672 614448 272678
rect 614396 272614 614448 272620
rect 617996 271318 618024 277780
rect 619100 275738 619128 277780
rect 619652 277766 620310 277794
rect 619088 275732 619140 275738
rect 619088 275674 619140 275680
rect 619180 275188 619232 275194
rect 619180 275130 619232 275136
rect 619192 274106 619220 275130
rect 619180 274100 619232 274106
rect 619180 274042 619232 274048
rect 617984 271312 618036 271318
rect 617984 271254 618036 271260
rect 619652 268530 619680 277766
rect 621492 271182 621520 277780
rect 622412 277766 622702 277794
rect 621480 271176 621532 271182
rect 621480 271118 621532 271124
rect 621664 271176 621716 271182
rect 621664 271118 621716 271124
rect 619640 268524 619692 268530
rect 619640 268466 619692 268472
rect 621676 267306 621704 271118
rect 621664 267300 621716 267306
rect 621664 267242 621716 267248
rect 622412 267034 622440 277766
rect 623884 275194 623912 277780
rect 623872 275188 623924 275194
rect 623872 275130 623924 275136
rect 625080 271153 625108 277780
rect 626184 275602 626212 277780
rect 626552 277766 627394 277794
rect 627932 277766 628590 277794
rect 629312 277766 629786 277794
rect 630692 277766 630982 277794
rect 626172 275596 626224 275602
rect 626172 275538 626224 275544
rect 625066 271144 625122 271153
rect 625066 271079 625122 271088
rect 626552 270230 626580 277766
rect 626540 270224 626592 270230
rect 626540 270166 626592 270172
rect 627932 270065 627960 277766
rect 627918 270056 627974 270065
rect 627918 269991 627974 270000
rect 629312 267073 629340 277766
rect 630692 269958 630720 277766
rect 632164 272542 632192 277780
rect 633360 275330 633388 277780
rect 633636 277766 634478 277794
rect 633348 275324 633400 275330
rect 633348 275266 633400 275272
rect 632152 272536 632204 272542
rect 632152 272478 632204 272484
rect 633636 270094 633664 277766
rect 635660 273873 635688 277780
rect 635646 273864 635702 273873
rect 635646 273799 635702 273808
rect 636856 271182 636884 277780
rect 637592 277766 638066 277794
rect 638972 277766 639262 277794
rect 636844 271176 636896 271182
rect 636844 271118 636896 271124
rect 633624 270088 633676 270094
rect 633624 270030 633676 270036
rect 630680 269952 630732 269958
rect 630680 269894 630732 269900
rect 637592 269793 637620 277766
rect 637578 269784 637634 269793
rect 637578 269719 637634 269728
rect 638972 268394 639000 277766
rect 640444 273086 640472 277780
rect 641640 275466 641668 277780
rect 641916 277766 642758 277794
rect 641628 275460 641680 275466
rect 641628 275402 641680 275408
rect 640432 273080 640484 273086
rect 640432 273022 640484 273028
rect 641916 269822 641944 277766
rect 643940 271590 643968 277780
rect 645136 272513 645164 277780
rect 645872 277766 646346 277794
rect 647252 277766 647542 277794
rect 645122 272504 645178 272513
rect 645122 272439 645178 272448
rect 643928 271584 643980 271590
rect 643928 271526 643980 271532
rect 641904 269816 641956 269822
rect 641904 269758 641956 269764
rect 638960 268388 639012 268394
rect 638960 268330 639012 268336
rect 629298 267064 629354 267073
rect 622400 267028 622452 267034
rect 629298 266999 629354 267008
rect 622400 266970 622452 266976
rect 613384 266756 613436 266762
rect 613384 266698 613436 266704
rect 575572 265804 575624 265810
rect 575572 265746 575624 265752
rect 554780 265668 554832 265674
rect 554780 265610 554832 265616
rect 558184 265668 558236 265674
rect 558184 265610 558236 265616
rect 554410 262168 554466 262177
rect 554410 262103 554466 262112
rect 554424 260914 554452 262103
rect 554412 260908 554464 260914
rect 554412 260850 554464 260856
rect 554318 259992 554374 260001
rect 554318 259927 554374 259936
rect 554332 259486 554360 259927
rect 554320 259480 554372 259486
rect 554320 259422 554372 259428
rect 553950 257816 554006 257825
rect 553950 257751 554006 257760
rect 553964 256766 553992 257751
rect 553952 256760 554004 256766
rect 553952 256702 554004 256708
rect 553674 255640 553730 255649
rect 553674 255575 553730 255584
rect 553490 251288 553546 251297
rect 553490 251223 553492 251232
rect 553544 251223 553546 251232
rect 553492 251194 553544 251200
rect 553688 249082 553716 255575
rect 554502 253464 554558 253473
rect 554502 253399 554504 253408
rect 554556 253399 554558 253408
rect 554504 253370 554556 253376
rect 555424 251252 555476 251258
rect 555424 251194 555476 251200
rect 553858 249112 553914 249121
rect 553676 249076 553728 249082
rect 553858 249047 553914 249056
rect 553676 249018 553728 249024
rect 553872 246362 553900 249047
rect 554410 246936 554466 246945
rect 554410 246871 554466 246880
rect 553860 246356 553912 246362
rect 553860 246298 553912 246304
rect 554424 245682 554452 246871
rect 554412 245676 554464 245682
rect 554412 245618 554464 245624
rect 554502 244760 554558 244769
rect 554502 244695 554558 244704
rect 554516 244322 554544 244695
rect 554504 244316 554556 244322
rect 554504 244258 554556 244264
rect 553950 242584 554006 242593
rect 553950 242519 554006 242528
rect 553964 241534 553992 242519
rect 553952 241528 554004 241534
rect 553952 241470 554004 241476
rect 553858 240408 553914 240417
rect 553858 240343 553914 240352
rect 553872 240174 553900 240343
rect 553860 240168 553912 240174
rect 553860 240110 553912 240116
rect 554320 238740 554372 238746
rect 554320 238682 554372 238688
rect 554332 238241 554360 238682
rect 554318 238232 554374 238241
rect 554318 238167 554374 238176
rect 554504 236088 554556 236094
rect 554502 236056 554504 236065
rect 554556 236056 554558 236065
rect 554502 235991 554558 236000
rect 554412 234592 554464 234598
rect 554412 234534 554464 234540
rect 554424 233889 554452 234534
rect 554410 233880 554466 233889
rect 554410 233815 554466 233824
rect 140792 231662 141174 231690
rect 141528 231662 141818 231690
rect 90364 230444 90416 230450
rect 90364 230386 90416 230392
rect 88248 230036 88300 230042
rect 88248 229978 88300 229984
rect 74448 229900 74500 229906
rect 74448 229842 74500 229848
rect 67548 229764 67600 229770
rect 67548 229706 67600 229712
rect 66168 228404 66220 228410
rect 66168 228346 66220 228352
rect 64788 225752 64840 225758
rect 64788 225694 64840 225700
rect 62946 222864 63002 222873
rect 62946 222799 63002 222808
rect 64604 221468 64656 221474
rect 64604 221410 64656 221416
rect 63132 220108 63184 220114
rect 63132 220050 63184 220056
rect 62764 218204 62816 218210
rect 62764 218146 62816 218152
rect 63144 217274 63172 220050
rect 64616 219434 64644 221410
rect 64800 219434 64828 225694
rect 63960 219428 64012 219434
rect 64616 219406 64736 219434
rect 64800 219428 64932 219434
rect 64800 219406 64880 219428
rect 63960 219370 64012 219376
rect 62270 217110 62344 217138
rect 63098 217246 63172 217274
rect 62270 216988 62298 217110
rect 63098 216988 63126 217246
rect 63972 217138 64000 219370
rect 64708 217274 64736 219406
rect 64880 219370 64932 219376
rect 66180 218074 66208 228346
rect 66444 220244 66496 220250
rect 66444 220186 66496 220192
rect 65616 218068 65668 218074
rect 65616 218010 65668 218016
rect 66168 218068 66220 218074
rect 66168 218010 66220 218016
rect 64708 217246 64782 217274
rect 63926 217110 64000 217138
rect 63926 216988 63954 217110
rect 64754 216988 64782 217246
rect 65628 217138 65656 218010
rect 66456 217274 66484 220186
rect 67560 219434 67588 229706
rect 73066 226944 73122 226953
rect 73066 226879 73122 226888
rect 69572 226160 69624 226166
rect 69572 226102 69624 226108
rect 68926 224224 68982 224233
rect 68926 224159 68982 224168
rect 68100 221740 68152 221746
rect 68100 221682 68152 221688
rect 67284 219406 67588 219434
rect 67284 217274 67312 219406
rect 68112 217274 68140 221682
rect 68940 217274 68968 224159
rect 69584 218618 69612 226102
rect 71412 221876 71464 221882
rect 71412 221818 71464 221824
rect 69754 220144 69810 220153
rect 69754 220079 69810 220088
rect 69572 218612 69624 218618
rect 69572 218554 69624 218560
rect 69768 217274 69796 220079
rect 70584 219020 70636 219026
rect 70584 218962 70636 218968
rect 65582 217110 65656 217138
rect 66410 217246 66484 217274
rect 67238 217246 67312 217274
rect 68066 217246 68140 217274
rect 68894 217246 68968 217274
rect 69722 217246 69796 217274
rect 65582 216988 65610 217110
rect 66410 216988 66438 217246
rect 67238 216988 67266 217246
rect 68066 216988 68094 217246
rect 68894 216988 68922 217246
rect 69722 216988 69750 217246
rect 70596 217138 70624 218962
rect 71424 217274 71452 221818
rect 72882 220416 72938 220425
rect 72882 220351 72938 220360
rect 72896 219434 72924 220351
rect 73080 219434 73108 226879
rect 72240 219428 72292 219434
rect 72896 219406 73016 219434
rect 73080 219428 73212 219434
rect 73080 219406 73160 219428
rect 72240 219370 72292 219376
rect 70550 217110 70624 217138
rect 71378 217246 71452 217274
rect 70550 216988 70578 217110
rect 71378 216988 71406 217246
rect 72252 217138 72280 219370
rect 72988 217274 73016 219406
rect 73160 219370 73212 219376
rect 74460 218074 74488 229842
rect 82084 228676 82136 228682
rect 82084 228618 82136 228624
rect 79966 228304 80022 228313
rect 79966 228239 80022 228248
rect 75828 227180 75880 227186
rect 75828 227122 75880 227128
rect 75552 218340 75604 218346
rect 75552 218282 75604 218288
rect 73896 218068 73948 218074
rect 73896 218010 73948 218016
rect 74448 218068 74500 218074
rect 74448 218010 74500 218016
rect 74724 218068 74776 218074
rect 74724 218010 74776 218016
rect 72988 217246 73062 217274
rect 72206 217110 72280 217138
rect 72206 216988 72234 217110
rect 73034 216988 73062 217246
rect 73908 217138 73936 218010
rect 74736 217138 74764 218010
rect 75564 217138 75592 218282
rect 75840 218074 75868 227122
rect 76564 223984 76616 223990
rect 76564 223926 76616 223932
rect 76380 220380 76432 220386
rect 76380 220322 76432 220328
rect 75828 218068 75880 218074
rect 75828 218010 75880 218016
rect 76392 217274 76420 220322
rect 76576 218890 76604 223926
rect 78588 223168 78640 223174
rect 78588 223110 78640 223116
rect 76564 218884 76616 218890
rect 76564 218826 76616 218832
rect 77208 218748 77260 218754
rect 77208 218690 77260 218696
rect 73862 217110 73936 217138
rect 74690 217110 74764 217138
rect 75518 217110 75592 217138
rect 76346 217246 76420 217274
rect 73862 216988 73890 217110
rect 74690 216988 74718 217110
rect 75518 216988 75546 217110
rect 76346 216988 76374 217246
rect 77220 217138 77248 218690
rect 78600 218074 78628 223110
rect 79692 218204 79744 218210
rect 79692 218146 79744 218152
rect 78036 218068 78088 218074
rect 78036 218010 78088 218016
rect 78588 218068 78640 218074
rect 78588 218010 78640 218016
rect 78864 218068 78916 218074
rect 78864 218010 78916 218016
rect 78048 217138 78076 218010
rect 78876 217138 78904 218010
rect 79704 217138 79732 218146
rect 79980 218074 80008 228239
rect 81348 223304 81400 223310
rect 81348 223246 81400 223252
rect 80520 219428 80572 219434
rect 80520 219370 80572 219376
rect 79968 218068 80020 218074
rect 79968 218010 80020 218016
rect 80532 217138 80560 219370
rect 81360 217274 81388 223246
rect 82096 218210 82124 228618
rect 86868 227316 86920 227322
rect 86868 227258 86920 227264
rect 83464 226296 83516 226302
rect 83464 226238 83516 226244
rect 82728 224392 82780 224398
rect 82728 224334 82780 224340
rect 82084 218204 82136 218210
rect 82084 218146 82136 218152
rect 82740 218074 82768 224334
rect 83004 220516 83056 220522
rect 83004 220458 83056 220464
rect 82176 218068 82228 218074
rect 82176 218010 82228 218016
rect 82728 218068 82780 218074
rect 82728 218010 82780 218016
rect 77174 217110 77248 217138
rect 78002 217110 78076 217138
rect 78830 217110 78904 217138
rect 79658 217110 79732 217138
rect 80486 217110 80560 217138
rect 81314 217246 81388 217274
rect 77174 216988 77202 217110
rect 78002 216988 78030 217110
rect 78830 216988 78858 217110
rect 79658 216988 79686 217110
rect 80486 216988 80514 217110
rect 81314 216988 81342 217246
rect 82188 217138 82216 218010
rect 83016 217274 83044 220458
rect 83476 218346 83504 226238
rect 85488 223576 85540 223582
rect 85488 223518 85540 223524
rect 85304 219156 85356 219162
rect 85304 219098 85356 219104
rect 83832 218884 83884 218890
rect 83832 218826 83884 218832
rect 83464 218340 83516 218346
rect 83464 218282 83516 218288
rect 82142 217110 82216 217138
rect 82970 217246 83044 217274
rect 82142 216988 82170 217110
rect 82970 216988 82998 217246
rect 83844 217138 83872 218826
rect 84660 218068 84712 218074
rect 84660 218010 84712 218016
rect 84672 217138 84700 218010
rect 85316 217274 85344 219098
rect 85500 218074 85528 223518
rect 86880 218074 86908 227258
rect 87972 222760 88024 222766
rect 87972 222702 88024 222708
rect 85488 218068 85540 218074
rect 85488 218010 85540 218016
rect 86316 218068 86368 218074
rect 86316 218010 86368 218016
rect 86868 218068 86920 218074
rect 86868 218010 86920 218016
rect 87144 218068 87196 218074
rect 87144 218010 87196 218016
rect 85316 217246 85482 217274
rect 83798 217110 83872 217138
rect 84626 217110 84700 217138
rect 83798 216988 83826 217110
rect 84626 216988 84654 217110
rect 85454 216988 85482 217246
rect 86328 217138 86356 218010
rect 87156 217138 87184 218010
rect 87984 217274 88012 222702
rect 88260 218074 88288 229978
rect 90376 229094 90404 230386
rect 118424 230308 118476 230314
rect 118424 230250 118476 230256
rect 111064 230172 111116 230178
rect 111064 230114 111116 230120
rect 103610 229800 103666 229809
rect 103610 229735 103666 229744
rect 92480 229220 92532 229226
rect 92480 229162 92532 229168
rect 90284 229066 90404 229094
rect 89628 227452 89680 227458
rect 89628 227394 89680 227400
rect 89444 223032 89496 223038
rect 89444 222974 89496 222980
rect 89456 218074 89484 222974
rect 88248 218068 88300 218074
rect 88248 218010 88300 218016
rect 88800 218068 88852 218074
rect 88800 218010 88852 218016
rect 89444 218068 89496 218074
rect 89444 218010 89496 218016
rect 86282 217110 86356 217138
rect 87110 217110 87184 217138
rect 87938 217246 88012 217274
rect 86282 216988 86310 217110
rect 87110 216988 87138 217110
rect 87938 216988 87966 217246
rect 88812 217138 88840 218010
rect 89640 217274 89668 227394
rect 90284 219434 90312 229066
rect 92492 225758 92520 229162
rect 97908 229084 97960 229090
rect 97908 229026 97960 229032
rect 96252 228676 96304 228682
rect 96252 228618 96304 228624
rect 93768 226024 93820 226030
rect 93768 225966 93820 225972
rect 92480 225752 92532 225758
rect 92480 225694 92532 225700
rect 92112 222896 92164 222902
rect 92112 222838 92164 222844
rect 91284 220788 91336 220794
rect 91284 220730 91336 220736
rect 90272 219428 90324 219434
rect 90272 219370 90324 219376
rect 90456 219428 90508 219434
rect 90456 219370 90508 219376
rect 88766 217110 88840 217138
rect 89594 217246 89668 217274
rect 88766 216988 88794 217110
rect 89594 216988 89622 217246
rect 90468 217138 90496 219370
rect 91296 217274 91324 220730
rect 92124 217274 92152 222838
rect 93780 218618 93808 225966
rect 95148 225888 95200 225894
rect 95148 225830 95200 225836
rect 92940 218612 92992 218618
rect 92940 218554 92992 218560
rect 93768 218612 93820 218618
rect 93768 218554 93820 218560
rect 90422 217110 90496 217138
rect 91250 217246 91324 217274
rect 92078 217246 92152 217274
rect 90422 216988 90450 217110
rect 91250 216988 91278 217246
rect 92078 216988 92106 217246
rect 92952 217138 92980 218554
rect 93768 218476 93820 218482
rect 93768 218418 93820 218424
rect 93780 217138 93808 218418
rect 95160 218074 95188 225830
rect 95424 221332 95476 221338
rect 95424 221274 95476 221280
rect 94596 218068 94648 218074
rect 94596 218010 94648 218016
rect 95148 218068 95200 218074
rect 95148 218010 95200 218016
rect 94608 217138 94636 218010
rect 95436 217274 95464 221274
rect 96264 217274 96292 228618
rect 97724 220652 97776 220658
rect 97724 220594 97776 220600
rect 97736 219434 97764 220594
rect 97736 219406 97856 219434
rect 97080 218068 97132 218074
rect 97080 218010 97132 218016
rect 92906 217110 92980 217138
rect 93734 217110 93808 217138
rect 94562 217110 94636 217138
rect 95390 217246 95464 217274
rect 96218 217246 96292 217274
rect 92906 216988 92934 217110
rect 93734 216988 93762 217110
rect 94562 216988 94590 217110
rect 95390 216988 95418 217246
rect 96218 216988 96246 217246
rect 97092 217138 97120 218010
rect 97828 217274 97856 219406
rect 97920 218090 97948 229026
rect 102048 228948 102100 228954
rect 102048 228890 102100 228896
rect 100668 227588 100720 227594
rect 100668 227530 100720 227536
rect 99288 222624 99340 222630
rect 99288 222566 99340 222572
rect 97920 218074 98040 218090
rect 99300 218074 99328 222566
rect 100392 218340 100444 218346
rect 100392 218282 100444 218288
rect 97920 218068 98052 218074
rect 97920 218062 98000 218068
rect 98000 218010 98052 218016
rect 98736 218068 98788 218074
rect 98736 218010 98788 218016
rect 99288 218068 99340 218074
rect 99288 218010 99340 218016
rect 99564 218068 99616 218074
rect 99564 218010 99616 218016
rect 97828 217246 97902 217274
rect 97046 217110 97120 217138
rect 97046 216988 97074 217110
rect 97874 216988 97902 217246
rect 98748 217138 98776 218010
rect 99576 217138 99604 218010
rect 100404 217138 100432 218282
rect 100680 218074 100708 227530
rect 101862 221504 101918 221513
rect 101862 221439 101918 221448
rect 101876 219434 101904 221439
rect 101876 219406 101996 219434
rect 100668 218068 100720 218074
rect 100668 218010 100720 218016
rect 101220 218068 101272 218074
rect 101220 218010 101272 218016
rect 101232 217138 101260 218010
rect 101968 217274 101996 219406
rect 102060 218090 102088 228890
rect 103428 225480 103480 225486
rect 103428 225422 103480 225428
rect 102060 218074 102180 218090
rect 103440 218074 103468 225422
rect 103624 224534 103652 229735
rect 107292 229084 107344 229090
rect 107292 229026 107344 229032
rect 107476 229084 107528 229090
rect 107476 229026 107528 229032
rect 107304 228818 107332 229026
rect 107108 228812 107160 228818
rect 107108 228754 107160 228760
rect 107292 228812 107344 228818
rect 107292 228754 107344 228760
rect 107120 228274 107148 228754
rect 107108 228268 107160 228274
rect 107108 228210 107160 228216
rect 107488 228138 107516 229026
rect 106188 228132 106240 228138
rect 106188 228074 106240 228080
rect 107476 228132 107528 228138
rect 107476 228074 107528 228080
rect 106004 225344 106056 225350
rect 106004 225286 106056 225292
rect 103612 224528 103664 224534
rect 103612 224470 103664 224476
rect 104808 224120 104860 224126
rect 104808 224062 104860 224068
rect 104532 222012 104584 222018
rect 104532 221954 104584 221960
rect 102060 218068 102192 218074
rect 102060 218062 102140 218068
rect 102140 218010 102192 218016
rect 102876 218068 102928 218074
rect 102876 218010 102928 218016
rect 103428 218068 103480 218074
rect 103428 218010 103480 218016
rect 103704 218068 103756 218074
rect 103704 218010 103756 218016
rect 101968 217246 102042 217274
rect 98702 217110 98776 217138
rect 99530 217110 99604 217138
rect 100358 217110 100432 217138
rect 101186 217110 101260 217138
rect 98702 216988 98730 217110
rect 99530 216988 99558 217110
rect 100358 216988 100386 217110
rect 101186 216988 101214 217110
rect 102014 216988 102042 217246
rect 102888 217138 102916 218010
rect 103716 217138 103744 218010
rect 104544 217274 104572 221954
rect 104820 218074 104848 224062
rect 105820 219496 105872 219502
rect 105820 219438 105872 219444
rect 105832 218346 105860 219438
rect 105820 218340 105872 218346
rect 105820 218282 105872 218288
rect 106016 218074 106044 225286
rect 104808 218068 104860 218074
rect 104808 218010 104860 218016
rect 105360 218068 105412 218074
rect 105360 218010 105412 218016
rect 106004 218068 106056 218074
rect 106004 218010 106056 218016
rect 102842 217110 102916 217138
rect 103670 217110 103744 217138
rect 104498 217246 104572 217274
rect 102842 216988 102870 217110
rect 103670 216988 103698 217110
rect 104498 216988 104526 217246
rect 105372 217138 105400 218010
rect 106200 217274 106228 228074
rect 110144 227724 110196 227730
rect 110144 227666 110196 227672
rect 106924 226908 106976 226914
rect 106924 226850 106976 226856
rect 106936 219298 106964 226850
rect 108304 225752 108356 225758
rect 108304 225694 108356 225700
rect 108316 225486 108344 225694
rect 108304 225480 108356 225486
rect 108304 225422 108356 225428
rect 108672 224528 108724 224534
rect 108672 224470 108724 224476
rect 107844 222148 107896 222154
rect 107844 222090 107896 222096
rect 106924 219292 106976 219298
rect 106924 219234 106976 219240
rect 107016 218476 107068 218482
rect 107016 218418 107068 218424
rect 105326 217110 105400 217138
rect 106154 217246 106228 217274
rect 105326 216988 105354 217110
rect 106154 216988 106182 217246
rect 107028 217138 107056 218418
rect 107856 217274 107884 222090
rect 108684 217274 108712 224470
rect 110156 218074 110184 227666
rect 111076 219434 111104 230114
rect 112996 228132 113048 228138
rect 112996 228074 113048 228080
rect 112812 223440 112864 223446
rect 112812 223382 112864 223388
rect 111248 219972 111300 219978
rect 111248 219914 111300 219920
rect 111260 219434 111288 219914
rect 110984 219406 111104 219434
rect 111168 219406 111288 219434
rect 110984 218074 111012 219406
rect 109500 218068 109552 218074
rect 109500 218010 109552 218016
rect 110144 218068 110196 218074
rect 110144 218010 110196 218016
rect 110328 218068 110380 218074
rect 110328 218010 110380 218016
rect 110972 218068 111024 218074
rect 110972 218010 111024 218016
rect 106982 217110 107056 217138
rect 107810 217246 107884 217274
rect 108638 217246 108712 217274
rect 106982 216988 107010 217110
rect 107810 216988 107838 217246
rect 108638 216988 108666 217246
rect 109512 217138 109540 218010
rect 110340 217138 110368 218010
rect 111168 217274 111196 219406
rect 112824 218074 112852 223382
rect 111984 218068 112036 218074
rect 111984 218010 112036 218016
rect 112812 218068 112864 218074
rect 112812 218010 112864 218016
rect 109466 217110 109540 217138
rect 110294 217110 110368 217138
rect 111122 217246 111196 217274
rect 109466 216988 109494 217110
rect 110294 216988 110322 217110
rect 111122 216988 111150 217246
rect 111996 217138 112024 218010
rect 113008 217274 113036 228074
rect 117228 225344 117280 225350
rect 117228 225286 117280 225292
rect 115848 224800 115900 224806
rect 115848 224742 115900 224748
rect 114468 221332 114520 221338
rect 114468 221274 114520 221280
rect 113640 218340 113692 218346
rect 113640 218282 113692 218288
rect 111950 217110 112024 217138
rect 112778 217246 113036 217274
rect 111950 216988 111978 217110
rect 112778 216988 112806 217246
rect 113652 217138 113680 218282
rect 114480 217274 114508 221274
rect 115860 218074 115888 224742
rect 116768 224664 116820 224670
rect 116768 224606 116820 224612
rect 116780 224262 116808 224606
rect 116768 224256 116820 224262
rect 116768 224198 116820 224204
rect 116952 224256 117004 224262
rect 116952 224198 117004 224204
rect 115296 218068 115348 218074
rect 115296 218010 115348 218016
rect 115848 218068 115900 218074
rect 115848 218010 115900 218016
rect 116124 218068 116176 218074
rect 116124 218010 116176 218016
rect 113606 217110 113680 217138
rect 114434 217246 114508 217274
rect 113606 216988 113634 217110
rect 114434 216988 114462 217246
rect 115308 217138 115336 218010
rect 116136 217138 116164 218010
rect 116964 217274 116992 224198
rect 117240 218074 117268 225286
rect 118148 224664 118200 224670
rect 118148 224606 118200 224612
rect 118160 224126 118188 224606
rect 118436 224262 118464 230250
rect 140044 229628 140096 229634
rect 140044 229570 140096 229576
rect 131120 229492 131172 229498
rect 131120 229434 131172 229440
rect 122932 229356 122984 229362
rect 122932 229298 122984 229304
rect 122748 227996 122800 228002
rect 122748 227938 122800 227944
rect 121092 226772 121144 226778
rect 121092 226714 121144 226720
rect 119988 226636 120040 226642
rect 119988 226578 120040 226584
rect 118792 224800 118844 224806
rect 118792 224742 118844 224748
rect 118608 224528 118660 224534
rect 118608 224470 118660 224476
rect 118620 224262 118648 224470
rect 118424 224256 118476 224262
rect 118424 224198 118476 224204
rect 118608 224256 118660 224262
rect 118608 224198 118660 224204
rect 117964 224120 118016 224126
rect 117964 224062 118016 224068
rect 118148 224120 118200 224126
rect 118804 224074 118832 224742
rect 118148 224062 118200 224068
rect 117976 223854 118004 224062
rect 118620 224046 118832 224074
rect 117964 223848 118016 223854
rect 117964 223790 118016 223796
rect 117780 221060 117832 221066
rect 117780 221002 117832 221008
rect 117228 218068 117280 218074
rect 117228 218010 117280 218016
rect 117792 217274 117820 221002
rect 117964 219428 118016 219434
rect 117964 219370 118016 219376
rect 117976 219162 118004 219370
rect 117964 219156 118016 219162
rect 117964 219098 118016 219104
rect 118620 217274 118648 224046
rect 120000 218074 120028 226578
rect 120264 218204 120316 218210
rect 120264 218146 120316 218152
rect 119436 218068 119488 218074
rect 119436 218010 119488 218016
rect 119988 218068 120040 218074
rect 119988 218010 120040 218016
rect 115262 217110 115336 217138
rect 116090 217110 116164 217138
rect 116918 217246 116992 217274
rect 117746 217246 117820 217274
rect 118574 217246 118648 217274
rect 115262 216988 115290 217110
rect 116090 216988 116118 217110
rect 116918 216988 116946 217246
rect 117746 216988 117774 217246
rect 118574 216988 118602 217246
rect 119448 217138 119476 218010
rect 120276 217138 120304 218146
rect 121104 217274 121132 226714
rect 122564 224936 122616 224942
rect 122564 224878 122616 224884
rect 122576 218074 122604 224878
rect 121920 218068 121972 218074
rect 121920 218010 121972 218016
rect 122564 218068 122616 218074
rect 122564 218010 122616 218016
rect 119402 217110 119476 217138
rect 120230 217110 120304 217138
rect 121058 217246 121132 217274
rect 119402 216988 119430 217110
rect 120230 216988 120258 217110
rect 121058 216988 121086 217246
rect 121932 217138 121960 218010
rect 122760 217274 122788 227938
rect 122944 223854 122972 229298
rect 125784 226908 125836 226914
rect 125784 226850 125836 226856
rect 125796 226506 125824 226850
rect 125784 226500 125836 226506
rect 125784 226442 125836 226448
rect 129372 226500 129424 226506
rect 129372 226442 129424 226448
rect 127440 225480 127492 225486
rect 127440 225422 127492 225428
rect 127452 225214 127480 225422
rect 127440 225208 127492 225214
rect 127440 225150 127492 225156
rect 128268 225208 128320 225214
rect 128268 225150 128320 225156
rect 126888 225072 126940 225078
rect 126888 225014 126940 225020
rect 126704 224528 126756 224534
rect 126704 224470 126756 224476
rect 122932 223848 122984 223854
rect 122932 223790 122984 223796
rect 125232 223848 125284 223854
rect 125232 223790 125284 223796
rect 123482 222864 123538 222873
rect 123482 222799 123538 222808
rect 123496 219434 123524 222799
rect 124404 219836 124456 219842
rect 124404 219778 124456 219784
rect 123484 219428 123536 219434
rect 123484 219370 123536 219376
rect 123576 219156 123628 219162
rect 123576 219098 123628 219104
rect 121886 217110 121960 217138
rect 122714 217246 122788 217274
rect 121886 216988 121914 217110
rect 122714 216988 122742 217246
rect 123588 217138 123616 219098
rect 124416 217274 124444 219778
rect 125244 217274 125272 223790
rect 126716 219434 126744 224470
rect 126900 219434 126928 225014
rect 126060 219428 126112 219434
rect 126716 219406 126836 219434
rect 126900 219428 127032 219434
rect 126900 219406 126980 219428
rect 126060 219370 126112 219376
rect 123542 217110 123616 217138
rect 124370 217246 124444 217274
rect 125198 217246 125272 217274
rect 123542 216988 123570 217110
rect 124370 216988 124398 217246
rect 125198 216988 125226 217246
rect 126072 217138 126100 219370
rect 126808 217274 126836 219406
rect 126980 219370 127032 219376
rect 128280 218210 128308 225150
rect 128544 220924 128596 220930
rect 128544 220866 128596 220872
rect 127716 218204 127768 218210
rect 127716 218146 127768 218152
rect 128268 218204 128320 218210
rect 128268 218146 128320 218152
rect 126808 217246 126882 217274
rect 126026 217110 126100 217138
rect 126026 216988 126054 217110
rect 126854 216988 126882 217246
rect 127728 217138 127756 218146
rect 128556 217274 128584 220866
rect 128728 219156 128780 219162
rect 128728 219098 128780 219104
rect 128740 218346 128768 219098
rect 128728 218340 128780 218346
rect 128728 218282 128780 218288
rect 129384 217274 129412 226442
rect 131132 224534 131160 229434
rect 140056 229094 140084 229570
rect 139964 229066 140084 229094
rect 135166 228032 135222 228041
rect 135166 227967 135222 227976
rect 133788 227860 133840 227866
rect 133788 227802 133840 227808
rect 131120 224528 131172 224534
rect 131120 224470 131172 224476
rect 131304 224528 131356 224534
rect 131304 224470 131356 224476
rect 131316 223854 131344 224470
rect 131304 223848 131356 223854
rect 131304 223790 131356 223796
rect 132408 223712 132460 223718
rect 132408 223654 132460 223660
rect 131028 219700 131080 219706
rect 131028 219642 131080 219648
rect 130200 219428 130252 219434
rect 130200 219370 130252 219376
rect 127682 217110 127756 217138
rect 128510 217246 128584 217274
rect 129338 217246 129412 217274
rect 127682 216988 127710 217110
rect 128510 216988 128538 217246
rect 129338 216988 129366 217246
rect 130212 217138 130240 219370
rect 131040 217274 131068 219642
rect 132420 219162 132448 223654
rect 133512 222488 133564 222494
rect 133512 222430 133564 222436
rect 131856 219156 131908 219162
rect 131856 219098 131908 219104
rect 132408 219156 132460 219162
rect 132408 219098 132460 219104
rect 130166 217110 130240 217138
rect 130994 217246 131068 217274
rect 130166 216988 130194 217110
rect 130994 216988 131022 217246
rect 131868 217138 131896 219098
rect 132776 219020 132828 219026
rect 132776 218962 132828 218968
rect 132788 217274 132816 218962
rect 133524 217274 133552 222430
rect 133800 219026 133828 227802
rect 134984 227044 135036 227050
rect 134984 226986 135036 226992
rect 134996 226681 135024 226986
rect 134982 226672 135038 226681
rect 134982 226607 135038 226616
rect 134984 223848 135036 223854
rect 134984 223790 135036 223796
rect 134996 219434 135024 223790
rect 135180 219434 135208 227967
rect 135444 227044 135496 227050
rect 135444 226986 135496 226992
rect 135456 226642 135484 226986
rect 135626 226672 135682 226681
rect 135444 226636 135496 226642
rect 135626 226607 135628 226616
rect 135444 226578 135496 226584
rect 135680 226607 135682 226616
rect 137560 226636 137612 226642
rect 135628 226578 135680 226584
rect 137560 226578 137612 226584
rect 137572 226522 137600 226578
rect 137204 226506 137600 226522
rect 137192 226500 137600 226506
rect 137244 226494 137600 226500
rect 139306 226536 139362 226545
rect 139306 226471 139362 226480
rect 137192 226442 137244 226448
rect 136836 226222 137692 226250
rect 136546 226128 136602 226137
rect 136546 226063 136602 226072
rect 134156 219428 134208 219434
rect 134156 219370 134208 219376
rect 134340 219428 134392 219434
rect 134996 219406 135116 219434
rect 135180 219428 135312 219434
rect 135180 219406 135260 219428
rect 134340 219370 134392 219376
rect 134168 219162 134196 219370
rect 134156 219156 134208 219162
rect 134156 219098 134208 219104
rect 133788 219020 133840 219026
rect 133788 218962 133840 218968
rect 131822 217110 131896 217138
rect 132650 217246 132816 217274
rect 133478 217246 133552 217274
rect 131822 216988 131850 217110
rect 132650 216988 132678 217246
rect 133478 216988 133506 217246
rect 134352 217138 134380 219370
rect 135088 217274 135116 219406
rect 135260 219370 135312 219376
rect 135812 219428 135864 219434
rect 135812 219370 135864 219376
rect 135824 219026 135852 219370
rect 136560 219026 136588 226063
rect 136836 225622 136864 226222
rect 137664 226166 137692 226222
rect 137468 226160 137520 226166
rect 137468 226102 137520 226108
rect 137652 226160 137704 226166
rect 137652 226102 137704 226108
rect 136824 225616 136876 225622
rect 136824 225558 136876 225564
rect 137008 225616 137060 225622
rect 137008 225558 137060 225564
rect 137020 225350 137048 225558
rect 137008 225344 137060 225350
rect 137008 225286 137060 225292
rect 137480 225078 137508 226102
rect 137468 225072 137520 225078
rect 137468 225014 137520 225020
rect 137284 221604 137336 221610
rect 137284 221546 137336 221552
rect 137468 221604 137520 221610
rect 137468 221546 137520 221552
rect 137296 221202 137324 221546
rect 137100 221196 137152 221202
rect 137100 221138 137152 221144
rect 137284 221196 137336 221202
rect 137284 221138 137336 221144
rect 137112 221082 137140 221138
rect 137480 221082 137508 221546
rect 138478 221232 138534 221241
rect 138478 221167 138534 221176
rect 137112 221054 137508 221082
rect 137652 219564 137704 219570
rect 137652 219506 137704 219512
rect 136916 219156 136968 219162
rect 136916 219098 136968 219104
rect 135812 219020 135864 219026
rect 135812 218962 135864 218968
rect 135996 219020 136048 219026
rect 135996 218962 136048 218968
rect 136548 219020 136600 219026
rect 136548 218962 136600 218968
rect 135088 217246 135162 217274
rect 134306 217110 134380 217138
rect 134306 216988 134334 217110
rect 135134 216988 135162 217246
rect 136008 217138 136036 218962
rect 136928 217274 136956 219098
rect 137664 217274 137692 219506
rect 138492 217274 138520 221167
rect 139320 217274 139348 226471
rect 139964 219434 139992 229066
rect 140792 228546 140820 231662
rect 140780 228540 140832 228546
rect 140780 228482 140832 228488
rect 140964 228540 141016 228546
rect 140964 228482 141016 228488
rect 140976 228274 141004 228482
rect 140964 228268 141016 228274
rect 140964 228210 141016 228216
rect 141148 228268 141200 228274
rect 141148 228210 141200 228216
rect 141160 228041 141188 228210
rect 141146 228032 141202 228041
rect 141146 227967 141202 227976
rect 141528 226166 141556 231662
rect 142158 227216 142214 227225
rect 142158 227151 142214 227160
rect 142172 226658 142200 227151
rect 142126 226630 142200 226658
rect 142126 226506 142154 226630
rect 142250 226536 142306 226545
rect 142114 226500 142166 226506
rect 142250 226471 142252 226480
rect 142114 226442 142166 226448
rect 142304 226471 142306 226480
rect 142252 226442 142304 226448
rect 142448 226386 142476 231676
rect 143092 227225 143120 231676
rect 143552 231662 143750 231690
rect 144012 231662 144394 231690
rect 145038 231662 145236 231690
rect 143078 227216 143134 227225
rect 143078 227151 143134 227160
rect 142356 226358 142476 226386
rect 141516 226160 141568 226166
rect 141700 226160 141752 226166
rect 141516 226102 141568 226108
rect 141698 226128 141700 226137
rect 141752 226128 141754 226137
rect 141698 226063 141754 226072
rect 142158 224632 142214 224641
rect 142158 224567 142214 224576
rect 142172 223990 142200 224567
rect 142160 223984 142212 223990
rect 141790 223952 141846 223961
rect 142160 223926 142212 223932
rect 141790 223887 141846 223896
rect 140778 219600 140834 219609
rect 140778 219535 140780 219544
rect 140832 219535 140834 219544
rect 140964 219564 141016 219570
rect 140780 219506 140832 219512
rect 140964 219506 141016 219512
rect 139952 219428 140004 219434
rect 139952 219370 140004 219376
rect 140136 219428 140188 219434
rect 140136 219370 140188 219376
rect 135962 217110 136036 217138
rect 136790 217246 136956 217274
rect 137618 217246 137692 217274
rect 138446 217246 138520 217274
rect 139274 217246 139348 217274
rect 135962 216988 135990 217110
rect 136790 216988 136818 217246
rect 137618 216988 137646 217246
rect 138446 216988 138474 217246
rect 139274 216988 139302 217246
rect 140148 217138 140176 219370
rect 140976 217274 141004 219506
rect 141804 217274 141832 223887
rect 142356 222358 142384 226358
rect 143170 225584 143226 225593
rect 143170 225519 143226 225528
rect 142620 224120 142672 224126
rect 142620 224062 142672 224068
rect 142632 223961 142660 224062
rect 142618 223952 142674 223961
rect 142618 223887 142674 223896
rect 142988 222488 143040 222494
rect 142986 222456 142988 222465
rect 143040 222456 143042 222465
rect 142986 222391 143042 222400
rect 142344 222352 142396 222358
rect 142344 222294 142396 222300
rect 142158 221912 142214 221921
rect 142158 221847 142214 221856
rect 142172 221762 142200 221847
rect 142126 221746 142200 221762
rect 142114 221740 142200 221746
rect 142166 221734 142200 221740
rect 142344 221740 142396 221746
rect 142114 221682 142166 221688
rect 142344 221682 142396 221688
rect 142356 221626 142384 221682
rect 142126 221598 142384 221626
rect 142126 221474 142154 221598
rect 142114 221468 142166 221474
rect 142114 221410 142166 221416
rect 142252 221468 142304 221474
rect 142252 221410 142304 221416
rect 142264 221354 142292 221410
rect 142126 221326 142292 221354
rect 142126 221202 142154 221326
rect 142250 221232 142306 221241
rect 142114 221196 142166 221202
rect 142250 221167 142252 221176
rect 142114 221138 142166 221144
rect 142304 221167 142306 221176
rect 142252 221138 142304 221144
rect 142158 220824 142214 220833
rect 142158 220759 142214 220768
rect 142172 220402 142200 220759
rect 142126 220374 142200 220402
rect 142126 220250 142154 220374
rect 142114 220244 142166 220250
rect 142114 220186 142166 220192
rect 142252 220244 142304 220250
rect 142252 220186 142304 220192
rect 142264 219881 142292 220186
rect 141974 219872 142030 219881
rect 141974 219807 142030 219816
rect 142250 219872 142306 219881
rect 142250 219807 142306 219816
rect 141988 219570 142016 219807
rect 142158 219600 142214 219609
rect 141976 219564 142028 219570
rect 142158 219535 142160 219544
rect 141976 219506 142028 219512
rect 142212 219535 142214 219544
rect 142160 219506 142212 219512
rect 142250 218784 142306 218793
rect 142250 218719 142252 218728
rect 142304 218719 142306 218728
rect 142252 218690 142304 218696
rect 143184 218618 143212 225519
rect 143552 225078 143580 231662
rect 143540 225072 143592 225078
rect 143540 225014 143592 225020
rect 143356 222488 143408 222494
rect 143356 222430 143408 222436
rect 142620 218612 142672 218618
rect 142620 218554 142672 218560
rect 143172 218612 143224 218618
rect 143172 218554 143224 218560
rect 140102 217110 140176 217138
rect 140930 217246 141004 217274
rect 141758 217246 141832 217274
rect 140102 216988 140130 217110
rect 140930 216988 140958 217246
rect 141758 216988 141786 217246
rect 142632 217138 142660 218554
rect 143368 217274 143396 222430
rect 144012 221474 144040 231662
rect 144644 230580 144696 230586
rect 144644 230522 144696 230528
rect 144656 229770 144684 230522
rect 144644 229764 144696 229770
rect 144644 229706 144696 229712
rect 144828 229764 144880 229770
rect 144828 229706 144880 229712
rect 144840 222494 144868 229706
rect 145208 223990 145236 231662
rect 145668 229809 145696 231676
rect 146326 231662 146524 231690
rect 145654 229800 145710 229809
rect 145654 229735 145710 229744
rect 146298 229256 146354 229265
rect 146298 229191 146300 229200
rect 146352 229191 146354 229200
rect 146300 229162 146352 229168
rect 145930 225312 145986 225321
rect 145930 225247 145986 225256
rect 145562 224088 145618 224097
rect 145562 224023 145618 224032
rect 145196 223984 145248 223990
rect 145196 223926 145248 223932
rect 144828 222488 144880 222494
rect 145012 222488 145064 222494
rect 144828 222430 144880 222436
rect 145010 222456 145012 222465
rect 145064 222456 145066 222465
rect 145010 222391 145066 222400
rect 144276 222352 144328 222358
rect 144276 222294 144328 222300
rect 144000 221468 144052 221474
rect 144000 221410 144052 221416
rect 144288 217274 144316 222294
rect 144460 221740 144512 221746
rect 144460 221682 144512 221688
rect 144472 221474 144500 221682
rect 144460 221468 144512 221474
rect 144460 221410 144512 221416
rect 145576 218754 145604 224023
rect 145748 219428 145800 219434
rect 145748 219370 145800 219376
rect 145760 218754 145788 219370
rect 145564 218748 145616 218754
rect 145564 218690 145616 218696
rect 145748 218748 145800 218754
rect 145748 218690 145800 218696
rect 145104 218612 145156 218618
rect 145104 218554 145156 218560
rect 143368 217246 143442 217274
rect 142586 217110 142660 217138
rect 142586 216988 142614 217110
rect 143414 216988 143442 217246
rect 144242 217246 144316 217274
rect 144242 216988 144270 217246
rect 145116 217138 145144 218554
rect 145944 217274 145972 225247
rect 146208 221740 146260 221746
rect 146208 221682 146260 221688
rect 146220 218618 146248 221682
rect 146496 220114 146524 231662
rect 146680 231662 146970 231690
rect 147232 231662 147614 231690
rect 147968 231662 148258 231690
rect 148428 231662 148902 231690
rect 149072 231662 149546 231690
rect 149808 231662 150190 231690
rect 150544 231662 150834 231690
rect 151096 231662 151478 231690
rect 151740 231662 152122 231690
rect 146680 229094 146708 231662
rect 146944 229628 146996 229634
rect 146944 229570 146996 229576
rect 146956 229226 146984 229570
rect 146944 229220 146996 229226
rect 146944 229162 146996 229168
rect 146588 229066 146708 229094
rect 147232 229094 147260 231662
rect 147968 229265 147996 231662
rect 147954 229256 148010 229265
rect 147954 229191 148010 229200
rect 147232 229066 147352 229094
rect 146588 221490 146616 229066
rect 146760 226160 146812 226166
rect 146760 226102 146812 226108
rect 146772 225434 146800 226102
rect 146942 225992 146998 226001
rect 146942 225927 146998 225936
rect 146956 225622 146984 225927
rect 146944 225616 146996 225622
rect 147128 225616 147180 225622
rect 146944 225558 146996 225564
rect 147126 225584 147128 225593
rect 147180 225584 147182 225593
rect 147126 225519 147182 225528
rect 146772 225406 147168 225434
rect 147140 225350 147168 225406
rect 146944 225344 146996 225350
rect 146944 225286 146996 225292
rect 147128 225344 147180 225350
rect 147128 225286 147180 225292
rect 146956 225078 146984 225286
rect 146944 225072 146996 225078
rect 146944 225014 146996 225020
rect 147324 224641 147352 229066
rect 147678 228576 147734 228585
rect 147678 228511 147734 228520
rect 147692 228426 147720 228511
rect 147646 228410 147720 228426
rect 147634 228404 147720 228410
rect 147686 228398 147720 228404
rect 147634 228346 147686 228352
rect 147310 224632 147366 224641
rect 147310 224567 147366 224576
rect 147680 223984 147732 223990
rect 147678 223952 147680 223961
rect 147732 223952 147734 223961
rect 147678 223887 147734 223896
rect 146588 221474 146708 221490
rect 146588 221468 146720 221474
rect 146588 221462 146668 221468
rect 146668 221410 146720 221416
rect 148428 220833 148456 231662
rect 148600 229764 148652 229770
rect 148600 229706 148652 229712
rect 148414 220824 148470 220833
rect 148414 220759 148470 220768
rect 146484 220108 146536 220114
rect 146484 220050 146536 220056
rect 147588 220108 147640 220114
rect 147588 220050 147640 220056
rect 146484 219428 146536 219434
rect 146484 219370 146536 219376
rect 146496 219162 146524 219370
rect 146484 219156 146536 219162
rect 146484 219098 146536 219104
rect 146944 219156 146996 219162
rect 146944 219098 146996 219104
rect 146956 218754 146984 219098
rect 146944 218748 146996 218754
rect 146944 218690 146996 218696
rect 146208 218612 146260 218618
rect 146208 218554 146260 218560
rect 146760 218612 146812 218618
rect 146760 218554 146812 218560
rect 145070 217110 145144 217138
rect 145898 217246 145972 217274
rect 145070 216988 145098 217110
rect 145898 216988 145926 217246
rect 146772 217138 146800 218554
rect 147600 217274 147628 220050
rect 148414 219328 148470 219337
rect 148382 219298 148414 219314
rect 148370 219292 148414 219298
rect 148422 219263 148470 219272
rect 148370 219234 148422 219240
rect 148232 218884 148284 218890
rect 148232 218826 148284 218832
rect 148416 218884 148468 218890
rect 148416 218826 148468 218832
rect 148244 218482 148272 218826
rect 148232 218476 148284 218482
rect 148232 218418 148284 218424
rect 146726 217110 146800 217138
rect 147554 217246 147628 217274
rect 146726 216988 146754 217110
rect 147554 216988 147582 217246
rect 148428 217138 148456 218826
rect 148612 218793 148640 229706
rect 149072 221921 149100 231662
rect 149808 228585 149836 231662
rect 150544 230586 150572 231662
rect 150532 230580 150584 230586
rect 150532 230522 150584 230528
rect 150900 230580 150952 230586
rect 150900 230522 150952 230528
rect 150912 229770 150940 230522
rect 150900 229764 150952 229770
rect 150900 229706 150952 229712
rect 149794 228576 149850 228585
rect 149794 228511 149850 228520
rect 150162 227216 150218 227225
rect 150162 227151 150164 227160
rect 150216 227151 150218 227160
rect 150348 227180 150400 227186
rect 150164 227122 150216 227128
rect 150348 227122 150400 227128
rect 149058 221912 149114 221921
rect 149058 221847 149114 221856
rect 149244 221876 149296 221882
rect 149244 221818 149296 221824
rect 149256 221762 149284 221818
rect 148980 221734 149284 221762
rect 148980 218890 149008 221734
rect 150360 219298 150388 227122
rect 150714 220824 150770 220833
rect 150714 220759 150770 220768
rect 150728 220386 150756 220759
rect 150716 220380 150768 220386
rect 150716 220322 150768 220328
rect 150900 220380 150952 220386
rect 150900 220322 150952 220328
rect 149244 219292 149296 219298
rect 149244 219234 149296 219240
rect 150348 219292 150400 219298
rect 150348 219234 150400 219240
rect 148968 218884 149020 218890
rect 148968 218826 149020 218832
rect 148598 218784 148654 218793
rect 148598 218719 148654 218728
rect 149256 217138 149284 219234
rect 149888 218884 149940 218890
rect 149888 218826 149940 218832
rect 149900 218482 149928 218826
rect 149888 218476 149940 218482
rect 149888 218418 149940 218424
rect 150072 218476 150124 218482
rect 150072 218418 150124 218424
rect 150084 217138 150112 218418
rect 150912 217138 150940 220322
rect 151096 220153 151124 231662
rect 151360 229764 151412 229770
rect 151360 229706 151412 229712
rect 151372 222494 151400 229706
rect 151740 226930 151768 231662
rect 151910 227488 151966 227497
rect 151910 227423 151966 227432
rect 151924 227322 151952 227423
rect 151912 227316 151964 227322
rect 151912 227258 151964 227264
rect 152280 227180 152332 227186
rect 151924 227140 152280 227168
rect 151924 227050 151952 227140
rect 152280 227122 152332 227128
rect 151912 227044 151964 227050
rect 151912 226986 151964 226992
rect 151740 226902 152136 226930
rect 151726 223816 151782 223825
rect 151726 223751 151782 223760
rect 151360 222488 151412 222494
rect 151360 222430 151412 222436
rect 151082 220144 151138 220153
rect 151082 220079 151138 220088
rect 151740 217138 151768 223751
rect 152108 221746 152136 226902
rect 152752 226386 152780 231676
rect 153396 229226 153424 231676
rect 153672 231662 154054 231690
rect 154592 231662 154698 231690
rect 153384 229220 153436 229226
rect 153384 229162 153436 229168
rect 153292 228540 153344 228546
rect 153292 228482 153344 228488
rect 152922 227488 152978 227497
rect 152922 227423 152978 227432
rect 152936 227322 152964 227423
rect 152924 227316 152976 227322
rect 152924 227258 152976 227264
rect 152568 226358 152780 226386
rect 152568 224369 152596 226358
rect 152832 226296 152884 226302
rect 152832 226238 152884 226244
rect 152844 226001 152872 226238
rect 153106 226128 153162 226137
rect 153106 226063 153162 226072
rect 152830 225992 152886 226001
rect 152830 225927 152886 225936
rect 152554 224360 152610 224369
rect 152554 224295 152610 224304
rect 152096 221740 152148 221746
rect 152096 221682 152148 221688
rect 152922 219328 152978 219337
rect 152556 219292 152608 219298
rect 153120 219298 153148 226063
rect 153304 225321 153332 228482
rect 153290 225312 153346 225321
rect 153290 225247 153346 225256
rect 153672 220561 153700 231662
rect 153844 229220 153896 229226
rect 153844 229162 153896 229168
rect 153658 220552 153714 220561
rect 153658 220487 153714 220496
rect 152922 219263 152978 219272
rect 153108 219292 153160 219298
rect 152556 219234 152608 219240
rect 152280 219156 152332 219162
rect 152280 219098 152332 219104
rect 152094 218920 152150 218929
rect 152292 218890 152320 219098
rect 152094 218855 152096 218864
rect 152148 218855 152150 218864
rect 152280 218884 152332 218890
rect 152096 218826 152148 218832
rect 152280 218826 152332 218832
rect 152568 217138 152596 219234
rect 152740 219020 152792 219026
rect 152740 218962 152792 218968
rect 152752 218754 152780 218962
rect 152936 218754 152964 219263
rect 153108 219234 153160 219240
rect 153384 219292 153436 219298
rect 153384 219234 153436 219240
rect 152740 218748 152792 218754
rect 152740 218690 152792 218696
rect 152924 218748 152976 218754
rect 152924 218690 152976 218696
rect 153396 217138 153424 219234
rect 153856 218929 153884 229162
rect 154592 227225 154620 231662
rect 154578 227216 154634 227225
rect 154578 227151 154634 227160
rect 155328 226953 155356 231676
rect 155972 229906 156000 231676
rect 156156 231662 156630 231690
rect 155960 229900 156012 229906
rect 155960 229842 156012 229848
rect 155866 228032 155922 228041
rect 155866 227967 155922 227976
rect 155314 226944 155370 226953
rect 155314 226879 155370 226888
rect 154578 224224 154634 224233
rect 154578 224159 154634 224168
rect 154592 223990 154620 224159
rect 154580 223984 154632 223990
rect 154580 223926 154632 223932
rect 155038 222592 155094 222601
rect 155038 222527 155094 222536
rect 154212 222488 154264 222494
rect 154212 222430 154264 222436
rect 153842 218920 153898 218929
rect 153842 218855 153898 218864
rect 154224 217138 154252 222430
rect 155052 217138 155080 222527
rect 155880 217274 155908 227967
rect 156156 220833 156184 231662
rect 156328 229900 156380 229906
rect 156328 229842 156380 229848
rect 156142 220824 156198 220833
rect 156142 220759 156198 220768
rect 156340 218754 156368 229842
rect 157260 224954 157288 231676
rect 157628 231662 157918 231690
rect 158272 231662 158562 231690
rect 158824 231662 159206 231690
rect 157430 228576 157486 228585
rect 157430 228511 157486 228520
rect 157444 228410 157472 228511
rect 157432 228404 157484 228410
rect 157432 228346 157484 228352
rect 157628 226250 157656 231662
rect 158272 230722 158300 231662
rect 158260 230716 158312 230722
rect 158260 230658 158312 230664
rect 157982 228984 158038 228993
rect 157982 228919 158038 228928
rect 157800 228404 157852 228410
rect 157800 228346 157852 228352
rect 157812 228041 157840 228346
rect 157798 228032 157854 228041
rect 157798 227967 157854 227976
rect 157444 226222 157656 226250
rect 157444 226166 157472 226222
rect 157432 226160 157484 226166
rect 157616 226160 157668 226166
rect 157432 226102 157484 226108
rect 157614 226128 157616 226137
rect 157668 226128 157670 226137
rect 157614 226063 157670 226072
rect 157076 224926 157288 224954
rect 156880 223984 156932 223990
rect 156880 223926 156932 223932
rect 156892 223825 156920 223926
rect 156878 223816 156934 223825
rect 156878 223751 156934 223760
rect 156880 223304 156932 223310
rect 156878 223272 156880 223281
rect 156932 223272 156934 223281
rect 156878 223207 156934 223216
rect 157076 223174 157104 224926
rect 157338 224632 157394 224641
rect 157338 224567 157394 224576
rect 157352 224482 157380 224567
rect 157306 224454 157380 224482
rect 157306 224398 157334 224454
rect 157294 224392 157346 224398
rect 157294 224334 157346 224340
rect 157432 224392 157484 224398
rect 157432 224334 157484 224340
rect 157444 224233 157472 224334
rect 157430 224224 157486 224233
rect 157430 224159 157486 224168
rect 157432 223304 157484 223310
rect 157430 223272 157432 223281
rect 157484 223272 157486 223281
rect 157430 223207 157486 223216
rect 157064 223168 157116 223174
rect 157064 223110 157116 223116
rect 157248 223168 157300 223174
rect 157248 223110 157300 223116
rect 157260 222601 157288 223110
rect 157246 222592 157302 222601
rect 157246 222527 157302 222536
rect 157338 220552 157394 220561
rect 157338 220487 157340 220496
rect 157392 220487 157394 220496
rect 157524 220516 157576 220522
rect 157340 220458 157392 220464
rect 157524 220458 157576 220464
rect 156328 218748 156380 218754
rect 156328 218690 156380 218696
rect 156696 218748 156748 218754
rect 156696 218690 156748 218696
rect 148382 217110 148456 217138
rect 149210 217110 149284 217138
rect 150038 217110 150112 217138
rect 150866 217110 150940 217138
rect 151694 217110 151768 217138
rect 152522 217110 152596 217138
rect 153350 217110 153424 217138
rect 154178 217110 154252 217138
rect 155006 217110 155080 217138
rect 155834 217246 155908 217274
rect 148382 216988 148410 217110
rect 149210 216988 149238 217110
rect 150038 216988 150066 217110
rect 150866 216988 150894 217110
rect 151694 216988 151722 217110
rect 152522 216988 152550 217110
rect 153350 216988 153378 217110
rect 154178 216988 154206 217110
rect 155006 216988 155034 217110
rect 155834 216988 155862 217246
rect 156708 217138 156736 218690
rect 157246 218648 157302 218657
rect 157246 218583 157302 218592
rect 157260 218482 157288 218583
rect 157248 218476 157300 218482
rect 157248 218418 157300 218424
rect 157536 217138 157564 220458
rect 157996 218618 158024 228919
rect 158824 228585 158852 231662
rect 158810 228576 158866 228585
rect 158810 228511 158866 228520
rect 159638 227488 159694 227497
rect 159638 227423 159640 227432
rect 159692 227423 159694 227432
rect 159640 227394 159692 227400
rect 159836 223310 159864 231676
rect 160480 228313 160508 231676
rect 161124 230450 161152 231676
rect 161112 230444 161164 230450
rect 161112 230386 161164 230392
rect 161296 230444 161348 230450
rect 161296 230386 161348 230392
rect 160466 228304 160522 228313
rect 160466 228239 160522 228248
rect 161308 227746 161336 230386
rect 160664 227718 161336 227746
rect 160008 227452 160060 227458
rect 160008 227394 160060 227400
rect 159824 223304 159876 223310
rect 159824 223246 159876 223252
rect 158350 223136 158406 223145
rect 158350 223071 158406 223080
rect 157984 218612 158036 218618
rect 157984 218554 158036 218560
rect 157706 218512 157762 218521
rect 157706 218447 157708 218456
rect 157760 218447 157762 218456
rect 157708 218418 157760 218424
rect 158364 217138 158392 223071
rect 160020 218618 160048 227394
rect 159180 218612 159232 218618
rect 159180 218554 159232 218560
rect 160008 218612 160060 218618
rect 160008 218554 160060 218560
rect 159192 217138 159220 218554
rect 160664 218482 160692 227718
rect 161202 226128 161258 226137
rect 161202 226063 161258 226072
rect 161216 225894 161244 226063
rect 161204 225888 161256 225894
rect 161204 225830 161256 225836
rect 160928 223304 160980 223310
rect 160928 223246 160980 223252
rect 160940 222766 160968 223246
rect 161204 223168 161256 223174
rect 161204 223110 161256 223116
rect 161388 223168 161440 223174
rect 161388 223110 161440 223116
rect 161216 222766 161244 223110
rect 160928 222760 160980 222766
rect 160928 222702 160980 222708
rect 161204 222760 161256 222766
rect 161204 222702 161256 222708
rect 161400 218618 161428 223110
rect 161768 220561 161796 231676
rect 162136 231662 162426 231690
rect 162964 231662 163070 231690
rect 161940 226296 161992 226302
rect 161940 226238 161992 226244
rect 161952 225894 161980 226238
rect 161940 225888 161992 225894
rect 161940 225830 161992 225836
rect 162136 224954 162164 231662
rect 162308 226296 162360 226302
rect 162308 226238 162360 226244
rect 162320 226137 162348 226238
rect 162306 226128 162362 226137
rect 162306 226063 162362 226072
rect 162306 225584 162362 225593
rect 162306 225519 162362 225528
rect 162320 225078 162348 225519
rect 162308 225072 162360 225078
rect 162308 225014 162360 225020
rect 162492 225072 162544 225078
rect 162492 225014 162544 225020
rect 161952 224926 162164 224954
rect 161952 223582 161980 224926
rect 161940 223576 161992 223582
rect 161940 223518 161992 223524
rect 162124 223576 162176 223582
rect 162124 223518 162176 223524
rect 162136 223038 162164 223518
rect 162124 223032 162176 223038
rect 162124 222974 162176 222980
rect 162124 221876 162176 221882
rect 162124 221818 162176 221824
rect 162136 221474 162164 221818
rect 162308 221740 162360 221746
rect 162308 221682 162360 221688
rect 162320 221474 162348 221682
rect 162124 221468 162176 221474
rect 162124 221410 162176 221416
rect 162308 221468 162360 221474
rect 162308 221410 162360 221416
rect 162308 220788 162360 220794
rect 162308 220730 162360 220736
rect 161754 220552 161810 220561
rect 161754 220487 161810 220496
rect 161938 220552 161994 220561
rect 162320 220522 162348 220730
rect 161938 220487 161994 220496
rect 162308 220516 162360 220522
rect 161952 220402 161980 220487
rect 162308 220458 162360 220464
rect 161768 220386 161980 220402
rect 161756 220380 161980 220386
rect 161808 220374 161980 220380
rect 161756 220322 161808 220328
rect 162308 219292 162360 219298
rect 162308 219234 162360 219240
rect 162320 218754 162348 219234
rect 162308 218748 162360 218754
rect 162308 218690 162360 218696
rect 160836 218612 160888 218618
rect 160836 218554 160888 218560
rect 161388 218612 161440 218618
rect 161388 218554 161440 218560
rect 160652 218476 160704 218482
rect 160652 218418 160704 218424
rect 159638 218240 159694 218249
rect 159638 218175 159640 218184
rect 159692 218175 159694 218184
rect 159640 218146 159692 218152
rect 160008 218068 160060 218074
rect 160008 218010 160060 218016
rect 160020 217138 160048 218010
rect 160848 217138 160876 218554
rect 161664 218476 161716 218482
rect 161664 218418 161716 218424
rect 161676 217138 161704 218418
rect 162504 217274 162532 225014
rect 162964 224641 162992 231662
rect 163700 229226 163728 231676
rect 163688 229220 163740 229226
rect 163688 229162 163740 229168
rect 163872 229220 163924 229226
rect 163872 229162 163924 229168
rect 163884 228993 163912 229162
rect 163870 228984 163926 228993
rect 163870 228919 163926 228928
rect 164344 227322 164372 231676
rect 164528 231662 165002 231690
rect 164332 227316 164384 227322
rect 164332 227258 164384 227264
rect 162950 224632 163006 224641
rect 162950 224567 163006 224576
rect 163962 224496 164018 224505
rect 163962 224431 164018 224440
rect 162676 221740 162728 221746
rect 162676 221682 162728 221688
rect 162688 218482 162716 221682
rect 162858 220552 162914 220561
rect 162858 220487 162860 220496
rect 162912 220487 162914 220496
rect 162860 220458 162912 220464
rect 163976 219298 164004 224431
rect 164528 223310 164556 231662
rect 165436 230580 165488 230586
rect 165436 230522 165488 230528
rect 165448 228682 165476 230522
rect 165436 228676 165488 228682
rect 165436 228618 165488 228624
rect 165436 227316 165488 227322
rect 165436 227258 165488 227264
rect 164516 223304 164568 223310
rect 164516 223246 164568 223252
rect 164148 223168 164200 223174
rect 165068 223168 165120 223174
rect 164148 223110 164200 223116
rect 165066 223136 165068 223145
rect 165120 223136 165122 223145
rect 162860 219292 162912 219298
rect 162860 219234 162912 219240
rect 163964 219292 164016 219298
rect 163964 219234 164016 219240
rect 162676 218476 162728 218482
rect 162676 218418 162728 218424
rect 162872 218249 162900 219234
rect 163320 218476 163372 218482
rect 163320 218418 163372 218424
rect 162858 218240 162914 218249
rect 162858 218175 162914 218184
rect 156662 217110 156736 217138
rect 157490 217110 157564 217138
rect 158318 217110 158392 217138
rect 159146 217110 159220 217138
rect 159974 217110 160048 217138
rect 160802 217110 160876 217138
rect 161630 217110 161704 217138
rect 162458 217246 162532 217274
rect 156662 216988 156690 217110
rect 157490 216988 157518 217110
rect 158318 216988 158346 217110
rect 159146 216988 159174 217110
rect 159974 216988 160002 217110
rect 160802 216988 160830 217110
rect 161630 216988 161658 217110
rect 162458 216988 162486 217246
rect 163332 217138 163360 218418
rect 164160 217138 164188 223110
rect 165066 223071 165122 223080
rect 165448 219298 165476 227258
rect 165632 222873 165660 231676
rect 166276 230042 166304 231676
rect 166644 231662 166934 231690
rect 167196 231662 167578 231690
rect 167840 231662 168222 231690
rect 166264 230036 166316 230042
rect 166264 229978 166316 229984
rect 166448 230036 166500 230042
rect 166448 229978 166500 229984
rect 166460 229226 166488 229978
rect 166448 229220 166500 229226
rect 166448 229162 166500 229168
rect 166446 228848 166502 228857
rect 166446 228783 166448 228792
rect 166500 228783 166502 228792
rect 166448 228754 166500 228760
rect 166446 228440 166502 228449
rect 166446 228375 166502 228384
rect 166460 225162 166488 228375
rect 166644 227497 166672 231662
rect 166908 229220 166960 229226
rect 166908 229162 166960 229168
rect 166920 228954 166948 229162
rect 166908 228948 166960 228954
rect 166908 228890 166960 228896
rect 166630 227488 166686 227497
rect 166630 227423 166686 227432
rect 166816 227452 166868 227458
rect 166816 227394 166868 227400
rect 166828 226370 166856 227394
rect 166816 226364 166868 226370
rect 166816 226306 166868 226312
rect 166632 226296 166684 226302
rect 166632 226238 166684 226244
rect 166644 225434 166672 226238
rect 166816 226024 166868 226030
rect 166814 225992 166816 226001
rect 166954 226024 167006 226030
rect 166868 225992 166870 226001
rect 166954 225966 167006 225972
rect 166814 225927 166870 225936
rect 166966 225842 166994 225966
rect 166920 225814 166994 225842
rect 166920 225593 166948 225814
rect 166906 225584 166962 225593
rect 166906 225519 166962 225528
rect 166644 225406 166856 225434
rect 166460 225134 166672 225162
rect 166448 225072 166500 225078
rect 166446 225040 166448 225049
rect 166500 225040 166502 225049
rect 166446 224975 166502 224984
rect 166446 223136 166502 223145
rect 166446 223071 166502 223080
rect 166460 222902 166488 223071
rect 166448 222896 166500 222902
rect 165618 222864 165674 222873
rect 166448 222838 166500 222844
rect 165618 222799 165674 222808
rect 166262 219328 166318 219337
rect 164976 219292 165028 219298
rect 164976 219234 165028 219240
rect 165436 219292 165488 219298
rect 165436 219234 165488 219240
rect 165804 219292 165856 219298
rect 166644 219314 166672 225134
rect 166828 225078 166856 225406
rect 166998 225312 167054 225321
rect 166998 225247 167054 225256
rect 167012 225078 167040 225247
rect 166816 225072 166868 225078
rect 166816 225014 166868 225020
rect 167000 225072 167052 225078
rect 167000 225014 167052 225020
rect 166954 223032 167006 223038
rect 166460 219298 166672 219314
rect 166262 219263 166318 219272
rect 166448 219292 166672 219298
rect 165804 219234 165856 219240
rect 164988 217138 165016 219234
rect 165816 217138 165844 219234
rect 166078 218920 166134 218929
rect 166078 218855 166080 218864
rect 166132 218855 166134 218864
rect 166080 218826 166132 218832
rect 166276 218482 166304 219263
rect 166500 219286 166672 219292
rect 166828 222980 166954 222986
rect 166828 222974 167006 222980
rect 166828 222958 166994 222974
rect 166448 219234 166500 219240
rect 166828 218906 166856 222958
rect 167196 220658 167224 231662
rect 167642 229256 167698 229265
rect 167642 229191 167698 229200
rect 167368 225072 167420 225078
rect 167366 225040 167368 225049
rect 167420 225040 167422 225049
rect 167366 224975 167422 224984
rect 167184 220652 167236 220658
rect 167184 220594 167236 220600
rect 167656 219434 167684 229191
rect 167840 223582 167868 231662
rect 168196 229084 168248 229090
rect 168196 229026 168248 229032
rect 168208 228857 168236 229026
rect 168194 228848 168250 228857
rect 168012 228812 168064 228818
rect 168194 228783 168250 228792
rect 168012 228754 168064 228760
rect 168024 228449 168052 228754
rect 168010 228440 168066 228449
rect 168010 228375 168066 228384
rect 168852 227186 168880 231676
rect 169036 231662 169510 231690
rect 169864 231662 170154 231690
rect 170416 231662 170798 231690
rect 168840 227180 168892 227186
rect 168840 227122 168892 227128
rect 169036 226001 169064 231662
rect 169576 227180 169628 227186
rect 169576 227122 169628 227128
rect 169206 226128 169262 226137
rect 169206 226063 169262 226072
rect 169022 225992 169078 226001
rect 169022 225927 169078 225936
rect 167828 223576 167880 223582
rect 167828 223518 167880 223524
rect 168288 223576 168340 223582
rect 168288 223518 168340 223524
rect 167288 219406 167684 219434
rect 167092 219156 167144 219162
rect 167092 219098 167144 219104
rect 167104 218929 167132 219098
rect 166460 218878 166856 218906
rect 167090 218920 167146 218929
rect 166954 218884 167006 218890
rect 166264 218476 166316 218482
rect 166264 218418 166316 218424
rect 166460 218210 166488 218878
rect 167090 218855 167146 218864
rect 166954 218826 167006 218832
rect 166966 218770 166994 218826
rect 166828 218742 166994 218770
rect 166448 218204 166500 218210
rect 166448 218146 166500 218152
rect 166632 218204 166684 218210
rect 166632 218146 166684 218152
rect 166644 217138 166672 218146
rect 166828 218074 166856 218742
rect 167288 218618 167316 219406
rect 167276 218612 167328 218618
rect 167276 218554 167328 218560
rect 167000 218476 167052 218482
rect 167000 218418 167052 218424
rect 167012 218210 167040 218418
rect 167000 218204 167052 218210
rect 167000 218146 167052 218152
rect 168104 218204 168156 218210
rect 168104 218146 168156 218152
rect 166816 218068 166868 218074
rect 166816 218010 166868 218016
rect 167460 218068 167512 218074
rect 167460 218010 167512 218016
rect 167472 217138 167500 218010
rect 168116 217274 168144 218146
rect 168300 218074 168328 223518
rect 169220 219434 169248 226063
rect 168944 219406 169248 219434
rect 168944 219298 168972 219406
rect 169114 219328 169170 219337
rect 168932 219292 168984 219298
rect 169114 219263 169116 219272
rect 168932 219234 168984 219240
rect 169168 219263 169170 219272
rect 169116 219234 169168 219240
rect 169588 218074 169616 227122
rect 169864 225321 169892 231662
rect 169850 225312 169906 225321
rect 169850 225247 169906 225256
rect 170416 223145 170444 231662
rect 170770 224496 170826 224505
rect 170826 224454 171134 224482
rect 170770 224431 170826 224440
rect 171106 224398 171134 224454
rect 170956 224392 171008 224398
rect 170956 224334 171008 224340
rect 171094 224392 171146 224398
rect 171094 224334 171146 224340
rect 170968 224233 170996 224334
rect 171428 224233 171456 231676
rect 172072 230586 172100 231676
rect 172060 230580 172112 230586
rect 172060 230522 172112 230528
rect 172426 229256 172482 229265
rect 172244 229220 172296 229226
rect 172426 229191 172428 229200
rect 172244 229162 172296 229168
rect 172480 229191 172482 229200
rect 172428 229162 172480 229168
rect 172256 228954 172284 229162
rect 172426 228984 172482 228993
rect 172244 228948 172296 228954
rect 172426 228919 172482 228928
rect 172244 228890 172296 228896
rect 170954 224224 171010 224233
rect 170954 224159 171010 224168
rect 171414 224224 171470 224233
rect 171414 224159 171470 224168
rect 170402 223136 170458 223145
rect 170402 223071 170458 223080
rect 171230 222320 171286 222329
rect 171230 222255 171286 222264
rect 171244 222170 171272 222255
rect 171060 222154 171272 222170
rect 171048 222148 171272 222154
rect 171100 222142 171272 222148
rect 171048 222090 171100 222096
rect 171046 221912 171102 221921
rect 171046 221847 171102 221856
rect 171506 221912 171562 221921
rect 171506 221847 171508 221856
rect 170772 220652 170824 220658
rect 170772 220594 170824 220600
rect 169944 218612 169996 218618
rect 169944 218554 169996 218560
rect 168288 218068 168340 218074
rect 168288 218010 168340 218016
rect 169116 218068 169168 218074
rect 169116 218010 169168 218016
rect 169576 218068 169628 218074
rect 169576 218010 169628 218016
rect 168116 217246 168282 217274
rect 163286 217110 163360 217138
rect 164114 217110 164188 217138
rect 164942 217110 165016 217138
rect 165770 217110 165844 217138
rect 166598 217110 166672 217138
rect 167426 217110 167500 217138
rect 163286 216988 163314 217110
rect 164114 216988 164142 217110
rect 164942 216988 164970 217110
rect 165770 216988 165798 217110
rect 166598 216988 166626 217110
rect 167426 216988 167454 217110
rect 168254 216988 168282 217246
rect 169128 217138 169156 218010
rect 169956 217138 169984 218554
rect 170784 217274 170812 220594
rect 171060 218210 171088 221847
rect 171560 221847 171562 221856
rect 171508 221818 171560 221824
rect 172440 219434 172468 228919
rect 172716 220794 172744 231676
rect 172992 231662 173374 231690
rect 172992 222018 173020 231662
rect 174004 229090 174032 231676
rect 173992 229084 174044 229090
rect 173992 229026 174044 229032
rect 174648 227594 174676 231676
rect 174820 229084 174872 229090
rect 174820 229026 174872 229032
rect 174636 227588 174688 227594
rect 174636 227530 174688 227536
rect 174832 224210 174860 229026
rect 175292 228954 175320 231676
rect 175476 231662 175950 231690
rect 175280 228948 175332 228954
rect 175280 228890 175332 228896
rect 175188 227452 175240 227458
rect 175188 227394 175240 227400
rect 174556 224182 174860 224210
rect 172980 222012 173032 222018
rect 172980 221954 173032 221960
rect 172704 220788 172756 220794
rect 172704 220730 172756 220736
rect 173348 220788 173400 220794
rect 173348 220730 173400 220736
rect 173360 219978 173388 220730
rect 173532 220516 173584 220522
rect 173532 220458 173584 220464
rect 173544 219978 173572 220458
rect 173348 219972 173400 219978
rect 173348 219914 173400 219920
rect 173532 219972 173584 219978
rect 173532 219914 173584 219920
rect 172348 219406 172468 219434
rect 171048 218204 171100 218210
rect 171048 218146 171100 218152
rect 171600 218204 171652 218210
rect 171600 218146 171652 218152
rect 169082 217110 169156 217138
rect 169910 217110 169984 217138
rect 170738 217246 170812 217274
rect 169082 216988 169110 217110
rect 169910 216988 169938 217110
rect 170738 216988 170766 217246
rect 171612 217138 171640 218146
rect 172348 217274 172376 219406
rect 174556 218346 174584 224182
rect 174912 222216 174964 222222
rect 174912 222158 174964 222164
rect 174544 218340 174596 218346
rect 174544 218282 174596 218288
rect 173256 218068 173308 218074
rect 173256 218010 173308 218016
rect 174084 218068 174136 218074
rect 174084 218010 174136 218016
rect 172348 217246 172422 217274
rect 171566 217110 171640 217138
rect 171566 216988 171594 217110
rect 172394 216988 172422 217246
rect 173268 217138 173296 218010
rect 174096 217138 174124 218010
rect 174924 217274 174952 222158
rect 175200 218074 175228 227394
rect 175476 222630 175504 231662
rect 176108 230580 176160 230586
rect 176108 230522 176160 230528
rect 175646 228984 175702 228993
rect 175646 228919 175648 228928
rect 175700 228919 175702 228928
rect 175648 228890 175700 228896
rect 176120 225894 176148 230522
rect 176580 229906 176608 231676
rect 177040 231662 177238 231690
rect 177408 231662 177882 231690
rect 178052 231662 178526 231690
rect 176568 229900 176620 229906
rect 176568 229842 176620 229848
rect 176476 226024 176528 226030
rect 176476 225966 176528 225972
rect 176108 225888 176160 225894
rect 176108 225830 176160 225836
rect 176488 225842 176516 225966
rect 176488 225814 176700 225842
rect 176672 225758 176700 225814
rect 176476 225752 176528 225758
rect 176476 225694 176528 225700
rect 176660 225752 176712 225758
rect 176660 225694 176712 225700
rect 176488 225593 176516 225694
rect 177040 225593 177068 231662
rect 177212 225888 177264 225894
rect 177212 225830 177264 225836
rect 176474 225584 176530 225593
rect 176474 225519 176530 225528
rect 177026 225584 177082 225593
rect 177026 225519 177082 225528
rect 177224 225321 177252 225830
rect 176474 225312 176530 225321
rect 176474 225247 176530 225256
rect 177210 225312 177266 225321
rect 177210 225247 177266 225256
rect 176108 223032 176160 223038
rect 176108 222974 176160 222980
rect 176292 223032 176344 223038
rect 176292 222974 176344 222980
rect 176120 222766 176148 222974
rect 176108 222760 176160 222766
rect 176108 222702 176160 222708
rect 175464 222624 175516 222630
rect 175464 222566 175516 222572
rect 176304 222222 176332 222974
rect 176292 222216 176344 222222
rect 176292 222158 176344 222164
rect 176108 222080 176160 222086
rect 176106 222048 176108 222057
rect 176160 222048 176162 222057
rect 176106 221983 176162 221992
rect 176292 222012 176344 222018
rect 176292 221954 176344 221960
rect 176304 218346 176332 221954
rect 176292 218340 176344 218346
rect 176292 218282 176344 218288
rect 176488 218210 176516 225247
rect 177408 224954 177436 231662
rect 177580 229900 177632 229906
rect 177580 229842 177632 229848
rect 177592 224954 177620 229842
rect 177040 224926 177436 224954
rect 177500 224926 177620 224954
rect 177040 222057 177068 224926
rect 177500 224210 177528 224926
rect 177224 224182 177528 224210
rect 177026 222048 177082 222057
rect 177026 221983 177082 221992
rect 175740 218204 175792 218210
rect 175740 218146 175792 218152
rect 176476 218204 176528 218210
rect 176476 218146 176528 218152
rect 175188 218068 175240 218074
rect 175188 218010 175240 218016
rect 173222 217110 173296 217138
rect 174050 217110 174124 217138
rect 174878 217246 174952 217274
rect 173222 216988 173250 217110
rect 174050 216988 174078 217110
rect 174878 216988 174906 217246
rect 175752 217138 175780 218146
rect 177224 218074 177252 224182
rect 178052 221513 178080 231662
rect 179156 229362 179184 231676
rect 179144 229356 179196 229362
rect 179144 229298 179196 229304
rect 179800 228682 179828 231676
rect 179984 231662 180458 231690
rect 179788 228676 179840 228682
rect 179788 228618 179840 228624
rect 179052 227588 179104 227594
rect 179052 227530 179104 227536
rect 178684 226024 178736 226030
rect 178682 225992 178684 226001
rect 178736 225992 178738 226001
rect 178682 225927 178738 225936
rect 178224 222148 178276 222154
rect 178224 222090 178276 222096
rect 178038 221504 178094 221513
rect 178038 221439 178094 221448
rect 177396 220652 177448 220658
rect 177396 220594 177448 220600
rect 176568 218068 176620 218074
rect 176568 218010 176620 218016
rect 177212 218068 177264 218074
rect 177212 218010 177264 218016
rect 176580 217138 176608 218010
rect 177408 217274 177436 220594
rect 177580 218612 177632 218618
rect 177580 218554 177632 218560
rect 177592 218074 177620 218554
rect 177580 218068 177632 218074
rect 177580 218010 177632 218016
rect 178236 217274 178264 222090
rect 179064 217274 179092 227530
rect 179984 222329 180012 231662
rect 181088 230586 181116 231676
rect 181076 230580 181128 230586
rect 181076 230522 181128 230528
rect 181732 230042 181760 231676
rect 181720 230036 181772 230042
rect 181720 229978 181772 229984
rect 181352 229356 181404 229362
rect 181352 229298 181404 229304
rect 180614 228984 180670 228993
rect 180614 228919 180670 228928
rect 179970 222320 180026 222329
rect 179970 222255 180026 222264
rect 180628 222170 180656 228919
rect 181364 228834 181392 229298
rect 181720 229084 181772 229090
rect 181720 229026 181772 229032
rect 181364 228806 181484 228834
rect 181260 228744 181312 228750
rect 181258 228712 181260 228721
rect 181312 228712 181314 228721
rect 181258 228647 181314 228656
rect 181074 228032 181130 228041
rect 181074 227967 181076 227976
rect 181128 227967 181130 227976
rect 181076 227938 181128 227944
rect 180444 222142 180656 222170
rect 180444 219434 180472 222142
rect 180616 222012 180668 222018
rect 180616 221954 180668 221960
rect 180628 221241 180656 221954
rect 180614 221232 180670 221241
rect 180614 221167 180670 221176
rect 180890 221232 180946 221241
rect 180890 221167 180946 221176
rect 180904 221066 180932 221167
rect 180754 221060 180806 221066
rect 180754 221002 180806 221008
rect 180892 221060 180944 221066
rect 180892 221002 180944 221008
rect 180766 220946 180794 221002
rect 180766 220918 180840 220946
rect 180812 220833 180840 220918
rect 180798 220824 180854 220833
rect 180798 220759 180854 220768
rect 181456 219434 181484 228806
rect 181732 228041 181760 229026
rect 181902 228984 181958 228993
rect 181902 228919 181904 228928
rect 181956 228919 181958 228928
rect 181904 228890 181956 228896
rect 181902 228712 181958 228721
rect 181902 228647 181958 228656
rect 181916 228138 181944 228647
rect 181904 228132 181956 228138
rect 181904 228074 181956 228080
rect 181718 228032 181774 228041
rect 181718 227967 181774 227976
rect 182376 227730 182404 231676
rect 182652 231662 183034 231690
rect 183678 231662 183876 231690
rect 182364 227724 182416 227730
rect 182364 227666 182416 227672
rect 181628 222148 181680 222154
rect 181628 222090 181680 222096
rect 181640 219434 181668 222090
rect 182652 220794 182680 231662
rect 183282 225176 183338 225185
rect 183282 225111 183338 225120
rect 182640 220788 182692 220794
rect 182640 220730 182692 220736
rect 183100 220788 183152 220794
rect 183100 220730 183152 220736
rect 180444 219406 180748 219434
rect 179880 218204 179932 218210
rect 179880 218146 179932 218152
rect 175706 217110 175780 217138
rect 176534 217110 176608 217138
rect 177362 217246 177436 217274
rect 178190 217246 178264 217274
rect 179018 217246 179092 217274
rect 175706 216988 175734 217110
rect 176534 216988 176562 217110
rect 177362 216988 177390 217246
rect 178190 216988 178218 217246
rect 179018 216988 179046 217246
rect 179892 217138 179920 218146
rect 180720 217274 180748 219406
rect 181364 219406 181484 219434
rect 181548 219406 181668 219434
rect 181364 218074 181392 219406
rect 181352 218068 181404 218074
rect 181352 218010 181404 218016
rect 181548 217274 181576 219406
rect 182364 218068 182416 218074
rect 182364 218010 182416 218016
rect 179846 217110 179920 217138
rect 180674 217246 180748 217274
rect 181502 217246 181576 217274
rect 179846 216988 179874 217110
rect 180674 216988 180702 217246
rect 181502 216988 181530 217246
rect 182376 217138 182404 218010
rect 183112 217274 183140 220730
rect 183296 218074 183324 225111
rect 183848 224262 183876 231662
rect 184308 230178 184336 231676
rect 184296 230172 184348 230178
rect 184296 230114 184348 230120
rect 184204 230036 184256 230042
rect 184204 229978 184256 229984
rect 183836 224256 183888 224262
rect 183836 224198 183888 224204
rect 184216 220794 184244 229978
rect 184952 228002 184980 231676
rect 185136 231662 185610 231690
rect 185872 231662 186254 231690
rect 184940 227996 184992 228002
rect 184940 227938 184992 227944
rect 184846 225720 184902 225729
rect 184846 225655 184902 225664
rect 184664 224256 184716 224262
rect 184664 224198 184716 224204
rect 184204 220788 184256 220794
rect 184204 220730 184256 220736
rect 184676 218074 184704 224198
rect 183284 218068 183336 218074
rect 183284 218010 183336 218016
rect 184020 218068 184072 218074
rect 184020 218010 184072 218016
rect 184664 218068 184716 218074
rect 184664 218010 184716 218016
rect 183112 217246 183186 217274
rect 182330 217110 182404 217138
rect 182330 216988 182358 217110
rect 183158 216988 183186 217246
rect 184032 217138 184060 218010
rect 184860 217274 184888 225655
rect 185136 221338 185164 231662
rect 185492 227724 185544 227730
rect 185492 227666 185544 227672
rect 185504 225486 185532 227666
rect 185674 225992 185730 226001
rect 185674 225927 185730 225936
rect 185688 225758 185716 225927
rect 185676 225752 185728 225758
rect 185676 225694 185728 225700
rect 185492 225480 185544 225486
rect 185492 225422 185544 225428
rect 185674 225448 185730 225457
rect 185674 225383 185730 225392
rect 185688 225214 185716 225383
rect 185676 225208 185728 225214
rect 185676 225150 185728 225156
rect 185676 225072 185728 225078
rect 185676 225014 185728 225020
rect 185688 224913 185716 225014
rect 185674 224904 185730 224913
rect 185674 224839 185730 224848
rect 185872 223446 185900 231662
rect 186136 227996 186188 228002
rect 186136 227938 186188 227944
rect 186148 224954 186176 227938
rect 186148 224926 186268 224954
rect 185860 223440 185912 223446
rect 185860 223382 185912 223388
rect 185768 221468 185820 221474
rect 185768 221410 185820 221416
rect 185124 221332 185176 221338
rect 185124 221274 185176 221280
rect 185780 221066 185808 221410
rect 185768 221060 185820 221066
rect 185768 221002 185820 221008
rect 185952 221060 186004 221066
rect 185952 221002 186004 221008
rect 185964 220833 185992 221002
rect 185950 220824 186006 220833
rect 185950 220759 186006 220768
rect 186240 219434 186268 224926
rect 186884 224398 186912 231676
rect 187528 227730 187556 231676
rect 187896 231662 188186 231690
rect 187516 227724 187568 227730
rect 187516 227666 187568 227672
rect 187148 226024 187200 226030
rect 187148 225966 187200 225972
rect 187332 226024 187384 226030
rect 187332 225966 187384 225972
rect 187160 225570 187188 225966
rect 187344 225729 187372 225966
rect 187516 225752 187568 225758
rect 187330 225720 187386 225729
rect 187516 225694 187568 225700
rect 187330 225655 187386 225664
rect 187160 225542 187372 225570
rect 187344 225486 187372 225542
rect 187332 225480 187384 225486
rect 187332 225422 187384 225428
rect 187332 225208 187384 225214
rect 187528 225185 187556 225694
rect 187332 225150 187384 225156
rect 187514 225176 187570 225185
rect 187056 225072 187108 225078
rect 187056 225014 187108 225020
rect 187068 224913 187096 225014
rect 187054 224904 187110 224913
rect 187054 224839 187110 224848
rect 186872 224392 186924 224398
rect 186872 224334 186924 224340
rect 186148 219406 186268 219434
rect 185768 219156 185820 219162
rect 185768 219098 185820 219104
rect 185584 218612 185636 218618
rect 185584 218554 185636 218560
rect 185596 218346 185624 218554
rect 185780 218346 185808 219098
rect 185584 218340 185636 218346
rect 185584 218282 185636 218288
rect 185768 218340 185820 218346
rect 185768 218282 185820 218288
rect 186148 218074 186176 219406
rect 185676 218068 185728 218074
rect 185676 218010 185728 218016
rect 186136 218068 186188 218074
rect 186136 218010 186188 218016
rect 186504 218068 186556 218074
rect 186504 218010 186556 218016
rect 183986 217110 184060 217138
rect 184814 217246 184888 217274
rect 183986 216988 184014 217110
rect 184814 216988 184842 217246
rect 185688 217138 185716 218010
rect 186516 217138 186544 218010
rect 187344 217274 187372 225150
rect 187514 225111 187570 225120
rect 187896 221066 187924 231662
rect 188816 224670 188844 231676
rect 189460 230314 189488 231676
rect 189448 230308 189500 230314
rect 189448 230250 189500 230256
rect 189724 230036 189776 230042
rect 189724 229978 189776 229984
rect 188804 224664 188856 224670
rect 188804 224606 188856 224612
rect 188988 224392 189040 224398
rect 188988 224334 189040 224340
rect 187884 221060 187936 221066
rect 187884 221002 187936 221008
rect 188160 221060 188212 221066
rect 188160 221002 188212 221008
rect 188172 217274 188200 221002
rect 189000 217274 189028 224334
rect 189736 219434 189764 229978
rect 190104 226778 190132 231676
rect 190762 231662 191144 231690
rect 190920 230308 190972 230314
rect 190920 230250 190972 230256
rect 190932 229770 190960 230250
rect 190920 229764 190972 229770
rect 190920 229706 190972 229712
rect 190550 228848 190606 228857
rect 190550 228783 190552 228792
rect 190604 228783 190606 228792
rect 190736 228812 190788 228818
rect 190552 228754 190604 228760
rect 190736 228754 190788 228760
rect 190748 228002 190776 228754
rect 190920 228268 190972 228274
rect 190920 228210 190972 228216
rect 190932 228002 190960 228210
rect 190736 227996 190788 228002
rect 190736 227938 190788 227944
rect 190920 227996 190972 228002
rect 190920 227938 190972 227944
rect 191116 226914 191144 231662
rect 191104 226908 191156 226914
rect 191104 226850 191156 226856
rect 190092 226772 190144 226778
rect 190092 226714 190144 226720
rect 191392 224806 191420 231676
rect 191564 230172 191616 230178
rect 191564 230114 191616 230120
rect 191576 229906 191604 230114
rect 191564 229900 191616 229906
rect 191564 229842 191616 229848
rect 191564 227724 191616 227730
rect 191564 227666 191616 227672
rect 191380 224800 191432 224806
rect 191380 224742 191432 224748
rect 190460 220788 190512 220794
rect 190460 220730 190512 220736
rect 190472 219706 190500 220730
rect 190460 219700 190512 219706
rect 190460 219642 190512 219648
rect 190644 219700 190696 219706
rect 190644 219642 190696 219648
rect 189736 219406 190316 219434
rect 190288 218074 190316 219406
rect 189816 218068 189868 218074
rect 189816 218010 189868 218016
rect 190276 218068 190328 218074
rect 190276 218010 190328 218016
rect 185642 217110 185716 217138
rect 186470 217110 186544 217138
rect 187298 217246 187372 217274
rect 188126 217246 188200 217274
rect 188954 217246 189028 217274
rect 185642 216988 185670 217110
rect 186470 216988 186498 217110
rect 187298 216988 187326 217246
rect 188126 216988 188154 217246
rect 188954 216988 188982 217246
rect 189828 217138 189856 218010
rect 190656 217274 190684 219642
rect 191576 219434 191604 227666
rect 192036 222766 192064 231676
rect 192680 229090 192708 231676
rect 192668 229084 192720 229090
rect 192668 229026 192720 229032
rect 192852 229084 192904 229090
rect 192852 229026 192904 229032
rect 192864 228857 192892 229026
rect 192850 228848 192906 228857
rect 192850 228783 192906 228792
rect 192484 224800 192536 224806
rect 192484 224742 192536 224748
rect 192024 222760 192076 222766
rect 192024 222702 192076 222708
rect 192300 222760 192352 222766
rect 192300 222702 192352 222708
rect 191484 219406 191604 219434
rect 191484 217274 191512 219406
rect 192312 218346 192340 222702
rect 192300 218340 192352 218346
rect 192300 218282 192352 218288
rect 192496 217274 192524 224742
rect 193324 219842 193352 231676
rect 193968 224942 193996 231676
rect 194612 229090 194640 231676
rect 194888 231662 195270 231690
rect 195440 231662 195914 231690
rect 194600 229084 194652 229090
rect 194600 229026 194652 229032
rect 194888 225457 194916 231662
rect 195440 226001 195468 231662
rect 195612 229084 195664 229090
rect 195612 229026 195664 229032
rect 195426 225992 195482 226001
rect 195426 225927 195482 225936
rect 194874 225448 194930 225457
rect 194874 225383 194930 225392
rect 195624 224954 195652 229026
rect 195796 226772 195848 226778
rect 195796 226714 195848 226720
rect 195808 225486 195836 226714
rect 195796 225480 195848 225486
rect 195796 225422 195848 225428
rect 193956 224936 194008 224942
rect 193956 224878 194008 224884
rect 194508 224936 194560 224942
rect 195624 224926 195928 224954
rect 194508 224878 194560 224884
rect 193312 219836 193364 219842
rect 193312 219778 193364 219784
rect 193128 219292 193180 219298
rect 193128 219234 193180 219240
rect 189782 217110 189856 217138
rect 190610 217246 190684 217274
rect 191438 217246 191512 217274
rect 192266 217246 192524 217274
rect 189782 216988 189810 217110
rect 190610 216988 190638 217246
rect 191438 216988 191466 217246
rect 192266 216988 192294 217246
rect 193140 217138 193168 219234
rect 193772 218340 193824 218346
rect 193772 218282 193824 218288
rect 193784 218074 193812 218282
rect 194520 218074 194548 224878
rect 195612 224664 195664 224670
rect 195612 224606 195664 224612
rect 195244 221332 195296 221338
rect 195244 221274 195296 221280
rect 195428 221332 195480 221338
rect 195428 221274 195480 221280
rect 195256 221066 195284 221274
rect 195244 221060 195296 221066
rect 195244 221002 195296 221008
rect 195440 220930 195468 221274
rect 195428 220924 195480 220930
rect 195428 220866 195480 220872
rect 194782 220824 194838 220833
rect 194782 220759 194784 220768
rect 194836 220759 194838 220768
rect 194784 220730 194836 220736
rect 195428 219972 195480 219978
rect 195428 219914 195480 219920
rect 195440 219706 195468 219914
rect 195428 219700 195480 219706
rect 195428 219642 195480 219648
rect 195058 219328 195114 219337
rect 195058 219263 195114 219272
rect 195428 219292 195480 219298
rect 195072 219162 195100 219263
rect 195428 219234 195480 219240
rect 195060 219156 195112 219162
rect 195060 219098 195112 219104
rect 195244 219156 195296 219162
rect 195244 219098 195296 219104
rect 195256 218618 195284 219098
rect 195440 218618 195468 219234
rect 195244 218612 195296 218618
rect 195244 218554 195296 218560
rect 195428 218612 195480 218618
rect 195428 218554 195480 218560
rect 193772 218068 193824 218074
rect 193772 218010 193824 218016
rect 193956 218068 194008 218074
rect 193956 218010 194008 218016
rect 194508 218068 194560 218074
rect 194508 218010 194560 218016
rect 194784 218068 194836 218074
rect 194784 218010 194836 218016
rect 193968 217138 193996 218010
rect 194796 217138 194824 218010
rect 195624 217274 195652 224606
rect 195900 218074 195928 224926
rect 196544 224534 196572 231676
rect 196992 230172 197044 230178
rect 196992 230114 197044 230120
rect 197004 224954 197032 230114
rect 197188 229498 197216 231676
rect 197464 231662 197846 231690
rect 198016 231662 198490 231690
rect 198936 231662 199134 231690
rect 199488 231662 199778 231690
rect 197176 229492 197228 229498
rect 197176 229434 197228 229440
rect 197464 226642 197492 231662
rect 198016 228290 198044 231662
rect 197740 228262 198044 228290
rect 197452 226636 197504 226642
rect 197452 226578 197504 226584
rect 197004 224926 197124 224954
rect 196532 224528 196584 224534
rect 196532 224470 196584 224476
rect 196070 220824 196126 220833
rect 196070 220759 196072 220768
rect 196124 220759 196126 220768
rect 196072 220730 196124 220736
rect 196070 219328 196126 219337
rect 196070 219263 196072 219272
rect 196124 219263 196126 219272
rect 196072 219234 196124 219240
rect 197096 218074 197124 224926
rect 197740 220794 197768 228262
rect 197912 228132 197964 228138
rect 197912 228074 197964 228080
rect 197728 220788 197780 220794
rect 197728 220730 197780 220736
rect 197268 219700 197320 219706
rect 197268 219642 197320 219648
rect 195888 218068 195940 218074
rect 195888 218010 195940 218016
rect 196440 218068 196492 218074
rect 196440 218010 196492 218016
rect 197084 218068 197136 218074
rect 197084 218010 197136 218016
rect 193094 217110 193168 217138
rect 193922 217110 193996 217138
rect 194750 217110 194824 217138
rect 195578 217246 195652 217274
rect 193094 216988 193122 217110
rect 193922 216988 193950 217110
rect 194750 216988 194778 217110
rect 195578 216988 195606 217246
rect 196452 217138 196480 218010
rect 197280 217274 197308 219642
rect 197924 219434 197952 228074
rect 198936 220930 198964 231662
rect 199488 226778 199516 231662
rect 200212 229492 200264 229498
rect 200212 229434 200264 229440
rect 200224 228002 200252 229434
rect 200212 227996 200264 228002
rect 200212 227938 200264 227944
rect 200408 227866 200436 231676
rect 200776 231662 201066 231690
rect 200776 229498 200804 231662
rect 200764 229492 200816 229498
rect 200764 229434 200816 229440
rect 200580 228540 200632 228546
rect 200580 228482 200632 228488
rect 200764 228540 200816 228546
rect 200764 228482 200816 228488
rect 200592 228002 200620 228482
rect 200776 228274 200804 228482
rect 200764 228268 200816 228274
rect 200764 228210 200816 228216
rect 201408 228268 201460 228274
rect 201408 228210 201460 228216
rect 200580 227996 200632 228002
rect 200580 227938 200632 227944
rect 200396 227860 200448 227866
rect 200396 227802 200448 227808
rect 200028 226908 200080 226914
rect 200028 226850 200080 226856
rect 199476 226772 199528 226778
rect 199476 226714 199528 226720
rect 199384 225480 199436 225486
rect 199384 225422 199436 225428
rect 198924 220924 198976 220930
rect 198924 220866 198976 220872
rect 198096 220788 198148 220794
rect 198096 220730 198148 220736
rect 197912 219428 197964 219434
rect 197912 219370 197964 219376
rect 198108 217274 198136 220730
rect 199396 219298 199424 225422
rect 199752 219428 199804 219434
rect 199752 219370 199804 219376
rect 199384 219292 199436 219298
rect 199384 219234 199436 219240
rect 198924 218068 198976 218074
rect 198924 218010 198976 218016
rect 196406 217110 196480 217138
rect 197234 217246 197308 217274
rect 198062 217246 198136 217274
rect 196406 216988 196434 217110
rect 197234 216988 197262 217246
rect 198062 216988 198090 217246
rect 198936 217138 198964 218010
rect 199764 217138 199792 219370
rect 200040 218074 200068 226850
rect 201040 225616 201092 225622
rect 200500 225564 201040 225570
rect 200500 225558 201092 225564
rect 200500 225542 201080 225558
rect 200500 225486 200528 225542
rect 200488 225480 200540 225486
rect 201040 225480 201092 225486
rect 200488 225422 200540 225428
rect 200684 225440 201040 225468
rect 200684 225298 200712 225440
rect 201040 225422 201092 225428
rect 200592 225270 200712 225298
rect 200592 225214 200620 225270
rect 200580 225208 200632 225214
rect 200580 225150 200632 225156
rect 201224 224528 201276 224534
rect 201224 224470 201276 224476
rect 201236 219434 201264 224470
rect 201236 219406 201356 219434
rect 200580 219020 200632 219026
rect 200580 218962 200632 218968
rect 200028 218068 200080 218074
rect 200028 218010 200080 218016
rect 200592 217138 200620 218962
rect 201328 217274 201356 219406
rect 201420 219042 201448 228210
rect 201696 223718 201724 231676
rect 202340 230314 202368 231676
rect 202892 231662 202998 231690
rect 203444 231662 203642 231690
rect 202328 230308 202380 230314
rect 202328 230250 202380 230256
rect 202892 225298 202920 231662
rect 202524 225270 202920 225298
rect 202524 225214 202552 225270
rect 202512 225208 202564 225214
rect 202512 225150 202564 225156
rect 202696 225208 202748 225214
rect 202696 225150 202748 225156
rect 201684 223712 201736 223718
rect 201684 223654 201736 223660
rect 201420 219026 201540 219042
rect 201420 219020 201552 219026
rect 201420 219014 201500 219020
rect 201500 218962 201552 218968
rect 202708 218074 202736 225150
rect 203248 221196 203300 221202
rect 203248 221138 203300 221144
rect 203260 220930 203288 221138
rect 203248 220924 203300 220930
rect 203248 220866 203300 220872
rect 203444 219570 203472 231662
rect 203708 230308 203760 230314
rect 203708 230250 203760 230256
rect 203432 219564 203484 219570
rect 203432 219506 203484 219512
rect 203340 219428 203392 219434
rect 203340 219370 203392 219376
rect 203352 219162 203380 219370
rect 203340 219156 203392 219162
rect 203340 219098 203392 219104
rect 203720 218074 203748 230250
rect 204272 223854 204300 231676
rect 204916 228138 204944 231676
rect 204904 228132 204956 228138
rect 204904 228074 204956 228080
rect 205364 228132 205416 228138
rect 205364 228074 205416 228080
rect 205376 223938 205404 228074
rect 205560 226506 205588 231676
rect 205744 231662 206218 231690
rect 206388 231662 206862 231690
rect 205548 226500 205600 226506
rect 205548 226442 205600 226448
rect 205376 223910 205496 223938
rect 204260 223848 204312 223854
rect 204260 223790 204312 223796
rect 205272 223848 205324 223854
rect 205272 223790 205324 223796
rect 203892 223440 203944 223446
rect 203892 223382 203944 223388
rect 202236 218068 202288 218074
rect 202236 218010 202288 218016
rect 202696 218068 202748 218074
rect 202696 218010 202748 218016
rect 203064 218068 203116 218074
rect 203064 218010 203116 218016
rect 203708 218068 203760 218074
rect 203708 218010 203760 218016
rect 201328 217246 201402 217274
rect 198890 217110 198964 217138
rect 199718 217110 199792 217138
rect 200546 217110 200620 217138
rect 198890 216988 198918 217110
rect 199718 216988 199746 217110
rect 200546 216988 200574 217110
rect 201374 216988 201402 217246
rect 202248 217138 202276 218010
rect 203076 217138 203104 218010
rect 203904 217274 203932 223382
rect 204904 221604 204956 221610
rect 204904 221546 204956 221552
rect 205088 221604 205140 221610
rect 205088 221546 205140 221552
rect 204916 221066 204944 221546
rect 205100 221202 205128 221546
rect 205088 221196 205140 221202
rect 205088 221138 205140 221144
rect 204904 221060 204956 221066
rect 204904 221002 204956 221008
rect 204536 220108 204588 220114
rect 204536 220050 204588 220056
rect 204720 220108 204772 220114
rect 204720 220050 204772 220056
rect 204548 219570 204576 220050
rect 204732 219842 204760 220050
rect 204720 219836 204772 219842
rect 204720 219778 204772 219784
rect 204536 219564 204588 219570
rect 204536 219506 204588 219512
rect 205284 219434 205312 223790
rect 204916 219406 205312 219434
rect 204916 219026 204944 219406
rect 204904 219020 204956 219026
rect 204904 218962 204956 218968
rect 204720 218068 204772 218074
rect 204720 218010 204772 218016
rect 202202 217110 202276 217138
rect 203030 217110 203104 217138
rect 203858 217246 203932 217274
rect 202202 216988 202230 217110
rect 203030 216988 203058 217110
rect 203858 216988 203886 217246
rect 204732 217138 204760 218010
rect 205468 217274 205496 223910
rect 205744 220250 205772 231662
rect 206008 221196 206060 221202
rect 206008 221138 206060 221144
rect 205732 220244 205784 220250
rect 205732 220186 205784 220192
rect 206020 218074 206048 221138
rect 206388 220930 206416 231662
rect 207492 222766 207520 231676
rect 207768 231662 208150 231690
rect 207768 225350 207796 231662
rect 207756 225344 207808 225350
rect 207756 225286 207808 225292
rect 208032 225344 208084 225350
rect 208032 225286 208084 225292
rect 207480 222760 207532 222766
rect 207480 222702 207532 222708
rect 206376 220924 206428 220930
rect 206376 220866 206428 220872
rect 207204 219700 207256 219706
rect 207204 219642 207256 219648
rect 206376 219020 206428 219026
rect 206376 218962 206428 218968
rect 206008 218068 206060 218074
rect 206008 218010 206060 218016
rect 205468 217246 205542 217274
rect 204686 217110 204760 217138
rect 204686 216988 204714 217110
rect 205514 216988 205542 217246
rect 206388 217138 206416 218962
rect 207216 217274 207244 219642
rect 208044 217274 208072 225286
rect 208780 222358 208808 231676
rect 209424 224126 209452 231676
rect 210068 229634 210096 231676
rect 210056 229628 210108 229634
rect 210056 229570 210108 229576
rect 210240 229628 210292 229634
rect 210240 229570 210292 229576
rect 209412 224120 209464 224126
rect 209412 224062 209464 224068
rect 209688 224120 209740 224126
rect 209688 224062 209740 224068
rect 209504 222760 209556 222766
rect 209504 222702 209556 222708
rect 208768 222352 208820 222358
rect 208768 222294 208820 222300
rect 209516 219434 209544 222702
rect 209700 219450 209728 224062
rect 210252 222766 210280 229570
rect 210712 228002 210740 231676
rect 211356 229094 211384 231676
rect 211172 229066 211384 229094
rect 211632 231662 212014 231690
rect 210700 227996 210752 228002
rect 210700 227938 210752 227944
rect 210240 222760 210292 222766
rect 210240 222702 210292 222708
rect 210976 222352 211028 222358
rect 210976 222294 211028 222300
rect 209700 219434 209820 219450
rect 208860 219428 208912 219434
rect 209516 219406 209636 219434
rect 209700 219428 209832 219434
rect 209700 219422 209780 219428
rect 208860 219370 208912 219376
rect 206342 217110 206416 217138
rect 207170 217246 207244 217274
rect 207998 217246 208072 217274
rect 206342 216988 206370 217110
rect 207170 216988 207198 217246
rect 207998 216988 208026 217246
rect 208872 217138 208900 219370
rect 209608 217274 209636 219406
rect 209780 219370 209832 219376
rect 209792 219339 209820 219370
rect 210988 218074 211016 222294
rect 211172 219570 211200 229066
rect 211632 221066 211660 231662
rect 212172 228404 212224 228410
rect 212172 228346 212224 228352
rect 212184 228002 212212 228346
rect 212172 227996 212224 228002
rect 212172 227938 212224 227944
rect 212172 226772 212224 226778
rect 212172 226714 212224 226720
rect 211620 221060 211672 221066
rect 211620 221002 211672 221008
rect 211344 220244 211396 220250
rect 211344 220186 211396 220192
rect 211160 219564 211212 219570
rect 211160 219506 211212 219512
rect 210516 218068 210568 218074
rect 210516 218010 210568 218016
rect 210976 218068 211028 218074
rect 210976 218010 211028 218016
rect 209608 217246 209682 217274
rect 208826 217110 208900 217138
rect 208826 216988 208854 217110
rect 209654 216988 209682 217246
rect 210528 217138 210556 218010
rect 211356 217274 211384 220186
rect 212184 217274 212212 226714
rect 212644 223854 212672 231676
rect 213288 227050 213316 231676
rect 213946 231662 214144 231690
rect 214116 229094 214144 231662
rect 214300 231662 214590 231690
rect 214300 229094 214328 231662
rect 215220 230450 215248 231676
rect 215208 230444 215260 230450
rect 215208 230386 215260 230392
rect 214024 229066 214144 229094
rect 214208 229066 214328 229094
rect 213276 227044 213328 227050
rect 213276 226986 213328 226992
rect 213184 226500 213236 226506
rect 213184 226442 213236 226448
rect 212632 223848 212684 223854
rect 212632 223790 212684 223796
rect 213196 218754 213224 226442
rect 213828 222760 213880 222766
rect 213828 222702 213880 222708
rect 213184 218748 213236 218754
rect 213184 218690 213236 218696
rect 213552 218748 213604 218754
rect 213552 218690 213604 218696
rect 213564 218482 213592 218690
rect 213552 218476 213604 218482
rect 213552 218418 213604 218424
rect 213000 218068 213052 218074
rect 213000 218010 213052 218016
rect 210482 217110 210556 217138
rect 211310 217246 211384 217274
rect 212138 217246 212212 217274
rect 210482 216988 210510 217110
rect 211310 216988 211338 217246
rect 212138 216988 212166 217246
rect 213012 217138 213040 218010
rect 213840 217274 213868 222702
rect 214024 220114 214052 229066
rect 214208 221610 214236 229066
rect 215864 226166 215892 231676
rect 216232 231662 216522 231690
rect 215852 226160 215904 226166
rect 215852 226102 215904 226108
rect 215944 223848 215996 223854
rect 215944 223790 215996 223796
rect 214748 222624 214800 222630
rect 214748 222566 214800 222572
rect 214380 222488 214432 222494
rect 214380 222430 214432 222436
rect 214392 222170 214420 222430
rect 214760 222358 214788 222566
rect 214748 222352 214800 222358
rect 214748 222294 214800 222300
rect 214932 222284 214984 222290
rect 214932 222226 214984 222232
rect 214944 222170 214972 222226
rect 214392 222142 214972 222170
rect 214196 221604 214248 221610
rect 214196 221546 214248 221552
rect 214656 221604 214708 221610
rect 214656 221546 214708 221552
rect 214012 220108 214064 220114
rect 214012 220050 214064 220056
rect 214668 217274 214696 221546
rect 215956 218890 215984 223790
rect 216232 222290 216260 231662
rect 216496 226160 216548 226166
rect 216496 226102 216548 226108
rect 216220 222284 216272 222290
rect 216220 222226 216272 222232
rect 215944 218884 215996 218890
rect 215944 218826 215996 218832
rect 216312 218476 216364 218482
rect 216312 218418 216364 218424
rect 215484 218068 215536 218074
rect 215484 218010 215536 218016
rect 212966 217110 213040 217138
rect 213794 217246 213868 217274
rect 214622 217246 214696 217274
rect 212966 216988 212994 217110
rect 213794 216988 213822 217246
rect 214622 216988 214650 217246
rect 215496 217138 215524 218010
rect 216324 217138 216352 218418
rect 216508 218074 216536 226102
rect 217152 223990 217180 231676
rect 217796 226506 217824 231676
rect 218440 228002 218468 231676
rect 218624 231662 219098 231690
rect 218428 227996 218480 228002
rect 218428 227938 218480 227944
rect 217784 226500 217836 226506
rect 217784 226442 217836 226448
rect 217140 223984 217192 223990
rect 217140 223926 217192 223932
rect 217324 223984 217376 223990
rect 217324 223926 217376 223932
rect 217140 220108 217192 220114
rect 217140 220050 217192 220056
rect 216496 218068 216548 218074
rect 216496 218010 216548 218016
rect 217152 217274 217180 220050
rect 217336 218754 217364 223926
rect 218624 220386 218652 231662
rect 219348 228540 219400 228546
rect 219348 228482 219400 228488
rect 218612 220380 218664 220386
rect 218612 220322 218664 220328
rect 217968 218884 218020 218890
rect 217968 218826 218020 218832
rect 217324 218748 217376 218754
rect 217324 218690 217376 218696
rect 215450 217110 215524 217138
rect 216278 217110 216352 217138
rect 217106 217246 217180 217274
rect 215450 216988 215478 217110
rect 216278 216988 216306 217110
rect 217106 216988 217134 217246
rect 217980 217138 218008 218826
rect 219360 218754 219388 228482
rect 219728 222494 219756 231676
rect 220372 229226 220400 231676
rect 220360 229220 220412 229226
rect 220360 229162 220412 229168
rect 221016 226370 221044 231676
rect 221004 226364 221056 226370
rect 221004 226306 221056 226312
rect 221660 222902 221688 231676
rect 222016 226636 222068 226642
rect 222016 226578 222068 226584
rect 221832 226500 221884 226506
rect 221832 226442 221884 226448
rect 221648 222896 221700 222902
rect 221648 222838 221700 222844
rect 219716 222488 219768 222494
rect 219716 222430 219768 222436
rect 220084 222488 220136 222494
rect 220084 222430 220136 222436
rect 220096 218890 220124 222430
rect 220452 222352 220504 222358
rect 220452 222294 220504 222300
rect 220084 218884 220136 218890
rect 220084 218826 220136 218832
rect 218796 218748 218848 218754
rect 218796 218690 218848 218696
rect 219348 218748 219400 218754
rect 219348 218690 219400 218696
rect 219624 218748 219676 218754
rect 219624 218690 219676 218696
rect 218808 217138 218836 218690
rect 219636 217138 219664 218690
rect 220464 217274 220492 222294
rect 220912 218748 220964 218754
rect 220912 218690 220964 218696
rect 220924 218482 220952 218690
rect 220912 218476 220964 218482
rect 220912 218418 220964 218424
rect 221096 218476 221148 218482
rect 221096 218418 221148 218424
rect 221108 218210 221136 218418
rect 221844 218210 221872 226442
rect 221096 218204 221148 218210
rect 221096 218146 221148 218152
rect 221280 218204 221332 218210
rect 221280 218146 221332 218152
rect 221832 218204 221884 218210
rect 221832 218146 221884 218152
rect 217934 217110 218008 217138
rect 218762 217110 218836 217138
rect 219590 217110 219664 217138
rect 220418 217246 220492 217274
rect 217934 216988 217962 217110
rect 218762 216988 218790 217110
rect 219590 216988 219618 217110
rect 220418 216988 220446 217246
rect 221292 217138 221320 218146
rect 222028 217274 222056 226578
rect 222304 223174 222332 231676
rect 222476 226296 222528 226302
rect 222476 226238 222528 226244
rect 222488 225622 222516 226238
rect 222476 225616 222528 225622
rect 222476 225558 222528 225564
rect 222948 223854 222976 231676
rect 223396 230444 223448 230450
rect 223396 230386 223448 230392
rect 222936 223848 222988 223854
rect 222936 223790 222988 223796
rect 222292 223168 222344 223174
rect 222292 223110 222344 223116
rect 223408 218210 223436 230386
rect 223592 225078 223620 231676
rect 224236 229094 224264 231676
rect 224052 229066 224264 229094
rect 224512 231662 224894 231690
rect 223580 225072 223632 225078
rect 223580 225014 223632 225020
rect 224052 223310 224080 229066
rect 224224 226024 224276 226030
rect 224224 225966 224276 225972
rect 224236 225622 224264 225966
rect 224224 225616 224276 225622
rect 224224 225558 224276 225564
rect 224040 223304 224092 223310
rect 224040 223246 224092 223252
rect 224224 223168 224276 223174
rect 224224 223110 224276 223116
rect 224236 218482 224264 223110
rect 224512 221746 224540 231662
rect 225524 226302 225552 231676
rect 226168 228410 226196 231676
rect 226812 229094 226840 231676
rect 226720 229066 226840 229094
rect 226156 228404 226208 228410
rect 226156 228346 226208 228352
rect 226340 228404 226392 228410
rect 226340 228346 226392 228352
rect 226156 227996 226208 228002
rect 226156 227938 226208 227944
rect 225696 227860 225748 227866
rect 225696 227802 225748 227808
rect 225512 226296 225564 226302
rect 225512 226238 225564 226244
rect 224868 225072 224920 225078
rect 224868 225014 224920 225020
rect 224500 221740 224552 221746
rect 224500 221682 224552 221688
rect 224224 218476 224276 218482
rect 224224 218418 224276 218424
rect 224592 218476 224644 218482
rect 224592 218418 224644 218424
rect 222936 218204 222988 218210
rect 222936 218146 222988 218152
rect 223396 218204 223448 218210
rect 223396 218146 223448 218152
rect 223764 218204 223816 218210
rect 223764 218146 223816 218152
rect 222028 217246 222102 217274
rect 221246 217110 221320 217138
rect 221246 216988 221274 217110
rect 222074 216988 222102 217246
rect 222948 217138 222976 218146
rect 223776 217138 223804 218146
rect 224604 217138 224632 218418
rect 224880 218210 224908 225014
rect 225420 219428 225472 219434
rect 225420 219370 225472 219376
rect 224868 218204 224920 218210
rect 224868 218146 224920 218152
rect 225432 217138 225460 219370
rect 225708 218482 225736 227802
rect 226168 219434 226196 227938
rect 226352 227866 226380 228346
rect 226340 227860 226392 227866
rect 226340 227802 226392 227808
rect 226720 223582 226748 229066
rect 227456 227322 227484 231676
rect 227444 227316 227496 227322
rect 227444 227258 227496 227264
rect 226892 227044 226944 227050
rect 226892 226986 226944 226992
rect 226708 223576 226760 223582
rect 226708 223518 226760 223524
rect 226156 219428 226208 219434
rect 226156 219370 226208 219376
rect 226904 219298 226932 226986
rect 228100 223990 228128 231676
rect 228744 227186 228772 231676
rect 229296 231662 229402 231690
rect 229664 231662 230046 231690
rect 228732 227180 228784 227186
rect 228732 227122 228784 227128
rect 229054 227044 229106 227050
rect 229054 226986 229106 226992
rect 229066 226930 229094 226986
rect 229020 226902 229094 226930
rect 229020 226506 229048 226902
rect 229008 226500 229060 226506
rect 229008 226442 229060 226448
rect 228732 226296 228784 226302
rect 228732 226238 228784 226244
rect 228088 223984 228140 223990
rect 228088 223926 228140 223932
rect 227076 221740 227128 221746
rect 227076 221682 227128 221688
rect 226892 219292 226944 219298
rect 226892 219234 226944 219240
rect 225696 218476 225748 218482
rect 225696 218418 225748 218424
rect 226248 218476 226300 218482
rect 226248 218418 226300 218424
rect 226260 217138 226288 218418
rect 227088 217138 227116 221682
rect 228548 219428 228600 219434
rect 228548 219370 228600 219376
rect 228560 218754 228588 219370
rect 228548 218748 228600 218754
rect 228548 218690 228600 218696
rect 227904 218204 227956 218210
rect 227904 218146 227956 218152
rect 227916 217138 227944 218146
rect 228744 217274 228772 226238
rect 229296 220522 229324 231662
rect 229664 221882 229692 231662
rect 230676 229362 230704 231676
rect 231124 229492 231176 229498
rect 231124 229434 231176 229440
rect 230664 229356 230716 229362
rect 230664 229298 230716 229304
rect 229652 221876 229704 221882
rect 229652 221818 229704 221824
rect 230388 221876 230440 221882
rect 230388 221818 230440 221824
rect 229284 220516 229336 220522
rect 229284 220458 229336 220464
rect 229744 220380 229796 220386
rect 229744 220322 229796 220328
rect 229376 219292 229428 219298
rect 229376 219234 229428 219240
rect 229388 218346 229416 219234
rect 229376 218340 229428 218346
rect 229376 218282 229428 218288
rect 229560 218340 229612 218346
rect 229560 218282 229612 218288
rect 222902 217110 222976 217138
rect 223730 217110 223804 217138
rect 224558 217110 224632 217138
rect 225386 217110 225460 217138
rect 226214 217110 226288 217138
rect 227042 217110 227116 217138
rect 227870 217110 227944 217138
rect 228698 217246 228772 217274
rect 222902 216988 222930 217110
rect 223730 216988 223758 217110
rect 224558 216988 224586 217110
rect 225386 216988 225414 217110
rect 226214 216988 226242 217110
rect 227042 216988 227070 217110
rect 227870 216988 227898 217110
rect 228698 216988 228726 217246
rect 229572 217138 229600 218282
rect 229756 218210 229784 220322
rect 229928 218884 229980 218890
rect 229928 218826 229980 218832
rect 229940 218482 229968 218826
rect 229928 218476 229980 218482
rect 229928 218418 229980 218424
rect 229744 218204 229796 218210
rect 229744 218146 229796 218152
rect 230400 217138 230428 221818
rect 231136 218346 231164 229434
rect 231320 228682 231348 231676
rect 231308 228676 231360 228682
rect 231308 228618 231360 228624
rect 231964 227458 231992 231676
rect 232148 231662 232622 231690
rect 231952 227452 232004 227458
rect 231952 227394 232004 227400
rect 231308 223984 231360 223990
rect 231308 223926 231360 223932
rect 231124 218340 231176 218346
rect 231124 218282 231176 218288
rect 231320 217274 231348 223926
rect 231952 222896 232004 222902
rect 231952 222838 232004 222844
rect 229526 217110 229600 217138
rect 230354 217110 230428 217138
rect 231182 217246 231348 217274
rect 229526 216988 229554 217110
rect 230354 216988 230382 217110
rect 231182 216988 231210 217246
rect 231964 217138 231992 222838
rect 232148 221474 232176 231662
rect 233252 227322 233280 231676
rect 233240 227316 233292 227322
rect 233240 227258 233292 227264
rect 232504 226500 232556 226506
rect 232504 226442 232556 226448
rect 232136 221468 232188 221474
rect 232136 221410 232188 221416
rect 232516 219434 232544 226442
rect 233896 226030 233924 231676
rect 234080 231662 234554 231690
rect 234816 231662 235198 231690
rect 233884 226024 233936 226030
rect 233884 225966 233936 225972
rect 234080 220658 234108 231662
rect 234528 227316 234580 227322
rect 234528 227258 234580 227264
rect 234344 225616 234396 225622
rect 234344 225558 234396 225564
rect 234356 224954 234384 225558
rect 234356 224926 234476 224954
rect 234068 220652 234120 220658
rect 234068 220594 234120 220600
rect 232504 219428 232556 219434
rect 232504 219370 232556 219376
rect 233700 219428 233752 219434
rect 233700 219370 233752 219376
rect 232872 218340 232924 218346
rect 232872 218282 232924 218288
rect 232884 217138 232912 218282
rect 233712 217138 233740 219370
rect 234448 217274 234476 224926
rect 234540 219434 234568 227258
rect 234816 223038 234844 231662
rect 235828 229770 235856 231676
rect 235816 229764 235868 229770
rect 235816 229706 235868 229712
rect 236472 227594 236500 231676
rect 236920 229764 236972 229770
rect 236920 229706 236972 229712
rect 236460 227588 236512 227594
rect 236460 227530 236512 227536
rect 235908 227180 235960 227186
rect 235908 227122 235960 227128
rect 234804 223032 234856 223038
rect 234804 222974 234856 222980
rect 235172 223032 235224 223038
rect 235172 222974 235224 222980
rect 234540 219428 234672 219434
rect 234540 219406 234620 219428
rect 234620 219370 234672 219376
rect 234804 219428 234856 219434
rect 234804 219370 234856 219376
rect 234816 218346 234844 219370
rect 235184 219298 235212 222974
rect 235172 219292 235224 219298
rect 235172 219234 235224 219240
rect 234804 218340 234856 218346
rect 234804 218282 234856 218288
rect 235920 218210 235948 227122
rect 236932 218210 236960 229706
rect 237116 228954 237144 231676
rect 237576 231662 237774 231690
rect 237104 228948 237156 228954
rect 237104 228890 237156 228896
rect 237576 222018 237604 231662
rect 238404 223174 238432 231676
rect 239048 225894 239076 231676
rect 239404 228676 239456 228682
rect 239404 228618 239456 228624
rect 239036 225888 239088 225894
rect 239036 225830 239088 225836
rect 238668 223848 238720 223854
rect 238668 223790 238720 223796
rect 238392 223168 238444 223174
rect 238392 223110 238444 223116
rect 237564 222012 237616 222018
rect 237564 221954 237616 221960
rect 237104 221060 237156 221066
rect 237104 221002 237156 221008
rect 235356 218204 235408 218210
rect 235356 218146 235408 218152
rect 235908 218204 235960 218210
rect 235908 218146 235960 218152
rect 236184 218204 236236 218210
rect 236184 218146 236236 218152
rect 236920 218204 236972 218210
rect 236920 218146 236972 218152
rect 234448 217246 234522 217274
rect 231964 217110 232038 217138
rect 232010 216988 232038 217110
rect 232838 217110 232912 217138
rect 233666 217110 233740 217138
rect 232838 216988 232866 217110
rect 233666 216988 233694 217110
rect 234494 216988 234522 217246
rect 235368 217138 235396 218146
rect 236196 217138 236224 218146
rect 237116 217274 237144 221002
rect 237840 219292 237892 219298
rect 237840 219234 237892 219240
rect 235322 217110 235396 217138
rect 236150 217110 236224 217138
rect 236978 217246 237144 217274
rect 235322 216988 235350 217110
rect 236150 216988 236178 217110
rect 236978 216988 237006 217246
rect 237852 217138 237880 219234
rect 238680 217274 238708 223790
rect 239416 219298 239444 228618
rect 239692 224262 239720 231676
rect 240152 231662 240350 231690
rect 239680 224256 239732 224262
rect 239680 224198 239732 224204
rect 240152 222154 240180 231662
rect 240980 229906 241008 231676
rect 240968 229900 241020 229906
rect 240968 229842 241020 229848
rect 241624 228818 241652 231676
rect 241612 228812 241664 228818
rect 241612 228754 241664 228760
rect 242268 225486 242296 231676
rect 242716 227792 242768 227798
rect 242716 227734 242768 227740
rect 242256 225480 242308 225486
rect 242256 225422 242308 225428
rect 241980 224256 242032 224262
rect 241980 224198 242032 224204
rect 240140 222148 240192 222154
rect 240140 222090 240192 222096
rect 241152 221468 241204 221474
rect 241152 221410 241204 221416
rect 240324 220516 240376 220522
rect 240324 220458 240376 220464
rect 239404 219292 239456 219298
rect 239404 219234 239456 219240
rect 239496 218476 239548 218482
rect 239496 218418 239548 218424
rect 237806 217110 237880 217138
rect 238634 217246 238708 217274
rect 237806 216988 237834 217110
rect 238634 216988 238662 217246
rect 239508 217138 239536 218418
rect 240336 217274 240364 220458
rect 241164 217274 241192 221410
rect 241992 217274 242020 224198
rect 239462 217110 239536 217138
rect 240290 217246 240364 217274
rect 241118 217246 241192 217274
rect 241946 217246 242020 217274
rect 242728 217274 242756 227734
rect 242912 225758 242940 231676
rect 243280 231662 243570 231690
rect 243832 231662 244214 231690
rect 244476 231662 244858 231690
rect 245120 231662 245502 231690
rect 242900 225752 242952 225758
rect 242900 225694 242952 225700
rect 243280 223038 243308 231662
rect 243452 226024 243504 226030
rect 243452 225966 243504 225972
rect 243268 223032 243320 223038
rect 243268 222974 243320 222980
rect 243464 218618 243492 225966
rect 243832 224398 243860 231662
rect 243820 224392 243872 224398
rect 243820 224334 243872 224340
rect 243636 222012 243688 222018
rect 243636 221954 243688 221960
rect 243452 218612 243504 218618
rect 243452 218554 243504 218560
rect 243648 217274 243676 221954
rect 244476 219978 244504 231662
rect 245120 221338 245148 231662
rect 246132 230042 246160 231676
rect 246120 230036 246172 230042
rect 246120 229978 246172 229984
rect 245660 229900 245712 229906
rect 245660 229842 245712 229848
rect 245672 227798 245700 229842
rect 246304 228812 246356 228818
rect 246304 228754 246356 228760
rect 245660 227792 245712 227798
rect 245660 227734 245712 227740
rect 245292 223168 245344 223174
rect 245292 223110 245344 223116
rect 245108 221332 245160 221338
rect 245108 221274 245160 221280
rect 244464 219972 244516 219978
rect 244464 219914 244516 219920
rect 244464 218068 244516 218074
rect 244464 218010 244516 218016
rect 242728 217246 242802 217274
rect 239462 216988 239490 217110
rect 240290 216988 240318 217246
rect 241118 216988 241146 217246
rect 241946 216988 241974 217246
rect 242774 216988 242802 217246
rect 243602 217246 243676 217274
rect 243602 216988 243630 217246
rect 244476 217138 244504 218010
rect 245304 217274 245332 223110
rect 246120 219292 246172 219298
rect 246120 219234 246172 219240
rect 244430 217110 244504 217138
rect 245258 217246 245332 217274
rect 244430 216988 244458 217110
rect 245258 216988 245286 217246
rect 246132 217138 246160 219234
rect 246316 219162 246344 228754
rect 246776 224806 246804 231676
rect 247420 224942 247448 231676
rect 248064 227662 248092 231676
rect 248052 227656 248104 227662
rect 248052 227598 248104 227604
rect 248236 227452 248288 227458
rect 248236 227394 248288 227400
rect 247408 224936 247460 224942
rect 247408 224878 247460 224884
rect 246764 224800 246816 224806
rect 246764 224742 246816 224748
rect 247592 224800 247644 224806
rect 247592 224742 247644 224748
rect 246948 224392 247000 224398
rect 246948 224334 247000 224340
rect 246304 219156 246356 219162
rect 246304 219098 246356 219104
rect 246960 217274 246988 224334
rect 247604 218074 247632 224742
rect 248248 218074 248276 227394
rect 248708 226030 248736 231676
rect 248892 231662 249366 231690
rect 249904 231662 250010 231690
rect 248696 226024 248748 226030
rect 248696 225966 248748 225972
rect 248892 224670 248920 231662
rect 249708 225888 249760 225894
rect 249708 225830 249760 225836
rect 248880 224664 248932 224670
rect 248880 224606 248932 224612
rect 249064 224664 249116 224670
rect 249064 224606 249116 224612
rect 249076 218210 249104 224606
rect 249064 218204 249116 218210
rect 249064 218146 249116 218152
rect 249432 218204 249484 218210
rect 249432 218146 249484 218152
rect 247592 218068 247644 218074
rect 247592 218010 247644 218016
rect 247776 218068 247828 218074
rect 247776 218010 247828 218016
rect 248236 218068 248288 218074
rect 248236 218010 248288 218016
rect 248604 218068 248656 218074
rect 248604 218010 248656 218016
rect 246086 217110 246160 217138
rect 246914 217246 246988 217274
rect 246086 216988 246114 217110
rect 246914 216988 246942 217246
rect 247788 217138 247816 218010
rect 248616 217138 248644 218010
rect 249444 217138 249472 218146
rect 249720 218074 249748 225830
rect 249904 219842 249932 231662
rect 250640 229090 250668 231676
rect 251284 230178 251312 231676
rect 251272 230172 251324 230178
rect 251272 230114 251324 230120
rect 251732 230036 251784 230042
rect 251732 229978 251784 229984
rect 250628 229084 250680 229090
rect 250628 229026 250680 229032
rect 251088 228948 251140 228954
rect 251088 228890 251140 228896
rect 250904 223032 250956 223038
rect 250904 222974 250956 222980
rect 249892 219836 249944 219842
rect 249892 219778 249944 219784
rect 250916 219434 250944 222974
rect 250916 219406 251036 219434
rect 249708 218068 249760 218074
rect 249708 218010 249760 218016
rect 250260 218068 250312 218074
rect 250260 218010 250312 218016
rect 250272 217138 250300 218010
rect 251008 217274 251036 219406
rect 251100 218090 251128 228890
rect 251744 218210 251772 229978
rect 251928 226914 251956 231676
rect 252572 228274 252600 231676
rect 252756 231662 253230 231690
rect 252560 228268 252612 228274
rect 252560 228210 252612 228216
rect 252468 227588 252520 227594
rect 252468 227530 252520 227536
rect 251916 226908 251968 226914
rect 251916 226850 251968 226856
rect 251732 218204 251784 218210
rect 251732 218146 251784 218152
rect 251100 218074 251220 218090
rect 252480 218074 252508 227530
rect 252756 220794 252784 231662
rect 253860 228818 253888 231676
rect 253848 228812 253900 228818
rect 253848 228754 253900 228760
rect 254504 225214 254532 231676
rect 254872 231662 255162 231690
rect 254492 225208 254544 225214
rect 254492 225150 254544 225156
rect 254872 223446 254900 231662
rect 255136 228812 255188 228818
rect 255136 228754 255188 228760
rect 254860 223440 254912 223446
rect 254860 223382 254912 223388
rect 252744 220788 252796 220794
rect 252744 220730 252796 220736
rect 253572 220788 253624 220794
rect 253572 220730 253624 220736
rect 252744 218612 252796 218618
rect 252744 218554 252796 218560
rect 251100 218068 251232 218074
rect 251100 218062 251180 218068
rect 251180 218010 251232 218016
rect 251916 218068 251968 218074
rect 251916 218010 251968 218016
rect 252468 218068 252520 218074
rect 252468 218010 252520 218016
rect 251008 217246 251082 217274
rect 247742 217110 247816 217138
rect 248570 217110 248644 217138
rect 249398 217110 249472 217138
rect 250226 217110 250300 217138
rect 247742 216988 247770 217110
rect 248570 216988 248598 217110
rect 249398 216988 249426 217110
rect 250226 216988 250254 217110
rect 251054 216988 251082 217246
rect 251928 217138 251956 218010
rect 252756 217138 252784 218554
rect 253584 217274 253612 220730
rect 254400 220652 254452 220658
rect 254400 220594 254452 220600
rect 251882 217110 251956 217138
rect 252710 217110 252784 217138
rect 253538 217246 253612 217274
rect 251882 216988 251910 217110
rect 252710 216988 252738 217110
rect 253538 216988 253566 217246
rect 254412 217138 254440 220594
rect 255148 217274 255176 228754
rect 255792 224534 255820 231676
rect 256436 230314 256464 231676
rect 256424 230308 256476 230314
rect 256424 230250 256476 230256
rect 257080 228138 257108 231676
rect 257264 231662 257738 231690
rect 258184 231662 258382 231690
rect 257068 228132 257120 228138
rect 257068 228074 257120 228080
rect 255964 227792 256016 227798
rect 255964 227734 256016 227740
rect 255780 224528 255832 224534
rect 255780 224470 255832 224476
rect 255976 221082 256004 227734
rect 255884 221054 256004 221082
rect 255884 219026 255912 221054
rect 256056 220924 256108 220930
rect 256056 220866 256108 220872
rect 255872 219020 255924 219026
rect 255872 218962 255924 218968
rect 255148 217246 255222 217274
rect 254366 217110 254440 217138
rect 254366 216988 254394 217110
rect 255194 216988 255222 217246
rect 256068 217138 256096 220866
rect 256884 219972 256936 219978
rect 256884 219914 256936 219920
rect 256896 217138 256924 219914
rect 257264 219706 257292 231662
rect 258184 229094 258212 231662
rect 258184 229066 258396 229094
rect 257712 225752 257764 225758
rect 257712 225694 257764 225700
rect 257252 219700 257304 219706
rect 257252 219642 257304 219648
rect 257724 217274 257752 225694
rect 258368 221202 258396 229066
rect 259012 227798 259040 231676
rect 259276 229084 259328 229090
rect 259276 229026 259328 229032
rect 259000 227792 259052 227798
rect 259000 227734 259052 227740
rect 258724 221876 258776 221882
rect 258724 221818 258776 221824
rect 258736 221610 258764 221818
rect 258540 221604 258592 221610
rect 258540 221546 258592 221552
rect 258724 221604 258776 221610
rect 258724 221546 258776 221552
rect 258552 221338 258580 221546
rect 258540 221332 258592 221338
rect 258540 221274 258592 221280
rect 258356 221196 258408 221202
rect 258356 221138 258408 221144
rect 259288 219162 259316 229026
rect 259656 224126 259684 231676
rect 259644 224120 259696 224126
rect 259644 224062 259696 224068
rect 260104 223440 260156 223446
rect 260104 223382 260156 223388
rect 258540 219156 258592 219162
rect 258540 219098 258592 219104
rect 259276 219156 259328 219162
rect 259276 219098 259328 219104
rect 259460 219156 259512 219162
rect 259460 219098 259512 219104
rect 256022 217110 256096 217138
rect 256850 217110 256924 217138
rect 257678 217246 257752 217274
rect 256022 216988 256050 217110
rect 256850 216988 256878 217110
rect 257678 216988 257706 217246
rect 258552 217138 258580 219098
rect 259276 219020 259328 219026
rect 259276 218962 259328 218968
rect 258506 217110 258580 217138
rect 259288 217138 259316 218962
rect 259472 218618 259500 219098
rect 259460 218612 259512 218618
rect 259460 218554 259512 218560
rect 260116 217138 260144 223382
rect 260300 222630 260328 231676
rect 260944 225350 260972 231676
rect 261392 230308 261444 230314
rect 261392 230250 261444 230256
rect 260932 225344 260984 225350
rect 260932 225286 260984 225292
rect 260288 222624 260340 222630
rect 260288 222566 260340 222572
rect 261024 222148 261076 222154
rect 261024 222090 261076 222096
rect 261036 217138 261064 222090
rect 261404 220930 261432 230250
rect 261588 229634 261616 231676
rect 261576 229628 261628 229634
rect 261576 229570 261628 229576
rect 262232 226778 262260 231676
rect 262220 226772 262272 226778
rect 262220 226714 262272 226720
rect 261852 224528 261904 224534
rect 261852 224470 261904 224476
rect 261392 220924 261444 220930
rect 261392 220866 261444 220872
rect 261864 217138 261892 224470
rect 262876 222766 262904 231676
rect 263060 231662 263534 231690
rect 263888 231662 264178 231690
rect 262864 222760 262916 222766
rect 262864 222702 262916 222708
rect 263060 220250 263088 231662
rect 263888 224670 263916 231662
rect 264808 226166 264836 231676
rect 265176 231662 265466 231690
rect 265728 231662 266110 231690
rect 264796 226160 264848 226166
rect 264796 226102 264848 226108
rect 264152 224936 264204 224942
rect 264152 224878 264204 224884
rect 263876 224664 263928 224670
rect 263876 224606 263928 224612
rect 263508 222760 263560 222766
rect 263508 222702 263560 222708
rect 263048 220244 263100 220250
rect 263048 220186 263100 220192
rect 263324 220244 263376 220250
rect 263324 220186 263376 220192
rect 262680 218068 262732 218074
rect 262680 218010 262732 218016
rect 262692 217138 262720 218010
rect 263336 217274 263364 220186
rect 263520 218090 263548 222702
rect 264164 218754 264192 224878
rect 264796 223304 264848 223310
rect 264796 223246 264848 223252
rect 264152 218748 264204 218754
rect 264152 218690 264204 218696
rect 263520 218074 263640 218090
rect 264808 218074 264836 223246
rect 265176 220114 265204 231662
rect 265728 221338 265756 231662
rect 266740 226506 266768 231676
rect 267384 228546 267412 231676
rect 267372 228540 267424 228546
rect 267372 228482 267424 228488
rect 267556 228540 267608 228546
rect 267556 228482 267608 228488
rect 266728 226500 266780 226506
rect 266728 226442 266780 226448
rect 266268 226160 266320 226166
rect 266268 226102 266320 226108
rect 265716 221332 265768 221338
rect 265716 221274 265768 221280
rect 265164 220108 265216 220114
rect 265164 220050 265216 220056
rect 265992 218748 266044 218754
rect 265992 218690 266044 218696
rect 263520 218068 263652 218074
rect 263520 218062 263600 218068
rect 263600 218010 263652 218016
rect 264336 218068 264388 218074
rect 264336 218010 264388 218016
rect 264796 218068 264848 218074
rect 264796 218010 264848 218016
rect 265164 218068 265216 218074
rect 265164 218010 265216 218016
rect 263336 217246 263502 217274
rect 259288 217110 259362 217138
rect 260116 217110 260190 217138
rect 258506 216988 258534 217110
rect 259334 216988 259362 217110
rect 260162 216988 260190 217110
rect 260990 217110 261064 217138
rect 261818 217110 261892 217138
rect 262646 217110 262720 217138
rect 260990 216988 261018 217110
rect 261818 216988 261846 217110
rect 262646 216988 262674 217110
rect 263474 216988 263502 217246
rect 264348 217138 264376 218010
rect 265176 217138 265204 218010
rect 266004 217274 266032 218690
rect 266280 218074 266308 226102
rect 266268 218068 266320 218074
rect 266268 218010 266320 218016
rect 266820 218068 266872 218074
rect 266820 218010 266872 218016
rect 264302 217110 264376 217138
rect 265130 217110 265204 217138
rect 265958 217246 266032 217274
rect 264302 216988 264330 217110
rect 265130 216988 265158 217110
rect 265958 216988 265986 217246
rect 266832 217138 266860 218010
rect 267568 217274 267596 228482
rect 267694 226024 267746 226030
rect 267660 225972 267694 225978
rect 267660 225966 267746 225972
rect 267660 225950 267734 225966
rect 267660 218090 267688 225950
rect 268028 222358 268056 231676
rect 268672 222494 268700 231676
rect 269316 224942 269344 231676
rect 269960 226642 269988 231676
rect 270132 227724 270184 227730
rect 270132 227666 270184 227672
rect 269948 226636 270000 226642
rect 269948 226578 270000 226584
rect 269304 224936 269356 224942
rect 269304 224878 269356 224884
rect 269028 223576 269080 223582
rect 269028 223518 269080 223524
rect 268660 222488 268712 222494
rect 268660 222430 268712 222436
rect 268016 222352 268068 222358
rect 268016 222294 268068 222300
rect 267832 221876 267884 221882
rect 267832 221818 267884 221824
rect 267844 218618 267872 221818
rect 267832 218612 267884 218618
rect 267832 218554 267884 218560
rect 267660 218074 267734 218090
rect 269040 218074 269068 223518
rect 269304 218204 269356 218210
rect 269304 218146 269356 218152
rect 267660 218068 267746 218074
rect 267660 218062 267694 218068
rect 267694 218010 267746 218016
rect 268476 218068 268528 218074
rect 268476 218010 268528 218016
rect 269028 218068 269080 218074
rect 269028 218010 269080 218016
rect 267568 217246 267642 217274
rect 266786 217110 266860 217138
rect 266786 216988 266814 217110
rect 267614 216988 267642 217246
rect 268488 217138 268516 218010
rect 269316 217138 269344 218146
rect 270144 217274 270172 227666
rect 270604 225078 270632 231676
rect 271248 227050 271276 231676
rect 271892 230450 271920 231676
rect 271880 230444 271932 230450
rect 271880 230386 271932 230392
rect 272536 228002 272564 231676
rect 272720 231662 273194 231690
rect 272524 227996 272576 228002
rect 272524 227938 272576 227944
rect 271236 227044 271288 227050
rect 271236 226986 271288 226992
rect 271788 227044 271840 227050
rect 271788 226986 271840 226992
rect 270592 225072 270644 225078
rect 270592 225014 270644 225020
rect 271604 224664 271656 224670
rect 271604 224606 271656 224612
rect 271616 218074 271644 224606
rect 270960 218068 271012 218074
rect 270960 218010 271012 218016
rect 271604 218068 271656 218074
rect 271604 218010 271656 218016
rect 268442 217110 268516 217138
rect 269270 217110 269344 217138
rect 270098 217246 270172 217274
rect 268442 216988 268470 217110
rect 269270 216988 269298 217110
rect 270098 216988 270126 217246
rect 270972 217138 271000 218010
rect 271800 217274 271828 226986
rect 272432 226908 272484 226914
rect 272432 226850 272484 226856
rect 272444 218482 272472 226850
rect 272720 221746 272748 231662
rect 273824 228410 273852 231676
rect 274008 231662 274482 231690
rect 273812 228404 273864 228410
rect 273812 228346 273864 228352
rect 274008 221882 274036 231662
rect 274180 230444 274232 230450
rect 274180 230386 274232 230392
rect 273996 221876 274048 221882
rect 273996 221818 274048 221824
rect 272708 221740 272760 221746
rect 272708 221682 272760 221688
rect 273444 221332 273496 221338
rect 273444 221274 273496 221280
rect 272616 218612 272668 218618
rect 272616 218554 272668 218560
rect 272432 218476 272484 218482
rect 272432 218418 272484 218424
rect 270926 217110 271000 217138
rect 271754 217246 271828 217274
rect 270926 216988 270954 217110
rect 271754 216988 271782 217246
rect 272628 217138 272656 218554
rect 273456 217274 273484 221274
rect 274192 219434 274220 230386
rect 275112 226302 275140 231676
rect 275296 231662 275770 231690
rect 276124 231662 276414 231690
rect 275100 226296 275152 226302
rect 275100 226238 275152 226244
rect 275100 221740 275152 221746
rect 275100 221682 275152 221688
rect 273916 219406 274220 219434
rect 273916 218210 273944 219406
rect 274272 218884 274324 218890
rect 274272 218826 274324 218832
rect 273904 218204 273956 218210
rect 273904 218146 273956 218152
rect 272582 217110 272656 217138
rect 273410 217246 273484 217274
rect 272582 216988 272610 217110
rect 273410 216988 273438 217246
rect 274284 217138 274312 218826
rect 275112 217274 275140 221682
rect 275296 221610 275324 231662
rect 275836 225004 275888 225010
rect 275836 224946 275888 224952
rect 275284 221604 275336 221610
rect 275284 221546 275336 221552
rect 274238 217110 274312 217138
rect 275066 217246 275140 217274
rect 275848 217274 275876 224946
rect 276124 220386 276152 231662
rect 276848 230172 276900 230178
rect 276848 230114 276900 230120
rect 276860 225010 276888 230114
rect 277044 229498 277072 231676
rect 277032 229492 277084 229498
rect 277032 229434 277084 229440
rect 277216 228268 277268 228274
rect 277216 228210 277268 228216
rect 276848 225004 276900 225010
rect 276848 224946 276900 224952
rect 276112 220380 276164 220386
rect 276112 220322 276164 220328
rect 277228 218074 277256 228210
rect 277688 222902 277716 231676
rect 278332 227322 278360 231676
rect 278320 227316 278372 227322
rect 278320 227258 278372 227264
rect 278504 226296 278556 226302
rect 278504 226238 278556 226244
rect 277676 222896 277728 222902
rect 277676 222838 277728 222844
rect 278320 221604 278372 221610
rect 278320 221546 278372 221552
rect 276756 218068 276808 218074
rect 276756 218010 276808 218016
rect 277216 218068 277268 218074
rect 277216 218010 277268 218016
rect 277584 218068 277636 218074
rect 277584 218010 277636 218016
rect 275848 217246 275922 217274
rect 274238 216988 274266 217110
rect 275066 216988 275094 217246
rect 275894 216988 275922 217246
rect 276768 217138 276796 218010
rect 277596 217138 277624 218010
rect 278332 217274 278360 221546
rect 278516 218074 278544 226238
rect 278976 223990 279004 231676
rect 279252 231662 279634 231690
rect 278964 223984 279016 223990
rect 278964 223926 279016 223932
rect 279252 219502 279280 231662
rect 280264 227186 280292 231676
rect 280448 231662 280922 231690
rect 280252 227180 280304 227186
rect 280252 227122 280304 227128
rect 280448 221066 280476 231662
rect 280712 227316 280764 227322
rect 280712 227258 280764 227264
rect 280436 221060 280488 221066
rect 280436 221002 280488 221008
rect 280068 220380 280120 220386
rect 280068 220322 280120 220328
rect 279240 219496 279292 219502
rect 279240 219438 279292 219444
rect 279240 218476 279292 218482
rect 279240 218418 279292 218424
rect 278504 218068 278556 218074
rect 278504 218010 278556 218016
rect 278332 217246 278406 217274
rect 276722 217110 276796 217138
rect 277550 217110 277624 217138
rect 276722 216988 276750 217110
rect 277550 216988 277578 217110
rect 278378 216988 278406 217246
rect 279252 217138 279280 218418
rect 280080 217274 280108 220322
rect 280724 218890 280752 227258
rect 281552 225622 281580 231676
rect 282196 229770 282224 231676
rect 282184 229764 282236 229770
rect 282184 229706 282236 229712
rect 282840 229094 282868 231676
rect 282380 229066 282868 229094
rect 283024 231662 283498 231690
rect 281540 225616 281592 225622
rect 281540 225558 281592 225564
rect 282380 223854 282408 229066
rect 282736 225004 282788 225010
rect 282736 224946 282788 224952
rect 282552 224256 282604 224262
rect 282552 224198 282604 224204
rect 282368 223848 282420 223854
rect 282368 223790 282420 223796
rect 280896 220108 280948 220114
rect 280896 220050 280948 220056
rect 280712 218884 280764 218890
rect 280712 218826 280764 218832
rect 280908 217274 280936 220050
rect 281080 218884 281132 218890
rect 281080 218826 281132 218832
rect 281092 218482 281120 218826
rect 281080 218476 281132 218482
rect 281080 218418 281132 218424
rect 282564 218074 282592 224198
rect 281724 218068 281776 218074
rect 281724 218010 281776 218016
rect 282552 218068 282604 218074
rect 282552 218010 282604 218016
rect 279206 217110 279280 217138
rect 280034 217246 280108 217274
rect 280862 217246 280936 217274
rect 279206 216988 279234 217110
rect 280034 216988 280062 217246
rect 280862 216988 280890 217246
rect 281736 217138 281764 218010
rect 282748 217274 282776 224946
rect 283024 220522 283052 231662
rect 284128 228682 284156 231676
rect 284116 228676 284168 228682
rect 284116 228618 284168 228624
rect 284116 228404 284168 228410
rect 284116 228346 284168 228352
rect 283380 222896 283432 222902
rect 283380 222838 283432 222844
rect 283012 220516 283064 220522
rect 283012 220458 283064 220464
rect 283392 217274 283420 222838
rect 281690 217110 281764 217138
rect 282518 217246 282776 217274
rect 283346 217246 283420 217274
rect 284128 217274 284156 228346
rect 284772 226914 284800 231676
rect 285048 231662 285430 231690
rect 285692 231662 286074 231690
rect 286244 231662 286718 231690
rect 284760 226908 284812 226914
rect 284760 226850 284812 226856
rect 285048 224126 285076 231662
rect 285312 229764 285364 229770
rect 285312 229706 285364 229712
rect 285324 225010 285352 229706
rect 285692 229094 285720 231662
rect 286244 229094 286272 231662
rect 287348 229906 287376 231676
rect 287624 231662 288006 231690
rect 287336 229900 287388 229906
rect 287336 229842 287388 229848
rect 285692 229066 285904 229094
rect 285496 225616 285548 225622
rect 285496 225558 285548 225564
rect 285312 225004 285364 225010
rect 285312 224946 285364 224952
rect 285036 224120 285088 224126
rect 285036 224062 285088 224068
rect 285508 218074 285536 225558
rect 285680 224936 285732 224942
rect 285680 224878 285732 224884
rect 285692 224262 285720 224878
rect 285680 224256 285732 224262
rect 285680 224198 285732 224204
rect 285876 222018 285904 229066
rect 286060 229066 286272 229094
rect 285864 222012 285916 222018
rect 285864 221954 285916 221960
rect 286060 221626 286088 229066
rect 286692 224120 286744 224126
rect 286692 224062 286744 224068
rect 285876 221598 286088 221626
rect 285876 221474 285904 221598
rect 285864 221468 285916 221474
rect 285864 221410 285916 221416
rect 286048 221468 286100 221474
rect 286048 221410 286100 221416
rect 285864 219428 285916 219434
rect 285864 219370 285916 219376
rect 285036 218068 285088 218074
rect 285036 218010 285088 218016
rect 285496 218068 285548 218074
rect 285496 218010 285548 218016
rect 284128 217246 284202 217274
rect 281690 216988 281718 217110
rect 282518 216988 282546 217246
rect 283346 216988 283374 217246
rect 284174 216988 284202 217246
rect 285048 217138 285076 218010
rect 285876 217138 285904 219370
rect 286060 219298 286088 221410
rect 286048 219292 286100 219298
rect 286048 219234 286100 219240
rect 286704 217274 286732 224062
rect 287624 223174 287652 231662
rect 288164 228132 288216 228138
rect 288164 228074 288216 228080
rect 287612 223168 287664 223174
rect 287612 223110 287664 223116
rect 288176 219434 288204 228074
rect 288636 224398 288664 231676
rect 289280 224806 289308 231676
rect 289924 229094 289952 231676
rect 289832 229066 289952 229094
rect 289268 224800 289320 224806
rect 289268 224742 289320 224748
rect 288624 224392 288676 224398
rect 288624 224334 288676 224340
rect 289636 224392 289688 224398
rect 289636 224334 289688 224340
rect 288348 224256 288400 224262
rect 288348 224198 288400 224204
rect 288176 219406 288296 219434
rect 287520 218068 287572 218074
rect 287520 218010 287572 218016
rect 285002 217110 285076 217138
rect 285830 217110 285904 217138
rect 286658 217246 286732 217274
rect 285002 216988 285030 217110
rect 285830 216988 285858 217110
rect 286658 216988 286686 217246
rect 287532 217138 287560 218010
rect 288268 217274 288296 219406
rect 288360 218090 288388 224198
rect 288360 218074 288480 218090
rect 289648 218074 289676 224334
rect 289832 221474 289860 229066
rect 290568 225894 290596 231676
rect 291212 228954 291240 231676
rect 291200 228948 291252 228954
rect 291200 228890 291252 228896
rect 291856 227458 291884 231676
rect 292500 230042 292528 231676
rect 292488 230036 292540 230042
rect 292488 229978 292540 229984
rect 292396 228676 292448 228682
rect 292396 228618 292448 228624
rect 291844 227452 291896 227458
rect 291844 227394 291896 227400
rect 291844 226432 291896 226438
rect 291844 226374 291896 226380
rect 290556 225888 290608 225894
rect 290556 225830 290608 225836
rect 290832 223168 290884 223174
rect 290832 223110 290884 223116
rect 289820 221468 289872 221474
rect 289820 221410 289872 221416
rect 290004 221468 290056 221474
rect 290004 221410 290056 221416
rect 288360 218068 288492 218074
rect 288360 218062 288440 218068
rect 288440 218010 288492 218016
rect 289176 218068 289228 218074
rect 289176 218010 289228 218016
rect 289636 218068 289688 218074
rect 289636 218010 289688 218016
rect 288268 217246 288342 217274
rect 287486 217110 287560 217138
rect 287486 216988 287514 217110
rect 288314 216988 288342 217246
rect 289188 217138 289216 218010
rect 290016 217274 290044 221410
rect 290844 217274 290872 223110
rect 291856 219162 291884 226374
rect 291844 219156 291896 219162
rect 291844 219098 291896 219104
rect 291660 218476 291712 218482
rect 291660 218418 291712 218424
rect 289142 217110 289216 217138
rect 289970 217246 290044 217274
rect 290798 217246 290872 217274
rect 289142 216988 289170 217110
rect 289970 216988 289998 217246
rect 290798 216988 290826 217246
rect 291672 217138 291700 218418
rect 292408 217274 292436 228618
rect 293144 227594 293172 231676
rect 293328 231662 293802 231690
rect 293132 227588 293184 227594
rect 293132 227530 293184 227536
rect 293328 220794 293356 231662
rect 293776 227452 293828 227458
rect 293776 227394 293828 227400
rect 293316 220788 293368 220794
rect 293316 220730 293368 220736
rect 293592 220788 293644 220794
rect 293592 220730 293644 220736
rect 293604 219026 293632 220730
rect 293592 219020 293644 219026
rect 293592 218962 293644 218968
rect 293788 218074 293816 227394
rect 294432 223038 294460 231676
rect 295076 226438 295104 231676
rect 295720 228818 295748 231676
rect 295904 231662 296378 231690
rect 296732 231662 297022 231690
rect 295708 228812 295760 228818
rect 295708 228754 295760 228760
rect 295064 226432 295116 226438
rect 295064 226374 295116 226380
rect 294972 225888 295024 225894
rect 294972 225830 295024 225836
rect 294420 223032 294472 223038
rect 294420 222974 294472 222980
rect 294144 219156 294196 219162
rect 294144 219098 294196 219104
rect 293316 218068 293368 218074
rect 293316 218010 293368 218016
rect 293776 218068 293828 218074
rect 293776 218010 293828 218016
rect 292408 217246 292482 217274
rect 291626 217110 291700 217138
rect 291626 216988 291654 217110
rect 292454 216988 292482 217246
rect 293328 217138 293356 218010
rect 294156 217138 294184 219098
rect 294984 217274 295012 225830
rect 295904 219978 295932 231662
rect 296444 227180 296496 227186
rect 296444 227122 296496 227128
rect 295892 219972 295944 219978
rect 295892 219914 295944 219920
rect 296456 218074 296484 227122
rect 296732 220658 296760 231662
rect 297652 230314 297680 231676
rect 297640 230308 297692 230314
rect 297640 230250 297692 230256
rect 296904 230036 296956 230042
rect 296904 229978 296956 229984
rect 296916 222766 296944 229978
rect 298296 229090 298324 231676
rect 298284 229084 298336 229090
rect 298284 229026 298336 229032
rect 298008 223576 298060 223582
rect 298008 223518 298060 223524
rect 296904 222760 296956 222766
rect 296904 222702 296956 222708
rect 296720 220652 296772 220658
rect 296720 220594 296772 220600
rect 296628 220516 296680 220522
rect 296628 220458 296680 220464
rect 295800 218068 295852 218074
rect 295800 218010 295852 218016
rect 296444 218068 296496 218074
rect 296444 218010 296496 218016
rect 293282 217110 293356 217138
rect 294110 217110 294184 217138
rect 294938 217246 295012 217274
rect 293282 216988 293310 217110
rect 294110 216988 294138 217110
rect 294938 216988 294966 217246
rect 295812 217138 295840 218010
rect 296640 217274 296668 220458
rect 296812 219972 296864 219978
rect 296812 219914 296864 219920
rect 296824 218618 296852 219914
rect 296812 218612 296864 218618
rect 296812 218554 296864 218560
rect 298020 218074 298048 223518
rect 298940 223446 298968 231676
rect 299296 227588 299348 227594
rect 299296 227530 299348 227536
rect 298928 223440 298980 223446
rect 298928 223382 298980 223388
rect 299112 218204 299164 218210
rect 299112 218146 299164 218152
rect 297456 218068 297508 218074
rect 297456 218010 297508 218016
rect 298008 218068 298060 218074
rect 298008 218010 298060 218016
rect 298284 218068 298336 218074
rect 298284 218010 298336 218016
rect 295766 217110 295840 217138
rect 296594 217246 296668 217274
rect 295766 216988 295794 217110
rect 296594 216988 296622 217246
rect 297468 217138 297496 218010
rect 298296 217138 298324 218010
rect 299124 217138 299152 218146
rect 299308 218074 299336 227530
rect 299584 225758 299612 231676
rect 299952 231662 300242 231690
rect 299572 225752 299624 225758
rect 299572 225694 299624 225700
rect 299952 220794 299980 231662
rect 300124 229900 300176 229906
rect 300124 229842 300176 229848
rect 300136 223582 300164 229842
rect 300872 224534 300900 231676
rect 301056 231662 301530 231690
rect 301700 231662 302174 231690
rect 302528 231662 302818 231690
rect 300860 224528 300912 224534
rect 300860 224470 300912 224476
rect 300124 223576 300176 223582
rect 300124 223518 300176 223524
rect 300308 223032 300360 223038
rect 300308 222974 300360 222980
rect 299940 220788 299992 220794
rect 299940 220730 299992 220736
rect 299940 220652 299992 220658
rect 299940 220594 299992 220600
rect 299296 218068 299348 218074
rect 299296 218010 299348 218016
rect 299952 217274 299980 220594
rect 300320 218210 300348 222974
rect 301056 220250 301084 231662
rect 301700 222154 301728 231662
rect 302528 230042 302556 231662
rect 302884 230308 302936 230314
rect 302884 230250 302936 230256
rect 302516 230036 302568 230042
rect 302516 229978 302568 229984
rect 302148 223440 302200 223446
rect 302148 223382 302200 223388
rect 301688 222148 301740 222154
rect 301688 222090 301740 222096
rect 301044 220244 301096 220250
rect 301044 220186 301096 220192
rect 301504 219428 301556 219434
rect 301504 219370 301556 219376
rect 301516 219026 301544 219370
rect 301504 219020 301556 219026
rect 301504 218962 301556 218968
rect 300768 218748 300820 218754
rect 300768 218690 300820 218696
rect 300308 218204 300360 218210
rect 300308 218146 300360 218152
rect 297422 217110 297496 217138
rect 298250 217110 298324 217138
rect 299078 217110 299152 217138
rect 299906 217246 299980 217274
rect 297422 216988 297450 217110
rect 298250 216988 298278 217110
rect 299078 216988 299106 217110
rect 299906 216988 299934 217246
rect 300780 217138 300808 218690
rect 302160 218074 302188 223382
rect 302896 218618 302924 230250
rect 303448 226166 303476 231676
rect 303436 226160 303488 226166
rect 303436 226102 303488 226108
rect 304092 226030 304120 231676
rect 304080 226024 304132 226030
rect 304080 225966 304132 225972
rect 303252 224528 303304 224534
rect 303252 224470 303304 224476
rect 302884 218612 302936 218618
rect 302884 218554 302936 218560
rect 301596 218068 301648 218074
rect 301596 218010 301648 218016
rect 302148 218068 302200 218074
rect 302148 218010 302200 218016
rect 302424 218068 302476 218074
rect 302424 218010 302476 218016
rect 301608 217138 301636 218010
rect 302436 217138 302464 218010
rect 303264 217274 303292 224470
rect 304736 223310 304764 231676
rect 305380 230314 305408 231676
rect 305368 230308 305420 230314
rect 305368 230250 305420 230256
rect 305644 230036 305696 230042
rect 305644 229978 305696 229984
rect 304908 225752 304960 225758
rect 304908 225694 304960 225700
rect 304724 223304 304776 223310
rect 304724 223246 304776 223252
rect 303712 221876 303764 221882
rect 303712 221818 303764 221824
rect 303724 218074 303752 221818
rect 304080 218204 304132 218210
rect 304080 218146 304132 218152
rect 303712 218068 303764 218074
rect 303712 218010 303764 218016
rect 300734 217110 300808 217138
rect 301562 217110 301636 217138
rect 302390 217110 302464 217138
rect 303218 217246 303292 217274
rect 300734 216988 300762 217110
rect 301562 216988 301590 217110
rect 302390 216988 302418 217110
rect 303218 216988 303246 217246
rect 304092 217138 304120 218146
rect 304920 217274 304948 225694
rect 305656 218210 305684 229978
rect 306024 223582 306052 231676
rect 306668 227730 306696 231676
rect 307312 228546 307340 231676
rect 307956 230450 307984 231676
rect 307944 230444 307996 230450
rect 307944 230386 307996 230392
rect 307852 230308 307904 230314
rect 307852 230250 307904 230256
rect 307300 228540 307352 228546
rect 307300 228482 307352 228488
rect 307668 228540 307720 228546
rect 307668 228482 307720 228488
rect 306656 227724 306708 227730
rect 306656 227666 306708 227672
rect 306012 223576 306064 223582
rect 306012 223518 306064 223524
rect 306288 223304 306340 223310
rect 306288 223246 306340 223252
rect 305644 218204 305696 218210
rect 305644 218146 305696 218152
rect 306300 218074 306328 223246
rect 306748 220788 306800 220794
rect 306748 220730 306800 220736
rect 306760 219026 306788 220730
rect 306748 219020 306800 219026
rect 306748 218962 306800 218968
rect 307392 218612 307444 218618
rect 307392 218554 307444 218560
rect 305736 218068 305788 218074
rect 305736 218010 305788 218016
rect 306288 218068 306340 218074
rect 306288 218010 306340 218016
rect 306564 218068 306616 218074
rect 306564 218010 306616 218016
rect 304046 217110 304120 217138
rect 304874 217246 304948 217274
rect 304046 216988 304074 217110
rect 304874 216988 304902 217246
rect 305748 217138 305776 218010
rect 306576 217138 306604 218010
rect 307404 217138 307432 218554
rect 307680 218074 307708 228482
rect 307864 224398 307892 230250
rect 308600 227050 308628 231676
rect 308588 227044 308640 227050
rect 308588 226986 308640 226992
rect 308772 227044 308824 227050
rect 308772 226986 308824 226992
rect 307852 224392 307904 224398
rect 307852 224334 307904 224340
rect 308784 218074 308812 226986
rect 308956 224392 309008 224398
rect 308956 224334 309008 224340
rect 307668 218068 307720 218074
rect 307668 218010 307720 218016
rect 308220 218068 308272 218074
rect 308220 218010 308272 218016
rect 308772 218068 308824 218074
rect 308772 218010 308824 218016
rect 308232 217138 308260 218010
rect 308968 217274 308996 224334
rect 309244 221338 309272 231676
rect 309888 224670 309916 231676
rect 310546 231662 310744 231690
rect 309876 224664 309928 224670
rect 309876 224606 309928 224612
rect 309876 222012 309928 222018
rect 309876 221954 309928 221960
rect 309232 221332 309284 221338
rect 309232 221274 309284 221280
rect 309888 217274 309916 221954
rect 310716 219978 310744 231662
rect 310900 231662 311190 231690
rect 310900 221746 310928 231662
rect 311820 228274 311848 231676
rect 312096 231662 312478 231690
rect 311808 228268 311860 228274
rect 311808 228210 311860 228216
rect 312096 227322 312124 231662
rect 312544 230444 312596 230450
rect 312544 230386 312596 230392
rect 312084 227316 312136 227322
rect 312084 227258 312136 227264
rect 310888 221740 310940 221746
rect 310888 221682 310940 221688
rect 311532 221740 311584 221746
rect 311532 221682 311584 221688
rect 310704 219972 310756 219978
rect 310704 219914 310756 219920
rect 310704 218204 310756 218210
rect 310704 218146 310756 218152
rect 308968 217246 309042 217274
rect 305702 217110 305776 217138
rect 306530 217110 306604 217138
rect 307358 217110 307432 217138
rect 308186 217110 308260 217138
rect 305702 216988 305730 217110
rect 306530 216988 306558 217110
rect 307358 216988 307386 217110
rect 308186 216988 308214 217110
rect 309014 216988 309042 217246
rect 309842 217246 309916 217274
rect 309842 216988 309870 217246
rect 310716 217138 310744 218146
rect 311544 217274 311572 221682
rect 311808 220244 311860 220250
rect 311808 220186 311860 220192
rect 311820 219162 311848 220186
rect 311808 219156 311860 219162
rect 311808 219098 311860 219104
rect 312556 218890 312584 230386
rect 313108 230178 313136 231676
rect 313292 231662 313766 231690
rect 313936 231662 314410 231690
rect 313096 230172 313148 230178
rect 313096 230114 313148 230120
rect 313096 226024 313148 226030
rect 313096 225966 313148 225972
rect 312544 218884 312596 218890
rect 312544 218826 312596 218832
rect 312360 218068 312412 218074
rect 312360 218010 312412 218016
rect 310670 217110 310744 217138
rect 311498 217246 311572 217274
rect 310670 216988 310698 217110
rect 311498 216988 311526 217246
rect 312372 217138 312400 218010
rect 313108 217274 313136 225966
rect 313292 221610 313320 231662
rect 313280 221604 313332 221610
rect 313280 221546 313332 221552
rect 313936 220386 313964 231662
rect 315040 226302 315068 231676
rect 315684 230450 315712 231676
rect 315672 230444 315724 230450
rect 315672 230386 315724 230392
rect 315304 230172 315356 230178
rect 315304 230114 315356 230120
rect 315028 226296 315080 226302
rect 315028 226238 315080 226244
rect 314476 221604 314528 221610
rect 314476 221546 314528 221552
rect 313924 220380 313976 220386
rect 313924 220322 313976 220328
rect 314016 218884 314068 218890
rect 314016 218826 314068 218832
rect 313108 217246 313182 217274
rect 312326 217110 312400 217138
rect 312326 216988 312354 217110
rect 313154 216988 313182 217246
rect 314028 217138 314056 218826
rect 314488 218074 314516 221546
rect 315316 218210 315344 230114
rect 316328 224942 316356 231676
rect 316316 224936 316368 224942
rect 316316 224878 316368 224884
rect 315856 224800 315908 224806
rect 315856 224742 315908 224748
rect 315672 219156 315724 219162
rect 315672 219098 315724 219104
rect 315304 218204 315356 218210
rect 315304 218146 315356 218152
rect 314476 218068 314528 218074
rect 314476 218010 314528 218016
rect 314844 218068 314896 218074
rect 314844 218010 314896 218016
rect 314856 217138 314884 218010
rect 315684 217138 315712 219098
rect 315868 218074 315896 224742
rect 316972 222902 317000 231676
rect 317524 231662 317630 231690
rect 317328 226296 317380 226302
rect 317328 226238 317380 226244
rect 316960 222896 317012 222902
rect 316960 222838 317012 222844
rect 317144 222896 317196 222902
rect 317144 222838 317196 222844
rect 317156 218074 317184 222838
rect 315856 218068 315908 218074
rect 315856 218010 315908 218016
rect 316500 218068 316552 218074
rect 316500 218010 316552 218016
rect 317144 218068 317196 218074
rect 317144 218010 317196 218016
rect 316512 217138 316540 218010
rect 317340 217274 317368 226238
rect 317524 220114 317552 231662
rect 318260 229770 318288 231676
rect 318248 229764 318300 229770
rect 318248 229706 318300 229712
rect 317972 228812 318024 228818
rect 317972 228754 318024 228760
rect 317512 220108 317564 220114
rect 317512 220050 317564 220056
rect 317984 219162 318012 228754
rect 318904 225622 318932 231676
rect 318892 225616 318944 225622
rect 318892 225558 318944 225564
rect 319548 224126 319576 231676
rect 319812 228948 319864 228954
rect 319812 228890 319864 228896
rect 319536 224120 319588 224126
rect 319536 224062 319588 224068
rect 318156 220108 318208 220114
rect 318156 220050 318208 220056
rect 317972 219156 318024 219162
rect 317972 219098 318024 219104
rect 318168 217274 318196 220050
rect 318984 218068 319036 218074
rect 318984 218010 319036 218016
rect 313982 217110 314056 217138
rect 314810 217110 314884 217138
rect 315638 217110 315712 217138
rect 316466 217110 316540 217138
rect 317294 217246 317368 217274
rect 318122 217246 318196 217274
rect 313982 216988 314010 217110
rect 314810 216988 314838 217110
rect 315638 216988 315666 217110
rect 316466 216988 316494 217110
rect 317294 216988 317322 217246
rect 318122 216988 318150 217246
rect 318996 217138 319024 218010
rect 319824 217274 319852 228890
rect 320192 228410 320220 231676
rect 320376 231662 320850 231690
rect 320180 228404 320232 228410
rect 320180 228346 320232 228352
rect 319996 224664 320048 224670
rect 319996 224606 320048 224612
rect 320008 218074 320036 224606
rect 320376 220794 320404 231662
rect 321480 228138 321508 231676
rect 321756 231662 322138 231690
rect 322400 231662 322782 231690
rect 321468 228132 321520 228138
rect 321468 228074 321520 228080
rect 321376 227724 321428 227730
rect 321376 227666 321428 227672
rect 320364 220788 320416 220794
rect 320364 220730 320416 220736
rect 320640 219156 320692 219162
rect 320640 219098 320692 219104
rect 319996 218068 320048 218074
rect 319996 218010 320048 218016
rect 318950 217110 319024 217138
rect 319778 217246 319852 217274
rect 318950 216988 318978 217110
rect 319778 216988 319806 217246
rect 320652 217138 320680 219098
rect 321388 217274 321416 227666
rect 321756 221474 321784 231662
rect 322400 224262 322428 231662
rect 323412 230314 323440 231676
rect 323688 231662 324070 231690
rect 323400 230308 323452 230314
rect 323400 230250 323452 230256
rect 322848 225616 322900 225622
rect 322848 225558 322900 225564
rect 322388 224256 322440 224262
rect 322388 224198 322440 224204
rect 321744 221468 321796 221474
rect 321744 221410 321796 221416
rect 322860 218074 322888 225558
rect 323688 223174 323716 231662
rect 324044 229764 324096 229770
rect 324044 229706 324096 229712
rect 323676 223168 323728 223174
rect 323676 223110 323728 223116
rect 323124 220380 323176 220386
rect 323124 220322 323176 220328
rect 322296 218068 322348 218074
rect 322296 218010 322348 218016
rect 322848 218068 322900 218074
rect 322848 218010 322900 218016
rect 321388 217246 321462 217274
rect 320606 217110 320680 217138
rect 320606 216988 320634 217110
rect 321434 216988 321462 217246
rect 322308 217138 322336 218010
rect 323136 217274 323164 220322
rect 324056 219434 324084 229706
rect 324700 219434 324728 231676
rect 325344 227458 325372 231676
rect 325332 227452 325384 227458
rect 325332 227394 325384 227400
rect 325424 226160 325476 226166
rect 325424 226102 325476 226108
rect 323964 219406 324084 219434
rect 324608 219406 324728 219434
rect 323964 217274 323992 219406
rect 324608 218482 324636 219406
rect 324596 218476 324648 218482
rect 324596 218418 324648 218424
rect 325436 218074 325464 226102
rect 325988 225894 326016 231676
rect 326632 228682 326660 231676
rect 326620 228676 326672 228682
rect 326620 228618 326672 228624
rect 326896 228404 326948 228410
rect 326896 228346 326948 228352
rect 326344 227316 326396 227322
rect 326344 227258 326396 227264
rect 325976 225888 326028 225894
rect 325976 225830 326028 225836
rect 326356 219434 326384 227258
rect 325608 219428 325660 219434
rect 325608 219370 325660 219376
rect 326344 219428 326396 219434
rect 326344 219370 326396 219376
rect 324780 218068 324832 218074
rect 324780 218010 324832 218016
rect 325424 218068 325476 218074
rect 325424 218010 325476 218016
rect 322262 217110 322336 217138
rect 323090 217246 323164 217274
rect 323918 217246 323992 217274
rect 322262 216988 322290 217110
rect 323090 216988 323118 217246
rect 323918 216988 323946 217246
rect 324792 217138 324820 218010
rect 325620 217138 325648 219370
rect 326908 218074 326936 228346
rect 327276 220250 327304 231676
rect 327552 231662 327934 231690
rect 327552 220522 327580 231662
rect 328564 227594 328592 231676
rect 328552 227588 328604 227594
rect 328552 227530 328604 227536
rect 329208 227186 329236 231676
rect 329852 229906 329880 231676
rect 330036 231662 330510 231690
rect 329840 229900 329892 229906
rect 329840 229842 329892 229848
rect 329196 227180 329248 227186
rect 329196 227122 329248 227128
rect 329748 227180 329800 227186
rect 329748 227122 329800 227128
rect 329104 223576 329156 223582
rect 329104 223518 329156 223524
rect 327540 220516 327592 220522
rect 327540 220458 327592 220464
rect 328092 220516 328144 220522
rect 328092 220458 328144 220464
rect 327264 220244 327316 220250
rect 327264 220186 327316 220192
rect 327264 219292 327316 219298
rect 327264 219234 327316 219240
rect 326436 218068 326488 218074
rect 326436 218010 326488 218016
rect 326896 218068 326948 218074
rect 326896 218010 326948 218016
rect 326448 217138 326476 218010
rect 327276 217274 327304 219234
rect 328104 217274 328132 220458
rect 329116 218890 329144 223518
rect 329564 220788 329616 220794
rect 329564 220730 329616 220736
rect 329576 219026 329604 220730
rect 329564 219020 329616 219026
rect 329564 218962 329616 218968
rect 329104 218884 329156 218890
rect 329104 218826 329156 218832
rect 328920 218068 328972 218074
rect 328920 218010 328972 218016
rect 324746 217110 324820 217138
rect 325574 217110 325648 217138
rect 326402 217110 326476 217138
rect 327230 217246 327304 217274
rect 328058 217246 328132 217274
rect 324746 216988 324774 217110
rect 325574 216988 325602 217110
rect 326402 216988 326430 217110
rect 327230 216988 327258 217246
rect 328058 216988 328086 217246
rect 328932 217138 328960 218010
rect 329760 217274 329788 227122
rect 330036 220658 330064 231662
rect 331140 223446 331168 231676
rect 331324 231662 331798 231690
rect 331968 231662 332442 231690
rect 331128 223440 331180 223446
rect 331128 223382 331180 223388
rect 330484 223168 330536 223174
rect 330484 223110 330536 223116
rect 330024 220652 330076 220658
rect 330024 220594 330076 220600
rect 330496 218074 330524 223110
rect 331324 223038 331352 231662
rect 331312 223032 331364 223038
rect 331312 222974 331364 222980
rect 331404 222148 331456 222154
rect 331404 222090 331456 222096
rect 330668 218204 330720 218210
rect 330668 218146 330720 218152
rect 330484 218068 330536 218074
rect 330484 218010 330536 218016
rect 330680 217274 330708 218146
rect 331416 217274 331444 222090
rect 331968 220794 331996 231662
rect 333072 224534 333100 231676
rect 333244 228676 333296 228682
rect 333244 228618 333296 228624
rect 333060 224528 333112 224534
rect 333060 224470 333112 224476
rect 331956 220788 332008 220794
rect 331956 220730 332008 220736
rect 332232 220244 332284 220250
rect 332232 220186 332284 220192
rect 332244 217274 332272 220186
rect 333256 218210 333284 228618
rect 333716 225758 333744 231676
rect 334084 231662 334374 231690
rect 333704 225752 333756 225758
rect 333704 225694 333756 225700
rect 333888 224528 333940 224534
rect 333888 224470 333940 224476
rect 333704 219020 333756 219026
rect 333704 218962 333756 218968
rect 333244 218204 333296 218210
rect 333244 218146 333296 218152
rect 333060 218068 333112 218074
rect 333060 218010 333112 218016
rect 328886 217110 328960 217138
rect 329714 217246 329788 217274
rect 330542 217246 330708 217274
rect 331370 217246 331444 217274
rect 332198 217246 332272 217274
rect 328886 216988 328914 217110
rect 329714 216988 329742 217246
rect 330542 216988 330570 217246
rect 331370 216988 331398 217246
rect 332198 216988 332226 217246
rect 333072 217138 333100 218010
rect 333716 217274 333744 218962
rect 333900 218074 333928 224470
rect 334084 221882 334112 231662
rect 335004 230042 335032 231676
rect 334992 230036 335044 230042
rect 334992 229978 335044 229984
rect 334256 229900 334308 229906
rect 334256 229842 334308 229848
rect 334268 226302 334296 229842
rect 335648 228546 335676 231676
rect 335636 228540 335688 228546
rect 335636 228482 335688 228488
rect 336292 227050 336320 231676
rect 336648 228540 336700 228546
rect 336648 228482 336700 228488
rect 336280 227044 336332 227050
rect 336280 226986 336332 226992
rect 336464 227044 336516 227050
rect 336464 226986 336516 226992
rect 334256 226296 334308 226302
rect 334256 226238 334308 226244
rect 335268 225752 335320 225758
rect 335268 225694 335320 225700
rect 334072 221876 334124 221882
rect 334072 221818 334124 221824
rect 335280 218074 335308 225694
rect 336476 219434 336504 226986
rect 336660 219434 336688 228482
rect 336936 223310 336964 231676
rect 337120 231662 337594 231690
rect 338238 231662 338436 231690
rect 336924 223304 336976 223310
rect 336924 223246 336976 223252
rect 337120 219434 337148 231662
rect 337936 223032 337988 223038
rect 337936 222974 337988 222980
rect 336384 219406 336504 219434
rect 336568 219406 336688 219434
rect 337028 219406 337148 219434
rect 336384 218074 336412 219406
rect 333888 218068 333940 218074
rect 333888 218010 333940 218016
rect 334716 218068 334768 218074
rect 334716 218010 334768 218016
rect 335268 218068 335320 218074
rect 335268 218010 335320 218016
rect 335544 218068 335596 218074
rect 335544 218010 335596 218016
rect 336372 218068 336424 218074
rect 336372 218010 336424 218016
rect 333716 217246 333882 217274
rect 333026 217110 333100 217138
rect 333026 216988 333054 217110
rect 333854 216988 333882 217246
rect 334728 217138 334756 218010
rect 335556 217138 335584 218010
rect 336568 217274 336596 219406
rect 337028 218754 337056 219406
rect 337200 218884 337252 218890
rect 337200 218826 337252 218832
rect 337016 218748 337068 218754
rect 337016 218690 337068 218696
rect 334682 217110 334756 217138
rect 335510 217110 335584 217138
rect 336338 217246 336596 217274
rect 334682 216988 334710 217110
rect 335510 216988 335538 217110
rect 336338 216988 336366 217246
rect 337212 217138 337240 218826
rect 337948 217274 337976 222974
rect 338408 222018 338436 231662
rect 338592 231662 338882 231690
rect 338396 222012 338448 222018
rect 338396 221954 338448 221960
rect 338592 221746 338620 231662
rect 339512 224398 339540 231676
rect 340156 230178 340184 231676
rect 340144 230172 340196 230178
rect 340144 230114 340196 230120
rect 340604 227452 340656 227458
rect 340604 227394 340656 227400
rect 340144 225888 340196 225894
rect 340144 225830 340196 225836
rect 339500 224392 339552 224398
rect 339500 224334 339552 224340
rect 338580 221740 338632 221746
rect 338580 221682 338632 221688
rect 338856 221468 338908 221474
rect 338856 221410 338908 221416
rect 338868 217274 338896 221410
rect 340156 219162 340184 225830
rect 340616 219434 340644 227394
rect 340800 226030 340828 231676
rect 340788 226024 340840 226030
rect 340788 225966 340840 225972
rect 341444 224806 341472 231676
rect 341628 231662 342102 231690
rect 341432 224800 341484 224806
rect 341432 224742 341484 224748
rect 341628 221746 341656 231662
rect 342076 224256 342128 224262
rect 342076 224198 342128 224204
rect 341616 221740 341668 221746
rect 341616 221682 341668 221688
rect 341340 221604 341392 221610
rect 341340 221546 341392 221552
rect 340616 219406 340736 219434
rect 340144 219156 340196 219162
rect 340144 219098 340196 219104
rect 340512 218748 340564 218754
rect 340512 218690 340564 218696
rect 339684 218068 339736 218074
rect 339684 218010 339736 218016
rect 337948 217246 338022 217274
rect 337166 217110 337240 217138
rect 337166 216988 337194 217110
rect 337994 216988 338022 217246
rect 338822 217246 338896 217274
rect 338822 216988 338850 217246
rect 339696 217138 339724 218010
rect 340524 217274 340552 218690
rect 340708 218074 340736 219406
rect 340696 218068 340748 218074
rect 340696 218010 340748 218016
rect 341352 217274 341380 221546
rect 339650 217110 339724 217138
rect 340478 217246 340552 217274
rect 341306 217246 341380 217274
rect 342088 217274 342116 224198
rect 342732 223582 342760 231676
rect 342720 223576 342772 223582
rect 342720 223518 342772 223524
rect 343376 222902 343404 231676
rect 343744 231662 344034 231690
rect 343548 223304 343600 223310
rect 343548 223246 343600 223252
rect 343364 222896 343416 222902
rect 343364 222838 343416 222844
rect 343560 218074 343588 223246
rect 343744 220114 343772 231662
rect 344664 228818 344692 231676
rect 345308 229906 345336 231676
rect 345664 230104 345716 230110
rect 345664 230046 345716 230052
rect 345296 229900 345348 229906
rect 345296 229842 345348 229848
rect 344652 228812 344704 228818
rect 344652 228754 344704 228760
rect 344652 224392 344704 224398
rect 344652 224334 344704 224340
rect 343732 220108 343784 220114
rect 343732 220050 343784 220056
rect 343824 219428 343876 219434
rect 343824 219370 343876 219376
rect 342996 218068 343048 218074
rect 342996 218010 343048 218016
rect 343548 218068 343600 218074
rect 343548 218010 343600 218016
rect 342088 217246 342162 217274
rect 339650 216988 339678 217110
rect 340478 216988 340506 217246
rect 341306 216988 341334 217246
rect 342134 216988 342162 217246
rect 343008 217138 343036 218010
rect 343836 217138 343864 219370
rect 344664 217274 344692 224334
rect 345480 220108 345532 220114
rect 345480 220050 345532 220056
rect 345492 217274 345520 220050
rect 345676 219162 345704 230046
rect 345952 228954 345980 231676
rect 345940 228948 345992 228954
rect 345940 228890 345992 228896
rect 346216 228812 346268 228818
rect 346216 228754 346268 228760
rect 345664 219156 345716 219162
rect 345664 219098 345716 219104
rect 342962 217110 343036 217138
rect 343790 217110 343864 217138
rect 344618 217246 344692 217274
rect 345446 217246 345520 217274
rect 346228 217274 346256 228754
rect 346596 227730 346624 231676
rect 346584 227724 346636 227730
rect 346584 227666 346636 227672
rect 347044 225888 347096 225894
rect 347044 225830 347096 225836
rect 347056 219434 347084 225830
rect 347240 224670 347268 231676
rect 347884 226030 347912 231676
rect 348160 231662 348542 231690
rect 347872 226024 347924 226030
rect 347872 225966 347924 225972
rect 347228 224664 347280 224670
rect 347228 224606 347280 224612
rect 347596 222896 347648 222902
rect 347596 222838 347648 222844
rect 347044 219428 347096 219434
rect 347044 219370 347096 219376
rect 347608 218074 347636 222838
rect 348160 220386 348188 231662
rect 349172 226166 349200 231676
rect 349160 226160 349212 226166
rect 349160 226102 349212 226108
rect 349068 226024 349120 226030
rect 349068 225966 349120 225972
rect 348148 220380 348200 220386
rect 348148 220322 348200 220328
rect 348792 218204 348844 218210
rect 348792 218146 348844 218152
rect 347136 218068 347188 218074
rect 347136 218010 347188 218016
rect 347596 218068 347648 218074
rect 347596 218010 347648 218016
rect 347964 218068 348016 218074
rect 347964 218010 348016 218016
rect 346228 217246 346302 217274
rect 342962 216988 342990 217110
rect 343790 216988 343818 217110
rect 344618 216988 344646 217246
rect 345446 216988 345474 217246
rect 346274 216988 346302 217246
rect 347148 217138 347176 218010
rect 347976 217138 348004 218010
rect 348804 217138 348832 218146
rect 349080 218074 349108 225966
rect 349816 225622 349844 231676
rect 350460 229770 350488 231676
rect 350448 229764 350500 229770
rect 350448 229706 350500 229712
rect 350540 229628 350592 229634
rect 350540 229570 350592 229576
rect 350172 228948 350224 228954
rect 350172 228890 350224 228896
rect 349804 225616 349856 225622
rect 349804 225558 349856 225564
rect 350184 218074 350212 228890
rect 350552 225026 350580 229570
rect 351104 228410 351132 231676
rect 351288 231662 351762 231690
rect 351288 229094 351316 231662
rect 351288 229066 351408 229094
rect 351092 228404 351144 228410
rect 351092 228346 351144 228352
rect 351184 225616 351236 225622
rect 351184 225558 351236 225564
rect 350368 224998 350580 225026
rect 349068 218068 349120 218074
rect 349068 218010 349120 218016
rect 349620 218068 349672 218074
rect 349620 218010 349672 218016
rect 350172 218068 350224 218074
rect 350172 218010 350224 218016
rect 349632 217138 349660 218010
rect 350368 217274 350396 224998
rect 351196 218210 351224 225558
rect 351380 220522 351408 229066
rect 352392 227322 352420 231676
rect 353036 230110 353064 231676
rect 353024 230104 353076 230110
rect 353024 230046 353076 230052
rect 352564 229900 352616 229906
rect 352564 229842 352616 229848
rect 352380 227316 352432 227322
rect 352380 227258 352432 227264
rect 351368 220516 351420 220522
rect 351368 220458 351420 220464
rect 352104 219428 352156 219434
rect 352104 219370 352156 219376
rect 351368 219020 351420 219026
rect 351368 218962 351420 218968
rect 351184 218204 351236 218210
rect 351184 218146 351236 218152
rect 351380 217274 351408 218962
rect 350368 217246 350442 217274
rect 347102 217110 347176 217138
rect 347930 217110 348004 217138
rect 348758 217110 348832 217138
rect 349586 217110 349660 217138
rect 347102 216988 347130 217110
rect 347930 216988 347958 217110
rect 348758 216988 348786 217110
rect 349586 216988 349614 217110
rect 350414 216988 350442 217246
rect 351242 217246 351408 217274
rect 351242 216988 351270 217246
rect 352116 217138 352144 219370
rect 352576 219162 352604 229842
rect 353680 227186 353708 231676
rect 353956 231662 354338 231690
rect 353668 227180 353720 227186
rect 353668 227122 353720 227128
rect 353956 222154 353984 231662
rect 354588 227180 354640 227186
rect 354588 227122 354640 227128
rect 353944 222148 353996 222154
rect 353944 222090 353996 222096
rect 352932 220380 352984 220386
rect 352932 220322 352984 220328
rect 352564 219156 352616 219162
rect 352564 219098 352616 219104
rect 352944 217274 352972 220322
rect 354404 219156 354456 219162
rect 354404 219098 354456 219104
rect 353760 218068 353812 218074
rect 353760 218010 353812 218016
rect 352070 217110 352144 217138
rect 352898 217246 352972 217274
rect 352070 216988 352098 217110
rect 352898 216988 352926 217246
rect 353772 217138 353800 218010
rect 354416 217274 354444 219098
rect 354600 218074 354628 227122
rect 354968 223174 354996 231676
rect 355612 228682 355640 231676
rect 355600 228676 355652 228682
rect 355600 228618 355652 228624
rect 355232 228404 355284 228410
rect 355232 228346 355284 228352
rect 354956 223168 355008 223174
rect 354956 223110 355008 223116
rect 355244 219026 355272 228346
rect 355508 227316 355560 227322
rect 355508 227258 355560 227264
rect 355520 219162 355548 227258
rect 356256 224534 356284 231676
rect 356900 225758 356928 231676
rect 356888 225752 356940 225758
rect 356888 225694 356940 225700
rect 356244 224528 356296 224534
rect 356244 224470 356296 224476
rect 357348 224528 357400 224534
rect 357348 224470 357400 224476
rect 357072 223168 357124 223174
rect 357072 223110 357124 223116
rect 355508 219156 355560 219162
rect 355508 219098 355560 219104
rect 355232 219020 355284 219026
rect 355232 218962 355284 218968
rect 355416 219020 355468 219026
rect 355416 218962 355468 218968
rect 354588 218068 354640 218074
rect 354588 218010 354640 218016
rect 354416 217246 354582 217274
rect 353726 217110 353800 217138
rect 353726 216988 353754 217110
rect 354554 216988 354582 217246
rect 355428 217138 355456 218962
rect 356244 218068 356296 218074
rect 356244 218010 356296 218016
rect 356256 217138 356284 218010
rect 357084 217274 357112 223110
rect 357360 218074 357388 224470
rect 357544 220250 357572 231676
rect 358188 229906 358216 231676
rect 358176 229900 358228 229906
rect 358176 229842 358228 229848
rect 358084 229288 358136 229294
rect 358084 229230 358136 229236
rect 357532 220244 357584 220250
rect 357532 220186 357584 220192
rect 358096 219434 358124 229230
rect 358832 228546 358860 231676
rect 359200 231662 359490 231690
rect 358820 228540 358872 228546
rect 358820 228482 358872 228488
rect 359200 223038 359228 231662
rect 359372 227588 359424 227594
rect 359372 227530 359424 227536
rect 359188 223032 359240 223038
rect 359188 222974 359240 222980
rect 357728 219406 358124 219434
rect 357728 218890 357756 219406
rect 358728 219156 358780 219162
rect 358728 219098 358780 219104
rect 357716 218884 357768 218890
rect 357716 218826 357768 218832
rect 357348 218068 357400 218074
rect 357348 218010 357400 218016
rect 357900 218068 357952 218074
rect 357900 218010 357952 218016
rect 355382 217110 355456 217138
rect 356210 217110 356284 217138
rect 357038 217246 357112 217274
rect 355382 216988 355410 217110
rect 356210 216988 356238 217110
rect 357038 216988 357066 217246
rect 357912 217138 357940 218010
rect 358740 217138 358768 219098
rect 359384 218074 359412 227530
rect 360120 227050 360148 231676
rect 360764 229294 360792 231676
rect 360752 229288 360804 229294
rect 360752 229230 360804 229236
rect 360936 229288 360988 229294
rect 360936 229230 360988 229236
rect 360108 227044 360160 227050
rect 360108 226986 360160 226992
rect 359556 221740 359608 221746
rect 359556 221682 359608 221688
rect 359372 218068 359424 218074
rect 359372 218010 359424 218016
rect 359568 217274 359596 221682
rect 360384 220244 360436 220250
rect 360384 220186 360436 220192
rect 360396 217274 360424 220186
rect 360948 219434 360976 229230
rect 361408 227458 361436 231676
rect 361592 231662 362066 231690
rect 362236 231662 362710 231690
rect 361396 227452 361448 227458
rect 361396 227394 361448 227400
rect 361212 227044 361264 227050
rect 361212 226986 361264 226992
rect 360856 219406 360976 219434
rect 360856 218754 360884 219406
rect 360844 218748 360896 218754
rect 360844 218690 360896 218696
rect 361224 217274 361252 226986
rect 361592 221610 361620 231662
rect 362236 221610 362264 231662
rect 363340 229294 363368 231676
rect 363328 229288 363380 229294
rect 363328 229230 363380 229236
rect 362868 228404 362920 228410
rect 362868 228346 362920 228352
rect 361580 221604 361632 221610
rect 361580 221546 361632 221552
rect 362224 221604 362276 221610
rect 362224 221546 362276 221552
rect 362040 221468 362092 221474
rect 362040 221410 362092 221416
rect 362052 217274 362080 221410
rect 362880 217274 362908 228346
rect 363984 223310 364012 231676
rect 364156 229900 364208 229906
rect 364156 229842 364208 229848
rect 363972 223304 364024 223310
rect 363972 223246 364024 223252
rect 364168 218074 364196 229842
rect 364628 224398 364656 231676
rect 364812 231662 365286 231690
rect 364616 224392 364668 224398
rect 364616 224334 364668 224340
rect 364812 224262 364840 231662
rect 365916 225894 365944 231676
rect 366560 228818 366588 231676
rect 366548 228812 366600 228818
rect 366548 228754 366600 228760
rect 366916 228540 366968 228546
rect 366916 228482 366968 228488
rect 366364 227792 366416 227798
rect 366364 227734 366416 227740
rect 365904 225888 365956 225894
rect 365904 225830 365956 225836
rect 364800 224256 364852 224262
rect 364800 224198 364852 224204
rect 364984 224256 365036 224262
rect 364984 224198 365036 224204
rect 364996 219162 365024 224198
rect 366376 219434 366404 227734
rect 366364 219428 366416 219434
rect 366364 219370 366416 219376
rect 364984 219156 365036 219162
rect 364984 219098 365036 219104
rect 366732 218884 366784 218890
rect 366732 218826 366784 218832
rect 365352 218340 365404 218346
rect 365352 218282 365404 218288
rect 364524 218204 364576 218210
rect 364524 218146 364576 218152
rect 363696 218068 363748 218074
rect 363696 218010 363748 218016
rect 364156 218068 364208 218074
rect 364156 218010 364208 218016
rect 357866 217110 357940 217138
rect 358694 217110 358768 217138
rect 359522 217246 359596 217274
rect 360350 217246 360424 217274
rect 361178 217246 361252 217274
rect 362006 217246 362080 217274
rect 362834 217246 362908 217274
rect 357866 216988 357894 217110
rect 358694 216988 358722 217110
rect 359522 216988 359550 217246
rect 360350 216988 360378 217246
rect 361178 216988 361206 217246
rect 362006 216988 362034 217246
rect 362834 216988 362862 217246
rect 363708 217138 363736 218010
rect 364536 217138 364564 218146
rect 365364 217138 365392 218282
rect 366180 218068 366232 218074
rect 366180 218010 366232 218016
rect 366192 217138 366220 218010
rect 366744 217274 366772 218826
rect 366928 218074 366956 228482
rect 367204 226030 367232 231676
rect 367388 231662 367862 231690
rect 367192 226024 367244 226030
rect 367192 225966 367244 225972
rect 367388 220114 367416 231662
rect 367652 225888 367704 225894
rect 367652 225830 367704 225836
rect 367376 220108 367428 220114
rect 367376 220050 367428 220056
rect 367664 218210 367692 225830
rect 368492 222902 368520 231676
rect 369136 228954 369164 231676
rect 369124 228948 369176 228954
rect 369124 228890 369176 228896
rect 369780 228682 369808 231676
rect 369768 228676 369820 228682
rect 369768 228618 369820 228624
rect 369124 227928 369176 227934
rect 369124 227870 369176 227876
rect 368480 222896 368532 222902
rect 368480 222838 368532 222844
rect 367836 220108 367888 220114
rect 367836 220050 367888 220056
rect 367652 218204 367704 218210
rect 367652 218146 367704 218152
rect 366916 218068 366968 218074
rect 366916 218010 366968 218016
rect 367848 217274 367876 220050
rect 369136 219026 369164 227870
rect 369768 227452 369820 227458
rect 369768 227394 369820 227400
rect 369124 219020 369176 219026
rect 369124 218962 369176 218968
rect 369492 218204 369544 218210
rect 369492 218146 369544 218152
rect 368664 218068 368716 218074
rect 368664 218010 368716 218016
rect 366744 217246 367002 217274
rect 363662 217110 363736 217138
rect 364490 217110 364564 217138
rect 365318 217110 365392 217138
rect 366146 217110 366220 217138
rect 363662 216988 363690 217110
rect 364490 216988 364518 217110
rect 365318 216988 365346 217110
rect 366146 216988 366174 217110
rect 366974 216988 367002 217246
rect 367802 217246 367876 217274
rect 367802 216988 367830 217246
rect 368676 217138 368704 218010
rect 369504 217138 369532 218146
rect 369780 218074 369808 227394
rect 370424 225622 370452 231676
rect 371068 229770 371096 231676
rect 371436 231662 371726 231690
rect 371056 229764 371108 229770
rect 371056 229706 371108 229712
rect 370964 229628 371016 229634
rect 370964 229570 371016 229576
rect 370412 225616 370464 225622
rect 370412 225558 370464 225564
rect 370504 223032 370556 223038
rect 370504 222974 370556 222980
rect 370516 218210 370544 222974
rect 370504 218204 370556 218210
rect 370504 218146 370556 218152
rect 370976 218074 371004 229570
rect 371148 220516 371200 220522
rect 371148 220458 371200 220464
rect 369768 218068 369820 218074
rect 369768 218010 369820 218016
rect 370320 218068 370372 218074
rect 370320 218010 370372 218016
rect 370964 218068 371016 218074
rect 370964 218010 371016 218016
rect 370332 217138 370360 218010
rect 371160 217274 371188 220458
rect 371436 220386 371464 231662
rect 372356 227322 372384 231676
rect 373000 227798 373028 231676
rect 372988 227792 373040 227798
rect 372988 227734 373040 227740
rect 373644 227322 373672 231676
rect 373816 228676 373868 228682
rect 373816 228618 373868 228624
rect 372344 227316 372396 227322
rect 372344 227258 372396 227264
rect 373632 227316 373684 227322
rect 373632 227258 373684 227264
rect 373264 227180 373316 227186
rect 373264 227122 373316 227128
rect 372528 225616 372580 225622
rect 372528 225558 372580 225564
rect 371424 220380 371476 220386
rect 371424 220322 371476 220328
rect 372540 218074 372568 225558
rect 373276 218346 373304 227122
rect 373632 219020 373684 219026
rect 373632 218962 373684 218968
rect 373264 218340 373316 218346
rect 373264 218282 373316 218288
rect 371976 218068 372028 218074
rect 371976 218010 372028 218016
rect 372528 218068 372580 218074
rect 372528 218010 372580 218016
rect 372804 218068 372856 218074
rect 372804 218010 372856 218016
rect 368630 217110 368704 217138
rect 369458 217110 369532 217138
rect 370286 217110 370360 217138
rect 371114 217246 371188 217274
rect 368630 216988 368658 217110
rect 369458 216988 369486 217110
rect 370286 216988 370314 217110
rect 371114 216988 371142 217246
rect 371988 217138 372016 218010
rect 372816 217138 372844 218010
rect 373644 217138 373672 218962
rect 373828 218074 373856 228618
rect 374288 224534 374316 231676
rect 374932 227594 374960 231676
rect 375576 227934 375604 231676
rect 375564 227928 375616 227934
rect 375564 227870 375616 227876
rect 374920 227588 374972 227594
rect 374920 227530 374972 227536
rect 374276 224528 374328 224534
rect 374276 224470 374328 224476
rect 375288 224392 375340 224398
rect 375288 224334 375340 224340
rect 375104 222896 375156 222902
rect 375104 222838 375156 222844
rect 375116 219434 375144 222838
rect 375300 219434 375328 224334
rect 376220 223174 376248 231676
rect 376576 228812 376628 228818
rect 376576 228754 376628 228760
rect 376208 223168 376260 223174
rect 376208 223110 376260 223116
rect 374460 219428 374512 219434
rect 375116 219406 375236 219434
rect 375300 219428 375432 219434
rect 375300 219406 375380 219428
rect 374460 219370 374512 219376
rect 373816 218068 373868 218074
rect 373816 218010 373868 218016
rect 374472 217138 374500 219370
rect 375208 217274 375236 219406
rect 375380 219370 375432 219376
rect 376588 218074 376616 228754
rect 376864 221746 376892 231676
rect 377232 231662 377522 231690
rect 377232 227050 377260 231662
rect 377404 230444 377456 230450
rect 377404 230386 377456 230392
rect 377220 227044 377272 227050
rect 377220 226986 377272 226992
rect 376852 221740 376904 221746
rect 376852 221682 376904 221688
rect 377416 220250 377444 230386
rect 378152 224262 378180 231676
rect 378796 230450 378824 231676
rect 378784 230444 378836 230450
rect 378784 230386 378836 230392
rect 378968 229152 379020 229158
rect 378968 229094 379020 229100
rect 378140 224256 378192 224262
rect 378140 224198 378192 224204
rect 377772 221604 377824 221610
rect 377772 221546 377824 221552
rect 377404 220244 377456 220250
rect 377404 220186 377456 220192
rect 376944 218204 376996 218210
rect 376944 218146 376996 218152
rect 376116 218068 376168 218074
rect 376116 218010 376168 218016
rect 376576 218068 376628 218074
rect 376576 218010 376628 218016
rect 375208 217246 375282 217274
rect 371942 217110 372016 217138
rect 372770 217110 372844 217138
rect 373598 217110 373672 217138
rect 374426 217110 374500 217138
rect 371942 216988 371970 217110
rect 372770 216988 372798 217110
rect 373598 216988 373626 217110
rect 374426 216988 374454 217110
rect 375254 216988 375282 217246
rect 376128 217138 376156 218010
rect 376956 217138 376984 218146
rect 377784 217274 377812 221546
rect 378980 219434 379008 229094
rect 379440 228410 379468 231676
rect 379428 228404 379480 228410
rect 379428 228346 379480 228352
rect 380084 225894 380112 231676
rect 380268 231662 380742 231690
rect 380072 225888 380124 225894
rect 380072 225830 380124 225836
rect 379336 225752 379388 225758
rect 379336 225694 379388 225700
rect 378796 219406 379008 219434
rect 378796 218890 378824 219406
rect 378784 218884 378836 218890
rect 378784 218826 378836 218832
rect 379152 218748 379204 218754
rect 379152 218690 379204 218696
rect 378600 218068 378652 218074
rect 378600 218010 378652 218016
rect 376082 217110 376156 217138
rect 376910 217110 376984 217138
rect 377738 217246 377812 217274
rect 376082 216988 376110 217110
rect 376910 216988 376938 217110
rect 377738 216988 377766 217246
rect 378612 217138 378640 218010
rect 379164 217274 379192 218690
rect 379348 218074 379376 225694
rect 380268 224346 380296 231662
rect 380440 230036 380492 230042
rect 380440 229978 380492 229984
rect 380452 229094 380480 229978
rect 381372 229906 381400 231676
rect 381360 229900 381412 229906
rect 381360 229842 381412 229848
rect 379900 224318 380296 224346
rect 380360 229066 380480 229094
rect 379900 221474 379928 224318
rect 380360 224210 380388 229066
rect 382016 228546 382044 231676
rect 382476 231662 382674 231690
rect 382004 228540 382056 228546
rect 382004 228482 382056 228488
rect 381728 228404 381780 228410
rect 381728 228346 381780 228352
rect 380084 224182 380388 224210
rect 379888 221468 379940 221474
rect 379888 221410 379940 221416
rect 380084 219026 380112 224182
rect 380256 219428 380308 219434
rect 380256 219370 380308 219376
rect 380072 219020 380124 219026
rect 380072 218962 380124 218968
rect 379336 218068 379388 218074
rect 379336 218010 379388 218016
rect 379164 217246 379422 217274
rect 378566 217110 378640 217138
rect 378566 216988 378594 217110
rect 379394 216988 379422 217246
rect 380268 217138 380296 219370
rect 381740 218074 381768 228346
rect 381912 227044 381964 227050
rect 381912 226986 381964 226992
rect 381084 218068 381136 218074
rect 381084 218010 381136 218016
rect 381728 218068 381780 218074
rect 381728 218010 381780 218016
rect 381096 217138 381124 218010
rect 381924 217274 381952 226986
rect 382476 220114 382504 231662
rect 382924 227316 382976 227322
rect 382924 227258 382976 227264
rect 382464 220108 382516 220114
rect 382464 220050 382516 220056
rect 382740 220108 382792 220114
rect 382740 220050 382792 220056
rect 382752 217274 382780 220050
rect 382936 218210 382964 227258
rect 383304 227186 383332 231676
rect 383948 229158 383976 231676
rect 384304 229900 384356 229906
rect 384304 229842 384356 229848
rect 383936 229152 383988 229158
rect 383936 229094 383988 229100
rect 383292 227180 383344 227186
rect 383292 227122 383344 227128
rect 384316 219434 384344 229842
rect 384592 223038 384620 231676
rect 384580 223032 384632 223038
rect 384580 222974 384632 222980
rect 385236 220522 385264 231676
rect 385880 227458 385908 231676
rect 386524 229770 386552 231676
rect 386512 229764 386564 229770
rect 386512 229706 386564 229712
rect 386972 229764 387024 229770
rect 386972 229706 387024 229712
rect 386984 229094 387012 229706
rect 387168 229094 387196 231676
rect 386984 229066 387104 229094
rect 387168 229066 387288 229094
rect 385868 227452 385920 227458
rect 385868 227394 385920 227400
rect 386328 227180 386380 227186
rect 386328 227122 386380 227128
rect 385224 220516 385276 220522
rect 385224 220458 385276 220464
rect 384304 219428 384356 219434
rect 384304 219370 384356 219376
rect 383568 219292 383620 219298
rect 383568 219234 383620 219240
rect 382924 218204 382976 218210
rect 382924 218146 382976 218152
rect 380222 217110 380296 217138
rect 381050 217110 381124 217138
rect 381878 217246 381952 217274
rect 382706 217246 382780 217274
rect 380222 216988 380250 217110
rect 381050 216988 381078 217110
rect 381878 216988 381906 217246
rect 382706 216988 382734 217246
rect 383580 217138 383608 219234
rect 384396 219020 384448 219026
rect 384396 218962 384448 218968
rect 384408 217138 384436 218962
rect 386052 218884 386104 218890
rect 386052 218826 386104 218832
rect 385224 218068 385276 218074
rect 385224 218010 385276 218016
rect 385236 217138 385264 218010
rect 386064 217138 386092 218826
rect 386340 218074 386368 227122
rect 387076 219298 387104 229066
rect 387260 228682 387288 229066
rect 387248 228676 387300 228682
rect 387248 228618 387300 228624
rect 387812 224398 387840 231676
rect 388088 231662 388470 231690
rect 388088 225622 388116 231662
rect 389100 230042 389128 231676
rect 389088 230036 389140 230042
rect 389088 229978 389140 229984
rect 389744 228818 389772 231676
rect 390020 231662 390402 231690
rect 389732 228812 389784 228818
rect 389732 228754 389784 228760
rect 388076 225616 388128 225622
rect 388076 225558 388128 225564
rect 388444 225616 388496 225622
rect 388444 225558 388496 225564
rect 387800 224392 387852 224398
rect 387800 224334 387852 224340
rect 387708 223032 387760 223038
rect 387708 222974 387760 222980
rect 387064 219292 387116 219298
rect 387064 219234 387116 219240
rect 386880 218204 386932 218210
rect 386880 218146 386932 218152
rect 386328 218068 386380 218074
rect 386328 218010 386380 218016
rect 386892 217138 386920 218146
rect 387720 217274 387748 222974
rect 388456 218210 388484 225558
rect 389088 224256 389140 224262
rect 389088 224198 389140 224204
rect 388444 218204 388496 218210
rect 388444 218146 388496 218152
rect 389100 218074 389128 224198
rect 390020 221610 390048 231662
rect 390284 228676 390336 228682
rect 390284 228618 390336 228624
rect 390008 221604 390060 221610
rect 390008 221546 390060 221552
rect 390100 220244 390152 220250
rect 390100 220186 390152 220192
rect 388536 218068 388588 218074
rect 388536 218010 388588 218016
rect 389088 218068 389140 218074
rect 389088 218010 389140 218016
rect 389364 218068 389416 218074
rect 389364 218010 389416 218016
rect 383534 217110 383608 217138
rect 384362 217110 384436 217138
rect 385190 217110 385264 217138
rect 386018 217110 386092 217138
rect 386846 217110 386920 217138
rect 387674 217246 387748 217274
rect 383534 216988 383562 217110
rect 384362 216988 384390 217110
rect 385190 216988 385218 217110
rect 386018 216988 386046 217110
rect 386846 216988 386874 217110
rect 387674 216988 387702 217246
rect 388548 217138 388576 218010
rect 389376 217138 389404 218010
rect 390112 217274 390140 220186
rect 390296 218074 390324 228618
rect 391032 222902 391060 231676
rect 391676 227322 391704 231676
rect 392136 231662 392334 231690
rect 391848 228404 391900 228410
rect 391848 228346 391900 228352
rect 391664 227316 391716 227322
rect 391664 227258 391716 227264
rect 391020 222896 391072 222902
rect 391020 222838 391072 222844
rect 391020 221468 391072 221474
rect 391020 221410 391072 221416
rect 390284 218068 390336 218074
rect 390284 218010 390336 218016
rect 391032 217274 391060 221410
rect 391860 217274 391888 228346
rect 392136 218754 392164 231662
rect 392964 228546 392992 231676
rect 392952 228540 393004 228546
rect 392952 228482 393004 228488
rect 393228 228540 393280 228546
rect 393228 228482 393280 228488
rect 392124 218748 392176 218754
rect 392124 218690 392176 218696
rect 393240 218074 393268 228482
rect 393608 225758 393636 231676
rect 394252 229906 394280 231676
rect 394804 231662 394910 231690
rect 394240 229900 394292 229906
rect 394240 229842 394292 229848
rect 393964 227792 394016 227798
rect 393964 227734 394016 227740
rect 393596 225752 393648 225758
rect 393596 225694 393648 225700
rect 393976 219026 394004 227734
rect 394608 225752 394660 225758
rect 394608 225694 394660 225700
rect 393964 219020 394016 219026
rect 393964 218962 394016 218968
rect 394332 218204 394384 218210
rect 394332 218146 394384 218152
rect 392676 218068 392728 218074
rect 392676 218010 392728 218016
rect 393228 218068 393280 218074
rect 393228 218010 393280 218016
rect 393504 218068 393556 218074
rect 393504 218010 393556 218016
rect 390112 217246 390186 217274
rect 388502 217110 388576 217138
rect 389330 217110 389404 217138
rect 388502 216988 388530 217110
rect 389330 216988 389358 217110
rect 390158 216988 390186 217246
rect 390986 217246 391060 217274
rect 391814 217246 391888 217274
rect 390986 216988 391014 217246
rect 391814 216988 391842 217246
rect 392688 217138 392716 218010
rect 393516 217138 393544 218010
rect 394344 217138 394372 218146
rect 394620 218074 394648 225694
rect 394804 220114 394832 231662
rect 395540 227798 395568 231676
rect 395528 227792 395580 227798
rect 395528 227734 395580 227740
rect 395988 227316 396040 227322
rect 395988 227258 396040 227264
rect 394792 220108 394844 220114
rect 394792 220050 394844 220056
rect 395804 218748 395856 218754
rect 395804 218690 395856 218696
rect 394608 218068 394660 218074
rect 394608 218010 394660 218016
rect 395160 218068 395212 218074
rect 395160 218010 395212 218016
rect 395172 217138 395200 218010
rect 395816 217274 395844 218690
rect 396000 218074 396028 227258
rect 396184 227050 396212 231676
rect 396828 229770 396856 231676
rect 396816 229764 396868 229770
rect 396816 229706 396868 229712
rect 397472 227798 397500 231676
rect 396632 227792 396684 227798
rect 396632 227734 396684 227740
rect 397460 227792 397512 227798
rect 397460 227734 397512 227740
rect 396172 227044 396224 227050
rect 396172 226986 396224 226992
rect 396644 218890 396672 227734
rect 398116 223038 398144 231676
rect 398760 227186 398788 231676
rect 398748 227180 398800 227186
rect 398748 227122 398800 227128
rect 398472 227044 398524 227050
rect 398472 226986 398524 226992
rect 398104 223032 398156 223038
rect 398104 222974 398156 222980
rect 397368 222896 397420 222902
rect 397368 222838 397420 222844
rect 396632 218884 396684 218890
rect 396632 218826 396684 218832
rect 397380 218074 397408 222838
rect 397644 220108 397696 220114
rect 397644 220050 397696 220056
rect 395988 218068 396040 218074
rect 395988 218010 396040 218016
rect 396816 218068 396868 218074
rect 396816 218010 396868 218016
rect 397368 218068 397420 218074
rect 397368 218010 397420 218016
rect 395816 217246 395982 217274
rect 392642 217110 392716 217138
rect 393470 217110 393544 217138
rect 394298 217110 394372 217138
rect 395126 217110 395200 217138
rect 392642 216988 392670 217110
rect 393470 216988 393498 217110
rect 394298 216988 394326 217110
rect 395126 216988 395154 217110
rect 395954 216988 395982 217246
rect 396828 217138 396856 218010
rect 397656 217274 397684 220050
rect 398484 217274 398512 226986
rect 399404 225622 399432 231676
rect 399852 229764 399904 229770
rect 399852 229706 399904 229712
rect 399392 225616 399444 225622
rect 399392 225558 399444 225564
rect 399864 219434 399892 229706
rect 400048 228682 400076 231676
rect 400416 231662 400706 231690
rect 400968 231662 401350 231690
rect 401704 231662 401994 231690
rect 400036 228676 400088 228682
rect 400036 228618 400088 228624
rect 400128 228540 400180 228546
rect 400128 228482 400180 228488
rect 400140 219434 400168 228482
rect 400416 221474 400444 231662
rect 400968 224262 400996 231662
rect 401416 228812 401468 228818
rect 401416 228754 401468 228760
rect 400956 224256 401008 224262
rect 400956 224198 401008 224204
rect 400404 221468 400456 221474
rect 400404 221410 400456 221416
rect 399300 219428 399352 219434
rect 399864 219406 400076 219434
rect 400140 219428 400272 219434
rect 400140 219406 400220 219428
rect 399300 219370 399352 219376
rect 396782 217110 396856 217138
rect 397610 217246 397684 217274
rect 398438 217246 398512 217274
rect 396782 216988 396810 217110
rect 397610 216988 397638 217246
rect 398438 216988 398466 217246
rect 399312 217138 399340 219370
rect 400048 217274 400076 219406
rect 400220 219370 400272 219376
rect 401428 218074 401456 228754
rect 401704 220250 401732 231662
rect 402624 228410 402652 231676
rect 402612 228404 402664 228410
rect 402612 228346 402664 228352
rect 403268 227798 403296 231676
rect 403912 228274 403940 231676
rect 404268 230376 404320 230382
rect 404268 230318 404320 230324
rect 403900 228268 403952 228274
rect 403900 228210 403952 228216
rect 402244 227792 402296 227798
rect 402244 227734 402296 227740
rect 403256 227792 403308 227798
rect 403256 227734 403308 227740
rect 404084 227792 404136 227798
rect 404084 227734 404136 227740
rect 401692 220244 401744 220250
rect 401692 220186 401744 220192
rect 401784 219020 401836 219026
rect 401784 218962 401836 218968
rect 400956 218068 401008 218074
rect 400956 218010 401008 218016
rect 401416 218068 401468 218074
rect 401416 218010 401468 218016
rect 400048 217246 400122 217274
rect 399266 217110 399340 217138
rect 399266 216988 399294 217110
rect 400094 216988 400122 217246
rect 400968 217138 400996 218010
rect 401796 217138 401824 218962
rect 402256 218210 402284 227734
rect 404096 219434 404124 227734
rect 404280 219434 404308 230318
rect 404556 225758 404584 231676
rect 404740 231662 405214 231690
rect 404544 225752 404596 225758
rect 404544 225694 404596 225700
rect 404740 219434 404768 231662
rect 405096 221468 405148 221474
rect 405096 221410 405148 221416
rect 403440 219428 403492 219434
rect 404096 219406 404216 219434
rect 404280 219428 404412 219434
rect 404280 219406 404360 219428
rect 403440 219370 403492 219376
rect 402612 218884 402664 218890
rect 402612 218826 402664 218832
rect 402244 218204 402296 218210
rect 402244 218146 402296 218152
rect 402624 217138 402652 218826
rect 403452 217138 403480 219370
rect 404188 217274 404216 219406
rect 404360 219370 404412 219376
rect 404556 219406 404768 219434
rect 404556 218754 404584 219406
rect 404544 218748 404596 218754
rect 404544 218690 404596 218696
rect 405108 217274 405136 221410
rect 405844 220114 405872 231676
rect 406488 227322 406516 231676
rect 406476 227316 406528 227322
rect 406476 227258 406528 227264
rect 406752 224936 406804 224942
rect 406752 224878 406804 224884
rect 405832 220108 405884 220114
rect 405832 220050 405884 220056
rect 405924 219496 405976 219502
rect 405924 219438 405976 219444
rect 405936 217274 405964 219438
rect 406764 217274 406792 224878
rect 407132 222902 407160 231676
rect 407776 228546 407804 231676
rect 408420 228818 408448 231676
rect 408696 231662 409078 231690
rect 408408 228812 408460 228818
rect 408408 228754 408460 228760
rect 407764 228540 407816 228546
rect 407764 228482 407816 228488
rect 407764 227928 407816 227934
rect 407764 227870 407816 227876
rect 407120 222896 407172 222902
rect 407120 222838 407172 222844
rect 407776 219026 407804 227870
rect 408696 227050 408724 231662
rect 408868 230240 408920 230246
rect 408868 230182 408920 230188
rect 408880 227798 408908 230182
rect 409708 229770 409736 231676
rect 409696 229764 409748 229770
rect 409696 229706 409748 229712
rect 409788 228404 409840 228410
rect 409788 228346 409840 228352
rect 408868 227792 408920 227798
rect 408868 227734 408920 227740
rect 409052 227792 409104 227798
rect 409052 227734 409104 227740
rect 408684 227044 408736 227050
rect 408684 226986 408736 226992
rect 408408 222896 408460 222902
rect 408408 222838 408460 222844
rect 407764 219020 407816 219026
rect 407764 218962 407816 218968
rect 407580 218204 407632 218210
rect 407580 218146 407632 218152
rect 404188 217246 404262 217274
rect 400922 217110 400996 217138
rect 401750 217110 401824 217138
rect 402578 217110 402652 217138
rect 403406 217110 403480 217138
rect 400922 216988 400950 217110
rect 401750 216988 401778 217110
rect 402578 216988 402606 217110
rect 403406 216988 403434 217110
rect 404234 216988 404262 217246
rect 405062 217246 405136 217274
rect 405890 217246 405964 217274
rect 406718 217246 406792 217274
rect 405062 216988 405090 217246
rect 405890 216988 405918 217246
rect 406718 216988 406746 217246
rect 407592 217138 407620 218146
rect 408420 217274 408448 222838
rect 409064 218890 409092 227734
rect 409052 218884 409104 218890
rect 409052 218826 409104 218832
rect 409800 218074 409828 228346
rect 410352 227798 410380 231676
rect 410996 230246 411024 231676
rect 410984 230240 411036 230246
rect 410984 230182 411036 230188
rect 411168 229764 411220 229770
rect 411168 229706 411220 229712
rect 410892 228676 410944 228682
rect 410892 228618 410944 228624
rect 410340 227792 410392 227798
rect 410340 227734 410392 227740
rect 409236 218068 409288 218074
rect 409236 218010 409288 218016
rect 409788 218068 409840 218074
rect 409788 218010 409840 218016
rect 410064 218068 410116 218074
rect 410064 218010 410116 218016
rect 407546 217110 407620 217138
rect 408374 217246 408448 217274
rect 407546 216988 407574 217110
rect 408374 216988 408402 217246
rect 409248 217138 409276 218010
rect 410076 217138 410104 218010
rect 410904 217274 410932 228618
rect 411180 218074 411208 229706
rect 411640 227934 411668 231676
rect 412284 230382 412312 231676
rect 412744 231662 412942 231690
rect 412272 230376 412324 230382
rect 412272 230318 412324 230324
rect 412456 229900 412508 229906
rect 412456 229842 412508 229848
rect 411628 227928 411680 227934
rect 411628 227870 411680 227876
rect 411904 227792 411956 227798
rect 411904 227734 411956 227740
rect 411720 218884 411772 218890
rect 411720 218826 411772 218832
rect 411168 218068 411220 218074
rect 411168 218010 411220 218016
rect 409202 217110 409276 217138
rect 410030 217110 410104 217138
rect 410858 217246 410932 217274
rect 409202 216988 409230 217110
rect 410030 216988 410058 217110
rect 410858 216988 410886 217246
rect 411732 217138 411760 218826
rect 411916 218210 411944 227734
rect 412468 218890 412496 229842
rect 412744 219502 412772 231662
rect 413572 227798 413600 231676
rect 413836 229084 413888 229090
rect 413836 229026 413888 229032
rect 413560 227792 413612 227798
rect 413560 227734 413612 227740
rect 412732 219496 412784 219502
rect 412732 219438 412784 219444
rect 412456 218884 412508 218890
rect 412456 218826 412508 218832
rect 412548 218748 412600 218754
rect 412548 218690 412600 218696
rect 411904 218204 411956 218210
rect 411904 218146 411956 218152
rect 412560 217138 412588 218690
rect 413848 218074 413876 229026
rect 414216 221474 414244 231676
rect 414860 224942 414888 231676
rect 415504 228410 415532 231676
rect 416148 228682 416176 231676
rect 416792 229094 416820 231676
rect 417436 229770 417464 231676
rect 417712 231662 418094 231690
rect 418264 231662 418738 231690
rect 417424 229764 417476 229770
rect 417424 229706 417476 229712
rect 417712 229094 417740 231662
rect 416792 229066 416912 229094
rect 416136 228676 416188 228682
rect 416136 228618 416188 228624
rect 415492 228404 415544 228410
rect 415492 228346 415544 228352
rect 416688 227792 416740 227798
rect 416688 227734 416740 227740
rect 414848 224936 414900 224942
rect 414848 224878 414900 224884
rect 416504 224256 416556 224262
rect 416504 224198 416556 224204
rect 414204 221468 414256 221474
rect 414204 221410 414256 221416
rect 415032 221060 415084 221066
rect 415032 221002 415084 221008
rect 414204 220788 414256 220794
rect 414204 220730 414256 220736
rect 413376 218068 413428 218074
rect 413376 218010 413428 218016
rect 413836 218068 413888 218074
rect 413836 218010 413888 218016
rect 413388 217138 413416 218010
rect 414216 217274 414244 220730
rect 415044 217274 415072 221002
rect 416516 219434 416544 224198
rect 416700 219434 416728 227734
rect 416884 222902 416912 229066
rect 417160 229066 417740 229094
rect 416872 222896 416924 222902
rect 416872 222838 416924 222844
rect 415860 219428 415912 219434
rect 416516 219406 416636 219434
rect 416700 219428 416832 219434
rect 416700 219406 416780 219428
rect 415860 219370 415912 219376
rect 411686 217110 411760 217138
rect 412514 217110 412588 217138
rect 413342 217110 413416 217138
rect 414170 217246 414244 217274
rect 414998 217246 415072 217274
rect 411686 216988 411714 217110
rect 412514 216988 412542 217110
rect 413342 216988 413370 217110
rect 414170 216988 414198 217246
rect 414998 216988 415026 217246
rect 415872 217138 415900 219370
rect 416608 217274 416636 219406
rect 416780 219370 416832 219376
rect 417160 218754 417188 229066
rect 418264 220794 418292 231662
rect 419368 229906 419396 231676
rect 419356 229900 419408 229906
rect 419356 229842 419408 229848
rect 419448 229288 419500 229294
rect 419448 229230 419500 229236
rect 418252 220788 418304 220794
rect 418252 220730 418304 220736
rect 417516 219428 417568 219434
rect 417516 219370 417568 219376
rect 417148 218748 417200 218754
rect 417148 218690 417200 218696
rect 416608 217246 416682 217274
rect 415826 217110 415900 217138
rect 415826 216988 415854 217110
rect 416654 216988 416682 217246
rect 417528 217138 417556 219370
rect 419172 219292 419224 219298
rect 419172 219234 419224 219240
rect 418344 218068 418396 218074
rect 418344 218010 418396 218016
rect 418356 217138 418384 218010
rect 419184 217138 419212 219234
rect 419460 218074 419488 229230
rect 420012 229158 420040 231676
rect 420000 229152 420052 229158
rect 420000 229094 420052 229100
rect 420184 229152 420236 229158
rect 420184 229094 420236 229100
rect 420196 221066 420224 229094
rect 420656 227798 420684 231676
rect 421024 231662 421314 231690
rect 420644 227792 420696 227798
rect 420644 227734 420696 227740
rect 420828 222896 420880 222902
rect 420828 222838 420880 222844
rect 420184 221060 420236 221066
rect 420184 221002 420236 221008
rect 420644 220856 420696 220862
rect 420644 220798 420696 220804
rect 420656 219434 420684 220798
rect 420656 219406 420776 219434
rect 419448 218068 419500 218074
rect 419448 218010 419500 218016
rect 420000 218068 420052 218074
rect 420000 218010 420052 218016
rect 420012 217138 420040 218010
rect 420748 217274 420776 219406
rect 420840 218090 420868 222838
rect 421024 219502 421052 231662
rect 421944 229158 421972 231676
rect 422312 231662 422602 231690
rect 422864 231662 423246 231690
rect 423784 231662 423890 231690
rect 421932 229152 421984 229158
rect 421932 229094 421984 229100
rect 422312 229094 422340 231662
rect 422220 229066 422340 229094
rect 422220 224262 422248 229066
rect 422208 224256 422260 224262
rect 422208 224198 422260 224204
rect 421656 220108 421708 220114
rect 421656 220050 421708 220056
rect 421012 219496 421064 219502
rect 421012 219438 421064 219444
rect 420840 218074 420960 218090
rect 420840 218068 420972 218074
rect 420840 218062 420920 218068
rect 420920 218010 420972 218016
rect 421668 217274 421696 220050
rect 422864 219434 422892 231662
rect 423312 224256 423364 224262
rect 423312 224198 423364 224204
rect 422680 219406 422892 219434
rect 422680 219298 422708 219406
rect 422668 219292 422720 219298
rect 422668 219234 422720 219240
rect 422484 218204 422536 218210
rect 422484 218146 422536 218152
rect 420748 217246 420822 217274
rect 417482 217110 417556 217138
rect 418310 217110 418384 217138
rect 419138 217110 419212 217138
rect 419966 217110 420040 217138
rect 417482 216988 417510 217110
rect 418310 216988 418338 217110
rect 419138 216988 419166 217110
rect 419966 216988 419994 217110
rect 420794 216988 420822 217246
rect 421622 217246 421696 217274
rect 421622 216988 421650 217246
rect 422496 217138 422524 218146
rect 423324 217274 423352 224198
rect 423784 220862 423812 231662
rect 424520 229294 424548 231676
rect 424508 229288 424560 229294
rect 424508 229230 424560 229236
rect 424324 229152 424376 229158
rect 424324 229094 424376 229100
rect 424336 224262 424364 229094
rect 424324 224256 424376 224262
rect 424324 224198 424376 224204
rect 425164 222902 425192 231676
rect 425440 231662 425822 231690
rect 425152 222896 425204 222902
rect 425152 222838 425204 222844
rect 424968 222148 425020 222154
rect 424968 222090 425020 222096
rect 423772 220856 423824 220862
rect 423772 220798 423824 220804
rect 424140 218068 424192 218074
rect 424140 218010 424192 218016
rect 422450 217110 422524 217138
rect 423278 217246 423352 217274
rect 422450 216988 422478 217110
rect 423278 216988 423306 217246
rect 424152 217138 424180 218010
rect 424980 217274 425008 222090
rect 425440 218210 425468 231662
rect 426452 223650 426480 231676
rect 426820 231662 427110 231690
rect 426440 223644 426492 223650
rect 426440 223586 426492 223592
rect 426820 220114 426848 231662
rect 427740 229158 427768 231676
rect 427728 229152 427780 229158
rect 427728 229094 427780 229100
rect 428384 229094 428412 231676
rect 428752 231662 429042 231690
rect 429304 231662 429686 231690
rect 429948 231662 430330 231690
rect 430684 231662 430974 231690
rect 431236 231662 431618 231690
rect 432064 231662 432262 231690
rect 432708 231662 432906 231690
rect 433550 231662 433748 231690
rect 428384 229066 428504 229094
rect 426992 223644 427044 223650
rect 426992 223586 427044 223592
rect 426808 220108 426860 220114
rect 426808 220050 426860 220056
rect 426624 218340 426676 218346
rect 426624 218282 426676 218288
rect 425428 218204 425480 218210
rect 425428 218146 425480 218152
rect 425796 218204 425848 218210
rect 425796 218146 425848 218152
rect 424106 217110 424180 217138
rect 424934 217246 425008 217274
rect 424106 216988 424134 217110
rect 424934 216988 424962 217246
rect 425808 217138 425836 218146
rect 426636 217138 426664 218282
rect 427004 218074 427032 223586
rect 427912 220108 427964 220114
rect 427912 220050 427964 220056
rect 427924 218074 427952 220050
rect 428280 219428 428332 219434
rect 428280 219370 428332 219376
rect 426992 218068 427044 218074
rect 426992 218010 427044 218016
rect 427452 218068 427504 218074
rect 427452 218010 427504 218016
rect 427912 218068 427964 218074
rect 427912 218010 427964 218016
rect 427464 217138 427492 218010
rect 428292 217138 428320 219370
rect 428476 218210 428504 229066
rect 428752 220114 428780 231662
rect 429304 222154 429332 231662
rect 429292 222148 429344 222154
rect 429292 222090 429344 222096
rect 428740 220108 428792 220114
rect 428740 220050 428792 220056
rect 429948 219434 429976 231662
rect 430684 219434 430712 231662
rect 431236 219434 431264 231662
rect 432064 219570 432092 231662
rect 432236 220244 432288 220250
rect 432236 220186 432288 220192
rect 432052 219564 432104 219570
rect 432052 219506 432104 219512
rect 432248 219434 432276 220186
rect 429580 219406 429976 219434
rect 430592 219406 430712 219434
rect 430776 219406 431264 219434
rect 431972 219406 432276 219434
rect 429580 218346 429608 219406
rect 429936 218748 429988 218754
rect 429936 218690 429988 218696
rect 429568 218340 429620 218346
rect 429568 218282 429620 218288
rect 428464 218204 428516 218210
rect 428464 218146 428516 218152
rect 429108 218068 429160 218074
rect 429108 218010 429160 218016
rect 429120 217138 429148 218010
rect 429948 217138 429976 218690
rect 430592 218074 430620 219406
rect 430580 218068 430632 218074
rect 430580 218010 430632 218016
rect 430776 217274 430804 219406
rect 431972 218090 432000 219406
rect 432708 218754 432736 231662
rect 433524 229832 433576 229838
rect 433524 229774 433576 229780
rect 433536 229094 433564 229774
rect 433720 229094 433748 231662
rect 434180 229838 434208 231676
rect 434168 229832 434220 229838
rect 434168 229774 434220 229780
rect 433536 229066 433656 229094
rect 433720 229066 433840 229094
rect 432696 218748 432748 218754
rect 432696 218690 432748 218696
rect 433248 218204 433300 218210
rect 433248 218146 433300 218152
rect 425762 217110 425836 217138
rect 426590 217110 426664 217138
rect 427418 217110 427492 217138
rect 428246 217110 428320 217138
rect 429074 217110 429148 217138
rect 429902 217110 429976 217138
rect 430730 217246 430804 217274
rect 431604 218062 432000 218090
rect 432420 218068 432472 218074
rect 425762 216988 425790 217110
rect 426590 216988 426618 217110
rect 427418 216988 427446 217110
rect 428246 216988 428274 217110
rect 429074 216988 429102 217110
rect 429902 216988 429930 217110
rect 430730 216988 430758 217246
rect 431604 217138 431632 218062
rect 432420 218010 432472 218016
rect 432432 217138 432460 218010
rect 433260 217138 433288 218146
rect 433628 217274 433656 229066
rect 433812 218074 433840 229066
rect 434824 220250 434852 231676
rect 435284 231662 435482 231690
rect 436126 231662 436324 231690
rect 434812 220244 434864 220250
rect 434812 220186 434864 220192
rect 434904 218340 434956 218346
rect 434904 218282 434956 218288
rect 433800 218068 433852 218074
rect 433800 218010 433852 218016
rect 433628 217246 434070 217274
rect 431558 217110 431632 217138
rect 432386 217110 432460 217138
rect 433214 217110 433288 217138
rect 431558 216988 431586 217110
rect 432386 216988 432414 217110
rect 433214 216988 433242 217110
rect 434042 216988 434070 217246
rect 434916 217138 434944 218282
rect 435284 218210 435312 231662
rect 436100 230376 436152 230382
rect 436100 230318 436152 230324
rect 435272 218204 435324 218210
rect 435272 218146 435324 218152
rect 435732 218068 435784 218074
rect 435732 218010 435784 218016
rect 435744 217138 435772 218010
rect 436112 217258 436140 230318
rect 436296 218074 436324 231662
rect 436756 230382 436784 231676
rect 436940 231662 437414 231690
rect 437768 231662 438058 231690
rect 436744 230376 436796 230382
rect 436744 230318 436796 230324
rect 436940 219434 436968 231662
rect 437768 219434 437796 231662
rect 438688 230382 438716 231676
rect 439332 230586 439360 231676
rect 439516 231662 439990 231690
rect 440344 231662 440634 231690
rect 439320 230580 439372 230586
rect 439320 230522 439372 230528
rect 439516 230466 439544 231662
rect 438964 230438 439544 230466
rect 438676 230376 438728 230382
rect 438676 230318 438728 230324
rect 438964 219434 438992 230438
rect 439320 230376 439372 230382
rect 439320 230318 439372 230324
rect 439332 219434 439360 230318
rect 436664 219406 436968 219434
rect 437492 219406 437796 219434
rect 438872 219406 438992 219434
rect 439056 219406 439360 219434
rect 436664 218346 436692 219406
rect 436652 218340 436704 218346
rect 436652 218282 436704 218288
rect 437492 218074 437520 219406
rect 438872 218074 438900 219406
rect 436284 218068 436336 218074
rect 436284 218010 436336 218016
rect 436560 218068 436612 218074
rect 436560 218010 436612 218016
rect 437480 218068 437532 218074
rect 437480 218010 437532 218016
rect 438216 218068 438268 218074
rect 438216 218010 438268 218016
rect 438860 218068 438912 218074
rect 438860 218010 438912 218016
rect 436100 217252 436152 217258
rect 436100 217194 436152 217200
rect 436572 217138 436600 218010
rect 437342 217252 437394 217258
rect 437342 217194 437394 217200
rect 434870 217110 434944 217138
rect 435698 217110 435772 217138
rect 436526 217110 436600 217138
rect 434870 216988 434898 217110
rect 435698 216988 435726 217110
rect 436526 216988 436554 217110
rect 437354 216988 437382 217194
rect 438228 217138 438256 218010
rect 439056 217274 439084 219406
rect 440344 218074 440372 231662
rect 440700 230444 440752 230450
rect 440700 230386 440752 230392
rect 439872 218068 439924 218074
rect 439872 218010 439924 218016
rect 440332 218068 440384 218074
rect 440332 218010 440384 218016
rect 438182 217110 438256 217138
rect 439010 217246 439084 217274
rect 438182 216988 438210 217110
rect 439010 216988 439038 217246
rect 439884 217138 439912 218010
rect 440712 217274 440740 230386
rect 441264 229158 441292 231676
rect 441908 230450 441936 231676
rect 442092 231662 442566 231690
rect 443104 231662 443210 231690
rect 441896 230444 441948 230450
rect 441896 230386 441948 230392
rect 442092 230330 442120 231662
rect 441724 230302 442120 230330
rect 441252 229152 441304 229158
rect 441252 229094 441304 229100
rect 441724 219434 441752 230302
rect 442080 229152 442132 229158
rect 442080 229094 442132 229100
rect 442092 229066 442304 229094
rect 441632 219406 441752 219434
rect 441632 218090 441660 219406
rect 439838 217110 439912 217138
rect 440666 217246 440740 217274
rect 441540 218062 441660 218090
rect 439838 216988 439866 217110
rect 440666 216988 440694 217246
rect 441540 217138 441568 218062
rect 442276 217274 442304 229066
rect 443104 217274 443132 231662
rect 443460 230444 443512 230450
rect 443460 230386 443512 230392
rect 443472 229094 443500 230386
rect 443840 230382 443868 231676
rect 443828 230376 443880 230382
rect 443828 230318 443880 230324
rect 444484 230110 444512 231676
rect 444668 231662 445142 231690
rect 444472 230104 444524 230110
rect 444472 230046 444524 230052
rect 444668 229094 444696 231662
rect 444840 230376 444892 230382
rect 444840 230318 444892 230324
rect 444852 229094 444880 230318
rect 445772 229094 445800 231676
rect 446416 230382 446444 231676
rect 446404 230376 446456 230382
rect 446404 230318 446456 230324
rect 447060 230246 447088 231676
rect 447244 231662 447718 231690
rect 447048 230240 447100 230246
rect 447048 230182 447100 230188
rect 443472 229066 443960 229094
rect 444668 229066 444788 229094
rect 444852 229066 445616 229094
rect 445772 229066 446444 229094
rect 443932 217274 443960 229066
rect 444760 217274 444788 229066
rect 445588 217274 445616 229066
rect 446416 217274 446444 229066
rect 447244 219434 447272 231662
rect 447600 230104 447652 230110
rect 447600 230046 447652 230052
rect 447612 219434 447640 230046
rect 448348 229094 448376 231676
rect 448992 229430 449020 231676
rect 449636 230382 449664 231676
rect 449164 230376 449216 230382
rect 449164 230318 449216 230324
rect 449624 230376 449676 230382
rect 449624 230318 449676 230324
rect 448980 229424 449032 229430
rect 448980 229366 449032 229372
rect 448348 229066 448652 229094
rect 447152 219406 447272 219434
rect 447336 219406 447640 219434
rect 442276 217246 442350 217274
rect 443104 217246 443178 217274
rect 443932 217246 444006 217274
rect 444760 217246 444834 217274
rect 445588 217246 445662 217274
rect 446416 217246 446490 217274
rect 447152 217258 447180 219406
rect 447336 217274 447364 219406
rect 441494 217110 441568 217138
rect 441494 216988 441522 217110
rect 442322 216988 442350 217246
rect 443150 216988 443178 217246
rect 443978 216988 444006 217246
rect 444806 216988 444834 217246
rect 445634 216988 445662 217246
rect 446462 216988 446490 217246
rect 447140 217252 447192 217258
rect 447140 217194 447192 217200
rect 447290 217246 447364 217274
rect 448624 217258 448652 229066
rect 449176 219434 449204 230318
rect 449900 230240 449952 230246
rect 449900 230182 449952 230188
rect 448992 219406 449204 219434
rect 449912 219434 449940 230182
rect 450280 229294 450308 231676
rect 450544 230376 450596 230382
rect 450544 230318 450596 230324
rect 450268 229288 450320 229294
rect 450268 229230 450320 229236
rect 450556 229094 450584 230318
rect 450924 229158 450952 231676
rect 451568 230246 451596 231676
rect 452226 231662 452608 231690
rect 451556 230240 451608 230246
rect 451556 230182 451608 230188
rect 451372 229424 451424 229430
rect 451372 229366 451424 229372
rect 450912 229152 450964 229158
rect 450912 229094 450964 229100
rect 450556 229066 450768 229094
rect 449912 219406 450584 219434
rect 448992 217274 449020 219406
rect 448106 217252 448158 217258
rect 447290 216988 447318 217246
rect 448106 217194 448158 217200
rect 448612 217252 448664 217258
rect 448612 217194 448664 217200
rect 448946 217246 449020 217274
rect 450556 217274 450584 219406
rect 450740 219298 450768 229066
rect 451384 224262 451412 229366
rect 451832 229288 451884 229294
rect 451832 229230 451884 229236
rect 451372 224256 451424 224262
rect 451372 224198 451424 224204
rect 451844 219434 451872 229230
rect 452200 224256 452252 224262
rect 452200 224198 452252 224204
rect 451476 219406 451872 219434
rect 450728 219292 450780 219298
rect 450728 219234 450780 219240
rect 451476 217274 451504 219406
rect 449762 217252 449814 217258
rect 448118 216988 448146 217194
rect 448946 216988 448974 217246
rect 450556 217246 450630 217274
rect 449762 217194 449814 217200
rect 449774 216988 449802 217194
rect 450602 216988 450630 217246
rect 451430 217246 451504 217274
rect 452212 217274 452240 224198
rect 452580 221474 452608 231662
rect 452856 230382 452884 231676
rect 452844 230376 452896 230382
rect 452844 230318 452896 230324
rect 453304 230240 453356 230246
rect 453304 230182 453356 230188
rect 452752 229152 452804 229158
rect 452752 229094 452804 229100
rect 452764 229066 453068 229094
rect 452568 221468 452620 221474
rect 452568 221410 452620 221416
rect 453040 217274 453068 229066
rect 453316 218074 453344 230182
rect 453500 229362 453528 231676
rect 454144 230246 454172 231676
rect 454802 231662 455092 231690
rect 454316 230376 454368 230382
rect 454316 230318 454368 230324
rect 454132 230240 454184 230246
rect 454132 230182 454184 230188
rect 453488 229356 453540 229362
rect 453488 229298 453540 229304
rect 454328 229094 454356 230318
rect 454328 229066 454724 229094
rect 453856 219292 453908 219298
rect 453856 219234 453908 219240
rect 453304 218068 453356 218074
rect 453304 218010 453356 218016
rect 452212 217246 452286 217274
rect 453040 217246 453114 217274
rect 451430 216988 451458 217246
rect 452258 216988 452286 217246
rect 453086 216988 453114 217246
rect 453868 217138 453896 219234
rect 454696 217274 454724 229066
rect 455064 218210 455092 231662
rect 455432 230382 455460 231676
rect 455420 230376 455472 230382
rect 455420 230318 455472 230324
rect 455236 230240 455288 230246
rect 455236 230182 455288 230188
rect 455248 220794 455276 230182
rect 455788 229356 455840 229362
rect 455788 229298 455840 229304
rect 455236 220788 455288 220794
rect 455236 220730 455288 220736
rect 455800 219434 455828 229298
rect 456076 224602 456104 231676
rect 456064 224596 456116 224602
rect 456064 224538 456116 224544
rect 456720 221610 456748 231676
rect 457168 230376 457220 230382
rect 457168 230318 457220 230324
rect 456708 221604 456760 221610
rect 456708 221546 456760 221552
rect 456708 221468 456760 221474
rect 456708 221410 456760 221416
rect 455800 219406 456380 219434
rect 455052 218204 455104 218210
rect 455052 218146 455104 218152
rect 455512 218068 455564 218074
rect 455512 218010 455564 218016
rect 454696 217246 454770 217274
rect 453868 217110 453942 217138
rect 453914 216988 453942 217110
rect 454742 216988 454770 217246
rect 455524 217138 455552 218010
rect 456352 217274 456380 219406
rect 456720 218074 456748 221410
rect 457180 219434 457208 230318
rect 457364 229770 457392 231676
rect 457352 229764 457404 229770
rect 457352 229706 457404 229712
rect 458008 223582 458036 231676
rect 458652 225826 458680 231676
rect 459310 231662 459508 231690
rect 458640 225820 458692 225826
rect 458640 225762 458692 225768
rect 457996 223576 458048 223582
rect 457996 223518 458048 223524
rect 458824 220788 458876 220794
rect 458824 220730 458876 220736
rect 457180 219406 458036 219434
rect 456708 218068 456760 218074
rect 456708 218010 456760 218016
rect 457168 218068 457220 218074
rect 457168 218010 457220 218016
rect 456352 217246 456426 217274
rect 455524 217110 455598 217138
rect 455570 216988 455598 217110
rect 456398 216988 456426 217246
rect 457180 217138 457208 218010
rect 458008 217274 458036 219406
rect 458836 217274 458864 220730
rect 459480 220250 459508 231662
rect 459652 224596 459704 224602
rect 459652 224538 459704 224544
rect 459468 220244 459520 220250
rect 459468 220186 459520 220192
rect 459664 217274 459692 224538
rect 459940 222902 459968 231676
rect 460584 224738 460612 231676
rect 461242 231662 461716 231690
rect 461886 231662 462176 231690
rect 461688 229094 461716 231662
rect 461688 229066 461992 229094
rect 460572 224732 460624 224738
rect 460572 224674 460624 224680
rect 460204 223576 460256 223582
rect 460204 223518 460256 223524
rect 459928 222896 459980 222902
rect 459928 222838 459980 222844
rect 460216 218754 460244 223518
rect 460204 218748 460256 218754
rect 460204 218690 460256 218696
rect 461308 218748 461360 218754
rect 461308 218690 461360 218696
rect 460480 218204 460532 218210
rect 460480 218146 460532 218152
rect 458008 217246 458082 217274
rect 458836 217246 458910 217274
rect 459664 217246 459738 217274
rect 457180 217110 457254 217138
rect 457226 216988 457254 217110
rect 458054 216988 458082 217246
rect 458882 216988 458910 217246
rect 459710 216988 459738 217246
rect 460492 217138 460520 218146
rect 461320 217138 461348 218690
rect 461964 218210 461992 229066
rect 462148 222154 462176 231662
rect 462516 224398 462544 231676
rect 462964 225820 463016 225826
rect 462964 225762 463016 225768
rect 462504 224392 462556 224398
rect 462504 224334 462556 224340
rect 462136 222148 462188 222154
rect 462136 222090 462188 222096
rect 462136 221604 462188 221610
rect 462136 221546 462188 221552
rect 461952 218204 462004 218210
rect 461952 218146 462004 218152
rect 462148 217274 462176 221546
rect 462976 217274 463004 225762
rect 463160 225418 463188 231676
rect 463804 230382 463832 231676
rect 464462 231662 465028 231690
rect 465106 231662 465488 231690
rect 465750 231662 465948 231690
rect 463792 230376 463844 230382
rect 463792 230318 463844 230324
rect 463884 229764 463936 229770
rect 463884 229706 463936 229712
rect 463148 225412 463200 225418
rect 463148 225354 463200 225360
rect 463148 224732 463200 224738
rect 463148 224674 463200 224680
rect 463160 218074 463188 224674
rect 463148 218068 463200 218074
rect 463148 218010 463200 218016
rect 463896 217274 463924 229706
rect 465000 219638 465028 231662
rect 465460 229770 465488 231662
rect 465724 230376 465776 230382
rect 465724 230318 465776 230324
rect 465448 229764 465500 229770
rect 465448 229706 465500 229712
rect 465736 220726 465764 230318
rect 465920 227662 465948 231662
rect 466104 231662 466394 231690
rect 465908 227656 465960 227662
rect 465908 227598 465960 227604
rect 466104 220862 466132 231662
rect 467024 229906 467052 231676
rect 467012 229900 467064 229906
rect 467012 229842 467064 229848
rect 467472 229764 467524 229770
rect 467472 229706 467524 229712
rect 467288 225412 467340 225418
rect 467288 225354 467340 225360
rect 467104 222896 467156 222902
rect 467104 222838 467156 222844
rect 466092 220856 466144 220862
rect 466092 220798 466144 220804
rect 465724 220720 465776 220726
rect 465724 220662 465776 220668
rect 465448 220244 465500 220250
rect 465448 220186 465500 220192
rect 464988 219632 465040 219638
rect 464988 219574 465040 219580
rect 464620 218068 464672 218074
rect 464620 218010 464672 218016
rect 462148 217246 462222 217274
rect 462976 217246 463050 217274
rect 460492 217110 460566 217138
rect 461320 217110 461394 217138
rect 460538 216988 460566 217110
rect 461366 216988 461394 217110
rect 462194 216988 462222 217246
rect 463022 216988 463050 217246
rect 463850 217246 463924 217274
rect 463850 216988 463878 217246
rect 464632 217138 464660 218010
rect 465460 217274 465488 220186
rect 466276 218204 466328 218210
rect 466276 218146 466328 218152
rect 465460 217246 465534 217274
rect 464632 217110 464706 217138
rect 464678 216988 464706 217110
rect 465506 216988 465534 217246
rect 466288 217138 466316 218146
rect 467116 217274 467144 222838
rect 467300 218074 467328 225354
rect 467484 222902 467512 229706
rect 467668 225622 467696 231676
rect 468312 230450 468340 231676
rect 468864 231662 468970 231690
rect 468300 230444 468352 230450
rect 468300 230386 468352 230392
rect 468864 230042 468892 231662
rect 469036 230444 469088 230450
rect 469036 230386 469088 230392
rect 468852 230036 468904 230042
rect 468852 229978 468904 229984
rect 467656 225616 467708 225622
rect 467656 225558 467708 225564
rect 467472 222896 467524 222902
rect 467472 222838 467524 222844
rect 468760 222148 468812 222154
rect 468760 222090 468812 222096
rect 467288 218068 467340 218074
rect 467288 218010 467340 218016
rect 467932 218068 467984 218074
rect 467932 218010 467984 218016
rect 467116 217246 467190 217274
rect 466288 217110 466362 217138
rect 466334 216988 466362 217110
rect 467162 216988 467190 217246
rect 467944 217138 467972 218010
rect 468772 217274 468800 222090
rect 469048 220250 469076 230386
rect 469600 229770 469628 231676
rect 469588 229764 469640 229770
rect 469588 229706 469640 229712
rect 469864 227656 469916 227662
rect 469864 227598 469916 227604
rect 469312 224392 469364 224398
rect 469312 224334 469364 224340
rect 469036 220244 469088 220250
rect 469036 220186 469088 220192
rect 468772 217246 468846 217274
rect 469324 217258 469352 224334
rect 469588 220720 469640 220726
rect 469588 220662 469640 220668
rect 469600 217274 469628 220662
rect 469876 218618 469904 227598
rect 470244 224398 470272 231676
rect 470888 230246 470916 231676
rect 470876 230240 470928 230246
rect 470876 230182 470928 230188
rect 471532 227934 471560 231676
rect 471888 230240 471940 230246
rect 471888 230182 471940 230188
rect 471520 227928 471572 227934
rect 471520 227870 471572 227876
rect 470232 224392 470284 224398
rect 470232 224334 470284 224340
rect 471900 222154 471928 230182
rect 472176 227050 472204 231676
rect 472834 231662 473032 231690
rect 472164 227044 472216 227050
rect 472164 226986 472216 226992
rect 471888 222148 471940 222154
rect 471888 222090 471940 222096
rect 470600 220856 470652 220862
rect 470600 220798 470652 220804
rect 469864 218612 469916 218618
rect 469864 218554 469916 218560
rect 470612 218074 470640 220798
rect 473004 220114 473032 231662
rect 473464 223582 473492 231676
rect 474122 231662 474504 231690
rect 474766 231662 475056 231690
rect 474004 229900 474056 229906
rect 474004 229842 474056 229848
rect 473452 223576 473504 223582
rect 473452 223518 473504 223524
rect 473728 222896 473780 222902
rect 473728 222838 473780 222844
rect 472992 220108 473044 220114
rect 472992 220050 473044 220056
rect 472072 219632 472124 219638
rect 472072 219574 472124 219580
rect 471244 218612 471296 218618
rect 471244 218554 471296 218560
rect 470600 218068 470652 218074
rect 470600 218010 470652 218016
rect 467944 217110 468018 217138
rect 467990 216988 468018 217110
rect 468818 216988 468846 217246
rect 469312 217252 469364 217258
rect 469600 217246 469674 217274
rect 469312 217194 469364 217200
rect 469646 216988 469674 217246
rect 470462 217252 470514 217258
rect 470462 217194 470514 217200
rect 470474 216988 470502 217194
rect 471256 217138 471284 218554
rect 472084 217274 472112 219574
rect 472900 218068 472952 218074
rect 472900 218010 472952 218016
rect 472084 217246 472158 217274
rect 471256 217110 471330 217138
rect 471302 216988 471330 217110
rect 472130 216988 472158 217246
rect 472912 217138 472940 218010
rect 473740 217274 473768 222838
rect 474016 220658 474044 229842
rect 474476 229094 474504 231662
rect 474476 229066 474780 229094
rect 474752 224262 474780 229066
rect 475028 227798 475056 231662
rect 475396 230382 475424 231676
rect 475384 230376 475436 230382
rect 475384 230318 475436 230324
rect 476040 230042 476068 231676
rect 476684 230178 476712 231676
rect 476672 230172 476724 230178
rect 476672 230114 476724 230120
rect 475384 230036 475436 230042
rect 475384 229978 475436 229984
rect 476028 230036 476080 230042
rect 476028 229978 476080 229984
rect 475016 227792 475068 227798
rect 475016 227734 475068 227740
rect 474740 224256 474792 224262
rect 474740 224198 474792 224204
rect 475396 220794 475424 229978
rect 476764 229764 476816 229770
rect 476764 229706 476816 229712
rect 476580 225616 476632 225622
rect 476580 225558 476632 225564
rect 475568 223576 475620 223582
rect 475568 223518 475620 223524
rect 475384 220788 475436 220794
rect 475384 220730 475436 220736
rect 474004 220652 474056 220658
rect 474004 220594 474056 220600
rect 475384 220652 475436 220658
rect 475384 220594 475436 220600
rect 474556 220244 474608 220250
rect 474556 220186 474608 220192
rect 474568 217274 474596 220186
rect 475396 217274 475424 220594
rect 475580 218618 475608 223518
rect 476212 220788 476264 220794
rect 476212 220730 476264 220736
rect 475568 218612 475620 218618
rect 475568 218554 475620 218560
rect 476224 217274 476252 220730
rect 476592 217274 476620 225558
rect 476776 220794 476804 229706
rect 477328 225622 477356 231676
rect 477986 231662 478552 231690
rect 478630 231662 478828 231690
rect 478328 230376 478380 230382
rect 478328 230318 478380 230324
rect 477316 225616 477368 225622
rect 477316 225558 477368 225564
rect 478340 222902 478368 230318
rect 478328 222896 478380 222902
rect 478328 222838 478380 222844
rect 477868 222148 477920 222154
rect 477868 222090 477920 222096
rect 476764 220788 476816 220794
rect 476764 220730 476816 220736
rect 477880 217274 477908 222090
rect 478524 220250 478552 231662
rect 478800 228682 478828 231662
rect 479260 229770 479288 231676
rect 479708 230172 479760 230178
rect 479708 230114 479760 230120
rect 479524 230036 479576 230042
rect 479524 229978 479576 229984
rect 479248 229764 479300 229770
rect 479248 229706 479300 229712
rect 478788 228676 478840 228682
rect 478788 228618 478840 228624
rect 479340 227928 479392 227934
rect 479340 227870 479392 227876
rect 478696 220788 478748 220794
rect 478696 220730 478748 220736
rect 478512 220244 478564 220250
rect 478512 220186 478564 220192
rect 478708 217274 478736 220730
rect 479352 219434 479380 227870
rect 479536 224534 479564 229978
rect 479720 228274 479748 230114
rect 479904 229294 479932 231676
rect 480548 230382 480576 231676
rect 480536 230376 480588 230382
rect 480536 230318 480588 230324
rect 479892 229288 479944 229294
rect 479892 229230 479944 229236
rect 479708 228268 479760 228274
rect 479708 228210 479760 228216
rect 481192 227186 481220 231676
rect 481548 230376 481600 230382
rect 481548 230318 481600 230324
rect 481180 227180 481232 227186
rect 481180 227122 481232 227128
rect 481180 227044 481232 227050
rect 481180 226986 481232 226992
rect 479524 224528 479576 224534
rect 479524 224470 479576 224476
rect 479708 224392 479760 224398
rect 479708 224334 479760 224340
rect 479352 219406 479564 219434
rect 479536 217274 479564 219406
rect 479720 219298 479748 224334
rect 479708 219292 479760 219298
rect 479708 219234 479760 219240
rect 480352 219292 480404 219298
rect 480352 219234 480404 219240
rect 473740 217246 473814 217274
rect 474568 217246 474642 217274
rect 475396 217246 475470 217274
rect 476224 217246 476298 217274
rect 476592 217246 477126 217274
rect 477880 217246 477954 217274
rect 478708 217246 478782 217274
rect 479536 217246 479610 217274
rect 472912 217110 472986 217138
rect 472958 216988 472986 217110
rect 473786 216988 473814 217246
rect 474614 216988 474642 217246
rect 475442 216988 475470 217246
rect 476270 216988 476298 217246
rect 477098 216988 477126 217246
rect 477926 216988 477954 217246
rect 478754 216988 478782 217246
rect 479582 216988 479610 217246
rect 480364 217138 480392 219234
rect 481192 217274 481220 226986
rect 481560 220386 481588 230318
rect 481836 229906 481864 231676
rect 481824 229900 481876 229906
rect 481824 229842 481876 229848
rect 482284 229288 482336 229294
rect 482284 229230 482336 229236
rect 482296 220522 482324 229230
rect 482480 228546 482508 231676
rect 483124 230042 483152 231676
rect 483112 230036 483164 230042
rect 483112 229978 483164 229984
rect 483768 229294 483796 231676
rect 484426 231662 484808 231690
rect 484780 230042 484808 231662
rect 484308 230036 484360 230042
rect 484308 229978 484360 229984
rect 484768 230036 484820 230042
rect 484768 229978 484820 229984
rect 484124 229764 484176 229770
rect 484124 229706 484176 229712
rect 483756 229288 483808 229294
rect 483756 229230 483808 229236
rect 484136 228682 484164 229706
rect 483572 228676 483624 228682
rect 483572 228618 483624 228624
rect 484124 228676 484176 228682
rect 484124 228618 484176 228624
rect 482468 228540 482520 228546
rect 482468 228482 482520 228488
rect 482928 227792 482980 227798
rect 482928 227734 482980 227740
rect 482940 222222 482968 227734
rect 482928 222216 482980 222222
rect 482928 222158 482980 222164
rect 482284 220516 482336 220522
rect 482284 220458 482336 220464
rect 481548 220380 481600 220386
rect 481548 220322 481600 220328
rect 482008 220108 482060 220114
rect 482008 220050 482060 220056
rect 482020 217274 482048 220050
rect 482940 218754 482968 222158
rect 483584 219162 483612 228618
rect 484320 221610 484348 229978
rect 485056 227322 485084 231676
rect 485044 227316 485096 227322
rect 485044 227258 485096 227264
rect 485700 224262 485728 231676
rect 486344 229770 486372 231676
rect 486332 229764 486384 229770
rect 486332 229706 486384 229712
rect 486792 229288 486844 229294
rect 486792 229230 486844 229236
rect 486608 224528 486660 224534
rect 486608 224470 486660 224476
rect 484584 224256 484636 224262
rect 484584 224198 484636 224204
rect 485688 224256 485740 224262
rect 485688 224198 485740 224204
rect 484308 221604 484360 221610
rect 484308 221546 484360 221552
rect 483756 221468 483808 221474
rect 483756 221410 483808 221416
rect 483572 219156 483624 219162
rect 483572 219098 483624 219104
rect 482928 218748 482980 218754
rect 482928 218690 482980 218696
rect 482836 218612 482888 218618
rect 482836 218554 482888 218560
rect 481192 217246 481266 217274
rect 482020 217246 482094 217274
rect 480364 217110 480438 217138
rect 480410 216988 480438 217110
rect 481238 216988 481266 217246
rect 482066 216988 482094 217246
rect 482848 217138 482876 218554
rect 483768 217274 483796 221410
rect 484596 219473 484624 224198
rect 486148 222896 486200 222902
rect 486148 222838 486200 222844
rect 484582 219464 484638 219473
rect 484582 219399 484638 219408
rect 484596 217274 484624 219399
rect 485320 218748 485372 218754
rect 485320 218690 485372 218696
rect 483722 217246 483796 217274
rect 484550 217246 484624 217274
rect 485332 217274 485360 218690
rect 485332 217246 485406 217274
rect 482848 217110 482922 217138
rect 482894 216988 482922 217110
rect 483722 216988 483750 217246
rect 484550 216988 484578 217246
rect 485378 216988 485406 217246
rect 486160 217138 486188 222838
rect 486620 220969 486648 224470
rect 486804 224398 486832 229230
rect 486792 224392 486844 224398
rect 486792 224334 486844 224340
rect 486988 222902 487016 231676
rect 487632 228410 487660 231676
rect 487620 228404 487672 228410
rect 487620 228346 487672 228352
rect 487804 228268 487856 228274
rect 487804 228210 487856 228216
rect 486976 222896 487028 222902
rect 486976 222838 487028 222844
rect 486606 220960 486662 220969
rect 486606 220895 486662 220904
rect 486620 217274 486648 220895
rect 487816 218113 487844 228210
rect 488276 220114 488304 231676
rect 488920 225894 488948 231676
rect 488908 225888 488960 225894
rect 488908 225830 488960 225836
rect 489184 225616 489236 225622
rect 489184 225558 489236 225564
rect 488264 220108 488316 220114
rect 488264 220050 488316 220056
rect 489196 219434 489224 225558
rect 489564 223310 489592 231676
rect 489920 229900 489972 229906
rect 489920 229842 489972 229848
rect 489932 225010 489960 229842
rect 489920 225004 489972 225010
rect 489920 224946 489972 224952
rect 489552 223304 489604 223310
rect 489552 223246 489604 223252
rect 490208 223174 490236 231676
rect 490852 230110 490880 231676
rect 490840 230104 490892 230110
rect 490840 230046 490892 230052
rect 490656 230036 490708 230042
rect 490656 229978 490708 229984
rect 490668 229634 490696 229978
rect 490656 229628 490708 229634
rect 490656 229570 490708 229576
rect 490564 228676 490616 228682
rect 490564 228618 490616 228624
rect 490196 223168 490248 223174
rect 490196 223110 490248 223116
rect 489460 220244 489512 220250
rect 489460 220186 489512 220192
rect 488724 219428 488776 219434
rect 488724 219370 488776 219376
rect 489184 219428 489236 219434
rect 489184 219370 489236 219376
rect 487802 218104 487858 218113
rect 488736 218074 488764 219370
rect 487802 218039 487858 218048
rect 488724 218068 488776 218074
rect 487816 217274 487844 218039
rect 488724 218010 488776 218016
rect 486620 217246 487062 217274
rect 487816 217246 487890 217274
rect 486160 217110 486234 217138
rect 486206 216988 486234 217110
rect 487034 216988 487062 217246
rect 487862 216988 487890 217246
rect 488736 217138 488764 218010
rect 489472 217274 489500 220186
rect 490576 219201 490604 228618
rect 491496 225758 491524 231676
rect 492154 231662 492352 231690
rect 491484 225752 491536 225758
rect 491484 225694 491536 225700
rect 491944 220516 491996 220522
rect 491944 220458 491996 220464
rect 490562 219192 490618 219201
rect 490288 219156 490340 219162
rect 490562 219127 490618 219136
rect 491114 219192 491170 219201
rect 491114 219127 491170 219136
rect 490288 219098 490340 219104
rect 490300 218929 490328 219098
rect 490286 218920 490342 218929
rect 490286 218855 490342 218864
rect 489472 217246 489546 217274
rect 488690 217110 488764 217138
rect 488690 216988 488718 217110
rect 489518 216988 489546 217246
rect 490300 217138 490328 218855
rect 491128 218657 491156 219127
rect 491114 218648 491170 218657
rect 491114 218583 491170 218592
rect 491128 217138 491156 218583
rect 491956 217274 491984 220458
rect 492324 220250 492352 231662
rect 492784 230382 492812 231676
rect 492772 230376 492824 230382
rect 492772 230318 492824 230324
rect 493428 230246 493456 231676
rect 494086 231662 494376 231690
rect 493968 230376 494020 230382
rect 493968 230318 494020 230324
rect 493416 230240 493468 230246
rect 493416 230182 493468 230188
rect 493784 230104 493836 230110
rect 493784 230046 493836 230052
rect 493796 228818 493824 230046
rect 493784 228812 493836 228818
rect 493784 228754 493836 228760
rect 492956 227180 493008 227186
rect 492956 227122 493008 227128
rect 492772 220380 492824 220386
rect 492772 220322 492824 220328
rect 492312 220244 492364 220250
rect 492312 220186 492364 220192
rect 491956 217246 492168 217274
rect 490300 217110 490374 217138
rect 491128 217110 491202 217138
rect 490346 216988 490374 217110
rect 491174 216988 491202 217110
rect 492002 216988 492030 217246
rect 492140 217161 492168 217246
rect 492126 217152 492182 217161
rect 492784 217138 492812 220322
rect 492968 219201 492996 227122
rect 493980 220522 494008 230318
rect 494348 230110 494376 231662
rect 494716 230382 494744 231676
rect 494704 230376 494756 230382
rect 494704 230318 494756 230324
rect 495164 230240 495216 230246
rect 495164 230182 495216 230188
rect 494336 230104 494388 230110
rect 494336 230046 494388 230052
rect 494612 228540 494664 228546
rect 494612 228482 494664 228488
rect 493968 220516 494020 220522
rect 493968 220458 494020 220464
rect 492954 219192 493010 219201
rect 492954 219127 493010 219136
rect 493598 219192 493654 219201
rect 493598 219127 493654 219136
rect 493612 217297 493640 219127
rect 494624 218210 494652 228482
rect 495176 225622 495204 230182
rect 495360 228682 495388 231676
rect 496004 229906 496032 231676
rect 496188 231662 496662 231690
rect 495992 229900 496044 229906
rect 495992 229842 496044 229848
rect 495348 228676 495400 228682
rect 495348 228618 495400 228624
rect 495164 225616 495216 225622
rect 495164 225558 495216 225564
rect 494796 225004 494848 225010
rect 494796 224946 494848 224952
rect 494808 219745 494836 224946
rect 496188 221882 496216 231662
rect 496360 230376 496412 230382
rect 496360 230318 496412 230324
rect 496176 221876 496228 221882
rect 496176 221818 496228 221824
rect 496084 221604 496136 221610
rect 496084 221546 496136 221552
rect 494794 219736 494850 219745
rect 494794 219671 494850 219680
rect 494612 218204 494664 218210
rect 494612 218146 494664 218152
rect 493598 217288 493654 217297
rect 494808 217274 494836 219671
rect 495256 218204 495308 218210
rect 495256 218146 495308 218152
rect 493598 217223 493654 217232
rect 494486 217246 494836 217274
rect 493612 217138 493640 217223
rect 492784 217110 492858 217138
rect 493612 217110 493686 217138
rect 492126 217087 492182 217096
rect 492830 216988 492858 217110
rect 493658 216988 493686 217110
rect 494486 216988 494514 217246
rect 495268 217138 495296 218146
rect 496096 217138 496124 221546
rect 496372 220386 496400 230318
rect 497292 227050 497320 231676
rect 497936 230314 497964 231676
rect 497924 230308 497976 230314
rect 497924 230250 497976 230256
rect 497464 229628 497516 229634
rect 497464 229570 497516 229576
rect 497280 227044 497332 227050
rect 497280 226986 497332 226992
rect 497476 224954 497504 229570
rect 498580 227186 498608 231676
rect 498752 227316 498804 227322
rect 498752 227258 498804 227264
rect 498568 227180 498620 227186
rect 498568 227122 498620 227128
rect 498764 224954 498792 227258
rect 497476 224926 497780 224954
rect 496912 224392 496964 224398
rect 496912 224334 496964 224340
rect 496360 220380 496412 220386
rect 496360 220322 496412 220328
rect 496924 218385 496952 224334
rect 497752 219201 497780 224926
rect 498672 224926 498792 224954
rect 497738 219192 497794 219201
rect 497738 219127 497794 219136
rect 496910 218376 496966 218385
rect 496910 218311 496966 218320
rect 496924 217138 496952 218311
rect 497556 218068 497608 218074
rect 497556 218010 497608 218016
rect 497568 217297 497596 218010
rect 497554 217288 497610 217297
rect 497752 217274 497780 219127
rect 498672 217569 498700 224926
rect 499224 224398 499252 231676
rect 499868 230382 499896 231676
rect 500052 231662 500526 231690
rect 501170 231662 501552 231690
rect 499856 230376 499908 230382
rect 499856 230318 499908 230324
rect 499672 230308 499724 230314
rect 499672 230250 499724 230256
rect 499684 230042 499712 230250
rect 499672 230036 499724 230042
rect 499672 229978 499724 229984
rect 499212 224392 499264 224398
rect 499212 224334 499264 224340
rect 499396 224256 499448 224262
rect 499396 224198 499448 224204
rect 498658 217560 498714 217569
rect 498658 217495 498714 217504
rect 498672 217274 498700 217495
rect 497752 217246 497826 217274
rect 497554 217223 497610 217232
rect 495268 217110 495342 217138
rect 496096 217110 496170 217138
rect 496924 217110 496998 217138
rect 495314 216988 495342 217110
rect 496142 216988 496170 217110
rect 496970 216988 496998 217110
rect 497798 216988 497826 217246
rect 498626 217246 498700 217274
rect 498626 216988 498654 217246
rect 499408 217138 499436 224198
rect 500052 221746 500080 231662
rect 501144 230376 501196 230382
rect 501144 230318 501196 230324
rect 500224 229764 500276 229770
rect 500224 229706 500276 229712
rect 500040 221740 500092 221746
rect 500040 221682 500092 221688
rect 500236 218385 500264 229706
rect 501156 227322 501184 230318
rect 501524 229094 501552 231662
rect 501800 229294 501828 231676
rect 501788 229288 501840 229294
rect 501788 229230 501840 229236
rect 501524 229066 501736 229094
rect 501512 228404 501564 228410
rect 501512 228346 501564 228352
rect 501144 227316 501196 227322
rect 501144 227258 501196 227264
rect 501524 224954 501552 228346
rect 501708 224954 501736 229066
rect 502444 228546 502472 231676
rect 503102 231662 503484 231690
rect 503260 230172 503312 230178
rect 503260 230114 503312 230120
rect 502432 228540 502484 228546
rect 502432 228482 502484 228488
rect 503272 226302 503300 230114
rect 503260 226296 503312 226302
rect 503260 226238 503312 226244
rect 502984 225888 503036 225894
rect 502984 225830 503036 225836
rect 501524 224926 501644 224954
rect 501708 224926 501828 224954
rect 501052 222896 501104 222902
rect 501052 222838 501104 222844
rect 501064 218482 501092 222838
rect 501052 218476 501104 218482
rect 501052 218418 501104 218424
rect 500038 218376 500094 218385
rect 500038 218311 500040 218320
rect 500092 218311 500094 218320
rect 500222 218376 500278 218385
rect 500222 218311 500278 218320
rect 500040 218282 500092 218288
rect 500236 217274 500264 218311
rect 500236 217246 500310 217274
rect 499408 217110 499482 217138
rect 499454 216988 499482 217110
rect 500282 216988 500310 217246
rect 501064 217138 501092 218418
rect 501616 217274 501644 224926
rect 501800 223038 501828 224926
rect 501788 223032 501840 223038
rect 501788 222974 501840 222980
rect 502708 220108 502760 220114
rect 502708 220050 502760 220056
rect 502720 219201 502748 220050
rect 502522 219192 502578 219201
rect 502522 219127 502578 219136
rect 502706 219192 502762 219201
rect 502996 219162 503024 225830
rect 503456 221610 503484 231662
rect 503732 230382 503760 231676
rect 504390 231662 504680 231690
rect 503720 230376 503772 230382
rect 503720 230318 503772 230324
rect 504364 230036 504416 230042
rect 504364 229978 504416 229984
rect 504376 229094 504404 229978
rect 504192 229066 504404 229094
rect 503444 221604 503496 221610
rect 503444 221546 503496 221552
rect 504192 220794 504220 229066
rect 504364 223304 504416 223310
rect 504364 223246 504416 223252
rect 504180 220788 504232 220794
rect 504180 220730 504232 220736
rect 502706 219127 502762 219136
rect 502984 219156 503036 219162
rect 502536 219026 502564 219127
rect 502524 219020 502576 219026
rect 502524 218962 502576 218968
rect 501616 217246 501966 217274
rect 501064 217110 501138 217138
rect 501110 216988 501138 217110
rect 501938 216988 501966 217246
rect 502720 217138 502748 219127
rect 502984 219098 503036 219104
rect 503536 219156 503588 219162
rect 503536 219098 503588 219104
rect 503548 217569 503576 219098
rect 503534 217560 503590 217569
rect 503534 217495 503590 217504
rect 503548 217138 503576 217495
rect 504376 217138 504404 223246
rect 504652 222902 504680 231662
rect 505020 229094 505048 231676
rect 505664 229770 505692 231676
rect 505652 229764 505704 229770
rect 505652 229706 505704 229712
rect 505020 229066 505140 229094
rect 505112 223310 505140 229066
rect 506020 228812 506072 228818
rect 506020 228754 506072 228760
rect 505100 223304 505152 223310
rect 505100 223246 505152 223252
rect 505652 223168 505704 223174
rect 505652 223110 505704 223116
rect 504640 222896 504692 222902
rect 504640 222838 504692 222844
rect 504640 219360 504692 219366
rect 504640 219302 504692 219308
rect 505284 219360 505336 219366
rect 505284 219302 505336 219308
rect 504652 218385 504680 219302
rect 505296 219201 505324 219302
rect 505098 219192 505154 219201
rect 505098 219127 505154 219136
rect 505282 219192 505338 219201
rect 505282 219127 505338 219136
rect 505112 219042 505140 219127
rect 505112 219014 505324 219042
rect 505296 218691 505324 219014
rect 505282 218682 505338 218691
rect 504822 218648 504878 218657
rect 505282 218617 505338 218626
rect 504822 218583 504878 218592
rect 504638 218376 504694 218385
rect 504638 218311 504694 218320
rect 504836 217841 504864 218583
rect 505664 218074 505692 223110
rect 505284 218068 505336 218074
rect 505284 218010 505336 218016
rect 505652 218068 505704 218074
rect 505652 218010 505704 218016
rect 504822 217832 504878 217841
rect 504822 217767 504878 217776
rect 505296 217138 505324 218010
rect 505468 217864 505520 217870
rect 505466 217832 505468 217841
rect 505520 217832 505522 217841
rect 505466 217767 505522 217776
rect 506032 217569 506060 228754
rect 506308 228410 506336 231676
rect 506966 231662 507348 231690
rect 506940 230376 506992 230382
rect 506940 230318 506992 230324
rect 506952 228834 506980 230318
rect 507124 229288 507176 229294
rect 507124 229230 507176 229236
rect 507136 228954 507164 229230
rect 507124 228948 507176 228954
rect 507124 228890 507176 228896
rect 506952 228806 507072 228834
rect 506296 228404 506348 228410
rect 506296 228346 506348 228352
rect 506848 225752 506900 225758
rect 506848 225694 506900 225700
rect 506018 217560 506074 217569
rect 506018 217495 506074 217504
rect 506032 217274 506060 217495
rect 506860 217274 506888 225694
rect 507044 220114 507072 228806
rect 507320 225758 507348 231662
rect 507596 229158 507624 231676
rect 507584 229152 507636 229158
rect 507584 229094 507636 229100
rect 507308 225752 507360 225758
rect 507308 225694 507360 225700
rect 508240 224534 508268 231676
rect 508228 224528 508280 224534
rect 508228 224470 508280 224476
rect 508884 224262 508912 231676
rect 509240 229900 509292 229906
rect 509240 229842 509292 229848
rect 509252 225010 509280 229842
rect 509528 229634 509556 231676
rect 509516 229628 509568 229634
rect 509516 229570 509568 229576
rect 510172 229094 510200 231676
rect 510172 229066 510384 229094
rect 510160 226296 510212 226302
rect 510160 226238 510212 226244
rect 509700 225616 509752 225622
rect 509700 225558 509752 225564
rect 509240 225004 509292 225010
rect 509712 224954 509740 225558
rect 509240 224946 509292 224952
rect 509436 224926 509740 224954
rect 508872 224256 508924 224262
rect 508872 224198 508924 224204
rect 508504 220516 508556 220522
rect 508504 220458 508556 220464
rect 507676 220244 507728 220250
rect 507676 220186 507728 220192
rect 507032 220108 507084 220114
rect 507032 220050 507084 220056
rect 507124 219224 507176 219230
rect 507124 219166 507176 219172
rect 507136 218346 507164 219166
rect 507308 219020 507360 219026
rect 507308 218962 507360 218968
rect 507320 218385 507348 218962
rect 507306 218376 507362 218385
rect 507124 218340 507176 218346
rect 507688 218346 507716 220186
rect 507306 218311 507362 218320
rect 507676 218340 507728 218346
rect 507124 218282 507176 218288
rect 507676 218282 507728 218288
rect 506032 217246 506106 217274
rect 506860 217246 506934 217274
rect 502720 217110 502794 217138
rect 503548 217110 503622 217138
rect 504376 217110 504450 217138
rect 502766 216988 502794 217110
rect 503594 216988 503622 217110
rect 504422 216988 504450 217110
rect 505250 217110 505324 217138
rect 505250 216988 505278 217110
rect 506078 216988 506106 217246
rect 506906 216988 506934 217246
rect 507688 217138 507716 218282
rect 508516 217841 508544 220458
rect 508502 217832 508558 217841
rect 508502 217767 508558 217776
rect 508516 217138 508544 217767
rect 509436 217274 509464 224926
rect 510172 218890 510200 226238
rect 510356 225622 510384 229066
rect 510816 226166 510844 231676
rect 511460 229974 511488 231676
rect 511448 229968 511500 229974
rect 511448 229910 511500 229916
rect 511264 229152 511316 229158
rect 511264 229094 511316 229100
rect 510804 226160 510856 226166
rect 510804 226102 510856 226108
rect 510344 225616 510396 225622
rect 510344 225558 510396 225564
rect 511276 220658 511304 229094
rect 512104 228682 512132 231676
rect 512762 231662 513144 231690
rect 511816 228676 511868 228682
rect 511816 228618 511868 228624
rect 512092 228676 512144 228682
rect 512092 228618 512144 228624
rect 511264 220652 511316 220658
rect 511264 220594 511316 220600
rect 510988 220380 511040 220386
rect 510988 220322 511040 220328
rect 511000 220017 511028 220322
rect 510986 220008 511042 220017
rect 510986 219943 511042 219952
rect 510160 218884 510212 218890
rect 510160 218826 510212 218832
rect 509390 217246 509464 217274
rect 510172 217274 510200 218826
rect 510172 217246 510246 217274
rect 507688 217110 507762 217138
rect 508516 217110 508590 217138
rect 507734 216988 507762 217110
rect 508562 216988 508590 217110
rect 509390 216988 509418 217246
rect 510218 216988 510246 217246
rect 511000 217138 511028 219943
rect 511828 217274 511856 228618
rect 512644 225004 512696 225010
rect 512644 224946 512696 224952
rect 512656 220017 512684 224946
rect 513116 223174 513144 231662
rect 513392 230246 513420 231676
rect 513380 230240 513432 230246
rect 513380 230182 513432 230188
rect 514036 227050 514064 231676
rect 514024 227044 514076 227050
rect 514024 226986 514076 226992
rect 514300 226908 514352 226914
rect 514300 226850 514352 226856
rect 513104 223168 513156 223174
rect 513104 223110 513156 223116
rect 513378 221912 513434 221921
rect 513378 221847 513380 221856
rect 513432 221847 513434 221856
rect 513380 221818 513432 221824
rect 512642 220008 512698 220017
rect 512642 219943 512698 219952
rect 512656 217274 512684 219943
rect 513392 217274 513420 221818
rect 514312 217274 514340 226850
rect 514680 224670 514708 231676
rect 515338 231662 515720 231690
rect 515404 230240 515456 230246
rect 515404 230182 515456 230188
rect 514668 224664 514720 224670
rect 514668 224606 514720 224612
rect 515416 221882 515444 230182
rect 515692 230110 515720 231662
rect 515876 231662 515982 231690
rect 515680 230104 515732 230110
rect 515680 230046 515732 230052
rect 515876 227594 515904 231662
rect 516612 230382 516640 231676
rect 516600 230376 516652 230382
rect 516600 230318 516652 230324
rect 517256 230246 517284 231676
rect 517428 230376 517480 230382
rect 517428 230318 517480 230324
rect 517244 230240 517296 230246
rect 517244 230182 517296 230188
rect 516784 229968 516836 229974
rect 516784 229910 516836 229916
rect 516048 229764 516100 229770
rect 516048 229706 516100 229712
rect 515864 227588 515916 227594
rect 515864 227530 515916 227536
rect 516060 227186 516088 229706
rect 515864 227180 515916 227186
rect 515864 227122 515916 227128
rect 516048 227180 516100 227186
rect 516048 227122 516100 227128
rect 515876 224954 515904 227122
rect 515876 224926 515996 224954
rect 516796 224942 516824 229910
rect 515404 221876 515456 221882
rect 515404 221818 515456 221824
rect 515968 221241 515996 224926
rect 516784 224936 516836 224942
rect 516784 224878 516836 224884
rect 516784 224392 516836 224398
rect 516784 224334 516836 224340
rect 515954 221232 516010 221241
rect 515954 221167 516010 221176
rect 515772 220788 515824 220794
rect 515772 220730 515824 220736
rect 515784 219570 515812 220730
rect 515220 219564 515272 219570
rect 515220 219506 515272 219512
rect 515772 219564 515824 219570
rect 515772 219506 515824 219512
rect 514482 219192 514538 219201
rect 514482 219127 514538 219136
rect 514758 219192 514814 219201
rect 514758 219127 514814 219136
rect 514496 217734 514524 219127
rect 514772 219042 514800 219127
rect 514772 219026 515076 219042
rect 514772 219020 515088 219026
rect 514772 219014 515036 219020
rect 515036 218962 515088 218968
rect 514760 218884 514812 218890
rect 514760 218826 514812 218832
rect 514772 218482 514800 218826
rect 514760 218476 514812 218482
rect 514760 218418 514812 218424
rect 514666 218342 514722 218351
rect 514666 218277 514722 218286
rect 514680 217870 514708 218277
rect 514668 217864 514720 217870
rect 514668 217806 514720 217812
rect 514484 217728 514536 217734
rect 514484 217670 514536 217676
rect 511828 217246 511902 217274
rect 512656 217246 512730 217274
rect 513392 217246 513558 217274
rect 514312 217246 514386 217274
rect 511000 217110 511074 217138
rect 511046 216988 511074 217110
rect 511874 216988 511902 217246
rect 512702 216988 512730 217246
rect 513530 216988 513558 217246
rect 514358 216988 514386 217246
rect 515232 217138 515260 219506
rect 515968 217274 515996 221167
rect 516600 219360 516652 219366
rect 516600 219302 516652 219308
rect 516612 219201 516640 219302
rect 516598 219192 516654 219201
rect 516598 219127 516654 219136
rect 515968 217246 516042 217274
rect 515186 217110 515260 217138
rect 515186 216988 515214 217110
rect 516014 216988 516042 217246
rect 516796 217138 516824 224334
rect 517440 220386 517468 230318
rect 517900 229090 517928 231676
rect 517888 229084 517940 229090
rect 517888 229026 517940 229032
rect 517796 227316 517848 227322
rect 517796 227258 517848 227264
rect 517808 221513 517836 227258
rect 518544 226030 518572 231676
rect 519188 230110 519216 231676
rect 519176 230104 519228 230110
rect 519176 230046 519228 230052
rect 518900 229764 518952 229770
rect 518900 229706 518952 229712
rect 518532 226024 518584 226030
rect 518532 225966 518584 225972
rect 518912 223446 518940 229706
rect 519832 228818 519860 231676
rect 520476 230382 520504 231676
rect 520464 230376 520516 230382
rect 520464 230318 520516 230324
rect 521120 229770 521148 231676
rect 521568 230376 521620 230382
rect 521568 230318 521620 230324
rect 521108 229764 521160 229770
rect 521108 229706 521160 229712
rect 520096 228948 520148 228954
rect 520096 228890 520148 228896
rect 519820 228812 519872 228818
rect 519820 228754 519872 228760
rect 518900 223440 518952 223446
rect 518900 223382 518952 223388
rect 519268 223032 519320 223038
rect 519268 222974 519320 222980
rect 518440 221740 518492 221746
rect 518440 221682 518492 221688
rect 517794 221504 517850 221513
rect 517794 221439 517850 221448
rect 517428 220380 517480 220386
rect 517428 220322 517480 220328
rect 517808 217274 517836 221439
rect 518452 220862 518480 221682
rect 518440 220856 518492 220862
rect 518440 220798 518492 220804
rect 517670 217246 517836 217274
rect 516796 217110 516870 217138
rect 516842 216988 516870 217110
rect 517670 216988 517698 217246
rect 518452 217138 518480 220798
rect 518808 219428 518860 219434
rect 518808 219370 518860 219376
rect 518820 218686 518848 219370
rect 518808 218680 518860 218686
rect 518808 218622 518860 218628
rect 519280 217138 519308 222974
rect 519542 220280 519598 220289
rect 519542 220215 519598 220224
rect 519556 219745 519584 220215
rect 519542 219736 519598 219745
rect 519542 219671 519598 219680
rect 519818 219736 519874 219745
rect 520108 219706 520136 228890
rect 520924 228540 520976 228546
rect 520924 228482 520976 228488
rect 519818 219671 519874 219680
rect 520096 219700 520148 219706
rect 519832 219434 519860 219671
rect 520096 219642 520148 219648
rect 519820 219428 519872 219434
rect 519820 219370 519872 219376
rect 519728 218748 519780 218754
rect 519728 218690 519780 218696
rect 519740 218210 519768 218690
rect 520108 218634 520136 219642
rect 520108 218606 520228 218634
rect 519728 218204 519780 218210
rect 519728 218146 519780 218152
rect 519912 218204 519964 218210
rect 519912 218146 519964 218152
rect 519924 217734 519952 218146
rect 519912 217728 519964 217734
rect 519912 217670 519964 217676
rect 520200 217274 520228 218606
rect 520154 217246 520228 217274
rect 520936 217274 520964 228482
rect 521580 220250 521608 230318
rect 521764 227322 521792 231676
rect 522422 231662 522896 231690
rect 522304 230240 522356 230246
rect 522304 230182 522356 230188
rect 521752 227316 521804 227322
rect 521752 227258 521804 227264
rect 521752 221604 521804 221610
rect 521752 221546 521804 221552
rect 521568 220244 521620 220250
rect 521568 220186 521620 220192
rect 520936 217246 521010 217274
rect 518452 217110 518526 217138
rect 519280 217110 519354 217138
rect 518498 216988 518526 217110
rect 519326 216988 519354 217110
rect 520154 216988 520182 217246
rect 520982 217122 521010 217246
rect 521764 217138 521792 221546
rect 522316 220522 522344 230182
rect 522868 221746 522896 231662
rect 523052 230042 523080 231676
rect 523040 230036 523092 230042
rect 523040 229978 523092 229984
rect 523696 223038 523724 231676
rect 524340 227458 524368 231676
rect 524984 229634 525012 231676
rect 525628 230330 525656 231676
rect 525628 230302 525748 230330
rect 525524 229900 525576 229906
rect 525524 229842 525576 229848
rect 524972 229628 525024 229634
rect 524972 229570 525024 229576
rect 525536 227730 525564 229842
rect 525524 227724 525576 227730
rect 525524 227666 525576 227672
rect 524328 227452 524380 227458
rect 524328 227394 524380 227400
rect 525064 227180 525116 227186
rect 525064 227122 525116 227128
rect 523960 223304 524012 223310
rect 523960 223246 524012 223252
rect 523684 223032 523736 223038
rect 523684 222974 523736 222980
rect 523776 222896 523828 222902
rect 523776 222838 523828 222844
rect 522856 221740 522908 221746
rect 522856 221682 522908 221688
rect 522304 220516 522356 220522
rect 522304 220458 522356 220464
rect 522580 220108 522632 220114
rect 522580 220050 522632 220056
rect 522592 219745 522620 220050
rect 522578 219736 522634 219745
rect 522578 219671 522634 219680
rect 522592 217138 522620 219671
rect 523788 217598 523816 222838
rect 523776 217592 523828 217598
rect 523776 217534 523828 217540
rect 523788 217274 523816 217534
rect 523466 217246 523816 217274
rect 523972 217274 524000 223246
rect 524418 219192 524474 219201
rect 524418 219127 524420 219136
rect 524472 219127 524474 219136
rect 524602 219192 524658 219201
rect 524602 219127 524658 219136
rect 524420 219098 524472 219104
rect 524616 218890 524644 219127
rect 525076 218890 525104 227122
rect 525720 224398 525748 230302
rect 526272 228954 526300 231676
rect 526916 230382 526944 231676
rect 526904 230376 526956 230382
rect 526904 230318 526956 230324
rect 526260 228948 526312 228954
rect 526260 228890 526312 228896
rect 525892 228404 525944 228410
rect 525892 228346 525944 228352
rect 525708 224392 525760 224398
rect 525708 224334 525760 224340
rect 525904 221610 525932 228346
rect 527560 225758 527588 231676
rect 527824 230376 527876 230382
rect 527824 230318 527876 230324
rect 526720 225752 526772 225758
rect 526720 225694 526772 225700
rect 527548 225752 527600 225758
rect 527548 225694 527600 225700
rect 525892 221604 525944 221610
rect 525892 221546 525944 221552
rect 524144 218884 524196 218890
rect 524144 218826 524196 218832
rect 524604 218884 524656 218890
rect 524604 218826 524656 218832
rect 525064 218884 525116 218890
rect 525064 218826 525116 218832
rect 524156 218385 524184 218826
rect 524142 218376 524198 218385
rect 524142 218311 524198 218320
rect 524602 218376 524658 218385
rect 524602 218311 524658 218320
rect 524616 218210 524644 218311
rect 524604 218204 524656 218210
rect 524604 218146 524656 218152
rect 524418 217832 524474 217841
rect 524418 217767 524474 217776
rect 524602 217832 524658 217841
rect 524602 217767 524658 217776
rect 524432 217462 524460 217767
rect 524616 217598 524644 217767
rect 524604 217592 524656 217598
rect 524604 217534 524656 217540
rect 524420 217456 524472 217462
rect 524420 217398 524472 217404
rect 525076 217274 525104 218826
rect 525904 217274 525932 221546
rect 526732 217274 526760 225694
rect 527548 220652 527600 220658
rect 527548 220594 527600 220600
rect 527560 218210 527588 220594
rect 527836 220114 527864 230318
rect 528204 225894 528232 231676
rect 528862 231662 529244 231690
rect 529506 231662 529796 231690
rect 529216 230314 529244 231662
rect 529204 230308 529256 230314
rect 529204 230250 529256 230256
rect 529020 230240 529072 230246
rect 529020 230182 529072 230188
rect 528192 225888 528244 225894
rect 528192 225830 528244 225836
rect 528376 224528 528428 224534
rect 528376 224470 528428 224476
rect 527824 220108 527876 220114
rect 527824 220050 527876 220056
rect 527548 218204 527600 218210
rect 527548 218146 527600 218152
rect 523972 217246 524322 217274
rect 525076 217246 525150 217274
rect 525904 217246 525978 217274
rect 526732 217246 526806 217274
rect 520970 217116 521022 217122
rect 521764 217110 521838 217138
rect 522592 217110 522666 217138
rect 520970 217058 521022 217064
rect 520982 216988 521010 217058
rect 521810 216988 521838 217110
rect 522638 216988 522666 217110
rect 523466 216988 523494 217246
rect 524294 216988 524322 217246
rect 525122 216988 525150 217246
rect 525950 216988 525978 217246
rect 526778 216988 526806 217246
rect 527560 217138 527588 218146
rect 528388 217870 528416 224470
rect 529032 223310 529060 230182
rect 529388 224256 529440 224262
rect 529388 224198 529440 224204
rect 529020 223304 529072 223310
rect 529020 223246 529072 223252
rect 529204 218612 529256 218618
rect 529204 218554 529256 218560
rect 529216 218346 529244 218554
rect 529204 218340 529256 218346
rect 529204 218282 529256 218288
rect 528376 217864 528428 217870
rect 528376 217806 528428 217812
rect 528388 217138 528416 217806
rect 529400 217274 529428 224198
rect 529768 222018 529796 231662
rect 529940 229764 529992 229770
rect 529940 229706 529992 229712
rect 529952 226302 529980 229706
rect 529940 226296 529992 226302
rect 529940 226238 529992 226244
rect 530136 224534 530164 231676
rect 530780 230178 530808 231676
rect 530768 230172 530820 230178
rect 530768 230114 530820 230120
rect 531424 228546 531452 231676
rect 531412 228540 531464 228546
rect 531412 228482 531464 228488
rect 531688 226160 531740 226166
rect 531688 226102 531740 226108
rect 530492 225616 530544 225622
rect 530492 225558 530544 225564
rect 530124 224528 530176 224534
rect 530124 224470 530176 224476
rect 530032 223440 530084 223446
rect 530032 223382 530084 223388
rect 529756 222012 529808 222018
rect 529756 221954 529808 221960
rect 530044 220017 530072 223382
rect 530030 220008 530086 220017
rect 530030 219943 530086 219952
rect 530306 220008 530362 220017
rect 530306 219943 530362 219952
rect 529572 218884 529624 218890
rect 529572 218826 529624 218832
rect 529584 218346 529612 218826
rect 529572 218340 529624 218346
rect 529572 218282 529624 218288
rect 529262 217246 529428 217274
rect 527560 217110 527634 217138
rect 528388 217110 528462 217138
rect 527606 216988 527634 217110
rect 528434 216988 528462 217110
rect 529262 216988 529290 217246
rect 530044 217138 530072 219943
rect 530320 218754 530348 219943
rect 530308 218748 530360 218754
rect 530308 218690 530360 218696
rect 530504 217258 530532 225558
rect 531320 224936 531372 224942
rect 531320 224878 531372 224884
rect 531332 219774 531360 224878
rect 531320 219768 531372 219774
rect 531320 219710 531372 219716
rect 531700 217274 531728 226102
rect 532068 225622 532096 231676
rect 532712 229770 532740 231676
rect 533370 231662 533752 231690
rect 532700 229764 532752 229770
rect 532700 229706 532752 229712
rect 532424 229628 532476 229634
rect 532424 229570 532476 229576
rect 532056 225616 532108 225622
rect 532056 225558 532108 225564
rect 532436 224806 532464 229570
rect 533528 228676 533580 228682
rect 533528 228618 533580 228624
rect 533540 224954 533568 228618
rect 533448 224926 533568 224954
rect 532424 224800 532476 224806
rect 532424 224742 532476 224748
rect 532608 219768 532660 219774
rect 532608 219710 532660 219716
rect 530492 217252 530544 217258
rect 530492 217194 530544 217200
rect 530906 217252 530958 217258
rect 531700 217246 531774 217274
rect 530906 217194 530958 217200
rect 530044 217110 530118 217138
rect 530090 216988 530118 217110
rect 530918 216988 530946 217194
rect 531746 216988 531774 217246
rect 532620 217138 532648 219710
rect 533448 217734 533476 224926
rect 533724 222902 533752 231662
rect 534000 228682 534028 231676
rect 534644 230450 534672 231676
rect 534632 230444 534684 230450
rect 534632 230386 534684 230392
rect 534724 230036 534776 230042
rect 534724 229978 534776 229984
rect 533988 228676 534040 228682
rect 533988 228618 534040 228624
rect 534736 223174 534764 229978
rect 535288 224262 535316 231676
rect 535932 227186 535960 231676
rect 536576 230178 536604 231676
rect 536564 230172 536616 230178
rect 536564 230114 536616 230120
rect 535920 227180 535972 227186
rect 535920 227122 535972 227128
rect 537220 227050 537248 231676
rect 537864 228410 537892 231676
rect 538508 229906 538536 231676
rect 538692 231662 539166 231690
rect 538496 229900 538548 229906
rect 538496 229842 538548 229848
rect 537852 228404 537904 228410
rect 537852 228346 537904 228352
rect 537484 227724 537536 227730
rect 537484 227666 537536 227672
rect 535644 227044 535696 227050
rect 535644 226986 535696 226992
rect 537208 227044 537260 227050
rect 537208 226986 537260 226992
rect 535656 224954 535684 226986
rect 535656 224926 535868 224954
rect 535276 224256 535328 224262
rect 535276 224198 535328 224204
rect 534448 223168 534500 223174
rect 534448 223110 534500 223116
rect 534724 223168 534776 223174
rect 534724 223110 534776 223116
rect 533712 222896 533764 222902
rect 533712 222838 533764 222844
rect 534170 219192 534226 219201
rect 533896 219156 533948 219162
rect 534170 219127 534226 219136
rect 533896 219098 533948 219104
rect 533908 218385 533936 219098
rect 534184 219042 534212 219127
rect 534184 219014 534304 219042
rect 534276 218890 534304 219014
rect 534264 218884 534316 218890
rect 534264 218826 534316 218832
rect 534080 218748 534132 218754
rect 534080 218690 534132 218696
rect 533710 218376 533766 218385
rect 533710 218311 533766 218320
rect 533894 218376 533950 218385
rect 533894 218311 533950 218320
rect 533436 217728 533488 217734
rect 533436 217670 533488 217676
rect 533448 217274 533476 217670
rect 533724 217598 533752 218311
rect 534092 218113 534120 218690
rect 534078 218104 534134 218113
rect 534078 218039 534134 218048
rect 534262 218104 534318 218113
rect 534262 218039 534318 218048
rect 534276 217598 534304 218039
rect 533712 217592 533764 217598
rect 533712 217534 533764 217540
rect 534264 217592 534316 217598
rect 534264 217534 534316 217540
rect 534460 217274 534488 223110
rect 535000 221876 535052 221882
rect 535000 221818 535052 221824
rect 535012 219366 535040 221818
rect 535000 219360 535052 219366
rect 535000 219302 535052 219308
rect 534630 219192 534686 219201
rect 534630 219127 534686 219136
rect 534644 218754 534672 219127
rect 534632 218748 534684 218754
rect 534632 218690 534684 218696
rect 532574 217110 532648 217138
rect 533402 217246 533476 217274
rect 534230 217246 534488 217274
rect 532574 216988 532602 217110
rect 533402 216988 533430 217246
rect 534230 216988 534258 217246
rect 535012 217138 535040 219302
rect 535840 217274 535868 224926
rect 536656 224664 536708 224670
rect 536656 224606 536708 224612
rect 535840 217246 535914 217274
rect 535886 217190 535914 217246
rect 535874 217184 535926 217190
rect 535012 217110 535086 217138
rect 535874 217126 535926 217132
rect 536668 217138 536696 224606
rect 537496 218754 537524 227666
rect 538692 221474 538720 231662
rect 544200 230444 544252 230450
rect 544200 230386 544252 230392
rect 541624 230308 541676 230314
rect 541624 230250 541676 230256
rect 540520 229084 540572 229090
rect 540520 229026 540572 229032
rect 538956 227588 539008 227594
rect 538956 227530 539008 227536
rect 538968 224954 538996 227530
rect 538876 224926 538996 224954
rect 540532 224954 540560 229026
rect 541440 226024 541492 226030
rect 541440 225966 541492 225972
rect 540532 224926 540836 224954
rect 538680 221468 538732 221474
rect 538680 221410 538732 221416
rect 538876 219314 538904 224926
rect 540060 220516 540112 220522
rect 540060 220458 540112 220464
rect 539140 220380 539192 220386
rect 539140 220322 539192 220328
rect 538416 219286 538904 219314
rect 537484 218748 537536 218754
rect 537484 218690 537536 218696
rect 537496 217274 537524 218690
rect 538416 217598 538444 219286
rect 538864 219156 538916 219162
rect 538864 219098 538916 219104
rect 538876 218482 538904 219098
rect 538864 218476 538916 218482
rect 538864 218418 538916 218424
rect 538404 217592 538456 217598
rect 538404 217534 538456 217540
rect 538416 217274 538444 217534
rect 537496 217246 537570 217274
rect 535058 216988 535086 217110
rect 535886 216988 535914 217126
rect 536668 217110 536742 217138
rect 536714 216988 536742 217110
rect 537542 216988 537570 217246
rect 538370 217246 538444 217274
rect 538370 216988 538398 217246
rect 539152 217138 539180 220322
rect 540072 217138 540100 220458
rect 540808 219910 540836 224926
rect 540796 219904 540848 219910
rect 540796 219846 540848 219852
rect 540808 217274 540836 219846
rect 541452 217274 541480 225966
rect 541636 224954 541664 230250
rect 543188 228812 543240 228818
rect 543188 228754 543240 228760
rect 541636 224926 541756 224954
rect 541728 220386 541756 224926
rect 543200 222194 543228 228754
rect 544212 226030 544240 230386
rect 549260 230172 549312 230178
rect 549260 230114 549312 230120
rect 547144 230036 547196 230042
rect 547144 229978 547196 229984
rect 545120 227316 545172 227322
rect 545120 227258 545172 227264
rect 544936 226296 544988 226302
rect 544936 226238 544988 226244
rect 544200 226024 544252 226030
rect 544200 225966 544252 225972
rect 543648 223304 543700 223310
rect 543648 223246 543700 223252
rect 543200 222166 543320 222194
rect 543292 221474 543320 222166
rect 543280 221468 543332 221474
rect 543280 221410 543332 221416
rect 542912 221264 542964 221270
rect 542912 221206 542964 221212
rect 542728 220652 542780 220658
rect 542728 220594 542780 220600
rect 541716 220380 541768 220386
rect 541716 220322 541768 220328
rect 542542 220280 542598 220289
rect 542542 220215 542598 220224
rect 542358 219192 542414 219201
rect 542358 219127 542414 219136
rect 542372 218482 542400 219127
rect 542556 219026 542584 220215
rect 542544 219020 542596 219026
rect 542544 218962 542596 218968
rect 542360 218476 542412 218482
rect 542360 218418 542412 218424
rect 542176 217728 542228 217734
rect 542176 217670 542228 217676
rect 542360 217728 542412 217734
rect 542360 217670 542412 217676
rect 542188 217462 542216 217670
rect 541992 217456 542044 217462
rect 541992 217398 542044 217404
rect 542176 217456 542228 217462
rect 542176 217398 542228 217404
rect 542004 217297 542032 217398
rect 542372 217326 542400 217670
rect 542360 217320 542412 217326
rect 541990 217288 542046 217297
rect 540808 217246 540882 217274
rect 541452 217246 541664 217274
rect 539152 217110 539226 217138
rect 539198 216988 539226 217110
rect 540026 217110 540100 217138
rect 540026 216988 540054 217110
rect 540854 216988 540882 217246
rect 541636 217138 541664 217246
rect 542360 217262 542412 217268
rect 541990 217223 542046 217232
rect 542740 217138 542768 220594
rect 542924 217598 542952 221206
rect 543292 220368 543320 221410
rect 543660 220658 543688 223246
rect 544948 220674 544976 226238
rect 545132 221882 545160 227258
rect 545120 221876 545172 221882
rect 545120 221818 545172 221824
rect 545132 221066 545160 221818
rect 547156 221746 547184 229978
rect 547880 227452 547932 227458
rect 547880 227394 547932 227400
rect 547420 223168 547472 223174
rect 547420 223110 547472 223116
rect 546592 221740 546644 221746
rect 546592 221682 546644 221688
rect 547144 221740 547196 221746
rect 547144 221682 547196 221688
rect 545120 221060 545172 221066
rect 545120 221002 545172 221008
rect 545764 221060 545816 221066
rect 545764 221002 545816 221008
rect 543648 220652 543700 220658
rect 544948 220646 545068 220674
rect 543648 220594 543700 220600
rect 545040 220561 545068 220646
rect 545026 220552 545082 220561
rect 545026 220487 545082 220496
rect 545302 220552 545358 220561
rect 545302 220487 545358 220496
rect 543108 220340 543320 220368
rect 542912 217592 542964 217598
rect 542912 217534 542964 217540
rect 543108 217308 543136 220340
rect 543370 220280 543426 220289
rect 543370 220215 543426 220224
rect 544200 220244 544252 220250
rect 543384 219201 543412 220215
rect 544200 220186 544252 220192
rect 543832 219360 543884 219366
rect 543832 219302 543884 219308
rect 544016 219360 544068 219366
rect 544016 219302 544068 219308
rect 543370 219192 543426 219201
rect 543370 219127 543426 219136
rect 543844 219026 543872 219302
rect 544028 219162 544056 219302
rect 544016 219156 544068 219162
rect 544016 219098 544068 219104
rect 543832 219020 543884 219026
rect 543832 218962 543884 218968
rect 543648 218476 543700 218482
rect 543648 218418 543700 218424
rect 543660 218113 543688 218418
rect 544014 218376 544070 218385
rect 544014 218311 544070 218320
rect 543462 218104 543518 218113
rect 543462 218039 543518 218048
rect 543646 218104 543702 218113
rect 543646 218039 543702 218048
rect 543476 217598 543504 218039
rect 544028 217682 544056 218311
rect 543706 217654 544056 217682
rect 543706 217598 543734 217654
rect 543464 217592 543516 217598
rect 543464 217534 543516 217540
rect 543694 217592 543746 217598
rect 543694 217534 543746 217540
rect 543832 217592 543884 217598
rect 543832 217534 543884 217540
rect 543108 217280 543366 217308
rect 543844 217297 543872 217534
rect 541636 217110 541710 217138
rect 541682 216988 541710 217110
rect 542510 217110 542768 217138
rect 542510 216988 542538 217110
rect 543338 216988 543366 217280
rect 543830 217288 543886 217297
rect 543830 217223 543886 217232
rect 544212 217138 544240 220186
rect 545040 217138 545068 220487
rect 545316 218890 545344 220487
rect 545304 218884 545356 218890
rect 545304 218826 545356 218832
rect 545776 217308 545804 221002
rect 545948 220652 546000 220658
rect 545948 220594 546000 220600
rect 546132 220652 546184 220658
rect 546132 220594 546184 220600
rect 545960 218482 545988 220594
rect 545948 218476 546000 218482
rect 545948 218418 546000 218424
rect 545776 217280 545850 217308
rect 544166 217110 544240 217138
rect 544994 217110 545068 217138
rect 544166 216988 544194 217110
rect 544994 216988 545022 217110
rect 545822 216988 545850 217280
rect 546144 217122 546172 220594
rect 546604 217138 546632 221682
rect 547432 218890 547460 223110
rect 547420 218884 547472 218890
rect 547420 218826 547472 218832
rect 547432 217138 547460 218826
rect 547892 217190 547920 227394
rect 549272 223038 549300 230114
rect 555436 230042 555464 251194
rect 558196 236094 558224 265610
rect 645872 261526 645900 277766
rect 647252 265674 647280 277766
rect 648724 277394 648752 277780
rect 648632 277366 648752 277394
rect 647240 265668 647292 265674
rect 647240 265610 647292 265616
rect 570604 261520 570656 261526
rect 570604 261462 570656 261468
rect 645860 261520 645912 261526
rect 645860 261462 645912 261468
rect 568580 260908 568632 260914
rect 568580 260850 568632 260856
rect 567844 259480 567896 259486
rect 567844 259422 567896 259428
rect 562324 256760 562376 256766
rect 562324 256702 562376 256708
rect 559564 253428 559616 253434
rect 559564 253370 559616 253376
rect 558184 236088 558236 236094
rect 558184 236030 558236 236036
rect 555424 230036 555476 230042
rect 555424 229978 555476 229984
rect 556804 229900 556856 229906
rect 556804 229842 556856 229848
rect 555608 229764 555660 229770
rect 555608 229706 555660 229712
rect 551560 228948 551612 228954
rect 551560 228890 551612 228896
rect 549904 224800 549956 224806
rect 549904 224742 549956 224748
rect 548064 223032 548116 223038
rect 548064 222974 548116 222980
rect 549260 223032 549312 223038
rect 549260 222974 549312 222980
rect 548076 221134 548104 222974
rect 549916 222194 549944 224742
rect 550640 224392 550692 224398
rect 550640 224334 550692 224340
rect 549916 222166 550128 222194
rect 548064 221128 548116 221134
rect 548064 221070 548116 221076
rect 548076 217308 548104 221070
rect 550100 219910 550128 222166
rect 550652 221270 550680 224334
rect 550364 221264 550416 221270
rect 550364 221206 550416 221212
rect 550640 221264 550692 221270
rect 550640 221206 550692 221212
rect 551284 221264 551336 221270
rect 551284 221206 551336 221212
rect 550376 221082 550404 221206
rect 550376 221054 550588 221082
rect 550560 220658 550588 221054
rect 551296 220814 551324 221206
rect 551296 220786 551416 220814
rect 550272 220652 550324 220658
rect 550272 220594 550324 220600
rect 550548 220652 550600 220658
rect 550548 220594 550600 220600
rect 548892 219904 548944 219910
rect 548892 219846 548944 219852
rect 550088 219904 550140 219910
rect 550088 219846 550140 219852
rect 548904 218890 548932 219846
rect 548248 218884 548300 218890
rect 548248 218826 548300 218832
rect 548892 218884 548944 218890
rect 548892 218826 548944 218832
rect 548260 218770 548288 218826
rect 548260 218742 548840 218770
rect 548812 218482 548840 218742
rect 548800 218476 548852 218482
rect 548800 218418 548852 218424
rect 548444 218062 549484 218090
rect 548444 217326 548472 218062
rect 549076 217456 549128 217462
rect 549260 217456 549312 217462
rect 549128 217404 549260 217410
rect 549076 217398 549312 217404
rect 549088 217382 549300 217398
rect 548432 217320 548484 217326
rect 548076 217280 548334 217308
rect 547880 217184 547932 217190
rect 546132 217116 546184 217122
rect 546604 217110 546678 217138
rect 547432 217110 547506 217138
rect 547880 217126 547932 217132
rect 546132 217058 546184 217064
rect 546650 216988 546678 217110
rect 547478 216988 547506 217110
rect 548306 216988 548334 217280
rect 548432 217262 548484 217268
rect 549456 217122 549484 218062
rect 550100 217172 550128 219846
rect 550284 217326 550312 220594
rect 551020 217926 551232 217954
rect 551020 217802 551048 217926
rect 551008 217796 551060 217802
rect 551008 217738 551060 217744
rect 551204 217734 551232 217926
rect 551192 217728 551244 217734
rect 550468 217654 550864 217682
rect 551192 217670 551244 217676
rect 550272 217320 550324 217326
rect 550272 217262 550324 217268
rect 549962 217144 550128 217172
rect 549122 217116 549174 217122
rect 549122 217058 549174 217064
rect 549444 217116 549496 217122
rect 549444 217058 549496 217064
rect 549134 216988 549162 217058
rect 549962 216988 549990 217144
rect 550468 217138 550496 217654
rect 550836 217308 550864 217654
rect 551008 217320 551060 217326
rect 550836 217280 551008 217308
rect 551008 217262 551060 217268
rect 551388 217190 551416 220786
rect 551572 217308 551600 228890
rect 554044 225888 554096 225894
rect 554044 225830 554096 225836
rect 553216 225752 553268 225758
rect 553216 225694 553268 225700
rect 553228 220998 553256 225694
rect 553584 222148 553636 222154
rect 553584 222090 553636 222096
rect 552848 220992 552900 220998
rect 552848 220934 552900 220940
rect 553216 220992 553268 220998
rect 553216 220934 553268 220940
rect 552480 220244 552532 220250
rect 552480 220186 552532 220192
rect 551744 217456 551796 217462
rect 551744 217398 551796 217404
rect 551572 217280 551646 217308
rect 550916 217184 550968 217190
rect 550376 217122 550496 217138
rect 550364 217116 550496 217122
rect 550416 217110 550496 217116
rect 550790 217132 550916 217138
rect 550790 217126 550968 217132
rect 551376 217184 551428 217190
rect 551376 217126 551428 217132
rect 550790 217110 550956 217126
rect 550364 217058 550416 217064
rect 550790 216988 550818 217110
rect 551618 216988 551646 217280
rect 551756 217190 551784 217398
rect 551744 217184 551796 217190
rect 552492 217138 552520 220186
rect 551744 217126 551796 217132
rect 552446 217110 552520 217138
rect 552860 217138 552888 220934
rect 553030 220280 553086 220289
rect 553030 220215 553086 220224
rect 553044 219178 553072 220215
rect 553596 220046 553624 222090
rect 553768 220652 553820 220658
rect 553768 220594 553820 220600
rect 553780 220046 553808 220594
rect 553216 220040 553268 220046
rect 553216 219982 553268 219988
rect 553584 220040 553636 220046
rect 553584 219982 553636 219988
rect 553768 220040 553820 220046
rect 553768 219982 553820 219988
rect 553228 219298 553256 219982
rect 553216 219292 553268 219298
rect 553216 219234 553268 219240
rect 553044 219162 553532 219178
rect 553044 219156 553544 219162
rect 553044 219150 553492 219156
rect 553492 219098 553544 219104
rect 553584 218884 553636 218890
rect 553584 218826 553636 218832
rect 553596 217818 553624 218826
rect 553504 217790 553624 217818
rect 553504 217462 553532 217790
rect 553492 217456 553544 217462
rect 553492 217398 553544 217404
rect 554056 217308 554084 225830
rect 555620 220658 555648 229706
rect 556528 224528 556580 224534
rect 556528 224470 556580 224476
rect 555790 222048 555846 222057
rect 555790 221983 555792 221992
rect 555844 221983 555846 221992
rect 555792 221954 555844 221960
rect 555608 220652 555660 220658
rect 555608 220594 555660 220600
rect 554964 220380 555016 220386
rect 554964 220322 555016 220328
rect 554056 217280 554130 217308
rect 552860 217110 553302 217138
rect 552446 216988 552474 217110
rect 553274 216988 553302 217110
rect 554102 216988 554130 217280
rect 554976 217138 555004 220322
rect 555804 217138 555832 221954
rect 554930 217110 555004 217138
rect 555758 217110 555832 217138
rect 556540 217138 556568 224470
rect 556816 222018 556844 229842
rect 558184 228540 558236 228546
rect 558184 228482 558236 228488
rect 558196 224954 558224 228482
rect 559012 225616 559064 225622
rect 559012 225558 559064 225564
rect 558196 224926 558316 224954
rect 556804 222012 556856 222018
rect 556804 221954 556856 221960
rect 558288 221746 558316 224926
rect 556712 221740 556764 221746
rect 556712 221682 556764 221688
rect 557816 221740 557868 221746
rect 557816 221682 557868 221688
rect 558276 221740 558328 221746
rect 558276 221682 558328 221688
rect 556724 220289 556752 221682
rect 556710 220280 556766 220289
rect 556710 220215 556766 220224
rect 556724 217308 556752 220215
rect 557264 218748 557316 218754
rect 557264 218690 557316 218696
rect 557276 217598 557304 218690
rect 557264 217592 557316 217598
rect 557264 217534 557316 217540
rect 557540 217592 557592 217598
rect 557540 217534 557592 217540
rect 557552 217326 557580 217534
rect 557540 217320 557592 217326
rect 556724 217280 557442 217308
rect 556540 217110 556614 217138
rect 554930 216988 554958 217110
rect 555758 216988 555786 217110
rect 556586 216988 556614 217110
rect 557414 216988 557442 217280
rect 557828 217308 557856 221682
rect 558000 220040 558052 220046
rect 558052 219988 558776 219994
rect 558000 219982 558776 219988
rect 558012 219966 558776 219982
rect 558748 219162 558776 219966
rect 558552 219156 558604 219162
rect 558552 219098 558604 219104
rect 558736 219156 558788 219162
rect 558736 219098 558788 219104
rect 558564 218385 558592 219098
rect 558366 218376 558422 218385
rect 558366 218311 558422 218320
rect 558550 218376 558606 218385
rect 558550 218311 558606 218320
rect 558380 217326 558408 218311
rect 558368 217320 558420 217326
rect 557828 217280 558270 217308
rect 557540 217262 557592 217268
rect 558242 216988 558270 217280
rect 559024 217308 559052 225558
rect 559576 220386 559604 253370
rect 561588 228676 561640 228682
rect 561588 228618 561640 228624
rect 560668 222896 560720 222902
rect 560668 222838 560720 222844
rect 560680 222329 560708 222838
rect 560666 222320 560722 222329
rect 560666 222255 560722 222264
rect 559840 220652 559892 220658
rect 559840 220594 559892 220600
rect 559564 220380 559616 220386
rect 559564 220322 559616 220328
rect 559024 217280 559098 217308
rect 558368 217262 558420 217268
rect 559070 216988 559098 217280
rect 559852 217138 559880 220594
rect 560680 217308 560708 222255
rect 561600 217308 561628 228618
rect 562336 226302 562364 256702
rect 566372 228404 566424 228410
rect 566372 228346 566424 228352
rect 563888 227180 563940 227186
rect 563888 227122 563940 227128
rect 562324 226296 562376 226302
rect 562324 226238 562376 226244
rect 562692 226024 562744 226030
rect 562692 225966 562744 225972
rect 562508 222692 562560 222698
rect 562508 222634 562560 222640
rect 561954 222320 562010 222329
rect 562520 222290 562548 222634
rect 562704 222329 562732 225966
rect 563900 224954 563928 227122
rect 565636 227044 565688 227050
rect 565636 226986 565688 226992
rect 563900 224926 564020 224954
rect 563796 224256 563848 224262
rect 563796 224198 563848 224204
rect 563808 222834 563836 224198
rect 563796 222828 563848 222834
rect 563796 222770 563848 222776
rect 563808 222714 563836 222770
rect 563808 222686 563928 222714
rect 562690 222320 562746 222329
rect 561954 222255 562010 222264
rect 562508 222284 562560 222290
rect 560680 217280 560754 217308
rect 559852 217110 559926 217138
rect 559898 216988 559926 217110
rect 560726 216988 560754 217280
rect 561554 217280 561628 217308
rect 561968 217308 561996 222255
rect 562690 222255 562746 222264
rect 562508 222226 562560 222232
rect 562888 222166 563192 222194
rect 562692 222012 562744 222018
rect 562692 221954 562744 221960
rect 562704 221626 562732 221954
rect 562888 221746 562916 222166
rect 563164 221898 563192 222166
rect 563704 222148 563756 222154
rect 563704 222090 563756 222096
rect 563426 222048 563482 222057
rect 563426 221983 563428 221992
rect 563480 221983 563482 221992
rect 563428 221954 563480 221960
rect 563164 221870 563284 221898
rect 563256 221762 563284 221870
rect 563716 221762 563744 222090
rect 562876 221740 562928 221746
rect 562876 221682 562928 221688
rect 563060 221740 563112 221746
rect 563256 221734 563744 221762
rect 563060 221682 563112 221688
rect 563072 221626 563100 221682
rect 562704 221598 563100 221626
rect 562520 220374 563100 220402
rect 562520 220289 562548 220374
rect 562506 220280 562562 220289
rect 562874 220280 562930 220289
rect 562506 220215 562562 220224
rect 562692 220244 562744 220250
rect 563072 220250 563100 220374
rect 562874 220215 562930 220224
rect 563060 220244 563112 220250
rect 562692 220186 562744 220192
rect 562704 218634 562732 220186
rect 562888 219026 562916 220215
rect 563060 220186 563112 220192
rect 563014 219156 563066 219162
rect 563066 219116 563560 219144
rect 563014 219098 563066 219104
rect 562876 219020 562928 219026
rect 563152 219020 563204 219026
rect 562876 218962 562928 218968
rect 563026 218980 563152 219008
rect 563026 218906 563054 218980
rect 563152 218962 563204 218968
rect 563336 219020 563388 219026
rect 563336 218962 563388 218968
rect 562888 218878 563054 218906
rect 562888 218754 562916 218878
rect 563348 218872 563376 218962
rect 563164 218844 563376 218872
rect 563164 218770 563192 218844
rect 562876 218748 562928 218754
rect 563072 218742 563192 218770
rect 563336 218748 563388 218754
rect 563072 218736 563100 218742
rect 562876 218690 562928 218696
rect 563026 218708 563100 218736
rect 563026 218634 563054 218708
rect 563336 218690 563388 218696
rect 562704 218606 563054 218634
rect 563348 217954 563376 218690
rect 563532 218226 563560 219116
rect 563072 217926 563376 217954
rect 563440 218198 563560 218226
rect 563072 217841 563100 217926
rect 563058 217832 563114 217841
rect 563058 217767 563114 217776
rect 563242 217832 563298 217841
rect 563242 217767 563298 217776
rect 562876 217320 562928 217326
rect 561968 217280 562410 217308
rect 561554 216988 561582 217280
rect 562382 216988 562410 217280
rect 563256 217308 563284 217767
rect 563440 217326 563468 218198
rect 563900 217546 563928 222686
rect 563716 217518 563928 217546
rect 563992 217546 564020 224926
rect 564808 223032 564860 223038
rect 564808 222974 564860 222980
rect 564820 222698 564848 222974
rect 564624 222692 564676 222698
rect 564624 222634 564676 222640
rect 564808 222692 564860 222698
rect 564808 222634 564860 222640
rect 564636 222290 564664 222634
rect 564624 222284 564676 222290
rect 564624 222226 564676 222232
rect 564346 217832 564402 217841
rect 564346 217767 564402 217776
rect 564530 217832 564586 217841
rect 564530 217767 564586 217776
rect 563992 217518 564066 217546
rect 562928 217280 563284 217308
rect 563428 217320 563480 217326
rect 562876 217262 562928 217268
rect 563428 217262 563480 217268
rect 563716 217138 563744 217518
rect 563210 217110 563744 217138
rect 563210 216988 563238 217110
rect 564038 216988 564066 217518
rect 564360 217462 564388 217767
rect 564164 217456 564216 217462
rect 564164 217398 564216 217404
rect 564348 217456 564400 217462
rect 564348 217398 564400 217404
rect 564176 217308 564204 217398
rect 564544 217308 564572 217767
rect 564176 217280 564572 217308
rect 564820 217138 564848 222634
rect 565648 222601 565676 226986
rect 566384 224954 566412 228346
rect 567568 226296 567620 226302
rect 567568 226238 567620 226244
rect 566384 224926 566504 224954
rect 565634 222592 565690 222601
rect 565634 222527 565690 222536
rect 565648 217308 565676 222527
rect 566476 217308 566504 224926
rect 566832 222964 566884 222970
rect 566832 222906 566884 222912
rect 566648 221740 566700 221746
rect 566648 221682 566700 221688
rect 566660 217308 566688 221682
rect 566844 220561 566872 222906
rect 567384 222420 567436 222426
rect 567384 222362 567436 222368
rect 567396 221746 567424 222362
rect 567384 221740 567436 221746
rect 567384 221682 567436 221688
rect 567580 220810 567608 226238
rect 567856 224262 567884 259422
rect 568592 229094 568620 260850
rect 570616 234598 570644 261462
rect 571340 249076 571392 249082
rect 571340 249018 571392 249024
rect 570604 234592 570656 234598
rect 570604 234534 570656 234540
rect 569960 230036 570012 230042
rect 569960 229978 570012 229984
rect 569972 229094 570000 229978
rect 571352 229094 571380 249018
rect 632704 246356 632756 246362
rect 632704 246298 632756 246304
rect 591304 245676 591356 245682
rect 591304 245618 591356 245624
rect 576124 242208 576176 242214
rect 576124 242150 576176 242156
rect 576136 238746 576164 242150
rect 577504 240168 577556 240174
rect 577504 240110 577556 240116
rect 576124 238740 576176 238746
rect 576124 238682 576176 238688
rect 568592 229066 568896 229094
rect 569972 229066 570644 229094
rect 571352 229066 571656 229094
rect 568868 224954 568896 229066
rect 568868 224926 569816 224954
rect 567844 224256 567896 224262
rect 567844 224198 567896 224204
rect 568948 224256 569000 224262
rect 568948 224198 569000 224204
rect 567752 221740 567804 221746
rect 567752 221682 567804 221688
rect 567764 220998 567792 221682
rect 567752 220992 567804 220998
rect 567752 220934 567804 220940
rect 567580 220782 567792 220810
rect 566830 220552 566886 220561
rect 566830 220487 566886 220496
rect 567014 220552 567070 220561
rect 567014 220487 567070 220496
rect 567028 219450 567056 220487
rect 567200 220380 567252 220386
rect 567200 220322 567252 220328
rect 567384 220380 567436 220386
rect 567384 220322 567436 220328
rect 566936 219422 567056 219450
rect 566936 219026 566964 219422
rect 567212 219026 567240 220322
rect 566924 219020 566976 219026
rect 566924 218962 566976 218968
rect 567200 219020 567252 219026
rect 567200 218962 567252 218968
rect 567200 218884 567252 218890
rect 567200 218826 567252 218832
rect 567212 218362 567240 218826
rect 567396 218482 567424 220322
rect 567764 220266 567792 220782
rect 567672 220238 567792 220266
rect 567672 219314 567700 220238
rect 567844 219428 568172 219434
rect 567896 219406 568120 219428
rect 567844 219370 567896 219376
rect 568120 219370 568172 219376
rect 567672 219286 567884 219314
rect 567658 219192 567714 219201
rect 567658 219127 567714 219136
rect 567672 218754 567700 219127
rect 567660 218748 567712 218754
rect 567660 218690 567712 218696
rect 567384 218476 567436 218482
rect 567384 218418 567436 218424
rect 567568 218476 567620 218482
rect 567568 218418 567620 218424
rect 567580 218362 567608 218418
rect 567212 218334 567608 218362
rect 567856 218054 567884 219286
rect 568028 219292 568080 219298
rect 568028 219234 568080 219240
rect 568040 219144 568068 219234
rect 568396 219156 568448 219162
rect 568040 219116 568396 219144
rect 568396 219098 568448 219104
rect 568120 218748 568172 218754
rect 568120 218690 568172 218696
rect 568132 218385 568160 218690
rect 568118 218376 568174 218385
rect 568118 218311 568174 218320
rect 567856 218026 567976 218054
rect 567948 217308 567976 218026
rect 565648 217280 565722 217308
rect 566476 217280 566550 217308
rect 566660 217280 567378 217308
rect 567948 217280 568206 217308
rect 564820 217110 564894 217138
rect 564866 216988 564894 217110
rect 565694 216988 565722 217280
rect 566522 216988 566550 217280
rect 567350 216988 567378 217280
rect 568178 216988 568206 217280
rect 568960 217138 568988 224198
rect 569316 222012 569368 222018
rect 569316 221954 569368 221960
rect 569592 222012 569644 222018
rect 569592 221954 569644 221960
rect 569328 221270 569356 221954
rect 569604 221746 569632 221954
rect 569592 221740 569644 221746
rect 569592 221682 569644 221688
rect 569132 221264 569184 221270
rect 569132 221206 569184 221212
rect 569316 221264 569368 221270
rect 569316 221206 569368 221212
rect 569144 220998 569172 221206
rect 569132 220992 569184 220998
rect 569132 220934 569184 220940
rect 569788 217308 569816 224926
rect 569960 222828 570012 222834
rect 569960 222770 570012 222776
rect 569972 221746 570000 222770
rect 569960 221740 570012 221746
rect 569960 221682 570012 221688
rect 570616 217308 570644 229066
rect 571628 227714 571656 229066
rect 571444 227686 571656 227714
rect 570800 219116 571196 219144
rect 570800 217326 570828 219116
rect 571168 219026 571196 219116
rect 570972 219020 571024 219026
rect 570972 218962 571024 218968
rect 571156 219020 571208 219026
rect 571156 218962 571208 218968
rect 570788 217320 570840 217326
rect 569788 217280 569862 217308
rect 570616 217280 570690 217308
rect 568960 217110 569034 217138
rect 569006 216988 569034 217110
rect 569834 216988 569862 217280
rect 570662 216988 570690 217280
rect 570788 217262 570840 217268
rect 570984 217138 571012 218962
rect 571444 218634 571472 227686
rect 576400 222964 576452 222970
rect 576400 222906 576452 222912
rect 574100 222692 574152 222698
rect 574100 222634 574152 222640
rect 571708 222556 571760 222562
rect 571708 222498 571760 222504
rect 572812 222556 572864 222562
rect 572812 222498 572864 222504
rect 571720 222034 571748 222498
rect 572304 222048 572360 222057
rect 571720 222006 572304 222034
rect 572304 221983 572360 221992
rect 572824 220386 572852 222498
rect 572352 220380 572404 220386
rect 572352 220322 572404 220328
rect 572812 220380 572864 220386
rect 572812 220322 572864 220328
rect 572364 219298 572392 220322
rect 572994 220280 573050 220289
rect 572994 220215 573050 220224
rect 573008 219434 573036 220215
rect 573008 219406 573128 219434
rect 572168 219292 572220 219298
rect 572168 219234 572220 219240
rect 572352 219292 572404 219298
rect 572352 219234 572404 219240
rect 572180 219042 572208 219234
rect 572352 219156 572404 219162
rect 572404 219116 572944 219144
rect 572352 219098 572404 219104
rect 572180 219014 572300 219042
rect 571156 218612 571208 218618
rect 571444 218606 571840 218634
rect 571156 218554 571208 218560
rect 571168 218346 571196 218554
rect 571614 218376 571670 218385
rect 571156 218340 571208 218346
rect 571614 218311 571670 218320
rect 571156 218282 571208 218288
rect 571628 218210 571656 218311
rect 571616 218204 571668 218210
rect 571616 218146 571668 218152
rect 571154 217832 571210 217841
rect 571154 217767 571210 217776
rect 571168 217326 571196 217767
rect 571812 217682 571840 218606
rect 571984 218612 572036 218618
rect 572036 218572 572208 218600
rect 571984 218554 572036 218560
rect 572180 218054 572208 218572
rect 572272 218226 572300 219014
rect 572916 218754 572944 219116
rect 573100 218890 573128 219406
rect 574112 219298 574140 222634
rect 575846 220280 575902 220289
rect 575846 220215 575902 220224
rect 573732 219292 573784 219298
rect 573732 219234 573784 219240
rect 574100 219292 574152 219298
rect 574100 219234 574152 219240
rect 573088 218884 573140 218890
rect 573088 218826 573140 218832
rect 572720 218748 572772 218754
rect 572720 218690 572772 218696
rect 572904 218748 572956 218754
rect 572904 218690 572956 218696
rect 572536 218612 572588 218618
rect 572536 218554 572588 218560
rect 572548 218346 572576 218554
rect 572732 218346 572760 218690
rect 572536 218340 572588 218346
rect 572536 218282 572588 218288
rect 572720 218340 572772 218346
rect 572720 218282 572772 218288
rect 573744 218226 573772 219234
rect 574848 218980 575612 219008
rect 574848 218346 574876 218980
rect 575584 218890 575612 218980
rect 575434 218884 575486 218890
rect 575434 218826 575486 218832
rect 575572 218884 575624 218890
rect 575572 218826 575624 218832
rect 575446 218498 575474 218826
rect 575860 218754 575888 220215
rect 576032 219156 576084 219162
rect 576032 219098 576084 219104
rect 575572 218748 575624 218754
rect 575572 218690 575624 218696
rect 575848 218748 575900 218754
rect 575848 218690 575900 218696
rect 575400 218470 575474 218498
rect 574836 218340 574888 218346
rect 574836 218282 574888 218288
rect 572272 218198 573588 218226
rect 573744 218198 574692 218226
rect 573560 218054 573588 218198
rect 574664 218054 574692 218198
rect 572180 218026 573496 218054
rect 573560 218026 574600 218054
rect 574664 218026 574876 218054
rect 572272 217926 573312 217954
rect 572272 217682 572300 217926
rect 571628 217654 571840 217682
rect 572180 217654 572300 217682
rect 571156 217320 571208 217326
rect 571156 217262 571208 217268
rect 570984 217110 571518 217138
rect 571490 216988 571518 217110
rect 571628 217036 571656 217654
rect 572180 217546 572208 217654
rect 571812 217518 572208 217546
rect 572720 217592 572772 217598
rect 572772 217552 572944 217580
rect 572720 217534 572772 217540
rect 571812 217462 571840 217518
rect 571800 217456 571852 217462
rect 571800 217398 571852 217404
rect 571984 217456 572036 217462
rect 571984 217398 572036 217404
rect 572536 217456 572588 217462
rect 572720 217456 572772 217462
rect 572588 217416 572720 217444
rect 572536 217398 572588 217404
rect 572720 217398 572772 217404
rect 571996 217190 572024 217398
rect 572916 217308 572944 217552
rect 573284 217462 573312 217926
rect 573272 217456 573324 217462
rect 573272 217398 573324 217404
rect 573468 217410 573496 218026
rect 574572 217841 574600 218026
rect 574374 217832 574430 217841
rect 574374 217767 574430 217776
rect 574558 217832 574614 217841
rect 574558 217767 574614 217776
rect 574388 217682 574416 217767
rect 574388 217654 574600 217682
rect 574572 217410 574600 217654
rect 573468 217382 574416 217410
rect 574572 217382 574692 217410
rect 573272 217320 573324 217326
rect 572916 217280 573272 217308
rect 573272 217262 573324 217268
rect 571984 217184 572036 217190
rect 573088 217184 573140 217190
rect 572732 217144 573088 217172
rect 572732 217138 572760 217144
rect 571984 217126 572036 217132
rect 572180 217110 572346 217138
rect 572456 217122 572760 217138
rect 573088 217126 573140 217132
rect 574192 217184 574244 217190
rect 574192 217126 574244 217132
rect 572180 217036 572208 217110
rect 571628 217008 572208 217036
rect 572318 216988 572346 217110
rect 572444 217116 572760 217122
rect 572496 217110 572760 217116
rect 572444 217058 572496 217064
rect 574204 213518 574232 217126
rect 574388 215150 574416 217382
rect 574664 216646 574692 217382
rect 574652 216640 574704 216646
rect 574652 216582 574704 216588
rect 574376 215144 574428 215150
rect 574376 215086 574428 215092
rect 574848 214742 574876 218026
rect 575204 217592 575256 217598
rect 575204 217534 575256 217540
rect 575216 217190 575244 217534
rect 575204 217184 575256 217190
rect 575204 217126 575256 217132
rect 574836 214736 574888 214742
rect 574836 214678 574888 214684
rect 574192 213512 574244 213518
rect 574192 213454 574244 213460
rect 575400 213246 575428 218470
rect 575584 215286 575612 218690
rect 575756 218476 575808 218482
rect 575756 218418 575808 218424
rect 575572 215280 575624 215286
rect 575572 215222 575624 215228
rect 575768 214470 575796 218418
rect 576044 217598 576072 219098
rect 576216 219020 576268 219026
rect 576216 218962 576268 218968
rect 576032 217592 576084 217598
rect 576032 217534 576084 217540
rect 575756 214464 575808 214470
rect 575756 214406 575808 214412
rect 576228 213654 576256 218962
rect 576412 214878 576440 222906
rect 576582 222048 576638 222057
rect 576582 221983 576638 221992
rect 576596 218482 576624 221983
rect 576584 218476 576636 218482
rect 576584 218418 576636 218424
rect 576860 216504 576912 216510
rect 576860 216446 576912 216452
rect 577318 216472 577374 216481
rect 576872 215294 576900 216446
rect 577318 216407 577374 216416
rect 577332 215937 577360 216407
rect 577318 215928 577374 215937
rect 577318 215863 577374 215872
rect 576872 215266 577084 215294
rect 577056 215121 577084 215266
rect 577042 215112 577098 215121
rect 577042 215047 577098 215056
rect 576400 214872 576452 214878
rect 576400 214814 576452 214820
rect 576216 213648 576268 213654
rect 575662 213616 575718 213625
rect 576216 213590 576268 213596
rect 575662 213551 575718 213560
rect 575676 213382 575704 213551
rect 575664 213376 575716 213382
rect 575664 213318 575716 213324
rect 575388 213240 575440 213246
rect 575388 213182 575440 213188
rect 577516 99142 577544 240110
rect 591316 235278 591344 245618
rect 624424 244316 624476 244322
rect 624424 244258 624476 244264
rect 591304 235272 591356 235278
rect 591304 235214 591356 235220
rect 593972 222420 594024 222426
rect 593972 222362 594024 222368
rect 582194 222320 582250 222329
rect 582194 222255 582250 222264
rect 577686 220552 577742 220561
rect 582208 220538 582236 222255
rect 593236 222148 593288 222154
rect 593236 222090 593288 222096
rect 593248 221134 593276 222090
rect 593236 221128 593288 221134
rect 593236 221070 593288 221076
rect 591960 220918 592356 220946
rect 591960 220862 591988 220918
rect 591948 220856 592000 220862
rect 591948 220798 592000 220804
rect 592132 220788 592184 220794
rect 592132 220730 592184 220736
rect 582378 220688 582434 220697
rect 582378 220623 582434 220632
rect 591854 220688 591910 220697
rect 591854 220623 591910 220632
rect 582392 220538 582420 220623
rect 582208 220510 582420 220538
rect 591868 220538 591896 220623
rect 591868 220510 592034 220538
rect 577686 220487 577742 220496
rect 577700 215014 577728 220487
rect 582194 220416 582250 220425
rect 582194 220351 582196 220360
rect 582248 220351 582250 220360
rect 582378 220416 582434 220425
rect 582378 220351 582380 220360
rect 582196 220322 582248 220328
rect 582432 220351 582434 220360
rect 591854 220416 591910 220425
rect 592006 220386 592034 220510
rect 592144 220425 592172 220730
rect 592328 220697 592356 220918
rect 592314 220688 592370 220697
rect 592314 220623 592370 220632
rect 592130 220416 592186 220425
rect 591854 220351 591856 220360
rect 582380 220322 582432 220328
rect 591908 220351 591910 220360
rect 591994 220380 592046 220386
rect 591856 220322 591908 220328
rect 592130 220351 592186 220360
rect 591994 220322 592046 220328
rect 577872 219292 577924 219298
rect 577872 219234 577924 219240
rect 577688 215008 577740 215014
rect 577688 214950 577740 214956
rect 577884 214606 577912 219234
rect 592130 219192 592186 219201
rect 592130 219127 592132 219136
rect 592184 219127 592186 219136
rect 592314 219192 592370 219201
rect 592314 219127 592370 219136
rect 592132 219098 592184 219104
rect 582932 218748 582984 218754
rect 582932 218690 582984 218696
rect 591948 218748 592000 218754
rect 591948 218690 592000 218696
rect 592132 218748 592184 218754
rect 592132 218690 592184 218696
rect 582944 218385 582972 218690
rect 591960 218385 591988 218690
rect 592144 218385 592172 218690
rect 582102 218376 582158 218385
rect 582102 218311 582158 218320
rect 582286 218376 582342 218385
rect 582286 218311 582342 218320
rect 582746 218376 582802 218385
rect 582746 218311 582802 218320
rect 582930 218376 582986 218385
rect 582930 218311 582986 218320
rect 591946 218376 592002 218385
rect 591946 218311 592002 218320
rect 592130 218376 592186 218385
rect 592130 218311 592186 218320
rect 582116 218210 582144 218311
rect 581920 218204 581972 218210
rect 581920 218146 581972 218152
rect 582104 218204 582156 218210
rect 582104 218146 582156 218152
rect 581932 218090 581960 218146
rect 582300 218090 582328 218311
rect 582760 218210 582788 218311
rect 582564 218204 582616 218210
rect 582564 218146 582616 218152
rect 582748 218204 582800 218210
rect 582748 218146 582800 218152
rect 591684 218198 592172 218226
rect 592328 218210 592356 219127
rect 581932 218062 582328 218090
rect 582576 218090 582604 218146
rect 582930 218104 582986 218113
rect 582576 218062 582930 218090
rect 582930 218039 582986 218048
rect 591684 217841 591712 218198
rect 591854 218104 591910 218113
rect 591854 218039 591910 218048
rect 582378 217832 582434 217841
rect 591670 217832 591726 217841
rect 582434 217790 582696 217818
rect 582378 217767 582434 217776
rect 582668 217054 582696 217790
rect 591868 217818 591896 218039
rect 592144 217977 592172 218198
rect 592316 218204 592368 218210
rect 592316 218146 592368 218152
rect 592130 217968 592186 217977
rect 592130 217903 592186 217912
rect 591868 217790 592632 217818
rect 591670 217767 591726 217776
rect 590106 217560 590162 217569
rect 590106 217495 590162 217504
rect 582656 217048 582708 217054
rect 582332 217016 582388 217025
rect 582388 216974 582512 217002
rect 582656 216990 582708 216996
rect 582332 216951 582388 216960
rect 582484 216918 582512 216974
rect 582472 216912 582524 216918
rect 582472 216854 582524 216860
rect 582564 216640 582616 216646
rect 582564 216582 582616 216588
rect 582576 216481 582604 216582
rect 582748 216504 582800 216510
rect 582378 216472 582434 216481
rect 582378 216407 582434 216416
rect 582562 216472 582618 216481
rect 582748 216446 582800 216452
rect 582562 216407 582618 216416
rect 582392 216306 582420 216407
rect 582380 216300 582432 216306
rect 582380 216242 582432 216248
rect 582760 216209 582788 216446
rect 582746 216200 582802 216209
rect 590120 216170 590148 217495
rect 591762 217288 591818 217297
rect 591762 217223 591818 217232
rect 592222 217288 592278 217297
rect 592222 217223 592278 217232
rect 591776 217054 591804 217223
rect 592236 217054 592264 217223
rect 592604 217054 592632 217790
rect 593512 217592 593564 217598
rect 593512 217534 593564 217540
rect 590292 217048 590344 217054
rect 590292 216990 590344 216996
rect 591764 217048 591816 217054
rect 591764 216990 591816 216996
rect 592224 217048 592276 217054
rect 592224 216990 592276 216996
rect 592592 217048 592644 217054
rect 592592 216990 592644 216996
rect 582746 216135 582802 216144
rect 590108 216164 590160 216170
rect 590108 216106 590160 216112
rect 590304 215626 590332 216990
rect 593524 216918 593552 217534
rect 590752 216912 590804 216918
rect 590752 216854 590804 216860
rect 593512 216912 593564 216918
rect 593512 216854 593564 216860
rect 590764 216034 590792 216854
rect 591764 216640 591816 216646
rect 591764 216582 591816 216588
rect 591776 216481 591804 216582
rect 592040 216504 592092 216510
rect 591762 216472 591818 216481
rect 591762 216407 591818 216416
rect 592038 216472 592040 216481
rect 592092 216472 592094 216481
rect 592038 216407 592094 216416
rect 592222 216336 592278 216345
rect 592222 216271 592224 216280
rect 592276 216271 592278 216280
rect 592224 216242 592276 216248
rect 590752 216028 590804 216034
rect 590752 215970 590804 215976
rect 590292 215620 590344 215626
rect 590292 215562 590344 215568
rect 577872 214600 577924 214606
rect 577872 214542 577924 214548
rect 578882 214024 578938 214033
rect 578882 213959 578938 213968
rect 578514 211712 578570 211721
rect 578514 211647 578516 211656
rect 578568 211647 578570 211656
rect 578516 211618 578568 211624
rect 578896 208350 578924 213959
rect 580448 211676 580500 211682
rect 580448 211618 580500 211624
rect 579252 209840 579304 209846
rect 579250 209808 579252 209817
rect 579304 209808 579306 209817
rect 579250 209743 579306 209752
rect 578884 208344 578936 208350
rect 578884 208286 578936 208292
rect 580460 207670 580488 211618
rect 593984 210202 594012 222362
rect 597560 222284 597612 222290
rect 597560 222226 597612 222232
rect 596456 222012 596508 222018
rect 596456 221954 596508 221960
rect 596640 222012 596692 222018
rect 596640 221954 596692 221960
rect 597192 222012 597244 222018
rect 597192 221954 597244 221960
rect 596468 221134 596496 221954
rect 596652 221474 596680 221954
rect 596824 221876 596876 221882
rect 596824 221818 596876 221824
rect 596836 221474 596864 221818
rect 596640 221468 596692 221474
rect 596640 221410 596692 221416
rect 596824 221468 596876 221474
rect 596824 221410 596876 221416
rect 596456 221128 596508 221134
rect 596456 221070 596508 221076
rect 597204 220998 597232 221954
rect 597572 221134 597600 222226
rect 607496 222148 607548 222154
rect 607496 222090 607548 222096
rect 607312 222012 607364 222018
rect 607312 221954 607364 221960
rect 606024 221876 606076 221882
rect 606024 221818 606076 221824
rect 599490 221776 599546 221785
rect 599490 221711 599546 221720
rect 601514 221776 601570 221785
rect 601514 221711 601570 221720
rect 602250 221776 602306 221785
rect 602250 221711 602306 221720
rect 597560 221128 597612 221134
rect 597560 221070 597612 221076
rect 597192 220992 597244 220998
rect 597192 220934 597244 220940
rect 596546 219192 596602 219201
rect 596546 219127 596602 219136
rect 599216 219156 599268 219162
rect 596560 218906 596588 219127
rect 599216 219098 599268 219104
rect 597006 218920 597062 218929
rect 596560 218878 597006 218906
rect 597006 218855 597062 218864
rect 596824 218612 596876 218618
rect 596824 218554 596876 218560
rect 596836 217598 596864 218554
rect 596824 217592 596876 217598
rect 596824 217534 596876 217540
rect 594798 217288 594854 217297
rect 594798 217223 594854 217232
rect 594812 210202 594840 217223
rect 595166 216744 595222 216753
rect 595166 216679 595222 216688
rect 595180 210202 595208 216679
rect 595904 216640 595956 216646
rect 595904 216582 595956 216588
rect 597558 216608 597614 216617
rect 595916 216345 595944 216582
rect 597558 216543 597614 216552
rect 596824 216504 596876 216510
rect 596824 216446 596876 216452
rect 595718 216336 595774 216345
rect 595718 216271 595774 216280
rect 595902 216336 595958 216345
rect 595902 216271 595958 216280
rect 595732 210202 595760 216271
rect 596364 216028 596416 216034
rect 596364 215970 596416 215976
rect 596376 210202 596404 215970
rect 596836 210202 596864 216446
rect 597572 210202 597600 216543
rect 599030 216336 599086 216345
rect 599030 216271 599086 216280
rect 597928 216164 597980 216170
rect 597928 216106 597980 216112
rect 597940 210202 597968 216106
rect 598480 215620 598532 215626
rect 598480 215562 598532 215568
rect 598492 210202 598520 215562
rect 599044 210202 599072 216271
rect 599228 215966 599256 219098
rect 599216 215960 599268 215966
rect 599216 215902 599268 215908
rect 599504 210202 599532 221711
rect 601528 221610 601556 221711
rect 601516 221604 601568 221610
rect 601516 221546 601568 221552
rect 600594 221232 600650 221241
rect 600594 221167 600650 221176
rect 600410 220688 600466 220697
rect 600410 220623 600466 220632
rect 600424 214334 600452 220623
rect 600412 214328 600464 214334
rect 600412 214270 600464 214276
rect 600608 210202 600636 221167
rect 600780 214328 600832 214334
rect 600780 214270 600832 214276
rect 593984 210174 594412 210202
rect 594812 210174 594964 210202
rect 595180 210174 595516 210202
rect 595732 210174 596068 210202
rect 596376 210174 596620 210202
rect 596836 210174 597172 210202
rect 597572 210174 597724 210202
rect 597940 210174 598276 210202
rect 598492 210174 598828 210202
rect 599044 210174 599380 210202
rect 599504 210174 599932 210202
rect 600484 210174 600636 210202
rect 600792 210202 600820 214270
rect 601792 213648 601844 213654
rect 601792 213590 601844 213596
rect 601240 213512 601292 213518
rect 601240 213454 601292 213460
rect 601252 210202 601280 213454
rect 601804 210202 601832 213590
rect 602264 210202 602292 221711
rect 603078 219192 603134 219201
rect 603078 219127 603134 219136
rect 603092 217870 603120 219127
rect 604460 218340 604512 218346
rect 604460 218282 604512 218288
rect 602896 217864 602948 217870
rect 602896 217806 602948 217812
rect 603080 217864 603132 217870
rect 603080 217806 603132 217812
rect 602908 212534 602936 217806
rect 604472 217734 604500 218282
rect 603448 217728 603500 217734
rect 603448 217670 603500 217676
rect 604460 217728 604512 217734
rect 604460 217670 604512 217676
rect 602908 212506 603120 212534
rect 603092 210202 603120 212506
rect 603460 210202 603488 217670
rect 604552 217320 604604 217326
rect 604552 217262 604604 217268
rect 604000 217184 604052 217190
rect 604000 217126 604052 217132
rect 604012 210202 604040 217126
rect 604564 210202 604592 217262
rect 605104 216912 605156 216918
rect 605104 216854 605156 216860
rect 605116 210202 605144 216854
rect 605840 216776 605892 216782
rect 605840 216718 605892 216724
rect 605852 210202 605880 216718
rect 606036 210338 606064 221818
rect 606668 221604 606720 221610
rect 606668 221546 606720 221552
rect 606036 210310 606156 210338
rect 606128 210202 606156 210310
rect 606680 210202 606708 221546
rect 607128 218476 607180 218482
rect 607128 218418 607180 218424
rect 607140 217326 607168 218418
rect 607128 217320 607180 217326
rect 607128 217262 607180 217268
rect 607324 214334 607352 221954
rect 607312 214328 607364 214334
rect 607312 214270 607364 214276
rect 607508 210202 607536 222090
rect 610532 221740 610584 221746
rect 610532 221682 610584 221688
rect 610072 221264 610124 221270
rect 610072 221206 610124 221212
rect 608692 221128 608744 221134
rect 608692 221070 608744 221076
rect 608704 214334 608732 221070
rect 608876 220992 608928 220998
rect 608876 220934 608928 220940
rect 607864 214328 607916 214334
rect 607864 214270 607916 214276
rect 608692 214328 608744 214334
rect 608692 214270 608744 214276
rect 607876 210202 607904 214270
rect 608888 210202 608916 220934
rect 609060 217456 609112 217462
rect 609060 217398 609112 217404
rect 600792 210174 601036 210202
rect 601252 210174 601588 210202
rect 601804 210174 602140 210202
rect 602264 210174 602692 210202
rect 603092 210174 603244 210202
rect 603460 210174 603796 210202
rect 604012 210174 604348 210202
rect 604564 210174 604900 210202
rect 605116 210174 605452 210202
rect 605852 210174 606004 210202
rect 606128 210174 606556 210202
rect 606680 210174 607108 210202
rect 607508 210174 607660 210202
rect 607876 210174 608212 210202
rect 608764 210174 608916 210202
rect 609072 210202 609100 217398
rect 609520 214328 609572 214334
rect 609520 214270 609572 214276
rect 609532 210202 609560 214270
rect 610084 210202 610112 221206
rect 610544 210202 610572 221682
rect 616878 221504 616934 221513
rect 616878 221439 616934 221448
rect 611634 220960 611690 220969
rect 611634 220895 611690 220904
rect 610806 220280 610862 220289
rect 610806 220215 610862 220224
rect 610820 219745 610848 220215
rect 610806 219736 610862 219745
rect 610806 219671 610862 219680
rect 611358 215928 611414 215937
rect 611358 215863 611414 215872
rect 611372 210202 611400 215863
rect 611648 210202 611676 220895
rect 614486 218648 614542 218657
rect 614486 218583 614542 218592
rect 613844 218068 613896 218074
rect 613844 218010 613896 218016
rect 612280 217864 612332 217870
rect 612280 217806 612332 217812
rect 612292 210202 612320 217806
rect 613384 215960 613436 215966
rect 613384 215902 613436 215908
rect 612832 213376 612884 213382
rect 612832 213318 612884 213324
rect 612844 210202 612872 213318
rect 613396 210202 613424 215902
rect 613856 215422 613884 218010
rect 614120 217048 614172 217054
rect 614120 216990 614172 216996
rect 613844 215416 613896 215422
rect 613844 215358 613896 215364
rect 614132 210202 614160 216990
rect 614500 210202 614528 218583
rect 615684 217728 615736 217734
rect 615684 217670 615736 217676
rect 615040 215416 615092 215422
rect 615040 215358 615092 215364
rect 615052 210202 615080 215358
rect 615696 210202 615724 217670
rect 616144 217320 616196 217326
rect 616144 217262 616196 217268
rect 616156 210202 616184 217262
rect 616892 214742 616920 221439
rect 620284 220788 620336 220794
rect 620284 220730 620336 220736
rect 620296 220250 620324 220730
rect 622676 220516 622728 220522
rect 622676 220458 622728 220464
rect 620100 220244 620152 220250
rect 620100 220186 620152 220192
rect 620284 220244 620336 220250
rect 620284 220186 620336 220192
rect 617062 220008 617118 220017
rect 617062 219943 617118 219952
rect 616696 214736 616748 214742
rect 616696 214678 616748 214684
rect 616880 214736 616932 214742
rect 616880 214678 616932 214684
rect 616708 214334 616736 214678
rect 616696 214328 616748 214334
rect 616696 214270 616748 214276
rect 617076 210202 617104 219943
rect 620112 219638 620140 220186
rect 621020 219768 621072 219774
rect 621020 219710 621072 219716
rect 618260 219632 618312 219638
rect 618260 219574 618312 219580
rect 620100 219632 620152 219638
rect 620100 219574 620152 219580
rect 617248 219496 617300 219502
rect 617248 219438 617300 219444
rect 609072 210174 609316 210202
rect 609532 210174 609868 210202
rect 610084 210174 610420 210202
rect 610544 210174 610972 210202
rect 611372 210174 611524 210202
rect 611648 210174 612076 210202
rect 612292 210174 612628 210202
rect 612844 210174 613180 210202
rect 613396 210174 613732 210202
rect 614132 210174 614284 210202
rect 614500 210174 614836 210202
rect 615052 210174 615388 210202
rect 615696 210174 615940 210202
rect 616156 210174 616492 210202
rect 617044 210174 617104 210202
rect 617260 210202 617288 219438
rect 617800 214736 617852 214742
rect 617800 214678 617852 214684
rect 617812 210202 617840 214678
rect 618272 210202 618300 219574
rect 618902 215656 618958 215665
rect 618902 215591 618958 215600
rect 618916 210202 618944 215591
rect 620558 215384 620614 215393
rect 620558 215319 620614 215328
rect 619640 215144 619692 215150
rect 619640 215086 619692 215092
rect 619652 210202 619680 215086
rect 620008 214464 620060 214470
rect 620008 214406 620060 214412
rect 620020 210202 620048 214406
rect 620572 210202 620600 215319
rect 621032 210202 621060 219710
rect 621664 215280 621716 215286
rect 621664 215222 621716 215228
rect 621676 210202 621704 215222
rect 622400 214872 622452 214878
rect 622400 214814 622452 214820
rect 622412 210202 622440 214814
rect 622688 210202 622716 220458
rect 623320 217592 623372 217598
rect 623320 217534 623372 217540
rect 623332 210202 623360 217534
rect 624436 214742 624464 244258
rect 628564 241528 628616 241534
rect 628564 241470 628616 241476
rect 626632 220652 626684 220658
rect 626632 220594 626684 220600
rect 625528 220108 625580 220114
rect 625528 220050 625580 220056
rect 625344 219904 625396 219910
rect 625344 219846 625396 219852
rect 624424 214736 624476 214742
rect 624424 214678 624476 214684
rect 624424 214328 624476 214334
rect 624424 214270 624476 214276
rect 623872 213240 623924 213246
rect 623872 213182 623924 213188
rect 623884 210202 623912 213182
rect 624436 210202 624464 214270
rect 625356 210202 625384 219846
rect 625540 219434 625568 220050
rect 617260 210174 617596 210202
rect 617812 210174 618148 210202
rect 618272 210174 618700 210202
rect 618916 210174 619252 210202
rect 619652 210174 619804 210202
rect 620020 210174 620356 210202
rect 620572 210174 620908 210202
rect 621032 210174 621460 210202
rect 621676 210174 622012 210202
rect 622412 210174 622564 210202
rect 622688 210174 623116 210202
rect 623332 210174 623668 210202
rect 623884 210174 624220 210202
rect 624436 210174 624772 210202
rect 625324 210174 625384 210202
rect 625448 219406 625568 219434
rect 625448 210202 625476 219406
rect 626446 218104 626502 218113
rect 626446 218039 626502 218048
rect 626080 215008 626132 215014
rect 626080 214950 626132 214956
rect 626092 210202 626120 214950
rect 626460 213926 626488 218039
rect 626644 214606 626672 220594
rect 628196 220380 628248 220386
rect 628196 220322 628248 220328
rect 628012 220244 628064 220250
rect 628012 220186 628064 220192
rect 626816 219632 626868 219638
rect 626816 219574 626868 219580
rect 626632 214600 626684 214606
rect 626632 214542 626684 214548
rect 626448 213920 626500 213926
rect 626448 213862 626500 213868
rect 626828 210202 626856 219574
rect 628024 214606 628052 220186
rect 627184 214600 627236 214606
rect 627184 214542 627236 214548
rect 628012 214600 628064 214606
rect 628012 214542 628064 214548
rect 627196 210202 627224 214542
rect 628208 210202 628236 220322
rect 628380 214464 628432 214470
rect 628380 214406 628432 214412
rect 625448 210174 625876 210202
rect 626092 210174 626428 210202
rect 626828 210174 626980 210202
rect 627196 210174 627532 210202
rect 628084 210174 628236 210202
rect 628392 210202 628420 214406
rect 628576 212770 628604 241470
rect 630954 219736 631010 219745
rect 630954 219671 631010 219680
rect 630770 219464 630826 219473
rect 630770 219399 630826 219408
rect 629942 218376 629998 218385
rect 629942 218311 629998 218320
rect 628840 214600 628892 214606
rect 628840 214542 628892 214548
rect 628564 212764 628616 212770
rect 628564 212706 628616 212712
rect 628852 210202 628880 214542
rect 629392 213920 629444 213926
rect 629392 213862 629444 213868
rect 629404 210202 629432 213862
rect 629956 210202 629984 218311
rect 630784 214606 630812 219399
rect 630772 214600 630824 214606
rect 630772 214542 630824 214548
rect 630968 210202 630996 219671
rect 631138 218648 631194 218657
rect 631138 218583 631194 218592
rect 628392 210174 628636 210202
rect 628852 210174 629188 210202
rect 629404 210174 629740 210202
rect 629956 210174 630292 210202
rect 630844 210174 630996 210202
rect 631152 210202 631180 218583
rect 631600 214600 631652 214606
rect 631600 214542 631652 214548
rect 631612 210202 631640 214542
rect 632716 212906 632744 246298
rect 648632 242214 648660 277366
rect 648620 242208 648672 242214
rect 648620 242150 648672 242156
rect 633624 235272 633676 235278
rect 633624 235214 633676 235220
rect 632704 212900 632756 212906
rect 632704 212842 632756 212848
rect 632704 212764 632756 212770
rect 632704 212706 632756 212712
rect 632716 210202 632744 212706
rect 633636 210202 633664 235214
rect 652036 232558 652064 378111
rect 652206 298480 652262 298489
rect 652206 298415 652262 298424
rect 652024 232552 652076 232558
rect 652024 232494 652076 232500
rect 640246 231432 640302 231441
rect 640246 231367 640302 231376
rect 639602 230072 639658 230081
rect 639602 230007 639658 230016
rect 638866 219192 638922 219201
rect 638866 219127 638922 219136
rect 636660 215348 636712 215354
rect 636660 215290 636712 215296
rect 633808 214736 633860 214742
rect 633808 214678 633860 214684
rect 631152 210174 631396 210202
rect 631612 210174 631948 210202
rect 632716 210174 633052 210202
rect 633604 210174 633664 210202
rect 633820 210202 633848 214678
rect 635556 213376 635608 213382
rect 635556 213318 635608 213324
rect 634360 212900 634412 212906
rect 634360 212842 634412 212848
rect 634372 210202 634400 212842
rect 635568 210202 635596 213318
rect 636672 210202 636700 215290
rect 638316 213920 638368 213926
rect 638316 213862 638368 213868
rect 637212 212764 637264 212770
rect 637212 212706 637264 212712
rect 637224 210202 637252 212706
rect 638328 210202 638356 213862
rect 638880 210202 638908 219127
rect 639616 215354 639644 230007
rect 640062 218920 640118 218929
rect 640062 218855 640118 218864
rect 639604 215348 639656 215354
rect 639604 215290 639656 215296
rect 640076 213926 640104 218855
rect 640064 213920 640116 213926
rect 640064 213862 640116 213868
rect 639972 213512 640024 213518
rect 639972 213454 640024 213460
rect 639984 210202 640012 213454
rect 640260 210202 640288 231367
rect 650642 223136 650698 223145
rect 650642 223071 650698 223080
rect 643190 220416 643246 220425
rect 643190 220351 643246 220360
rect 641442 220144 641498 220153
rect 641442 220079 641498 220088
rect 641456 212770 641484 220079
rect 642086 217288 642142 217297
rect 642086 217223 642142 217232
rect 642100 213518 642128 217223
rect 643006 215928 643062 215937
rect 643006 215863 643062 215872
rect 642088 213512 642140 213518
rect 642088 213454 642140 213460
rect 641628 213240 641680 213246
rect 641628 213182 641680 213188
rect 642178 213208 642234 213217
rect 641444 212764 641496 212770
rect 641444 212706 641496 212712
rect 641640 210202 641668 213182
rect 642178 213143 642234 213152
rect 642192 210202 642220 213143
rect 643020 210202 643048 215863
rect 633820 210174 634156 210202
rect 634372 210174 634708 210202
rect 635260 210174 635596 210202
rect 636364 210174 636700 210202
rect 636916 210174 637252 210202
rect 638020 210174 638356 210202
rect 638572 210174 638908 210202
rect 639676 210174 640012 210202
rect 640228 210174 640288 210202
rect 641332 210174 641668 210202
rect 641884 210174 642220 210202
rect 642988 210174 643048 210202
rect 643204 210202 643232 220351
rect 647240 220108 647292 220114
rect 647240 220050 647292 220056
rect 644938 217560 644994 217569
rect 644938 217495 644994 217504
rect 644952 210202 644980 217495
rect 646594 216200 646650 216209
rect 646594 216135 646650 216144
rect 645492 213648 645544 213654
rect 645492 213590 645544 213596
rect 645504 210202 645532 213590
rect 646608 210202 646636 216135
rect 647252 214690 647280 220050
rect 649906 218648 649962 218657
rect 649906 218583 649962 218592
rect 647252 214662 647556 214690
rect 647146 214568 647202 214577
rect 647146 214503 647202 214512
rect 647160 210202 647188 214503
rect 643204 210174 643540 210202
rect 644644 210174 644980 210202
rect 645196 210174 645532 210202
rect 646300 210174 646636 210202
rect 646852 210174 647188 210202
rect 647528 210202 647556 214662
rect 648528 213920 648580 213926
rect 648528 213862 648580 213868
rect 648540 210202 648568 213862
rect 649920 210202 649948 218583
rect 650656 213926 650684 223071
rect 652022 222864 652078 222873
rect 652022 222799 652078 222808
rect 651286 214840 651342 214849
rect 651286 214775 651342 214784
rect 650644 213920 650696 213926
rect 650644 213862 650696 213868
rect 650460 213512 650512 213518
rect 650460 213454 650512 213460
rect 650472 210202 650500 213454
rect 651300 210202 651328 214775
rect 651840 213784 651892 213790
rect 651840 213726 651892 213732
rect 651852 210202 651880 213726
rect 652036 213382 652064 222799
rect 652024 213376 652076 213382
rect 652024 213318 652076 213324
rect 647528 210174 647956 210202
rect 648508 210174 648568 210202
rect 649612 210174 649948 210202
rect 650164 210174 650500 210202
rect 651268 210174 651328 210202
rect 651820 210174 651880 210202
rect 581736 209840 581788 209846
rect 581736 209782 581788 209788
rect 581552 208616 581604 208622
rect 581552 208558 581604 208564
rect 580448 207664 580500 207670
rect 580448 207606 580500 207612
rect 579526 207496 579582 207505
rect 579582 207454 579752 207482
rect 579526 207431 579582 207440
rect 579526 205864 579582 205873
rect 579526 205799 579528 205808
rect 579580 205799 579582 205808
rect 579528 205770 579580 205776
rect 579724 204270 579752 207454
rect 581000 205828 581052 205834
rect 581000 205770 581052 205776
rect 579712 204264 579764 204270
rect 579712 204206 579764 204212
rect 578330 203280 578386 203289
rect 578330 203215 578386 203224
rect 578344 202910 578372 203215
rect 578332 202904 578384 202910
rect 578332 202846 578384 202852
rect 580264 202904 580316 202910
rect 580264 202846 580316 202852
rect 578790 200832 578846 200841
rect 578790 200767 578846 200776
rect 578804 200190 578832 200767
rect 578792 200184 578844 200190
rect 578792 200126 578844 200132
rect 580276 200054 580304 202846
rect 581012 202842 581040 205770
rect 581000 202836 581052 202842
rect 581000 202778 581052 202784
rect 581564 200114 581592 208558
rect 581748 206310 581776 209782
rect 652220 209574 652248 298415
rect 658936 233889 658964 390526
rect 659120 360097 659148 510614
rect 660316 405657 660344 550598
rect 661868 523048 661920 523054
rect 661868 522990 661920 522996
rect 661684 456816 661736 456822
rect 661684 456758 661736 456764
rect 660302 405648 660358 405657
rect 660302 405583 660358 405592
rect 659106 360088 659162 360097
rect 659106 360023 659162 360032
rect 661696 313585 661724 456758
rect 661880 406337 661908 522990
rect 662064 492017 662092 590650
rect 664456 579737 664484 709310
rect 665836 626113 665864 749362
rect 666296 705537 666324 776999
rect 666466 742792 666522 742801
rect 666466 742727 666522 742736
rect 666282 705528 666338 705537
rect 666282 705463 666338 705472
rect 666480 665417 666508 742727
rect 667216 671129 667244 803150
rect 667754 786720 667810 786729
rect 667754 786655 667810 786664
rect 667570 743200 667626 743209
rect 667570 743135 667626 743144
rect 667202 671120 667258 671129
rect 667202 671055 667258 671064
rect 667584 665961 667612 743135
rect 667768 710841 667796 786655
rect 668228 752321 668256 868119
rect 668584 789404 668636 789410
rect 668584 789346 668636 789352
rect 668398 783864 668454 783873
rect 668398 783799 668454 783808
rect 668214 752312 668270 752321
rect 668214 752247 668270 752256
rect 668214 733408 668270 733417
rect 668214 733343 668270 733352
rect 667754 710832 667810 710841
rect 667754 710767 667810 710776
rect 667754 688936 667810 688945
rect 667754 688871 667810 688880
rect 667570 665952 667626 665961
rect 667570 665887 667626 665896
rect 666466 665408 666522 665417
rect 666466 665343 666522 665352
rect 667204 629332 667256 629338
rect 667204 629274 667256 629280
rect 665822 626104 665878 626113
rect 665822 626039 665878 626048
rect 664628 603152 664680 603158
rect 664628 603094 664680 603100
rect 666466 603120 666522 603129
rect 664442 579728 664498 579737
rect 664442 579663 664498 579672
rect 663248 496868 663300 496874
rect 663248 496810 663300 496816
rect 662050 492008 662106 492017
rect 662050 491943 662106 491952
rect 663064 416832 663116 416838
rect 663064 416774 663116 416780
rect 661866 406328 661922 406337
rect 661866 406263 661922 406272
rect 661868 364404 661920 364410
rect 661868 364346 661920 364352
rect 661682 313576 661738 313585
rect 661682 313511 661738 313520
rect 661880 234161 661908 364346
rect 663076 268161 663104 416774
rect 663260 358601 663288 496810
rect 664640 494057 664668 603094
rect 666466 603055 666522 603064
rect 665824 576904 665876 576910
rect 665824 576846 665876 576852
rect 665836 494737 665864 576846
rect 666480 529961 666508 603055
rect 667216 534177 667244 629274
rect 667768 621217 667796 688871
rect 668228 662561 668256 733343
rect 668412 708801 668440 783799
rect 668398 708792 668454 708801
rect 668398 708727 668454 708736
rect 668398 693288 668454 693297
rect 668398 693223 668454 693232
rect 668214 662552 668270 662561
rect 668214 662487 668270 662496
rect 668214 654256 668270 654265
rect 668214 654191 668270 654200
rect 667754 621208 667810 621217
rect 667754 621143 667810 621152
rect 668228 574161 668256 654191
rect 668412 620265 668440 693223
rect 668596 670585 668624 789346
rect 668768 775600 668820 775606
rect 668768 775542 668820 775548
rect 668780 734369 668808 775542
rect 668950 773800 669006 773809
rect 668950 773735 669006 773744
rect 668766 734360 668822 734369
rect 668766 734295 668822 734304
rect 668766 731504 668822 731513
rect 668766 731439 668822 731448
rect 668582 670576 668638 670585
rect 668582 670511 668638 670520
rect 668780 664601 668808 731439
rect 668964 710025 668992 773735
rect 669240 755177 669268 879135
rect 671158 872264 671214 872273
rect 671158 872199 671214 872208
rect 670606 867912 670662 867921
rect 670606 867847 670662 867856
rect 669778 864240 669834 864249
rect 669778 864175 669834 864184
rect 669594 789440 669650 789449
rect 669594 789375 669650 789384
rect 669226 755168 669282 755177
rect 669226 755103 669282 755112
rect 669410 741160 669466 741169
rect 669410 741095 669466 741104
rect 668950 710016 669006 710025
rect 668950 709951 669006 709960
rect 669226 705120 669282 705129
rect 669226 705055 669282 705064
rect 668766 664592 668822 664601
rect 668766 664527 668822 664536
rect 669042 648680 669098 648689
rect 669042 648615 669098 648624
rect 668584 643136 668636 643142
rect 668584 643078 668636 643084
rect 668398 620256 668454 620265
rect 668398 620191 668454 620200
rect 668398 601760 668454 601769
rect 668398 601695 668454 601704
rect 668214 574152 668270 574161
rect 668214 574087 668270 574096
rect 668214 564496 668270 564505
rect 668214 564431 668270 564440
rect 667202 534168 667258 534177
rect 667202 534103 667258 534112
rect 666466 529952 666522 529961
rect 666466 529887 666522 529896
rect 665822 494728 665878 494737
rect 665822 494663 665878 494672
rect 664626 494048 664682 494057
rect 664626 493983 664682 493992
rect 668228 485217 668256 564431
rect 668412 526561 668440 601695
rect 668596 535945 668624 643078
rect 668858 593736 668914 593745
rect 668858 593671 668914 593680
rect 668582 535936 668638 535945
rect 668582 535871 668638 535880
rect 668872 528601 668900 593671
rect 669056 573209 669084 648615
rect 669042 573200 669098 573209
rect 669042 573135 669098 573144
rect 669042 559192 669098 559201
rect 669042 559127 669098 559136
rect 668858 528592 668914 528601
rect 668858 528527 668914 528536
rect 668398 526552 668454 526561
rect 668398 526487 668454 526496
rect 668214 485208 668270 485217
rect 668214 485143 668270 485152
rect 667204 484424 667256 484430
rect 667204 484366 667256 484372
rect 665824 470620 665876 470626
rect 665824 470562 665876 470568
rect 664444 404388 664496 404394
rect 664444 404330 664496 404336
rect 663246 358592 663302 358601
rect 663246 358527 663302 358536
rect 664456 271153 664484 404330
rect 665836 315489 665864 470562
rect 667216 360913 667244 484366
rect 669056 483177 669084 559127
rect 669042 483168 669098 483177
rect 669042 483103 669098 483112
rect 669240 456521 669268 705055
rect 669424 663649 669452 741095
rect 669608 709617 669636 789375
rect 669792 750961 669820 864175
rect 669964 815652 670016 815658
rect 669964 815594 670016 815600
rect 669778 750952 669834 750961
rect 669778 750887 669834 750896
rect 669778 738576 669834 738585
rect 669778 738511 669834 738520
rect 669594 709608 669650 709617
rect 669594 709543 669650 709552
rect 669594 695192 669650 695201
rect 669594 695127 669650 695136
rect 669410 663640 669466 663649
rect 669410 663575 669466 663584
rect 669608 620673 669636 695127
rect 669792 666233 669820 738511
rect 669976 673169 670004 815594
rect 670330 783048 670386 783057
rect 670330 782983 670386 782992
rect 670146 780736 670202 780745
rect 670146 780671 670202 780680
rect 670160 710433 670188 780671
rect 670146 710424 670202 710433
rect 670146 710359 670202 710368
rect 670344 707577 670372 782983
rect 670620 751777 670648 867847
rect 670974 778696 671030 778705
rect 670974 778631 671030 778640
rect 670606 751768 670662 751777
rect 670606 751703 670662 751712
rect 670790 750136 670846 750145
rect 670790 750071 670846 750080
rect 670804 727977 670832 750071
rect 670988 736934 671016 778631
rect 671172 752593 671200 872199
rect 671356 763065 671384 895630
rect 671342 763056 671398 763065
rect 671342 762991 671398 763000
rect 671632 758554 671660 935711
rect 671816 758713 671844 936663
rect 672644 930134 672672 937479
rect 672828 930134 672856 937751
rect 673012 937666 673040 939766
rect 672920 937638 673040 937666
rect 672920 934538 672948 937638
rect 673104 934697 673132 962503
rect 673090 934688 673146 934697
rect 673090 934623 673146 934632
rect 672920 934510 673132 934538
rect 673104 930617 673132 934510
rect 673380 932657 673408 962775
rect 674194 957128 674250 957137
rect 674194 957063 674250 957072
rect 673366 932648 673422 932657
rect 673366 932583 673422 932592
rect 673090 930608 673146 930617
rect 673090 930543 673146 930552
rect 674208 930209 674236 957063
rect 674392 933065 674420 966039
rect 675036 963254 675064 966709
rect 675206 966104 675262 966113
rect 675262 966062 675418 966090
rect 675206 966039 675262 966048
rect 675772 965161 675800 965435
rect 675758 965152 675814 965161
rect 675758 965087 675814 965096
rect 675206 963656 675262 963665
rect 675206 963591 675262 963600
rect 675220 963254 675248 963591
rect 675404 963393 675432 963595
rect 675390 963384 675446 963393
rect 675390 963319 675446 963328
rect 674944 963226 675064 963254
rect 675128 963226 675248 963254
rect 674944 962577 674972 963226
rect 674930 962568 674986 962577
rect 674930 962503 674986 962512
rect 674654 962160 674710 962169
rect 674654 962095 674710 962104
rect 674378 933056 674434 933065
rect 674378 932991 674434 933000
rect 674668 932249 674696 962095
rect 675128 961769 675156 963226
rect 675496 962849 675524 963016
rect 675482 962840 675538 962849
rect 675482 962775 675538 962784
rect 675404 962169 675432 962404
rect 675390 962160 675446 962169
rect 675390 962095 675446 962104
rect 675128 961741 675418 961769
rect 675206 959304 675262 959313
rect 675262 959262 675418 959290
rect 675206 959239 675262 959248
rect 675114 958760 675170 958769
rect 675170 958718 675418 958746
rect 675114 958695 675170 958704
rect 675772 957817 675800 958052
rect 675298 957808 675354 957817
rect 675298 957743 675354 957752
rect 675758 957808 675814 957817
rect 675758 957743 675814 957752
rect 675312 955482 675340 957743
rect 675496 957137 675524 957440
rect 675482 957128 675538 957137
rect 675482 957063 675538 957072
rect 675758 956448 675814 956457
rect 675758 956383 675814 956392
rect 675772 956216 675800 956383
rect 675312 955454 675524 955482
rect 675496 955060 675524 955454
rect 675022 954544 675078 954553
rect 675022 954479 675078 954488
rect 674838 953456 674894 953465
rect 674838 953391 674894 953400
rect 674654 932240 674710 932249
rect 674654 932175 674710 932184
rect 674194 930200 674250 930209
rect 674194 930135 674250 930144
rect 672184 930106 672672 930134
rect 672736 930106 672856 930134
rect 671986 928296 672042 928305
rect 671986 928231 672042 928240
rect 671802 758704 671858 758713
rect 671802 758639 671858 758648
rect 671632 758526 671752 758554
rect 671526 758296 671582 758305
rect 671526 758231 671582 758240
rect 671158 752584 671214 752593
rect 671158 752519 671214 752528
rect 671158 737080 671214 737089
rect 671158 737015 671214 737024
rect 670896 736906 671016 736934
rect 670896 728090 670924 736906
rect 671172 734210 671200 737015
rect 671344 735616 671396 735622
rect 671344 735558 671396 735564
rect 671172 734182 671292 734210
rect 671066 730552 671122 730561
rect 671066 730487 671122 730496
rect 670896 728062 671016 728090
rect 670790 727968 670846 727977
rect 670790 727903 670846 727912
rect 670790 712464 670846 712473
rect 670790 712399 670846 712408
rect 670330 707568 670386 707577
rect 670330 707503 670386 707512
rect 670606 699816 670662 699825
rect 670606 699751 670662 699760
rect 670330 687440 670386 687449
rect 670330 687375 670386 687384
rect 669962 673160 670018 673169
rect 669962 673095 670018 673104
rect 669778 666224 669834 666233
rect 669778 666159 669834 666168
rect 670148 656940 670200 656946
rect 670148 656882 670200 656888
rect 669962 648136 670018 648145
rect 669962 648071 670018 648080
rect 669778 645416 669834 645425
rect 669778 645351 669834 645360
rect 669594 620664 669650 620673
rect 669594 620599 669650 620608
rect 669792 574977 669820 645351
rect 669778 574968 669834 574977
rect 669778 574903 669834 574912
rect 669976 571713 670004 648071
rect 669962 571704 670018 571713
rect 669962 571639 670018 571648
rect 669410 570888 669466 570897
rect 669410 570823 669466 570832
rect 669424 500993 669452 570823
rect 669594 556200 669650 556209
rect 669594 556135 669650 556144
rect 669410 500984 669466 500993
rect 669410 500919 669466 500928
rect 669608 482361 669636 556135
rect 669778 553888 669834 553897
rect 669778 553823 669834 553832
rect 669792 483585 669820 553823
rect 670160 537849 670188 656882
rect 670344 618225 670372 687375
rect 670620 619449 670648 699751
rect 670804 667729 670832 712399
rect 670988 706761 671016 728062
rect 671080 727274 671108 730487
rect 671080 727246 671200 727274
rect 670974 706752 671030 706761
rect 670974 706687 671030 706696
rect 670974 685536 671030 685545
rect 670974 685471 671030 685480
rect 670790 667720 670846 667729
rect 670790 667655 670846 667664
rect 670988 666482 671016 685471
rect 670896 666454 671016 666482
rect 670896 661858 670924 666454
rect 671172 666346 671200 727246
rect 671080 666318 671200 666346
rect 671080 666262 671108 666318
rect 671068 666256 671120 666262
rect 671068 666198 671120 666204
rect 671264 666074 671292 734182
rect 671172 666046 671292 666074
rect 671172 662425 671200 666046
rect 671158 662416 671214 662425
rect 671158 662351 671214 662360
rect 670896 661830 671016 661858
rect 670988 627162 671016 661830
rect 671158 640520 671214 640529
rect 671158 640455 671214 640464
rect 670976 627156 671028 627162
rect 670976 627098 671028 627104
rect 670790 623928 670846 623937
rect 670790 623863 670846 623872
rect 670606 619440 670662 619449
rect 670606 619375 670662 619384
rect 670330 618216 670386 618225
rect 670330 618151 670386 618160
rect 670606 608016 670662 608025
rect 670606 607951 670662 607960
rect 670330 598088 670386 598097
rect 670330 598023 670386 598032
rect 670146 537840 670202 537849
rect 670146 537775 670202 537784
rect 669964 536852 670016 536858
rect 669964 536794 670016 536800
rect 669778 483576 669834 483585
rect 669778 483511 669834 483520
rect 669594 482352 669650 482361
rect 669594 482287 669650 482296
rect 669226 456512 669282 456521
rect 669226 456447 669282 456456
rect 668584 444440 668636 444446
rect 668584 444382 668636 444388
rect 667202 360904 667258 360913
rect 667202 360839 667258 360848
rect 667388 350600 667440 350606
rect 667388 350542 667440 350548
rect 667020 324352 667072 324358
rect 667020 324294 667072 324300
rect 665822 315480 665878 315489
rect 665822 315415 665878 315424
rect 664442 271144 664498 271153
rect 664442 271079 664498 271088
rect 663062 268152 663118 268161
rect 663062 268087 663118 268096
rect 661866 234152 661922 234161
rect 661866 234087 661922 234096
rect 658922 233880 658978 233889
rect 658922 233815 658978 233824
rect 662328 232416 662380 232422
rect 662328 232358 662380 232364
rect 661682 230344 661738 230353
rect 661682 230279 661738 230288
rect 660946 229800 661002 229809
rect 660946 229735 661002 229744
rect 652758 226400 652814 226409
rect 652758 226335 652814 226344
rect 652772 220114 652800 226335
rect 658922 225584 658978 225593
rect 658922 225519 658978 225528
rect 655518 225312 655574 225321
rect 655518 225247 655574 225256
rect 654782 225040 654838 225049
rect 654782 224975 654838 224984
rect 654232 221468 654284 221474
rect 654232 221410 654284 221416
rect 653034 220688 653090 220697
rect 653034 220623 653090 220632
rect 652760 220108 652812 220114
rect 652760 220050 652812 220056
rect 652852 215960 652904 215966
rect 652852 215902 652904 215908
rect 652864 210202 652892 215902
rect 653048 210202 653076 220623
rect 654046 216472 654102 216481
rect 654046 216407 654102 216416
rect 654060 216322 654088 216407
rect 654060 216294 654180 216322
rect 654152 213058 654180 216294
rect 654060 213042 654180 213058
rect 654048 213036 654180 213042
rect 654100 213030 654180 213036
rect 654048 212978 654100 212984
rect 654244 210202 654272 221410
rect 654796 215966 654824 224975
rect 655532 221474 655560 225247
rect 656622 223952 656678 223961
rect 656622 223887 656678 223896
rect 655704 221604 655756 221610
rect 655704 221546 655756 221552
rect 655520 221468 655572 221474
rect 655520 221410 655572 221416
rect 654784 215960 654836 215966
rect 654784 215902 654836 215908
rect 655716 213926 655744 221546
rect 655704 213920 655756 213926
rect 655704 213862 655756 213868
rect 654784 213036 654836 213042
rect 654784 212978 654836 212984
rect 654796 210202 654824 212978
rect 656636 210202 656664 223887
rect 658186 223680 658242 223689
rect 658186 223615 658242 223624
rect 658002 221504 658058 221513
rect 658002 221439 658058 221448
rect 656808 213920 656860 213926
rect 656808 213862 656860 213868
rect 656820 210202 656848 213862
rect 658016 213790 658044 221439
rect 658004 213784 658056 213790
rect 658004 213726 658056 213732
rect 658200 210202 658228 223615
rect 658740 214192 658792 214198
rect 658740 214134 658792 214140
rect 658752 210202 658780 214134
rect 658936 213246 658964 225519
rect 659290 224496 659346 224505
rect 659290 224431 659346 224440
rect 659304 221610 659332 224431
rect 659474 221776 659530 221785
rect 659474 221711 659530 221720
rect 659292 221604 659344 221610
rect 659292 221546 659344 221552
rect 659488 213654 659516 221711
rect 659658 215112 659714 215121
rect 659658 215047 659714 215056
rect 659476 213648 659528 213654
rect 659476 213590 659528 213596
rect 658924 213240 658976 213246
rect 658924 213182 658976 213188
rect 659672 212534 659700 215047
rect 660960 213926 660988 229735
rect 661696 214198 661724 230279
rect 662340 215294 662368 232358
rect 665088 232212 665140 232218
rect 665088 232154 665140 232160
rect 663062 231704 663118 231713
rect 663062 231639 663118 231648
rect 663076 215294 663104 231639
rect 664442 230888 664498 230897
rect 664442 230823 664498 230832
rect 663706 230616 663762 230625
rect 663706 230551 663762 230560
rect 662248 215266 662368 215294
rect 662984 215266 663104 215294
rect 661684 214192 661736 214198
rect 661684 214134 661736 214140
rect 662052 214056 662104 214062
rect 662052 213998 662104 214004
rect 660396 213920 660448 213926
rect 660396 213862 660448 213868
rect 660948 213920 661000 213926
rect 660948 213862 661000 213868
rect 652864 210174 652924 210202
rect 653048 210174 653476 210202
rect 654244 210174 654580 210202
rect 654796 210174 655132 210202
rect 656236 210174 656664 210202
rect 656788 210174 656848 210202
rect 657892 210174 658228 210202
rect 658444 210174 658780 210202
rect 659488 212506 659700 212534
rect 659488 210202 659516 212506
rect 660408 210202 660436 213862
rect 660948 213784 661000 213790
rect 660948 213726 661000 213732
rect 660960 210202 660988 213726
rect 661498 213480 661554 213489
rect 661498 213415 661554 213424
rect 661512 210202 661540 213415
rect 662064 210202 662092 213998
rect 659488 210174 659548 210202
rect 660100 210174 660436 210202
rect 660652 210174 660988 210202
rect 661204 210174 661540 210202
rect 661756 210174 662092 210202
rect 662248 210202 662276 215266
rect 662984 213790 663012 215266
rect 662972 213784 663024 213790
rect 662972 213726 663024 213732
rect 663156 213784 663208 213790
rect 663156 213726 663208 213732
rect 663168 210202 663196 213726
rect 663720 210202 663748 230551
rect 664258 220416 664314 220425
rect 664258 220351 664314 220360
rect 664272 219745 664300 220351
rect 664258 219736 664314 219745
rect 664258 219671 664314 219680
rect 664258 216744 664314 216753
rect 664258 216679 664314 216688
rect 664272 216209 664300 216679
rect 664258 216200 664314 216209
rect 664258 216135 664314 216144
rect 664456 213790 664484 230823
rect 664444 213784 664496 213790
rect 664444 213726 664496 213732
rect 664810 213752 664866 213761
rect 664810 213687 664866 213696
rect 664260 213036 664312 213042
rect 664260 212978 664312 212984
rect 664272 210202 664300 212978
rect 664824 210202 664852 213687
rect 665100 213042 665128 232154
rect 665822 231160 665878 231169
rect 665822 231095 665878 231104
rect 665836 214062 665864 231095
rect 666836 229696 666888 229702
rect 666836 229638 666888 229644
rect 666652 226500 666704 226506
rect 666652 226442 666704 226448
rect 666008 226092 666060 226098
rect 666008 226034 666060 226040
rect 665824 214056 665876 214062
rect 665824 213998 665876 214004
rect 666020 213382 666048 226034
rect 666664 223281 666692 226442
rect 666650 223272 666706 223281
rect 666650 223207 666706 223216
rect 666848 222873 666876 229638
rect 666834 222864 666890 222873
rect 666834 222799 666890 222808
rect 666650 221096 666706 221105
rect 666650 221031 666706 221040
rect 666008 213376 666060 213382
rect 666008 213318 666060 213324
rect 665088 213036 665140 213042
rect 665088 212978 665140 212984
rect 662248 210174 662308 210202
rect 662860 210174 663196 210202
rect 663412 210174 663748 210202
rect 663964 210174 664300 210202
rect 664516 210174 664852 210202
rect 632152 209568 632204 209574
rect 652208 209568 652260 209574
rect 632204 209516 632500 209522
rect 632152 209510 632500 209516
rect 652208 209510 652260 209516
rect 632164 209494 632500 209510
rect 589464 208344 589516 208350
rect 589464 208286 589516 208292
rect 589476 208049 589504 208286
rect 589462 208040 589518 208049
rect 589462 207975 589518 207984
rect 589464 207664 589516 207670
rect 589464 207606 589516 207612
rect 589476 206417 589504 207606
rect 589462 206408 589518 206417
rect 589462 206343 589518 206352
rect 581736 206304 581788 206310
rect 581736 206246 581788 206252
rect 589648 206304 589700 206310
rect 589648 206246 589700 206252
rect 589660 204785 589688 206246
rect 589646 204776 589702 204785
rect 589646 204711 589702 204720
rect 589464 204264 589516 204270
rect 589464 204206 589516 204212
rect 589476 203153 589504 204206
rect 589462 203144 589518 203153
rect 589462 203079 589518 203088
rect 589464 202836 589516 202842
rect 589464 202778 589516 202784
rect 589476 201521 589504 202778
rect 589462 201512 589518 201521
rect 589462 201447 589518 201456
rect 590384 200184 590436 200190
rect 590384 200126 590436 200132
rect 581564 200086 581684 200114
rect 580264 200048 580316 200054
rect 580264 199990 580316 199996
rect 579526 198928 579582 198937
rect 579526 198863 579582 198872
rect 579540 198762 579568 198863
rect 579528 198756 579580 198762
rect 579528 198698 579580 198704
rect 578514 196480 578570 196489
rect 578514 196415 578570 196424
rect 578528 196042 578556 196415
rect 578516 196036 578568 196042
rect 578516 195978 578568 195984
rect 579526 194984 579582 194993
rect 579526 194919 579582 194928
rect 579540 194614 579568 194919
rect 579528 194608 579580 194614
rect 579528 194550 579580 194556
rect 579526 192264 579582 192273
rect 579526 192199 579582 192208
rect 579540 191894 579568 192199
rect 579528 191888 579580 191894
rect 579528 191830 579580 191836
rect 579526 190768 579582 190777
rect 579526 190703 579582 190712
rect 579540 190534 579568 190703
rect 579528 190528 579580 190534
rect 579528 190470 579580 190476
rect 579526 188048 579582 188057
rect 579526 187983 579582 187992
rect 579540 187746 579568 187983
rect 579528 187740 579580 187746
rect 579528 187682 579580 187688
rect 579528 186312 579580 186318
rect 579526 186280 579528 186289
rect 579580 186280 579582 186289
rect 579526 186215 579582 186224
rect 579528 184884 579580 184890
rect 579528 184826 579580 184832
rect 579540 184385 579568 184826
rect 579526 184376 579582 184385
rect 579526 184311 579582 184320
rect 579528 182164 579580 182170
rect 579528 182106 579580 182112
rect 579540 181937 579568 182106
rect 579526 181928 579582 181937
rect 579526 181863 579582 181872
rect 578792 180804 578844 180810
rect 578792 180746 578844 180752
rect 578804 180169 578832 180746
rect 578790 180160 578846 180169
rect 578790 180095 578846 180104
rect 578792 178084 578844 178090
rect 578792 178026 578844 178032
rect 578804 175137 578832 178026
rect 579528 177948 579580 177954
rect 579528 177890 579580 177896
rect 579540 177721 579568 177890
rect 579526 177712 579582 177721
rect 579526 177647 579582 177656
rect 579988 175296 580040 175302
rect 579988 175238 580040 175244
rect 578790 175128 578846 175137
rect 578790 175063 578846 175072
rect 578424 174548 578476 174554
rect 578424 174490 578476 174496
rect 578436 173505 578464 174490
rect 578422 173496 578478 173505
rect 578422 173431 578478 173440
rect 580000 172922 580028 175238
rect 578240 172916 578292 172922
rect 578240 172858 578292 172864
rect 579988 172916 580040 172922
rect 579988 172858 580040 172864
rect 578252 171057 578280 172858
rect 580908 172576 580960 172582
rect 580908 172518 580960 172524
rect 579896 171148 579948 171154
rect 579632 171106 579896 171134
rect 578238 171048 578294 171057
rect 578238 170983 578294 170992
rect 578700 169788 578752 169794
rect 578700 169730 578752 169736
rect 578712 169289 578740 169730
rect 578698 169280 578754 169289
rect 578698 169215 578754 169224
rect 579632 168586 579660 171106
rect 579896 171090 579948 171096
rect 580920 169794 580948 172518
rect 580908 169788 580960 169794
rect 580908 169730 580960 169736
rect 579540 168558 579660 168586
rect 579540 166977 579568 168558
rect 579712 168428 579764 168434
rect 579712 168370 579764 168376
rect 579526 166968 579582 166977
rect 579526 166903 579582 166912
rect 578884 165572 578936 165578
rect 578884 165514 578936 165520
rect 578896 164529 578924 165514
rect 578882 164520 578938 164529
rect 578882 164455 578938 164464
rect 579724 162874 579752 168370
rect 579540 162846 579752 162874
rect 580908 162920 580960 162926
rect 580908 162862 580960 162868
rect 579540 162761 579568 162846
rect 579526 162752 579582 162761
rect 578424 162716 578476 162722
rect 579526 162687 579582 162696
rect 578424 162658 578476 162664
rect 578240 162580 578292 162586
rect 578240 162522 578292 162528
rect 578252 159905 578280 162522
rect 578238 159896 578294 159905
rect 578238 159831 578294 159840
rect 578436 158409 578464 162658
rect 580540 161492 580592 161498
rect 580540 161434 580592 161440
rect 578884 158772 578936 158778
rect 578884 158714 578936 158720
rect 578422 158400 578478 158409
rect 578422 158335 578478 158344
rect 578896 155961 578924 158714
rect 578882 155952 578938 155961
rect 578882 155887 578938 155896
rect 580552 154698 580580 161434
rect 580724 160132 580776 160138
rect 580724 160074 580776 160080
rect 578332 154692 578384 154698
rect 578332 154634 578384 154640
rect 580540 154692 580592 154698
rect 580540 154634 580592 154640
rect 578344 154057 578372 154634
rect 578330 154048 578386 154057
rect 578330 153983 578386 153992
rect 580736 152794 580764 160074
rect 580920 158778 580948 162862
rect 580908 158772 580960 158778
rect 580908 158714 580960 158720
rect 578240 152788 578292 152794
rect 578240 152730 578292 152736
rect 580724 152788 580776 152794
rect 580724 152730 580776 152736
rect 578252 151745 578280 152730
rect 580448 151836 580500 151842
rect 580448 151778 580500 151784
rect 578238 151736 578294 151745
rect 578238 151671 578294 151680
rect 578332 151088 578384 151094
rect 578332 151030 578384 151036
rect 578344 149705 578372 151030
rect 578330 149696 578386 149705
rect 578330 149631 578386 149640
rect 578884 149116 578936 149122
rect 578884 149058 578936 149064
rect 578700 147280 578752 147286
rect 578698 147248 578700 147257
rect 578752 147248 578754 147257
rect 578698 147183 578754 147192
rect 578608 140752 578660 140758
rect 578608 140694 578660 140700
rect 578620 140593 578648 140694
rect 578606 140584 578662 140593
rect 578606 140519 578662 140528
rect 578608 139324 578660 139330
rect 578608 139266 578660 139272
rect 578620 138825 578648 139266
rect 578606 138816 578662 138825
rect 578606 138751 578662 138760
rect 578700 137284 578752 137290
rect 578700 137226 578752 137232
rect 578712 134473 578740 137226
rect 578896 136649 578924 149058
rect 579252 144696 579304 144702
rect 579250 144664 579252 144673
rect 579304 144664 579306 144673
rect 579250 144599 579306 144608
rect 579528 143472 579580 143478
rect 579528 143414 579580 143420
rect 579540 143041 579568 143414
rect 579526 143032 579582 143041
rect 579526 142967 579582 142976
rect 580460 140758 580488 151778
rect 580448 140752 580500 140758
rect 580448 140694 580500 140700
rect 580264 139460 580316 139466
rect 580264 139402 580316 139408
rect 579068 137148 579120 137154
rect 579068 137090 579120 137096
rect 578882 136640 578938 136649
rect 578882 136575 578938 136584
rect 578698 134464 578754 134473
rect 578698 134399 578754 134408
rect 579080 132297 579108 137090
rect 579066 132288 579122 132297
rect 579066 132223 579122 132232
rect 578884 131300 578936 131306
rect 578884 131242 578936 131248
rect 578332 124160 578384 124166
rect 578332 124102 578384 124108
rect 578344 123593 578372 124102
rect 578330 123584 578386 123593
rect 578330 123519 578386 123528
rect 578700 118584 578752 118590
rect 578700 118526 578752 118532
rect 578712 118425 578740 118526
rect 578698 118416 578754 118425
rect 578698 118351 578754 118360
rect 578700 117224 578752 117230
rect 578700 117166 578752 117172
rect 578712 116929 578740 117166
rect 578698 116920 578754 116929
rect 578698 116855 578754 116864
rect 578896 110401 578924 131242
rect 579068 131164 579120 131170
rect 579068 131106 579120 131112
rect 579080 129713 579108 131106
rect 579066 129704 579122 129713
rect 579066 129639 579122 129648
rect 579160 128308 579212 128314
rect 579160 128250 579212 128256
rect 579172 127809 579200 128250
rect 579158 127800 579214 127809
rect 579158 127735 579214 127744
rect 579068 126268 579120 126274
rect 579068 126210 579120 126216
rect 579080 113174 579108 126210
rect 579528 125384 579580 125390
rect 579526 125352 579528 125361
rect 579580 125352 579582 125361
rect 579526 125287 579582 125296
rect 580276 124166 580304 139402
rect 580632 131776 580684 131782
rect 580632 131718 580684 131724
rect 580264 124160 580316 124166
rect 580264 124102 580316 124108
rect 580448 122868 580500 122874
rect 580448 122810 580500 122816
rect 579528 121440 579580 121446
rect 579528 121382 579580 121388
rect 579540 121145 579568 121382
rect 579526 121136 579582 121145
rect 579526 121071 579582 121080
rect 579252 114504 579304 114510
rect 579250 114472 579252 114481
rect 579304 114472 579306 114481
rect 579250 114407 579306 114416
rect 578988 113146 579108 113174
rect 578988 110514 579016 113146
rect 579160 113076 579212 113082
rect 579160 113018 579212 113024
rect 579172 112577 579200 113018
rect 579158 112568 579214 112577
rect 579158 112503 579214 112512
rect 578988 110486 579108 110514
rect 578882 110392 578938 110401
rect 578882 110327 578938 110336
rect 578884 108996 578936 109002
rect 578884 108938 578936 108944
rect 578896 108361 578924 108938
rect 578882 108352 578938 108361
rect 578882 108287 578938 108296
rect 578884 107636 578936 107642
rect 578884 107578 578936 107584
rect 578332 103352 578384 103358
rect 578330 103320 578332 103329
rect 578384 103320 578386 103329
rect 578330 103255 578386 103264
rect 578516 102128 578568 102134
rect 578516 102070 578568 102076
rect 578528 101697 578556 102070
rect 578514 101688 578570 101697
rect 578514 101623 578570 101632
rect 577504 99136 577556 99142
rect 577504 99078 577556 99084
rect 578332 97980 578384 97986
rect 578332 97922 578384 97928
rect 578344 97481 578372 97922
rect 578330 97472 578386 97481
rect 578330 97407 578386 97416
rect 577504 95940 577556 95946
rect 577504 95882 577556 95888
rect 576860 57248 576912 57254
rect 576860 57190 576912 57196
rect 574560 56160 574612 56166
rect 574560 56102 574612 56108
rect 574572 53990 574600 56102
rect 574928 56024 574980 56030
rect 574928 55966 574980 55972
rect 574744 55888 574796 55894
rect 574744 55830 574796 55836
rect 574756 54126 574784 55830
rect 574744 54120 574796 54126
rect 574744 54062 574796 54068
rect 574560 53984 574612 53990
rect 574560 53926 574612 53932
rect 574940 53854 574968 55966
rect 576872 54233 576900 57190
rect 577516 55049 577544 95882
rect 578332 86964 578384 86970
rect 578332 86906 578384 86912
rect 578344 86465 578372 86906
rect 578330 86456 578386 86465
rect 578330 86391 578386 86400
rect 578424 85468 578476 85474
rect 578424 85410 578476 85416
rect 578436 77897 578464 85410
rect 578896 80073 578924 107578
rect 579080 105913 579108 110486
rect 579066 105904 579122 105913
rect 579066 105839 579122 105848
rect 580264 104916 580316 104922
rect 580264 104858 580316 104864
rect 579252 99272 579304 99278
rect 579250 99240 579252 99249
rect 579304 99240 579306 99249
rect 579250 99175 579306 99184
rect 579436 95056 579488 95062
rect 579434 95024 579436 95033
rect 579488 95024 579490 95033
rect 579434 94959 579490 94968
rect 579528 93424 579580 93430
rect 579528 93366 579580 93372
rect 579540 93129 579568 93366
rect 579526 93120 579582 93129
rect 579526 93055 579582 93064
rect 579344 91996 579396 92002
rect 579344 91938 579396 91944
rect 579356 90953 579384 91938
rect 579528 91792 579580 91798
rect 579528 91734 579580 91740
rect 579342 90944 579398 90953
rect 579342 90879 579398 90888
rect 579540 88097 579568 91734
rect 579526 88088 579582 88097
rect 579526 88023 579582 88032
rect 579528 84040 579580 84046
rect 579526 84008 579528 84017
rect 579580 84008 579582 84017
rect 579526 83943 579582 83952
rect 579436 82476 579488 82482
rect 579436 82418 579488 82424
rect 579448 82249 579476 82418
rect 579434 82240 579490 82249
rect 579434 82175 579490 82184
rect 578882 80064 578938 80073
rect 578882 79999 578938 80008
rect 579068 79348 579120 79354
rect 579068 79290 579120 79296
rect 578422 77888 578478 77897
rect 578422 77823 578478 77832
rect 578332 77716 578384 77722
rect 578332 77658 578384 77664
rect 578344 75721 578372 77658
rect 578330 75712 578386 75721
rect 578330 75647 578386 75656
rect 578884 75200 578936 75206
rect 578884 75142 578936 75148
rect 578516 62076 578568 62082
rect 578516 62018 578568 62024
rect 578528 61849 578556 62018
rect 578514 61840 578570 61849
rect 578514 61775 578570 61784
rect 578896 60489 578924 75142
rect 578882 60480 578938 60489
rect 578882 60415 578938 60424
rect 579080 55078 579108 79290
rect 580276 77722 580304 104858
rect 580460 102134 580488 122810
rect 580644 117230 580672 131718
rect 580632 117224 580684 117230
rect 580632 117166 580684 117172
rect 581656 114510 581684 200086
rect 589464 200048 589516 200054
rect 589464 199990 589516 199996
rect 589476 199889 589504 199990
rect 589462 199880 589518 199889
rect 589462 199815 589518 199824
rect 589464 198756 589516 198762
rect 589464 198698 589516 198704
rect 589476 196625 589504 198698
rect 590396 198257 590424 200126
rect 590382 198248 590438 198257
rect 590382 198183 590438 198192
rect 589462 196616 589518 196625
rect 589462 196551 589518 196560
rect 589280 196036 589332 196042
rect 589280 195978 589332 195984
rect 589292 194993 589320 195978
rect 589278 194984 589334 194993
rect 589278 194919 589334 194928
rect 589464 194608 589516 194614
rect 589464 194550 589516 194556
rect 589476 193361 589504 194550
rect 589462 193352 589518 193361
rect 589462 193287 589518 193296
rect 589464 191888 589516 191894
rect 589464 191830 589516 191836
rect 589476 191729 589504 191830
rect 589462 191720 589518 191729
rect 589462 191655 589518 191664
rect 590568 190528 590620 190534
rect 590568 190470 590620 190476
rect 590580 190097 590608 190470
rect 590566 190088 590622 190097
rect 590566 190023 590622 190032
rect 589646 188456 589702 188465
rect 589646 188391 589702 188400
rect 589464 187740 589516 187746
rect 589464 187682 589516 187688
rect 589476 186833 589504 187682
rect 589462 186824 589518 186833
rect 589462 186759 589518 186768
rect 589660 186318 589688 188391
rect 589648 186312 589700 186318
rect 589648 186254 589700 186260
rect 589462 185192 589518 185201
rect 589462 185127 589518 185136
rect 589476 184890 589504 185127
rect 589464 184884 589516 184890
rect 589464 184826 589516 184832
rect 589462 183560 589518 183569
rect 589462 183495 589518 183504
rect 589476 182170 589504 183495
rect 589464 182164 589516 182170
rect 589464 182106 589516 182112
rect 590566 181928 590622 181937
rect 590566 181863 590622 181872
rect 590580 180810 590608 181863
rect 590568 180804 590620 180810
rect 590568 180746 590620 180752
rect 589646 180296 589702 180305
rect 589646 180231 589702 180240
rect 589462 178664 589518 178673
rect 589462 178599 589518 178608
rect 589476 178090 589504 178599
rect 589464 178084 589516 178090
rect 589464 178026 589516 178032
rect 589660 177954 589688 180231
rect 589648 177948 589700 177954
rect 589648 177890 589700 177896
rect 589646 177032 589702 177041
rect 589646 176967 589702 176976
rect 589462 175400 589518 175409
rect 589462 175335 589464 175344
rect 589516 175335 589518 175344
rect 589464 175306 589516 175312
rect 589660 174554 589688 176967
rect 666664 176497 666692 221031
rect 666836 209092 666888 209098
rect 666836 209034 666888 209040
rect 666650 176488 666706 176497
rect 666650 176423 666706 176432
rect 589648 174548 589700 174554
rect 589648 174490 589700 174496
rect 589462 173768 589518 173777
rect 589462 173703 589518 173712
rect 589476 172582 589504 173703
rect 589464 172576 589516 172582
rect 589464 172518 589516 172524
rect 589462 172136 589518 172145
rect 589462 172071 589518 172080
rect 589476 171154 589504 172071
rect 589464 171148 589516 171154
rect 589464 171090 589516 171096
rect 589462 170504 589518 170513
rect 589462 170439 589518 170448
rect 589476 169794 589504 170439
rect 582380 169788 582432 169794
rect 582380 169730 582432 169736
rect 589464 169788 589516 169794
rect 589464 169730 589516 169736
rect 582392 165578 582420 169730
rect 589462 168872 589518 168881
rect 589462 168807 589518 168816
rect 589476 168434 589504 168807
rect 589464 168428 589516 168434
rect 589464 168370 589516 168376
rect 589462 167240 589518 167249
rect 589462 167175 589518 167184
rect 589476 167074 589504 167175
rect 583760 167068 583812 167074
rect 583760 167010 583812 167016
rect 589464 167068 589516 167074
rect 589464 167010 589516 167016
rect 582380 165572 582432 165578
rect 582380 165514 582432 165520
rect 582472 164280 582524 164286
rect 582472 164222 582524 164228
rect 582484 162722 582512 164222
rect 582472 162716 582524 162722
rect 582472 162658 582524 162664
rect 583772 162586 583800 167010
rect 589462 165608 589518 165617
rect 589462 165543 589518 165552
rect 589476 164286 589504 165543
rect 589464 164280 589516 164286
rect 589464 164222 589516 164228
rect 589462 163976 589518 163985
rect 589462 163911 589518 163920
rect 589476 162926 589504 163911
rect 589464 162920 589516 162926
rect 589464 162862 589516 162868
rect 583760 162580 583812 162586
rect 583760 162522 583812 162528
rect 589462 162344 589518 162353
rect 589462 162279 589518 162288
rect 589476 161498 589504 162279
rect 589464 161492 589516 161498
rect 589464 161434 589516 161440
rect 589462 160712 589518 160721
rect 589462 160647 589518 160656
rect 589476 160138 589504 160647
rect 589464 160132 589516 160138
rect 589464 160074 589516 160080
rect 589830 159080 589886 159089
rect 589830 159015 589886 159024
rect 589844 158778 589872 159015
rect 587164 158772 587216 158778
rect 587164 158714 587216 158720
rect 589832 158772 589884 158778
rect 589832 158714 589884 158720
rect 585784 157412 585836 157418
rect 585784 157354 585836 157360
rect 584404 154624 584456 154630
rect 584404 154566 584456 154572
rect 583024 153264 583076 153270
rect 583024 153206 583076 153212
rect 583036 143478 583064 153206
rect 584416 144702 584444 154566
rect 585796 147286 585824 157354
rect 587176 151094 587204 158714
rect 589462 157448 589518 157457
rect 589462 157383 589464 157392
rect 589516 157383 589518 157392
rect 589464 157354 589516 157360
rect 589462 155816 589518 155825
rect 589462 155751 589518 155760
rect 589476 154630 589504 155751
rect 589464 154624 589516 154630
rect 589464 154566 589516 154572
rect 589462 154184 589518 154193
rect 589462 154119 589518 154128
rect 589476 153270 589504 154119
rect 589464 153264 589516 153270
rect 589464 153206 589516 153212
rect 589462 152552 589518 152561
rect 589462 152487 589518 152496
rect 589476 151842 589504 152487
rect 589464 151836 589516 151842
rect 589464 151778 589516 151784
rect 587164 151088 587216 151094
rect 587164 151030 587216 151036
rect 590014 150920 590070 150929
rect 590014 150855 590070 150864
rect 589462 149288 589518 149297
rect 589462 149223 589518 149232
rect 589476 149122 589504 149223
rect 589464 149116 589516 149122
rect 589464 149058 589516 149064
rect 588542 147656 588598 147665
rect 588542 147591 588598 147600
rect 585784 147280 585836 147286
rect 585784 147222 585836 147228
rect 585968 144968 586020 144974
rect 585968 144910 586020 144916
rect 584404 144696 584456 144702
rect 584404 144638 584456 144644
rect 584588 143608 584640 143614
rect 584588 143550 584640 143556
rect 583024 143472 583076 143478
rect 583024 143414 583076 143420
rect 583024 140820 583076 140826
rect 583024 140762 583076 140768
rect 583036 125390 583064 140762
rect 584404 135312 584456 135318
rect 584404 135254 584456 135260
rect 583024 125384 583076 125390
rect 583024 125326 583076 125332
rect 583208 124908 583260 124914
rect 583208 124850 583260 124856
rect 581828 122120 581880 122126
rect 581828 122062 581880 122068
rect 581644 114504 581696 114510
rect 581644 114446 581696 114452
rect 581644 111104 581696 111110
rect 581644 111046 581696 111052
rect 580448 102128 580500 102134
rect 580448 102070 580500 102076
rect 580448 100020 580500 100026
rect 580448 99962 580500 99968
rect 580460 86970 580488 99962
rect 581656 99278 581684 111046
rect 581840 109002 581868 122062
rect 583024 109744 583076 109750
rect 583024 109686 583076 109692
rect 581828 108996 581880 109002
rect 581828 108938 581880 108944
rect 581828 106344 581880 106350
rect 581828 106286 581880 106292
rect 581644 99272 581696 99278
rect 581644 99214 581696 99220
rect 581644 89004 581696 89010
rect 581644 88946 581696 88952
rect 580448 86964 580500 86970
rect 580448 86906 580500 86912
rect 580264 77716 580316 77722
rect 580264 77658 580316 77664
rect 579528 73160 579580 73166
rect 579526 73128 579528 73137
rect 579580 73128 579582 73137
rect 579526 73063 579582 73072
rect 579528 71256 579580 71262
rect 579526 71224 579528 71233
rect 579580 71224 579582 71233
rect 579526 71159 579582 71168
rect 579526 66328 579582 66337
rect 579526 66263 579528 66272
rect 579580 66263 579582 66272
rect 579528 66234 579580 66240
rect 579528 64864 579580 64870
rect 579528 64806 579580 64812
rect 579540 64569 579568 64806
rect 579526 64560 579582 64569
rect 579526 64495 579582 64504
rect 580264 58676 580316 58682
rect 580264 58618 580316 58624
rect 579528 57928 579580 57934
rect 579526 57896 579528 57905
rect 579580 57896 579582 57905
rect 579526 57831 579582 57840
rect 579528 56568 579580 56574
rect 579528 56510 579580 56516
rect 579540 56137 579568 56510
rect 579526 56128 579582 56137
rect 579526 56063 579582 56072
rect 579068 55072 579120 55078
rect 577502 55040 577558 55049
rect 579068 55014 579120 55020
rect 577502 54975 577558 54984
rect 580276 54262 580304 58618
rect 581656 55214 581684 88946
rect 581840 85474 581868 106286
rect 581828 85468 581880 85474
rect 581828 85410 581880 85416
rect 583036 84046 583064 109686
rect 583220 103358 583248 124850
rect 584416 118590 584444 135254
rect 584600 131170 584628 143550
rect 585980 137154 586008 144910
rect 587164 142452 587216 142458
rect 587164 142394 587216 142400
rect 585968 137148 586020 137154
rect 585968 137090 586020 137096
rect 585784 136672 585836 136678
rect 585784 136614 585836 136620
rect 584588 131164 584640 131170
rect 584588 131106 584640 131112
rect 585796 121446 585824 136614
rect 587176 128314 587204 142394
rect 588556 137290 588584 147591
rect 589462 146024 589518 146033
rect 589462 145959 589518 145968
rect 589476 144974 589504 145959
rect 589464 144968 589516 144974
rect 589464 144910 589516 144916
rect 589462 144392 589518 144401
rect 589462 144327 589518 144336
rect 589476 143614 589504 144327
rect 589464 143608 589516 143614
rect 589464 143550 589516 143556
rect 589830 142760 589886 142769
rect 589830 142695 589886 142704
rect 589844 142458 589872 142695
rect 589832 142452 589884 142458
rect 589832 142394 589884 142400
rect 590028 142154 590056 150855
rect 589936 142126 590056 142154
rect 589462 141128 589518 141137
rect 589462 141063 589518 141072
rect 589476 140826 589504 141063
rect 589464 140820 589516 140826
rect 589464 140762 589516 140768
rect 589462 139496 589518 139505
rect 589462 139431 589464 139440
rect 589516 139431 589518 139440
rect 589464 139402 589516 139408
rect 589936 139330 589964 142126
rect 589924 139324 589976 139330
rect 589924 139266 589976 139272
rect 589462 137864 589518 137873
rect 589462 137799 589518 137808
rect 588544 137284 588596 137290
rect 588544 137226 588596 137232
rect 589476 136678 589504 137799
rect 589464 136672 589516 136678
rect 589464 136614 589516 136620
rect 589462 136232 589518 136241
rect 589462 136167 589518 136176
rect 589476 135318 589504 136167
rect 589464 135312 589516 135318
rect 589464 135254 589516 135260
rect 590290 134600 590346 134609
rect 590290 134535 590346 134544
rect 588726 132968 588782 132977
rect 588726 132903 588782 132912
rect 587164 128308 587216 128314
rect 587164 128250 587216 128256
rect 587624 127220 587676 127226
rect 587624 127162 587676 127168
rect 587636 126274 587664 127162
rect 587624 126268 587676 126274
rect 587624 126210 587676 126216
rect 587348 121508 587400 121514
rect 587348 121450 587400 121456
rect 585784 121440 585836 121446
rect 585784 121382 585836 121388
rect 584588 118720 584640 118726
rect 584588 118662 584640 118668
rect 584404 118584 584456 118590
rect 584404 118526 584456 118532
rect 584404 113212 584456 113218
rect 584404 113154 584456 113160
rect 583208 103352 583260 103358
rect 583208 103294 583260 103300
rect 583024 84040 583076 84046
rect 583024 83982 583076 83988
rect 584416 82482 584444 113154
rect 584600 95062 584628 118662
rect 585968 117360 586020 117366
rect 585968 117302 586020 117308
rect 585784 116000 585836 116006
rect 585784 115942 585836 115948
rect 584588 95056 584640 95062
rect 584588 94998 584640 95004
rect 585796 92002 585824 115942
rect 585980 93430 586008 117302
rect 587164 100768 587216 100774
rect 587164 100710 587216 100716
rect 585968 93424 586020 93430
rect 585968 93366 586020 93372
rect 585784 91996 585836 92002
rect 585784 91938 585836 91944
rect 584404 82476 584456 82482
rect 584404 82418 584456 82424
rect 585784 79484 585836 79490
rect 585784 79426 585836 79432
rect 583022 77888 583078 77897
rect 583022 77823 583078 77832
rect 581644 55208 581696 55214
rect 581644 55150 581696 55156
rect 583036 54398 583064 77823
rect 584404 77308 584456 77314
rect 584404 77250 584456 77256
rect 584416 54942 584444 77250
rect 585796 71262 585824 79426
rect 587176 73166 587204 100710
rect 587360 97986 587388 121450
rect 588542 115016 588598 115025
rect 588542 114951 588598 114960
rect 587348 97980 587400 97986
rect 587348 97922 587400 97928
rect 588556 91798 588584 114951
rect 588740 113082 588768 132903
rect 590304 131782 590332 134535
rect 666848 133113 666876 209034
rect 667032 178809 667060 324294
rect 667204 310548 667256 310554
rect 667204 310490 667256 310496
rect 667018 178800 667074 178809
rect 667018 178735 667074 178744
rect 667216 134609 667244 310490
rect 667400 181393 667428 350542
rect 667572 338156 667624 338162
rect 667572 338098 667624 338104
rect 667584 186969 667612 338098
rect 668596 312905 668624 444382
rect 669976 403753 670004 536794
rect 670344 527785 670372 598023
rect 670620 529009 670648 607951
rect 670804 579057 670832 623863
rect 671172 621014 671200 640455
rect 671356 630674 671384 735558
rect 671540 713697 671568 758231
rect 671724 757897 671752 758526
rect 671710 757888 671766 757897
rect 671710 757823 671766 757832
rect 671710 757480 671766 757489
rect 671710 757415 671766 757424
rect 671526 713688 671582 713697
rect 671526 713623 671582 713632
rect 671526 713280 671582 713289
rect 671526 713215 671582 713224
rect 671540 712094 671568 713215
rect 671724 712881 671752 757415
rect 672000 732873 672028 928231
rect 672184 770681 672212 930106
rect 672538 873624 672594 873633
rect 672538 873559 672594 873568
rect 672354 784408 672410 784417
rect 672354 784343 672410 784352
rect 672170 770672 672226 770681
rect 672170 770607 672226 770616
rect 672170 733680 672226 733689
rect 672170 733615 672226 733624
rect 671986 732864 672042 732873
rect 671986 732799 672042 732808
rect 671710 712872 671766 712881
rect 671710 712807 671766 712816
rect 671540 712066 671660 712094
rect 671632 668545 671660 712066
rect 671986 688664 672042 688673
rect 671986 688599 672042 688608
rect 671618 668536 671674 668545
rect 671618 668471 671674 668480
rect 671802 668128 671858 668137
rect 671802 668063 671858 668072
rect 671526 667312 671582 667321
rect 671526 667247 671582 667256
rect 671540 649994 671568 667247
rect 671540 649966 671660 649994
rect 671632 630674 671660 649966
rect 671356 630646 671568 630674
rect 671632 630646 671752 630674
rect 671540 627881 671568 630646
rect 671526 627872 671582 627881
rect 671526 627807 671582 627816
rect 671724 627178 671752 630646
rect 671448 627150 671752 627178
rect 671448 623370 671476 627150
rect 671816 627042 671844 668063
rect 671632 627014 671844 627042
rect 671632 623529 671660 627014
rect 671802 624472 671858 624481
rect 671802 624407 671858 624416
rect 671618 623520 671674 623529
rect 671618 623455 671674 623464
rect 671448 623342 671568 623370
rect 671540 622713 671568 623342
rect 671816 623234 671844 624407
rect 671816 623206 671936 623234
rect 671710 623112 671766 623121
rect 671710 623047 671766 623056
rect 671526 622704 671582 622713
rect 671526 622639 671582 622648
rect 671080 620986 671200 621014
rect 670790 579048 670846 579057
rect 670790 578983 670846 578992
rect 670790 578640 670846 578649
rect 670790 578575 670846 578584
rect 670804 577946 670832 578575
rect 670712 577918 670832 577946
rect 670712 572714 670740 577918
rect 670882 577824 670938 577833
rect 670882 577759 670938 577768
rect 670896 572714 670924 577759
rect 671080 576201 671108 620986
rect 671436 616208 671488 616214
rect 671436 616150 671488 616156
rect 671250 594824 671306 594833
rect 671250 594759 671306 594768
rect 671066 576192 671122 576201
rect 671066 576127 671122 576136
rect 671264 572714 671292 594759
rect 671448 579873 671476 616150
rect 671434 579864 671490 579873
rect 671434 579799 671490 579808
rect 671434 579456 671490 579465
rect 671434 579391 671490 579400
rect 671448 572714 671476 579391
rect 671724 578241 671752 623047
rect 671908 616214 671936 623206
rect 672000 616842 672028 688599
rect 672184 661609 672212 733615
rect 672368 709209 672396 784343
rect 672552 754225 672580 873559
rect 672736 760345 672764 930106
rect 673366 929520 673422 929529
rect 673366 929455 673422 929464
rect 672998 870088 673054 870097
rect 672998 870023 673054 870032
rect 672722 760336 672778 760345
rect 672722 760271 672778 760280
rect 672722 759928 672778 759937
rect 672722 759863 672778 759872
rect 672538 754216 672594 754225
rect 672538 754151 672594 754160
rect 672538 738304 672594 738313
rect 672538 738239 672594 738248
rect 672552 736934 672580 738239
rect 672736 736934 672764 759863
rect 673012 755449 673040 870023
rect 673182 759112 673238 759121
rect 673182 759047 673238 759056
rect 672998 755440 673054 755449
rect 672998 755375 673054 755384
rect 672906 751360 672962 751369
rect 672906 751295 672962 751304
rect 672920 736934 672948 751295
rect 672552 736906 672672 736934
rect 672736 736906 672856 736934
rect 672920 736906 673040 736934
rect 672354 709200 672410 709209
rect 672354 709135 672410 709144
rect 672448 707260 672500 707266
rect 672448 707202 672500 707208
rect 672460 670313 672488 707202
rect 672446 670304 672502 670313
rect 672446 670239 672502 670248
rect 672446 668944 672502 668953
rect 672446 668879 672502 668888
rect 672170 661600 672226 661609
rect 672170 661535 672226 661544
rect 672460 640334 672488 668879
rect 672644 662425 672672 736906
rect 672828 715329 672856 736906
rect 673012 728142 673040 736906
rect 673000 728136 673052 728142
rect 673000 728078 673052 728084
rect 672814 715320 672870 715329
rect 672814 715255 672870 715264
rect 672814 714912 672870 714921
rect 672814 714847 672870 714856
rect 672828 669905 672856 714847
rect 673196 714513 673224 759047
rect 673380 732873 673408 929455
rect 674852 928792 674880 953391
rect 675036 934289 675064 954479
rect 675220 954366 675418 954394
rect 675220 951425 675248 954366
rect 675404 953465 675432 953768
rect 675390 953456 675446 953465
rect 675390 953391 675446 953400
rect 675312 952530 675418 952558
rect 675312 951810 675340 952530
rect 675312 951782 675524 951810
rect 675496 951538 675524 951782
rect 677506 951552 677562 951561
rect 675496 951510 676076 951538
rect 675206 951416 675262 951425
rect 675206 951351 675262 951360
rect 675850 951416 675906 951425
rect 675850 951351 675906 951360
rect 675206 951144 675262 951153
rect 675206 951079 675262 951088
rect 675022 934280 675078 934289
rect 675022 934215 675078 934224
rect 675220 933881 675248 951079
rect 675864 949482 675892 951351
rect 675852 949476 675904 949482
rect 675852 949418 675904 949424
rect 676048 948054 676076 951510
rect 677506 951487 677562 951496
rect 676036 948048 676088 948054
rect 676036 947990 676088 947996
rect 676218 941760 676274 941769
rect 676218 941695 676274 941704
rect 676232 939321 676260 941695
rect 676218 939312 676274 939321
rect 676218 939247 676274 939256
rect 676494 938088 676550 938097
rect 676048 938046 676494 938074
rect 676048 937825 676076 938046
rect 676494 938023 676550 938032
rect 676034 937816 676090 937825
rect 676034 937751 676090 937760
rect 675206 933872 675262 933881
rect 675206 933807 675262 933816
rect 677520 931161 677548 951487
rect 678242 950736 678298 950745
rect 678242 950671 678298 950680
rect 678256 935649 678284 950671
rect 682384 949476 682436 949482
rect 682384 949418 682436 949424
rect 681004 948048 681056 948054
rect 681004 947990 681056 947996
rect 678242 935640 678298 935649
rect 678242 935575 678298 935584
rect 681016 933609 681044 947990
rect 682396 935241 682424 949418
rect 683118 947336 683174 947345
rect 683118 947271 683174 947280
rect 683132 939729 683160 947271
rect 703694 940508 703722 940644
rect 704154 940508 704182 940644
rect 704614 940508 704642 940644
rect 705074 940508 705102 940644
rect 705534 940508 705562 940644
rect 705994 940508 706022 940644
rect 706454 940508 706482 940644
rect 706914 940508 706942 940644
rect 707374 940508 707402 940644
rect 707834 940508 707862 940644
rect 708294 940508 708322 940644
rect 708754 940508 708782 940644
rect 709214 940508 709242 940644
rect 683118 939720 683174 939729
rect 683118 939655 683174 939664
rect 682382 935232 682438 935241
rect 682382 935167 682438 935176
rect 681002 933600 681058 933609
rect 681002 933535 681058 933544
rect 677506 931152 677562 931161
rect 677506 931087 677562 931096
rect 683118 929112 683174 929121
rect 683118 929047 683174 929056
rect 683132 928810 683160 929047
rect 675852 928804 675904 928810
rect 674852 928764 675852 928792
rect 675852 928746 675904 928752
rect 683120 928804 683172 928810
rect 683120 928746 683172 928752
rect 675298 879200 675354 879209
rect 675298 879135 675354 879144
rect 675312 877418 675340 879135
rect 675404 877418 675432 877540
rect 675312 877390 675432 877418
rect 675312 876982 675432 877010
rect 675312 876874 675340 876982
rect 674944 876846 675340 876874
rect 675404 876860 675432 876982
rect 674944 870913 674972 876846
rect 675772 875945 675800 876248
rect 675758 875936 675814 875945
rect 675758 875871 675814 875880
rect 675404 874041 675432 874412
rect 675390 874032 675446 874041
rect 675390 873967 675446 873976
rect 675404 873633 675432 873868
rect 675390 873624 675446 873633
rect 675390 873559 675446 873568
rect 675114 873216 675170 873225
rect 675170 873174 675418 873202
rect 675114 873151 675170 873160
rect 675404 872273 675432 872576
rect 675390 872264 675446 872273
rect 675390 872199 675446 872208
rect 674930 870904 674986 870913
rect 674930 870839 674986 870848
rect 675114 870088 675170 870097
rect 675170 870046 675418 870074
rect 675114 870023 675170 870032
rect 674116 869502 675418 869530
rect 673918 864920 673974 864929
rect 673918 864855 673974 864864
rect 673734 779376 673790 779385
rect 673734 779311 673790 779320
rect 673550 777472 673606 777481
rect 673550 777407 673606 777416
rect 673366 732864 673422 732873
rect 673366 732799 673422 732808
rect 673564 732154 673592 777407
rect 673748 756254 673776 779311
rect 673932 772041 673960 864855
rect 673918 772032 673974 772041
rect 673918 771967 673974 771976
rect 674116 756254 674144 869502
rect 674668 868861 675340 868889
rect 674470 788080 674526 788089
rect 674470 788015 674526 788024
rect 674286 780056 674342 780065
rect 674286 779991 674342 780000
rect 673656 756226 673776 756254
rect 673932 756226 674144 756254
rect 673656 736930 673684 756226
rect 673932 752185 673960 756226
rect 673918 752176 673974 752185
rect 673918 752111 673974 752120
rect 673656 736902 673776 736930
rect 673552 732148 673604 732154
rect 673552 732090 673604 732096
rect 673366 730144 673422 730153
rect 673366 730079 673422 730088
rect 673380 728634 673408 730079
rect 673748 728770 673776 736902
rect 674012 732148 674064 732154
rect 674012 732090 674064 732096
rect 673656 728742 673776 728770
rect 673380 728606 673592 728634
rect 673366 728512 673422 728521
rect 673366 728447 673368 728456
rect 673420 728447 673422 728456
rect 673368 728418 673420 728424
rect 673564 728362 673592 728606
rect 673380 728334 673592 728362
rect 673182 714504 673238 714513
rect 673182 714439 673238 714448
rect 672998 714096 673054 714105
rect 672998 714031 673054 714040
rect 673012 707266 673040 714031
rect 673000 707260 673052 707266
rect 673000 707202 673052 707208
rect 673182 698320 673238 698329
rect 673182 698255 673238 698264
rect 672998 685808 673054 685817
rect 672998 685743 673054 685752
rect 672814 669896 672870 669905
rect 672814 669831 672870 669840
rect 672814 669488 672870 669497
rect 672814 669423 672870 669432
rect 672630 662416 672686 662425
rect 672630 662351 672686 662360
rect 672630 661192 672686 661201
rect 672630 661127 672686 661136
rect 672184 640306 672488 640334
rect 672184 635497 672212 640306
rect 672354 638752 672410 638761
rect 672354 638687 672410 638696
rect 672170 635488 672226 635497
rect 672170 635423 672226 635432
rect 672172 627156 672224 627162
rect 672172 627098 672224 627104
rect 672184 619857 672212 627098
rect 672170 619848 672226 619857
rect 672170 619783 672226 619792
rect 672000 616814 672212 616842
rect 672184 616729 672212 616814
rect 672170 616720 672226 616729
rect 672170 616655 672226 616664
rect 671896 616208 671948 616214
rect 671896 616150 671948 616156
rect 671986 614952 672042 614961
rect 671986 614887 672042 614896
rect 671710 578232 671766 578241
rect 671710 578167 671766 578176
rect 670712 572686 670832 572714
rect 670896 572686 671016 572714
rect 671264 572686 671384 572714
rect 671448 572686 671568 572714
rect 670804 535129 670832 572686
rect 670790 535120 670846 535129
rect 670790 535055 670846 535064
rect 670988 534970 671016 572686
rect 671158 569664 671214 569673
rect 671158 569599 671214 569608
rect 671172 563054 671200 569599
rect 671356 563122 671384 572686
rect 671540 563122 671568 572686
rect 670896 534942 671016 534970
rect 671080 563026 671200 563054
rect 671264 563094 671384 563122
rect 671448 563094 671568 563122
rect 670896 533089 670924 534942
rect 670882 533080 670938 533089
rect 671080 533066 671108 563026
rect 671264 533186 671292 563094
rect 671448 534721 671476 563094
rect 671710 555248 671766 555257
rect 671710 555183 671766 555192
rect 671434 534712 671490 534721
rect 671434 534647 671490 534656
rect 671434 534440 671490 534449
rect 671434 534375 671490 534384
rect 671252 533180 671304 533186
rect 671252 533122 671304 533128
rect 671080 533038 671292 533066
rect 670882 533015 670938 533024
rect 670884 532908 670936 532914
rect 670884 532850 670936 532856
rect 670606 529000 670662 529009
rect 670606 528935 670662 528944
rect 670330 527776 670386 527785
rect 670330 527711 670386 527720
rect 670896 524929 670924 532850
rect 671264 532794 671292 533038
rect 671448 532930 671476 534375
rect 671080 532766 671292 532794
rect 671356 532902 671476 532930
rect 670882 524920 670938 524929
rect 670882 524855 670938 524864
rect 671080 455054 671108 532766
rect 671356 490929 671384 532902
rect 671526 532808 671582 532817
rect 671526 532743 671582 532752
rect 671342 490920 671398 490929
rect 671342 490855 671398 490864
rect 671540 489297 671568 532743
rect 671526 489288 671582 489297
rect 671526 489223 671582 489232
rect 671724 486033 671752 555183
rect 671710 486024 671766 486033
rect 671710 485959 671766 485968
rect 672000 455433 672028 614887
rect 672170 604752 672226 604761
rect 672170 604687 672226 604696
rect 672184 576854 672212 604687
rect 672368 579562 672396 638687
rect 672644 630674 672672 661127
rect 672644 630646 672764 630674
rect 672538 604344 672594 604353
rect 672538 604279 672594 604288
rect 672552 582374 672580 604279
rect 672736 582374 672764 630646
rect 672828 627914 672856 669423
rect 673012 627914 673040 685743
rect 673196 630674 673224 698255
rect 673380 666505 673408 728334
rect 673656 727274 673684 728742
rect 673828 728612 673880 728618
rect 673828 728554 673880 728560
rect 673840 728249 673868 728554
rect 673826 728240 673882 728249
rect 673826 728175 673882 728184
rect 673826 727696 673882 727705
rect 673826 727631 673882 727640
rect 673840 727274 673868 727631
rect 673564 727246 673684 727274
rect 673748 727246 673868 727274
rect 673564 724169 673592 727246
rect 673550 724160 673606 724169
rect 673550 724095 673606 724104
rect 673550 689616 673606 689625
rect 673550 689551 673606 689560
rect 673366 666496 673422 666505
rect 673366 666431 673422 666440
rect 673368 666256 673420 666262
rect 673368 666198 673420 666204
rect 673380 660793 673408 666198
rect 673366 660784 673422 660793
rect 673366 660719 673422 660728
rect 673366 659968 673422 659977
rect 673366 659903 673422 659912
rect 673196 630646 673316 630674
rect 672828 627886 672948 627914
rect 673012 627886 673132 627914
rect 672920 626754 672948 627886
rect 672908 626748 672960 626754
rect 672908 626690 672960 626696
rect 673104 626618 673132 627886
rect 673092 626612 673144 626618
rect 673092 626554 673144 626560
rect 672908 626408 672960 626414
rect 672908 626350 672960 626356
rect 672920 621738 672948 626350
rect 673288 625002 673316 630646
rect 672828 621710 672948 621738
rect 673012 624974 673316 625002
rect 672828 618254 672856 621710
rect 673012 621625 673040 624974
rect 673182 622296 673238 622305
rect 673182 622231 673238 622240
rect 672998 621616 673054 621625
rect 672998 621551 673054 621560
rect 672828 618226 672948 618254
rect 672920 615777 672948 618226
rect 672906 615768 672962 615777
rect 672906 615703 672962 615712
rect 672460 582346 672580 582374
rect 672644 582346 672764 582374
rect 672460 579614 672488 582346
rect 672644 579614 672672 582346
rect 672460 579586 672580 579614
rect 672644 579586 672764 579614
rect 672356 579556 672408 579562
rect 672356 579498 672408 579504
rect 672552 577538 672580 579586
rect 672092 576826 672212 576854
rect 672276 577510 672580 577538
rect 672092 567194 672120 576826
rect 672276 571962 672304 577510
rect 672446 577008 672502 577017
rect 672446 576943 672502 576952
rect 672460 572762 672488 576943
rect 672448 572756 672500 572762
rect 672448 572698 672500 572704
rect 672736 572642 672764 579586
rect 673000 579556 673052 579562
rect 673000 579498 673052 579504
rect 673012 574569 673040 579498
rect 673196 577425 673224 622231
rect 673182 577416 673238 577425
rect 673182 577351 673238 577360
rect 672998 574560 673054 574569
rect 672998 574495 673054 574504
rect 672908 572756 672960 572762
rect 672908 572698 672960 572704
rect 672184 571934 672304 571962
rect 672552 572614 672764 572642
rect 672184 569242 672212 571934
rect 672184 569214 672488 569242
rect 672264 567316 672316 567322
rect 672264 567258 672316 567264
rect 672092 567166 672212 567194
rect 672184 538214 672212 567166
rect 672092 538186 672212 538214
rect 672092 531298 672120 538186
rect 672276 531457 672304 567258
rect 672460 538214 672488 569214
rect 672552 567746 672580 572614
rect 672552 567718 672672 567746
rect 672644 546281 672672 567718
rect 672920 567322 672948 572698
rect 672908 567316 672960 567322
rect 672908 567258 672960 567264
rect 672906 559056 672962 559065
rect 672906 558991 672962 559000
rect 672630 546272 672686 546281
rect 672630 546207 672686 546216
rect 672368 538186 672488 538214
rect 672368 533338 672396 538186
rect 672538 533488 672594 533497
rect 672538 533423 672594 533432
rect 672368 533310 672488 533338
rect 672262 531448 672318 531457
rect 672262 531383 672318 531392
rect 672460 531298 672488 533310
rect 672092 531270 672212 531298
rect 672184 530233 672212 531270
rect 672368 531270 672488 531298
rect 672170 530224 672226 530233
rect 672170 530159 672226 530168
rect 672368 529417 672396 531270
rect 672354 529408 672410 529417
rect 672354 529343 672410 529352
rect 672552 528554 672580 533423
rect 672722 531856 672778 531865
rect 672722 531791 672778 531800
rect 672736 528714 672764 531791
rect 672736 528686 672856 528714
rect 672552 528526 672764 528554
rect 672736 490113 672764 528526
rect 672828 495434 672856 528686
rect 672920 505094 672948 558991
rect 673182 548448 673238 548457
rect 673182 548383 673238 548392
rect 672920 505066 673132 505094
rect 672828 495406 672948 495434
rect 672722 490104 672778 490113
rect 672722 490039 672778 490048
rect 672446 489696 672502 489705
rect 672446 489631 672502 489640
rect 671986 455424 672042 455433
rect 671986 455359 672042 455368
rect 671068 455048 671120 455054
rect 671068 454990 671120 454996
rect 672264 453960 672316 453966
rect 672264 453902 672316 453908
rect 672276 453801 672304 453902
rect 672262 453792 672318 453801
rect 672262 453727 672318 453736
rect 671344 430636 671396 430642
rect 671344 430578 671396 430584
rect 669962 403744 670018 403753
rect 669962 403679 670018 403688
rect 670606 393544 670662 393553
rect 670606 393479 670662 393488
rect 669962 347304 670018 347313
rect 669962 347239 670018 347248
rect 668582 312896 668638 312905
rect 668582 312831 668638 312840
rect 668306 302288 668362 302297
rect 668306 302223 668362 302232
rect 667756 284368 667808 284374
rect 667756 284310 667808 284316
rect 667570 186960 667626 186969
rect 667570 186895 667626 186904
rect 667386 181384 667442 181393
rect 667386 181319 667442 181328
rect 667768 135969 667796 284310
rect 668124 235340 668176 235346
rect 668124 235282 668176 235288
rect 667940 230308 667992 230314
rect 667940 230250 667992 230256
rect 667952 224942 667980 230250
rect 667940 224936 667992 224942
rect 667940 224878 667992 224884
rect 667940 224664 667992 224670
rect 667940 224606 667992 224612
rect 667952 223961 667980 224606
rect 667938 223952 667994 223961
rect 667938 223887 667994 223896
rect 667940 219564 667992 219570
rect 667940 219506 667992 219512
rect 667952 192681 667980 219506
rect 667938 192672 667994 192681
rect 667938 192607 667994 192616
rect 667940 189440 667992 189446
rect 667938 189408 667940 189417
rect 667992 189408 667994 189417
rect 667938 189343 667994 189352
rect 668136 182889 668164 235282
rect 668320 229537 668348 302223
rect 668768 237448 668820 237454
rect 668768 237390 668820 237396
rect 668490 234560 668546 234569
rect 668490 234495 668546 234504
rect 668306 229528 668362 229537
rect 668306 229463 668362 229472
rect 668308 226636 668360 226642
rect 668308 226578 668360 226584
rect 668320 226409 668348 226578
rect 668306 226400 668362 226409
rect 668306 226335 668362 226344
rect 668306 225312 668362 225321
rect 668306 225247 668362 225256
rect 668320 225078 668348 225247
rect 668308 225072 668360 225078
rect 668308 225014 668360 225020
rect 668308 224936 668360 224942
rect 668308 224878 668360 224884
rect 668320 222194 668348 224878
rect 668228 222166 668348 222194
rect 668228 215294 668256 222166
rect 668228 215266 668348 215294
rect 668122 182880 668178 182889
rect 668122 182815 668178 182824
rect 667940 174752 667992 174758
rect 667938 174720 667940 174729
rect 667992 174720 667994 174729
rect 667938 174655 667994 174664
rect 668032 169720 668084 169726
rect 668030 169688 668032 169697
rect 668084 169688 668086 169697
rect 668030 169623 668086 169632
rect 667940 164960 667992 164966
rect 667938 164928 667940 164937
rect 667992 164928 667994 164937
rect 667938 164863 667994 164872
rect 668320 163305 668348 215266
rect 668306 163296 668362 163305
rect 668306 163231 668362 163240
rect 668504 148617 668532 234495
rect 668780 153513 668808 237390
rect 668950 236736 669006 236745
rect 668950 236671 669006 236680
rect 668964 160041 668992 236671
rect 669780 235544 669832 235550
rect 669780 235486 669832 235492
rect 669596 234252 669648 234258
rect 669596 234194 669648 234200
rect 669136 233640 669188 233646
rect 669136 233582 669188 233588
rect 669148 209774 669176 233582
rect 669320 230444 669372 230450
rect 669320 230386 669372 230392
rect 669332 230058 669360 230386
rect 669240 230030 669360 230058
rect 669240 219586 669268 230030
rect 669412 225480 669464 225486
rect 669412 225422 669464 225428
rect 669424 225049 669452 225422
rect 669410 225040 669466 225049
rect 669410 224975 669466 224984
rect 669412 224188 669464 224194
rect 669412 224130 669464 224136
rect 669424 223689 669452 224130
rect 669410 223680 669466 223689
rect 669410 223615 669466 223624
rect 669240 219570 669360 219586
rect 669240 219564 669372 219570
rect 669240 219558 669320 219564
rect 669320 219506 669372 219512
rect 669410 214160 669466 214169
rect 669410 214095 669466 214104
rect 669056 209746 669176 209774
rect 669056 202450 669084 209746
rect 669226 208312 669282 208321
rect 669226 208247 669282 208256
rect 669240 207369 669268 208247
rect 669226 207360 669282 207369
rect 669226 207295 669282 207304
rect 669226 202464 669282 202473
rect 669056 202422 669226 202450
rect 669226 202399 669282 202408
rect 669136 199368 669188 199374
rect 669134 199336 669136 199345
rect 669188 199336 669190 199345
rect 669134 199271 669190 199280
rect 669226 198792 669282 198801
rect 669226 198727 669282 198736
rect 669240 194426 669268 198727
rect 669424 197169 669452 214095
rect 669410 197160 669466 197169
rect 669410 197095 669466 197104
rect 669240 194398 669360 194426
rect 669136 194336 669188 194342
rect 669134 194304 669136 194313
rect 669188 194304 669190 194313
rect 669134 194239 669190 194248
rect 669332 194154 669360 194398
rect 669148 194126 669360 194154
rect 669148 187649 669176 194126
rect 669608 190454 669636 234194
rect 669332 190426 669636 190454
rect 669134 187640 669190 187649
rect 669134 187575 669190 187584
rect 669332 184906 669360 190426
rect 669240 184878 669360 184906
rect 669240 184521 669268 184878
rect 669226 184512 669282 184521
rect 669226 184447 669282 184456
rect 669792 174758 669820 235486
rect 669780 174752 669832 174758
rect 669780 174694 669832 174700
rect 669778 168192 669834 168201
rect 669778 168127 669834 168136
rect 669134 164248 669190 164257
rect 669134 164183 669190 164192
rect 668950 160032 669006 160041
rect 668950 159967 669006 159976
rect 668766 153504 668822 153513
rect 668766 153439 668822 153448
rect 668766 149152 668822 149161
rect 668766 149087 668822 149096
rect 668490 148608 668546 148617
rect 668490 148543 668546 148552
rect 668584 145580 668636 145586
rect 668584 145522 668636 145528
rect 668596 145353 668624 145522
rect 668582 145344 668638 145353
rect 668582 145279 668638 145288
rect 667940 136400 667992 136406
rect 667940 136342 667992 136348
rect 667754 135960 667810 135969
rect 667754 135895 667810 135904
rect 667952 135561 667980 136342
rect 667938 135552 667994 135561
rect 667938 135487 667994 135496
rect 667202 134600 667258 134609
rect 667202 134535 667258 134544
rect 666834 133104 666890 133113
rect 666834 133039 666890 133048
rect 590292 131776 590344 131782
rect 590292 131718 590344 131724
rect 589462 131336 589518 131345
rect 589462 131271 589464 131280
rect 589516 131271 589518 131280
rect 589464 131242 589516 131248
rect 589646 129704 589702 129713
rect 589646 129639 589702 129648
rect 589462 128072 589518 128081
rect 589462 128007 589518 128016
rect 589476 127226 589504 128007
rect 589464 127220 589516 127226
rect 589464 127162 589516 127168
rect 589660 124914 589688 129639
rect 668582 128344 668638 128353
rect 668582 128279 668638 128288
rect 590106 126440 590162 126449
rect 590106 126375 590162 126384
rect 589648 124908 589700 124914
rect 589648 124850 589700 124856
rect 589922 124808 589978 124817
rect 589922 124743 589978 124752
rect 589462 123176 589518 123185
rect 589462 123111 589518 123120
rect 589476 122874 589504 123111
rect 589464 122868 589516 122874
rect 589464 122810 589516 122816
rect 589278 121544 589334 121553
rect 589278 121479 589280 121488
rect 589332 121479 589334 121488
rect 589280 121450 589332 121456
rect 589462 119912 589518 119921
rect 589462 119847 589518 119856
rect 589476 118726 589504 119847
rect 589464 118720 589516 118726
rect 589464 118662 589516 118668
rect 589462 118280 589518 118289
rect 589462 118215 589518 118224
rect 589476 117366 589504 118215
rect 589464 117360 589516 117366
rect 589464 117302 589516 117308
rect 589462 116648 589518 116657
rect 589462 116583 589518 116592
rect 589476 116006 589504 116583
rect 589464 116000 589516 116006
rect 589464 115942 589516 115948
rect 589462 113384 589518 113393
rect 589462 113319 589518 113328
rect 589476 113218 589504 113319
rect 589464 113212 589516 113218
rect 589464 113154 589516 113160
rect 588728 113076 588780 113082
rect 588728 113018 588780 113024
rect 589370 111752 589426 111761
rect 589370 111687 589426 111696
rect 589384 109750 589412 111687
rect 589936 111110 589964 124743
rect 590120 122126 590148 126375
rect 667940 125588 667992 125594
rect 667940 125530 667992 125536
rect 590108 122120 590160 122126
rect 590108 122062 590160 122068
rect 667952 119241 667980 125530
rect 668596 120873 668624 128279
rect 668780 125769 668808 149087
rect 669148 138825 669176 164183
rect 669134 138816 669190 138825
rect 669134 138751 669190 138760
rect 668766 125760 668822 125769
rect 668766 125695 668822 125704
rect 669792 125594 669820 168127
rect 669976 136406 670004 347239
rect 670422 256728 670478 256737
rect 670422 256663 670478 256672
rect 670436 235929 670464 256663
rect 670422 235920 670478 235929
rect 670422 235855 670478 235864
rect 670330 233200 670386 233209
rect 670330 233135 670386 233144
rect 670146 232928 670202 232937
rect 670146 232863 670202 232872
rect 670160 164966 670188 232863
rect 670344 169726 670372 233135
rect 670620 211177 670648 393479
rect 671356 269793 671384 430578
rect 672460 401713 672488 489631
rect 672920 488481 672948 495406
rect 672906 488472 672962 488481
rect 672906 488407 672962 488416
rect 672630 488064 672686 488073
rect 672630 487999 672686 488008
rect 672446 401704 672502 401713
rect 672446 401639 672502 401648
rect 672446 400480 672502 400489
rect 672446 400415 672502 400424
rect 672262 393952 672318 393961
rect 672262 393887 672318 393896
rect 672276 376281 672304 393887
rect 672262 376272 672318 376281
rect 672262 376207 672318 376216
rect 672460 355881 672488 400415
rect 672644 400081 672672 487999
rect 673104 485774 673132 505066
rect 673012 485746 673132 485774
rect 673012 484809 673040 485746
rect 673196 485625 673224 548383
rect 673182 485616 673238 485625
rect 673182 485551 673238 485560
rect 672998 484800 673054 484809
rect 672998 484735 673054 484744
rect 673380 455954 673408 659903
rect 673564 636857 673592 689551
rect 673748 681057 673776 727246
rect 674024 726617 674052 732090
rect 674150 728136 674202 728142
rect 674150 728078 674202 728084
rect 674162 727977 674190 728078
rect 674148 727968 674204 727977
rect 674148 727903 674204 727912
rect 674300 726889 674328 779991
rect 674484 736934 674512 788015
rect 674668 757217 674696 868861
rect 675312 868850 675340 868861
rect 675404 868850 675432 868875
rect 675312 868822 675432 868850
rect 675298 868456 675354 868465
rect 675298 868391 675354 868400
rect 674838 868184 674894 868193
rect 674838 868119 674894 868128
rect 674852 867513 674880 868119
rect 674838 867504 674894 867513
rect 674838 867439 674894 867448
rect 675312 866266 675340 868391
rect 675496 867921 675524 868224
rect 675482 867912 675538 867921
rect 675482 867847 675538 867856
rect 675482 867504 675538 867513
rect 675482 867439 675538 867448
rect 675496 867035 675524 867439
rect 675312 866238 675432 866266
rect 675404 865844 675432 866238
rect 675404 864929 675432 865195
rect 675390 864920 675446 864929
rect 675390 864855 675446 864864
rect 675496 864249 675524 864552
rect 675482 864240 675538 864249
rect 675482 864175 675538 864184
rect 675312 863382 675432 863410
rect 675312 863342 675340 863382
rect 675128 863314 675340 863342
rect 675404 863328 675432 863382
rect 675128 801794 675156 863314
rect 675298 863152 675354 863161
rect 675298 863087 675354 863096
rect 675312 859754 675340 863087
rect 675220 859726 675340 859754
rect 675220 856994 675248 859726
rect 675220 856966 675340 856994
rect 675312 804554 675340 856966
rect 675036 801766 675156 801794
rect 675220 804526 675340 804554
rect 674838 796920 674894 796929
rect 674838 796855 674894 796864
rect 674852 784145 674880 796855
rect 675036 792134 675064 801766
rect 675220 796929 675248 804526
rect 675206 796920 675262 796929
rect 675206 796855 675262 796864
rect 675036 792106 675156 792134
rect 675128 789698 675156 792106
rect 675036 789670 675156 789698
rect 675036 785234 675064 789670
rect 675206 789440 675262 789449
rect 675206 789375 675262 789384
rect 675220 787693 675248 789375
rect 675404 788089 675432 788324
rect 675390 788080 675446 788089
rect 675390 788015 675446 788024
rect 675220 787665 675418 787693
rect 674944 785206 675064 785234
rect 675128 787018 675418 787046
rect 674944 784258 674972 785206
rect 674944 784230 675064 784258
rect 674838 784136 674894 784145
rect 674838 784071 674894 784080
rect 674838 778968 674894 778977
rect 674838 778903 674894 778912
rect 674852 776529 674880 778903
rect 674838 776520 674894 776529
rect 674838 776455 674894 776464
rect 674838 775840 674894 775849
rect 674838 775775 674894 775784
rect 674852 768233 674880 775775
rect 675036 774897 675064 784230
rect 675128 779714 675156 787018
rect 675298 786720 675354 786729
rect 675298 786655 675354 786664
rect 675312 785234 675340 786655
rect 675312 785206 675432 785234
rect 675404 785196 675432 785206
rect 675404 784417 675432 784652
rect 675390 784408 675446 784417
rect 675390 784343 675446 784352
rect 675298 784136 675354 784145
rect 675298 784071 675354 784080
rect 675128 779686 675248 779714
rect 675220 775418 675248 779686
rect 675128 775390 675248 775418
rect 675128 775146 675156 775390
rect 675128 775118 675248 775146
rect 675022 774888 675078 774897
rect 675022 774823 675078 774832
rect 674838 768224 674894 768233
rect 674838 768159 674894 768168
rect 675220 766601 675248 775118
rect 675312 770054 675340 784071
rect 675496 783873 675524 783972
rect 675482 783864 675538 783873
rect 675482 783799 675538 783808
rect 675496 783057 675524 783360
rect 675482 783048 675538 783057
rect 675482 782983 675538 782992
rect 675496 780745 675524 780844
rect 675482 780736 675538 780745
rect 675482 780671 675538 780680
rect 675496 780065 675524 780300
rect 675482 780056 675538 780065
rect 675482 779991 675538 780000
rect 675496 779385 675524 779688
rect 675482 779376 675538 779385
rect 675482 779311 675538 779320
rect 675496 778705 675524 779008
rect 675482 778696 675538 778705
rect 675482 778631 675538 778640
rect 675496 777481 675524 777852
rect 675482 777472 675538 777481
rect 675482 777407 675538 777416
rect 675496 776529 675524 776628
rect 675482 776520 675538 776529
rect 675482 776455 675538 776464
rect 675496 775849 675524 776016
rect 675482 775840 675538 775849
rect 675482 775775 675538 775784
rect 675666 775704 675722 775713
rect 675666 775639 675722 775648
rect 675680 775336 675708 775639
rect 675496 773809 675524 774180
rect 675482 773800 675538 773809
rect 675482 773735 675538 773744
rect 682382 772712 682438 772721
rect 682382 772647 682438 772656
rect 675312 770026 675892 770054
rect 675206 766592 675262 766601
rect 675206 766527 675262 766536
rect 674654 757208 674710 757217
rect 674654 757143 674710 757152
rect 675864 755857 675892 770026
rect 676126 768224 676182 768233
rect 676126 768159 676182 768168
rect 676140 766601 676168 768159
rect 676126 766592 676182 766601
rect 676126 766527 676182 766536
rect 676034 763056 676090 763065
rect 676034 762991 676090 763000
rect 676048 760753 676076 762991
rect 677046 761968 677102 761977
rect 677046 761903 677102 761912
rect 676770 761832 676826 761841
rect 676770 761767 676826 761776
rect 676034 760744 676090 760753
rect 676034 760679 676090 760688
rect 676034 757208 676090 757217
rect 676034 757143 676036 757152
rect 676088 757143 676090 757152
rect 676036 757114 676088 757120
rect 675850 755848 675906 755857
rect 675850 755783 675906 755792
rect 676784 755041 676812 761767
rect 676770 755032 676826 755041
rect 676770 754967 676826 754976
rect 677060 754633 677088 761903
rect 682396 757081 682424 772647
rect 683210 772032 683266 772041
rect 683210 771967 683266 771976
rect 683224 770054 683252 771967
rect 683394 770944 683450 770953
rect 683394 770879 683450 770888
rect 683224 770026 683344 770054
rect 683120 757172 683172 757178
rect 683120 757114 683172 757120
rect 682382 757072 682438 757081
rect 682382 757007 682438 757016
rect 677046 754624 677102 754633
rect 677046 754559 677102 754568
rect 683132 753001 683160 757114
rect 683316 756673 683344 770026
rect 683408 759370 683436 770879
rect 683578 770672 683634 770681
rect 683578 770607 683634 770616
rect 683592 759529 683620 770607
rect 703694 762076 703722 762212
rect 704154 762076 704182 762212
rect 704614 762076 704642 762212
rect 705074 762076 705102 762212
rect 705534 762076 705562 762212
rect 705994 762076 706022 762212
rect 706454 762076 706482 762212
rect 706914 762076 706942 762212
rect 707374 762076 707402 762212
rect 707834 762076 707862 762212
rect 708294 762076 708322 762212
rect 708754 762076 708782 762212
rect 709214 762076 709242 762212
rect 683578 759520 683634 759529
rect 683578 759455 683634 759464
rect 683408 759342 683528 759370
rect 683302 756664 683358 756673
rect 683302 756599 683358 756608
rect 683500 753817 683528 759342
rect 683486 753808 683542 753817
rect 683486 753743 683542 753752
rect 683118 752992 683174 753001
rect 683118 752927 683174 752936
rect 675128 743294 675418 743322
rect 675128 743209 675156 743294
rect 675114 743200 675170 743209
rect 675114 743135 675170 743144
rect 674930 742792 674986 742801
rect 674930 742727 674986 742736
rect 674944 741418 674972 742727
rect 675404 742529 675432 742696
rect 675390 742520 675446 742529
rect 675390 742455 675446 742464
rect 675312 742070 675432 742098
rect 675312 742030 675340 742070
rect 675128 742002 675340 742030
rect 675404 742016 675432 742070
rect 675128 741577 675156 742002
rect 675114 741568 675170 741577
rect 675114 741503 675170 741512
rect 674944 741390 675156 741418
rect 674930 741160 674986 741169
rect 674930 741095 674986 741104
rect 674944 739038 674972 741095
rect 675128 740194 675156 741390
rect 675128 740166 675418 740194
rect 675114 739664 675170 739673
rect 675170 739622 675418 739650
rect 675114 739599 675170 739608
rect 674944 739010 675340 739038
rect 675312 738970 675340 739010
rect 675404 738970 675432 739024
rect 675312 738942 675432 738970
rect 675022 738576 675078 738585
rect 675022 738511 675078 738520
rect 675036 738154 675064 738511
rect 675206 738372 675262 738381
rect 675262 738330 675418 738358
rect 675206 738307 675262 738316
rect 675036 738126 675340 738154
rect 675114 737080 675170 737089
rect 675114 737015 675170 737024
rect 674484 736906 674604 736934
rect 674286 726880 674342 726889
rect 674286 726815 674342 726824
rect 674576 726617 674604 736906
rect 675128 735333 675156 737015
rect 675312 735842 675340 738126
rect 675404 735842 675432 735896
rect 675312 735814 675432 735842
rect 675128 735305 675418 735333
rect 674760 734658 675418 734686
rect 674760 727705 674788 734658
rect 674930 734360 674986 734369
rect 674930 734295 674986 734304
rect 674944 731626 674972 734295
rect 675128 734017 675418 734045
rect 675128 733689 675156 734017
rect 675114 733680 675170 733689
rect 675114 733615 675170 733624
rect 675114 733408 675170 733417
rect 675114 733343 675170 733352
rect 675128 732850 675156 733343
rect 675128 732822 675418 732850
rect 675312 731734 675432 731762
rect 675312 731626 675340 731734
rect 674944 731598 675340 731626
rect 675404 731612 675432 731734
rect 675114 731504 675170 731513
rect 675114 731439 675170 731448
rect 675128 729178 675156 731439
rect 675312 730986 675418 731014
rect 675312 730153 675340 730986
rect 675482 730552 675538 730561
rect 675482 730487 675538 730496
rect 675496 730351 675524 730487
rect 675298 730144 675354 730153
rect 675298 730079 675354 730088
rect 675128 729150 675418 729178
rect 674746 727696 674802 727705
rect 674746 727631 674802 727640
rect 683486 726880 683542 726889
rect 683486 726815 683542 726824
rect 674010 726608 674066 726617
rect 674010 726543 674066 726552
rect 674562 726608 674618 726617
rect 674562 726543 674618 726552
rect 682382 725792 682438 725801
rect 682382 725727 682438 725736
rect 677322 724296 677378 724305
rect 677322 724231 677324 724240
rect 677376 724231 677378 724240
rect 677324 724202 677376 724208
rect 676034 718312 676090 718321
rect 676034 718247 676090 718256
rect 676048 715737 676076 718247
rect 676034 715728 676090 715737
rect 676034 715663 676090 715672
rect 682396 711657 682424 725727
rect 683118 725520 683174 725529
rect 683118 725455 683174 725464
rect 682382 711648 682438 711657
rect 682382 711583 682438 711592
rect 683132 708393 683160 725455
rect 683304 724260 683356 724266
rect 683304 724202 683356 724208
rect 683118 708384 683174 708393
rect 683118 708319 683174 708328
rect 683316 707985 683344 724202
rect 683302 707976 683358 707985
rect 683302 707911 683358 707920
rect 683500 707169 683528 726815
rect 683670 726472 683726 726481
rect 683670 726407 683726 726416
rect 683684 711249 683712 726407
rect 703694 717196 703722 717264
rect 704154 717196 704182 717264
rect 704614 717196 704642 717264
rect 705074 717196 705102 717264
rect 705534 717196 705562 717264
rect 705994 717196 706022 717264
rect 706454 717196 706482 717264
rect 706914 717196 706942 717264
rect 707374 717196 707402 717264
rect 707834 717196 707862 717264
rect 708294 717196 708322 717264
rect 708754 717196 708782 717264
rect 709214 717196 709242 717264
rect 683670 711240 683726 711249
rect 683670 711175 683726 711184
rect 683486 707160 683542 707169
rect 683486 707095 683542 707104
rect 674378 706344 674434 706353
rect 674378 706279 674434 706288
rect 674010 693016 674066 693025
rect 674010 692951 674066 692960
rect 673734 681048 673790 681057
rect 673734 680983 673790 680992
rect 673734 647864 673790 647873
rect 673734 647799 673790 647808
rect 673550 636848 673606 636857
rect 673550 636783 673606 636792
rect 673552 626748 673604 626754
rect 673552 626690 673604 626696
rect 673564 625161 673592 626690
rect 673550 625152 673606 625161
rect 673550 625087 673606 625096
rect 673550 603528 673606 603537
rect 673550 603463 673606 603472
rect 673564 598934 673592 603463
rect 673472 598906 673592 598934
rect 673472 591410 673500 598906
rect 673748 598890 673776 647799
rect 674024 621014 674052 692951
rect 674194 690160 674250 690169
rect 674194 690095 674250 690104
rect 674208 683114 674236 690095
rect 674208 683086 674328 683114
rect 674300 652202 674328 683086
rect 674116 652174 674328 652202
rect 674116 647234 674144 652174
rect 674392 652066 674420 706279
rect 674930 699816 674986 699825
rect 674930 699751 674986 699760
rect 674944 697694 674972 699751
rect 675128 698329 675418 698337
rect 675114 698320 675418 698329
rect 675170 698309 675418 698320
rect 675114 698255 675170 698264
rect 674944 697666 675418 697694
rect 675404 696833 675432 697035
rect 675390 696824 675446 696833
rect 675390 696759 675446 696768
rect 675128 695201 675418 695209
rect 675114 695192 675418 695201
rect 675170 695181 675418 695192
rect 675114 695127 675170 695136
rect 675680 694385 675708 694620
rect 675666 694376 675722 694385
rect 675666 694311 675722 694320
rect 674668 693994 675418 694022
rect 674668 656894 674696 693994
rect 675312 693382 675432 693410
rect 675312 693342 675340 693382
rect 675128 693314 675340 693342
rect 675404 693328 675432 693382
rect 674930 693288 674986 693297
rect 674930 693223 674986 693232
rect 674944 690894 674972 693223
rect 675128 693025 675156 693314
rect 675114 693016 675170 693025
rect 675114 692951 675170 692960
rect 674944 690866 675418 690894
rect 675404 690169 675432 690336
rect 675390 690160 675446 690169
rect 675390 690095 675446 690104
rect 675312 689710 675432 689738
rect 675312 689625 675340 689710
rect 675404 689656 675432 689710
rect 675298 689616 675354 689625
rect 675298 689551 675354 689560
rect 675128 689030 675418 689058
rect 674930 688936 674986 688945
rect 674930 688871 674986 688880
rect 674944 687154 674972 688871
rect 675128 688673 675156 689030
rect 675298 688936 675354 688945
rect 675298 688871 675354 688880
rect 675114 688664 675170 688673
rect 675114 688599 675170 688608
rect 674944 687126 675156 687154
rect 674838 686488 674894 686497
rect 674838 686423 674894 686432
rect 674852 683114 674880 686423
rect 675128 685998 675156 687126
rect 675312 687018 675340 688871
rect 675496 687449 675524 687820
rect 675482 687440 675538 687449
rect 675482 687375 675538 687384
rect 675312 686990 675524 687018
rect 675496 686664 675524 686990
rect 675128 685970 675418 685998
rect 675482 685808 675538 685817
rect 675482 685743 675538 685752
rect 675206 685536 675262 685545
rect 675206 685471 675262 685480
rect 675220 684570 675248 685471
rect 675496 685372 675524 685743
rect 675220 684542 675432 684570
rect 675404 684148 675432 684542
rect 674852 683086 675248 683114
rect 674668 656866 674880 656894
rect 674208 652038 674420 652066
rect 674208 648530 674236 652038
rect 674562 648952 674618 648961
rect 674562 648887 674618 648896
rect 674208 648502 674512 648530
rect 674116 647206 674328 647234
rect 674300 641866 674328 647206
rect 674484 645153 674512 648502
rect 674576 645854 674604 648887
rect 674852 648802 674880 656866
rect 675022 651536 675078 651545
rect 675022 651471 675078 651480
rect 674668 648774 674880 648802
rect 674668 647170 674696 648774
rect 674838 647592 674894 647601
rect 674838 647527 674894 647536
rect 674668 647142 674788 647170
rect 674576 645826 674696 645854
rect 674470 645144 674526 645153
rect 674470 645079 674526 645088
rect 674300 641838 674420 641866
rect 674194 641744 674250 641753
rect 674194 641679 674250 641688
rect 673932 620986 674052 621014
rect 673932 617409 673960 620986
rect 673918 617400 673974 617409
rect 673918 617335 673974 617344
rect 674010 599584 674066 599593
rect 674010 599519 674066 599528
rect 674024 599434 674052 599519
rect 673656 598862 673776 598890
rect 673840 599406 674052 599434
rect 673656 595649 673684 598862
rect 673642 595640 673698 595649
rect 673642 595575 673698 595584
rect 673840 595354 673868 599406
rect 674010 599312 674066 599321
rect 674010 599247 674066 599256
rect 674024 595377 674052 599247
rect 674208 598934 674236 641679
rect 674392 641186 674420 641838
rect 674300 641158 674420 641186
rect 674300 630674 674328 641158
rect 674668 640334 674696 645826
rect 674576 640306 674696 640334
rect 674300 630646 674420 630674
rect 674392 624889 674420 630646
rect 674378 624880 674434 624889
rect 674378 624815 674434 624824
rect 674378 606520 674434 606529
rect 674378 606455 674434 606464
rect 674392 605834 674420 606455
rect 674392 605806 674512 605834
rect 674208 598906 674328 598934
rect 673564 595326 673868 595354
rect 674010 595368 674066 595377
rect 673564 591546 673592 595326
rect 674010 595303 674066 595312
rect 674300 592929 674328 598906
rect 674286 592920 674342 592929
rect 674286 592855 674342 592864
rect 673918 591696 673974 591705
rect 673918 591631 673974 591640
rect 673564 591518 673868 591546
rect 673472 591382 673684 591410
rect 673656 528329 673684 591382
rect 673840 532545 673868 591518
rect 673932 582374 673960 591631
rect 674484 582374 674512 605806
rect 674576 596174 674604 640306
rect 674760 618633 674788 647142
rect 674852 647034 674880 647527
rect 674852 647006 674972 647034
rect 674944 644065 674972 647006
rect 675036 644314 675064 651471
rect 675220 650185 675248 683086
rect 683210 682680 683266 682689
rect 683210 682615 683266 682624
rect 676494 673160 676550 673169
rect 676494 673095 676550 673104
rect 676508 671129 676536 673095
rect 676494 671120 676550 671129
rect 676494 671055 676550 671064
rect 676494 670304 676550 670313
rect 676494 670239 676550 670248
rect 676508 669497 676536 670239
rect 676494 669488 676550 669497
rect 676494 669423 676550 669432
rect 676494 666224 676550 666233
rect 676494 666159 676550 666168
rect 676508 665417 676536 666159
rect 676494 665408 676550 665417
rect 676494 665343 676550 665352
rect 683224 664601 683252 682615
rect 683670 682408 683726 682417
rect 683670 682343 683726 682352
rect 683486 681048 683542 681057
rect 683486 680983 683542 680992
rect 683210 664592 683266 664601
rect 683210 664527 683266 664536
rect 683500 662969 683528 680983
rect 683684 667049 683712 682343
rect 703694 671908 703722 672044
rect 704154 671908 704182 672044
rect 704614 671908 704642 672044
rect 705074 671908 705102 672044
rect 705534 671908 705562 672044
rect 705994 671908 706022 672044
rect 706454 671908 706482 672044
rect 706914 671908 706942 672044
rect 707374 671908 707402 672044
rect 707834 671908 707862 672044
rect 708294 671908 708322 672044
rect 708754 671908 708782 672044
rect 709214 671908 709242 672044
rect 683670 667040 683726 667049
rect 683670 666975 683726 666984
rect 683486 662960 683542 662969
rect 683486 662895 683542 662904
rect 675390 654256 675446 654265
rect 675390 654191 675446 654200
rect 675404 654134 675432 654191
rect 675312 654106 675432 654134
rect 675312 653018 675340 654106
rect 675312 652990 675432 653018
rect 675404 652460 675432 652990
rect 675588 652905 675616 653140
rect 675574 652896 675630 652905
rect 675574 652831 675630 652840
rect 675404 651545 675432 651848
rect 675390 651536 675446 651545
rect 675390 651471 675446 651480
rect 675206 650176 675262 650185
rect 675206 650111 675262 650120
rect 675128 649998 675340 650026
rect 675128 645810 675156 649998
rect 675312 649994 675340 649998
rect 675404 649994 675432 650012
rect 675312 649966 675432 649994
rect 675404 648961 675432 649468
rect 675390 648952 675446 648961
rect 675390 648887 675446 648896
rect 675496 648689 675524 648788
rect 675482 648680 675538 648689
rect 675482 648615 675538 648624
rect 675496 647873 675524 648176
rect 675482 647864 675538 647873
rect 675482 647799 675538 647808
rect 675298 647248 675354 647257
rect 675298 647183 675354 647192
rect 675312 646105 675340 647183
rect 675298 646096 675354 646105
rect 675298 646031 675354 646040
rect 675482 645824 675538 645833
rect 675128 645782 675482 645810
rect 675482 645759 675538 645768
rect 675496 645425 675524 645660
rect 675758 645552 675814 645561
rect 675758 645487 675814 645496
rect 675482 645416 675538 645425
rect 675482 645351 675538 645360
rect 675772 645116 675800 645487
rect 675772 644337 675800 644475
rect 675298 644328 675354 644337
rect 675036 644286 675298 644314
rect 675298 644263 675354 644272
rect 675758 644328 675814 644337
rect 675758 644263 675814 644272
rect 674930 644056 674986 644065
rect 674930 643991 674986 644000
rect 675114 643784 675170 643793
rect 675114 643719 675170 643728
rect 675128 641594 675156 643719
rect 675496 643521 675524 643824
rect 675482 643512 675538 643521
rect 675482 643447 675538 643456
rect 675312 642621 675418 642649
rect 675312 641753 675340 642621
rect 675298 641744 675354 641753
rect 675298 641679 675354 641688
rect 675128 641566 675340 641594
rect 675312 641458 675340 641566
rect 675312 641430 675418 641458
rect 674930 640792 674986 640801
rect 674930 640727 674986 640736
rect 674944 631417 674972 640727
rect 675404 640529 675432 640795
rect 675390 640520 675446 640529
rect 675390 640455 675446 640464
rect 675404 639826 675432 640152
rect 675220 639798 675432 639826
rect 674930 631408 674986 631417
rect 674930 631343 674986 631352
rect 674746 618624 674802 618633
rect 674746 618559 674802 618568
rect 674838 603120 674894 603129
rect 674838 603055 674894 603064
rect 674852 601089 674880 603055
rect 675022 601760 675078 601769
rect 675022 601695 675078 601704
rect 674838 601080 674894 601089
rect 674838 601015 674894 601024
rect 675036 600545 675064 601695
rect 675022 600536 675078 600545
rect 675022 600471 675078 600480
rect 675022 599040 675078 599049
rect 675022 598975 675078 598984
rect 675036 596873 675064 598975
rect 675022 596864 675078 596873
rect 675022 596799 675078 596808
rect 675220 596174 675248 639798
rect 675496 638761 675524 638928
rect 675482 638752 675538 638761
rect 675482 638687 675538 638696
rect 675390 638072 675446 638081
rect 675390 638007 675446 638016
rect 675404 637574 675432 638007
rect 677506 637936 677562 637945
rect 677506 637871 677562 637880
rect 675758 637664 675814 637673
rect 675758 637599 675814 637608
rect 674576 596146 674696 596174
rect 674668 592657 674696 596146
rect 675128 596146 675248 596174
rect 675312 637546 675432 637574
rect 674930 595504 674986 595513
rect 674930 595439 674986 595448
rect 674654 592648 674710 592657
rect 674654 592583 674710 592592
rect 674944 592034 674972 595439
rect 675128 592498 675156 596146
rect 675312 595898 675340 637546
rect 675772 631417 675800 637599
rect 675758 631408 675814 631417
rect 675758 631343 675814 631352
rect 675850 627872 675906 627881
rect 675850 627807 675906 627816
rect 675864 626618 675892 627807
rect 675852 626612 675904 626618
rect 675852 626554 675904 626560
rect 676496 626612 676548 626618
rect 676496 626554 676548 626560
rect 676508 625705 676536 626554
rect 676494 625696 676550 625705
rect 676494 625631 676550 625640
rect 677520 622033 677548 637871
rect 683394 636848 683450 636857
rect 683394 636783 683450 636792
rect 683210 635488 683266 635497
rect 683210 635423 683266 635432
rect 683224 624481 683252 635423
rect 683408 634814 683436 636783
rect 683408 634786 683620 634814
rect 683394 624880 683450 624889
rect 683394 624815 683450 624824
rect 683210 624472 683266 624481
rect 683210 624407 683266 624416
rect 677506 622024 677562 622033
rect 677506 621959 677562 621968
rect 676494 621616 676550 621625
rect 676494 621551 676550 621560
rect 676508 621217 676536 621551
rect 676494 621208 676550 621217
rect 676494 621143 676550 621152
rect 683408 617137 683436 624815
rect 683592 617953 683620 634786
rect 703694 626892 703722 627028
rect 704154 626892 704182 627028
rect 704614 626892 704642 627028
rect 705074 626892 705102 627028
rect 705534 626892 705562 627028
rect 705994 626892 706022 627028
rect 706454 626892 706482 627028
rect 706914 626892 706942 627028
rect 707374 626892 707402 627028
rect 707834 626892 707862 627028
rect 708294 626892 708322 627028
rect 708754 626892 708782 627028
rect 709214 626892 709242 627028
rect 683578 617944 683634 617953
rect 683578 617879 683634 617888
rect 683394 617128 683450 617137
rect 683394 617063 683450 617072
rect 675482 608288 675538 608297
rect 675482 608223 675538 608232
rect 675496 608124 675524 608223
rect 675482 608016 675538 608025
rect 675482 607951 675538 607960
rect 675496 607479 675524 607951
rect 675496 606529 675524 606832
rect 675482 606520 675538 606529
rect 675482 606455 675538 606464
rect 675496 604761 675524 604996
rect 675482 604752 675538 604761
rect 675482 604687 675538 604696
rect 675496 604353 675524 604452
rect 675482 604344 675538 604353
rect 675482 604279 675538 604288
rect 675496 603537 675524 603772
rect 675482 603528 675538 603537
rect 675482 603463 675538 603472
rect 675496 602857 675524 603160
rect 675482 602848 675538 602857
rect 675482 602783 675538 602792
rect 675482 601080 675538 601089
rect 675482 601015 675538 601024
rect 675496 600644 675524 601015
rect 675482 600536 675538 600545
rect 675482 600471 675538 600480
rect 675496 600100 675524 600471
rect 675496 599321 675524 599488
rect 675482 599312 675538 599321
rect 675482 599247 675538 599256
rect 675666 599176 675722 599185
rect 675666 599111 675722 599120
rect 675680 598808 675708 599111
rect 675482 598088 675538 598097
rect 675482 598023 675538 598032
rect 675496 597652 675524 598023
rect 675482 596864 675538 596873
rect 675482 596799 675538 596808
rect 675496 596428 675524 596799
rect 675220 595870 675340 595898
rect 675220 592634 675248 595870
rect 675404 595513 675432 595816
rect 675390 595504 675446 595513
rect 675390 595439 675446 595448
rect 675496 594833 675524 595136
rect 675482 594824 675538 594833
rect 675482 594759 675538 594768
rect 675404 593745 675432 593980
rect 675390 593736 675446 593745
rect 675390 593671 675446 593680
rect 683302 592920 683358 592929
rect 683302 592855 683358 592864
rect 675220 592606 676168 592634
rect 675128 592470 675984 592498
rect 675758 592376 675814 592385
rect 675758 592311 675814 592320
rect 675574 592104 675630 592113
rect 675574 592039 675630 592048
rect 674944 592006 675064 592034
rect 673932 582346 674052 582374
rect 674024 545737 674052 582346
rect 674392 582346 674512 582374
rect 674194 552120 674250 552129
rect 674194 552055 674250 552064
rect 674010 545728 674066 545737
rect 674010 545663 674066 545672
rect 674010 535392 674066 535401
rect 674010 535327 674066 535336
rect 674024 534177 674052 535327
rect 674010 534168 674066 534177
rect 674010 534103 674066 534112
rect 673826 532536 673882 532545
rect 673826 532471 673882 532480
rect 673642 528320 673698 528329
rect 673642 528255 673698 528264
rect 674208 483993 674236 552055
rect 674392 547097 674420 582346
rect 675036 563054 675064 592006
rect 675588 586265 675616 592039
rect 675574 586256 675630 586265
rect 675574 586191 675630 586200
rect 675772 576609 675800 592311
rect 675956 591394 675984 592470
rect 675944 591388 675996 591394
rect 675944 591330 675996 591336
rect 676140 591258 676168 592606
rect 679624 591388 679676 591394
rect 679624 591330 679676 591336
rect 676128 591252 676180 591258
rect 676128 591194 676180 591200
rect 676034 582992 676090 583001
rect 676034 582927 676090 582936
rect 676048 580281 676076 582927
rect 676034 580272 676090 580281
rect 676034 580207 676090 580216
rect 675758 576600 675814 576609
rect 675758 576535 675814 576544
rect 679636 571334 679664 591330
rect 682384 591252 682436 591258
rect 682384 591194 682436 591200
rect 682396 575657 682424 591194
rect 682382 575648 682438 575657
rect 682382 575583 682438 575592
rect 683316 573209 683344 592855
rect 683486 592648 683542 592657
rect 683486 592583 683542 592592
rect 683500 574025 683528 592583
rect 683762 591424 683818 591433
rect 683762 591359 683818 591368
rect 683486 574016 683542 574025
rect 683486 573951 683542 573960
rect 683302 573200 683358 573209
rect 683302 573135 683358 573144
rect 683776 572393 683804 591359
rect 703694 581740 703722 581876
rect 704154 581740 704182 581876
rect 704614 581740 704642 581876
rect 705074 581740 705102 581876
rect 705534 581740 705562 581876
rect 705994 581740 706022 581876
rect 706454 581740 706482 581876
rect 706914 581740 706942 581876
rect 707374 581740 707402 581876
rect 707834 581740 707862 581876
rect 708294 581740 708322 581876
rect 708754 581740 708782 581876
rect 709214 581740 709242 581876
rect 683762 572384 683818 572393
rect 683762 572319 683818 572328
rect 679624 571328 679676 571334
rect 679624 571270 679676 571276
rect 683120 571328 683172 571334
rect 683120 571270 683172 571276
rect 683132 570761 683160 571270
rect 683118 570752 683174 570761
rect 683118 570687 683174 570696
rect 675206 564496 675262 564505
rect 675206 564431 675262 564440
rect 674852 563026 675064 563054
rect 674654 558376 674710 558385
rect 674654 558311 674710 558320
rect 674378 547088 674434 547097
rect 674378 547023 674434 547032
rect 674470 535120 674526 535129
rect 674470 535055 674526 535064
rect 674484 534177 674512 535055
rect 674470 534168 674526 534177
rect 674470 534103 674526 534112
rect 674470 532264 674526 532273
rect 674470 532199 674526 532208
rect 674484 531457 674512 532199
rect 674470 531448 674526 531457
rect 674470 531383 674526 531392
rect 674668 484401 674696 558311
rect 674852 547369 674880 563026
rect 675220 562306 675248 564431
rect 675390 563136 675446 563145
rect 675390 563071 675446 563080
rect 675404 562904 675432 563071
rect 675220 562278 675418 562306
rect 675496 561241 675524 561612
rect 675482 561232 675538 561241
rect 675482 561167 675538 561176
rect 675312 559830 675432 559858
rect 675312 559790 675340 559830
rect 675036 559762 675340 559790
rect 675404 559776 675432 559830
rect 675036 548162 675064 559762
rect 675312 559218 675418 559246
rect 675312 559065 675340 559218
rect 675298 559056 675354 559065
rect 675298 558991 675354 559000
rect 675206 558784 675262 558793
rect 675206 558719 675262 558728
rect 675220 557954 675248 558719
rect 675404 558385 675432 558620
rect 675390 558376 675446 558385
rect 675390 558311 675446 558320
rect 675220 557926 675418 557954
rect 675206 556200 675262 556209
rect 675206 556135 675262 556144
rect 675220 553670 675248 556135
rect 675404 555257 675432 555492
rect 675390 555248 675446 555257
rect 675390 555183 675446 555192
rect 675772 554713 675800 554919
rect 675758 554704 675814 554713
rect 675758 554639 675814 554648
rect 675404 553897 675432 554268
rect 675390 553888 675446 553897
rect 675390 553823 675446 553832
rect 675220 553642 675340 553670
rect 675312 553602 675340 553642
rect 675404 553602 675432 553656
rect 675312 553574 675432 553602
rect 675206 553480 675262 553489
rect 675206 553415 675262 553424
rect 675220 551253 675248 553415
rect 675404 552129 675432 552432
rect 675390 552120 675446 552129
rect 675390 552055 675446 552064
rect 675220 551225 675418 551253
rect 675758 550760 675814 550769
rect 675758 550695 675814 550704
rect 675772 550596 675800 550695
rect 675404 549681 675432 549951
rect 675390 549672 675446 549681
rect 675390 549607 675446 549616
rect 675496 548457 675524 548760
rect 675482 548448 675538 548457
rect 675482 548383 675538 548392
rect 675036 548134 675340 548162
rect 675312 548026 675340 548134
rect 675312 547998 675432 548026
rect 675114 547904 675170 547913
rect 675114 547839 675170 547848
rect 675128 547754 675156 547839
rect 675036 547726 675156 547754
rect 674838 547360 674894 547369
rect 674838 547295 674894 547304
rect 674838 543824 674894 543833
rect 674838 543759 674894 543768
rect 674852 540974 674880 543759
rect 674852 540946 674972 540974
rect 674944 503849 674972 540946
rect 675036 538214 675064 547726
rect 675206 547632 675262 547641
rect 675206 547567 675262 547576
rect 675036 538186 675156 538214
rect 674930 503840 674986 503849
rect 674930 503775 674986 503784
rect 675128 503690 675156 538186
rect 675220 503826 675248 547567
rect 675404 540974 675432 547998
rect 675852 547664 675904 547670
rect 675852 547606 675904 547612
rect 678244 547664 678296 547670
rect 678244 547606 678296 547612
rect 675864 547369 675892 547606
rect 675850 547360 675906 547369
rect 675850 547295 675906 547304
rect 676402 546272 676458 546281
rect 676402 546207 676458 546216
rect 675312 540946 675432 540974
rect 675312 511994 675340 540946
rect 676034 537840 676090 537849
rect 676034 537775 676090 537784
rect 676048 535741 676076 537775
rect 676034 535732 676090 535741
rect 676034 535667 676090 535676
rect 675850 532536 675906 532545
rect 675850 532471 675906 532480
rect 675864 532302 675892 532471
rect 675852 532296 675904 532302
rect 675852 532238 675904 532244
rect 675758 529408 675814 529417
rect 675758 529343 675814 529352
rect 675942 529408 675998 529417
rect 675942 529343 675998 529352
rect 675772 528805 675800 529343
rect 675758 528796 675814 528805
rect 675758 528731 675814 528740
rect 675956 528601 675984 529343
rect 675942 528592 675998 528601
rect 675942 528527 675998 528536
rect 675852 518832 675904 518838
rect 675852 518774 675904 518780
rect 675864 511994 675892 518774
rect 675312 511966 675432 511994
rect 675220 503798 675340 503826
rect 675036 503662 675156 503690
rect 675036 503577 675064 503662
rect 675022 503568 675078 503577
rect 675022 503503 675078 503512
rect 675312 503418 675340 503798
rect 675036 503390 675340 503418
rect 675036 503305 675064 503390
rect 675022 503296 675078 503305
rect 675022 503231 675078 503240
rect 675404 502334 675432 511966
rect 675588 511966 675892 511994
rect 675588 502334 675616 511966
rect 675850 503840 675906 503849
rect 675850 503775 675906 503784
rect 675864 503674 675892 503775
rect 675852 503668 675904 503674
rect 675852 503610 675904 503616
rect 676034 503568 676090 503577
rect 676034 503503 676036 503512
rect 676088 503503 676090 503512
rect 676036 503474 676088 503480
rect 676034 503296 676090 503305
rect 676034 503231 676090 503240
rect 675312 502306 675432 502334
rect 675496 502306 675616 502334
rect 675852 502376 675904 502382
rect 675852 502318 675904 502324
rect 674930 500984 674986 500993
rect 674930 500919 674986 500928
rect 674654 484392 674710 484401
rect 674654 484327 674710 484336
rect 674194 483984 674250 483993
rect 674194 483919 674250 483928
rect 674746 464808 674802 464817
rect 674746 464743 674802 464752
rect 674760 456929 674788 464743
rect 673826 456920 673882 456929
rect 673826 456855 673882 456864
rect 674746 456920 674802 456929
rect 674746 456855 674802 456864
rect 673840 456074 673868 456855
rect 673946 456512 674002 456521
rect 673946 456447 673948 456456
rect 674000 456447 674002 456456
rect 673948 456418 674000 456424
rect 673828 456068 673880 456074
rect 673828 456010 673880 456016
rect 673380 455926 673500 455954
rect 673472 455870 673500 455926
rect 673460 455864 673512 455870
rect 673460 455806 673512 455812
rect 673596 455696 673652 455705
rect 673596 455631 673598 455640
rect 673650 455631 673652 455640
rect 673598 455602 673650 455608
rect 673504 455424 673560 455433
rect 673504 455359 673506 455368
rect 673558 455359 673560 455368
rect 673506 455330 673558 455336
rect 673388 455184 673440 455190
rect 673386 455152 673388 455161
rect 673440 455152 673442 455161
rect 673386 455087 673442 455096
rect 674944 454889 674972 500919
rect 675312 486441 675340 502306
rect 675298 486432 675354 486441
rect 675298 486367 675354 486376
rect 673162 454880 673218 454889
rect 673162 454815 673164 454824
rect 673216 454815 673218 454824
rect 674930 454880 674986 454889
rect 674930 454815 674986 454824
rect 673164 454786 673216 454792
rect 673046 454640 673098 454646
rect 673044 454608 673046 454617
rect 675496 454617 675524 502306
rect 675864 485774 675892 502318
rect 676048 500954 676076 503231
rect 676036 500948 676088 500954
rect 676036 500890 676088 500896
rect 676416 495434 676444 546207
rect 676588 532296 676640 532302
rect 676586 532264 676588 532273
rect 676640 532264 676642 532273
rect 676586 532199 676642 532208
rect 678256 531457 678284 547606
rect 683210 547088 683266 547097
rect 683210 547023 683266 547032
rect 679622 546544 679678 546553
rect 679622 546479 679678 546488
rect 678242 531448 678298 531457
rect 678242 531383 678298 531392
rect 679636 531049 679664 546479
rect 683224 531865 683252 547023
rect 683394 545728 683450 545737
rect 683394 545663 683450 545672
rect 683210 531856 683266 531865
rect 683210 531791 683266 531800
rect 679622 531040 679678 531049
rect 679622 530975 679678 530984
rect 683408 527785 683436 545663
rect 703694 536724 703722 536860
rect 704154 536724 704182 536860
rect 704614 536724 704642 536860
rect 705074 536724 705102 536860
rect 705534 536724 705562 536860
rect 705994 536724 706022 536860
rect 706454 536724 706482 536860
rect 706914 536724 706942 536860
rect 707374 536724 707402 536860
rect 707834 536724 707862 536860
rect 708294 536724 708322 536860
rect 708754 536724 708782 536860
rect 709214 536724 709242 536860
rect 683578 532264 683634 532273
rect 683578 532199 683634 532208
rect 683394 527776 683450 527785
rect 683394 527711 683450 527720
rect 683592 526561 683620 532199
rect 683578 526552 683634 526561
rect 683578 526487 683634 526496
rect 676862 525736 676918 525745
rect 676862 525671 676918 525680
rect 676876 502382 676904 525671
rect 677874 524512 677930 524521
rect 677874 524447 677930 524456
rect 677888 518838 677916 524447
rect 677876 518832 677928 518838
rect 677876 518774 677928 518780
rect 683210 503704 683266 503713
rect 679624 503668 679676 503674
rect 683210 503639 683266 503648
rect 679624 503610 679676 503616
rect 676864 502376 676916 502382
rect 676864 502318 676916 502324
rect 676416 495406 676812 495434
rect 676034 494048 676090 494057
rect 676034 493983 676090 493992
rect 676048 492726 676076 493983
rect 676036 492720 676088 492726
rect 676036 492662 676088 492668
rect 675680 485746 675892 485774
rect 673098 454608 673100 454617
rect 673044 454543 673100 454552
rect 675482 454608 675538 454617
rect 675482 454543 675538 454552
rect 672954 454368 673006 454374
rect 672952 454336 672954 454345
rect 675680 454345 675708 485746
rect 675850 481944 675906 481953
rect 675850 481879 675906 481888
rect 673006 454336 673008 454345
rect 672952 454271 673008 454280
rect 675666 454336 675722 454345
rect 675666 454271 675722 454280
rect 672816 454096 672868 454102
rect 672814 454064 672816 454073
rect 672868 454064 672870 454073
rect 672814 453999 672870 454008
rect 675864 453801 675892 481879
rect 676034 480720 676090 480729
rect 676034 480655 676090 480664
rect 676048 454073 676076 480655
rect 676784 455705 676812 495406
rect 677322 492416 677378 492425
rect 677322 492351 677378 492360
rect 676954 488880 677010 488889
rect 676954 488815 677010 488824
rect 676968 485797 676996 488815
rect 677336 487257 677364 492351
rect 677322 487248 677378 487257
rect 677322 487183 677378 487192
rect 679636 486849 679664 503610
rect 682384 503532 682436 503538
rect 682384 503474 682436 503480
rect 681004 500948 681056 500954
rect 681004 500890 681056 500896
rect 681016 487665 681044 500890
rect 681002 487656 681058 487665
rect 681002 487591 681058 487600
rect 679622 486840 679678 486849
rect 679622 486775 679678 486784
rect 676954 485788 677010 485797
rect 676954 485723 677010 485732
rect 682396 481545 682424 503474
rect 683224 482769 683252 503639
rect 683578 494728 683634 494737
rect 683578 494663 683634 494672
rect 683396 492720 683448 492726
rect 683396 492662 683448 492668
rect 683408 491745 683436 492662
rect 683394 491736 683450 491745
rect 683394 491671 683450 491680
rect 683592 491337 683620 494663
rect 703694 492796 703722 492864
rect 704154 492796 704182 492864
rect 704614 492796 704642 492864
rect 705074 492796 705102 492864
rect 705534 492796 705562 492864
rect 705994 492796 706022 492864
rect 706454 492796 706482 492864
rect 706914 492796 706942 492864
rect 707374 492796 707402 492864
rect 707834 492796 707862 492864
rect 708294 492796 708322 492864
rect 708754 492796 708782 492864
rect 709214 492796 709242 492864
rect 683578 491328 683634 491337
rect 683578 491263 683634 491272
rect 683210 482760 683266 482769
rect 683210 482695 683266 482704
rect 682382 481536 682438 481545
rect 682382 481471 682438 481480
rect 676770 455696 676826 455705
rect 676770 455631 676826 455640
rect 676034 454064 676090 454073
rect 676034 453999 676090 454008
rect 675850 453792 675906 453801
rect 675850 453727 675906 453736
rect 683118 406328 683174 406337
rect 683118 406263 683174 406272
rect 676034 405648 676090 405657
rect 676034 405583 676090 405592
rect 676048 403481 676076 405583
rect 676034 403472 676090 403481
rect 676034 403407 676090 403416
rect 683132 403345 683160 406263
rect 703694 404532 703722 404668
rect 704154 404532 704182 404668
rect 704614 404532 704642 404668
rect 705074 404532 705102 404668
rect 705534 404532 705562 404668
rect 705994 404532 706022 404668
rect 706454 404532 706482 404668
rect 706914 404532 706942 404668
rect 707374 404532 707402 404668
rect 707834 404532 707862 404668
rect 708294 404532 708322 404668
rect 708754 404532 708782 404668
rect 709214 404532 709242 404668
rect 683118 403336 683174 403345
rect 683118 403271 683174 403280
rect 674194 402248 674250 402257
rect 674194 402183 674250 402192
rect 672630 400072 672686 400081
rect 672630 400007 672686 400016
rect 673182 398848 673238 398857
rect 673182 398783 673238 398792
rect 672998 397216 673054 397225
rect 672998 397151 673054 397160
rect 672722 392592 672778 392601
rect 672722 392527 672778 392536
rect 672446 355872 672502 355881
rect 672446 355807 672502 355816
rect 672538 354648 672594 354657
rect 672538 354583 672594 354592
rect 672170 353424 672226 353433
rect 672170 353359 672226 353368
rect 671986 348936 672042 348945
rect 671986 348871 672042 348880
rect 672000 332353 672028 348871
rect 672184 340785 672212 353359
rect 672354 348528 672410 348537
rect 672354 348463 672410 348472
rect 672170 340776 672226 340785
rect 672170 340711 672226 340720
rect 671986 332344 672042 332353
rect 671986 332279 672042 332288
rect 672170 311264 672226 311273
rect 672170 311199 672226 311208
rect 671986 302016 672042 302025
rect 671986 301951 672042 301960
rect 671342 269784 671398 269793
rect 671342 269719 671398 269728
rect 671342 264072 671398 264081
rect 671342 264007 671398 264016
rect 671356 238241 671384 264007
rect 671710 262032 671766 262041
rect 671710 261967 671766 261976
rect 671526 257952 671582 257961
rect 671526 257887 671582 257896
rect 671540 241505 671568 257887
rect 671724 244769 671752 261967
rect 671710 244760 671766 244769
rect 671710 244695 671766 244704
rect 671526 241496 671582 241505
rect 671526 241431 671582 241440
rect 671342 238232 671398 238241
rect 671342 238167 671398 238176
rect 671252 237652 671304 237658
rect 671252 237594 671304 237600
rect 671068 235884 671120 235890
rect 671068 235826 671120 235832
rect 671080 234614 671108 235826
rect 671264 234614 671292 237594
rect 671436 237176 671488 237182
rect 671436 237118 671488 237124
rect 671080 234586 671200 234614
rect 671264 234586 671384 234614
rect 670792 234048 670844 234054
rect 670712 233996 670792 234002
rect 670712 233990 670844 233996
rect 670712 233974 670832 233990
rect 670712 215294 670740 233974
rect 671172 233209 671200 234586
rect 671158 233200 671214 233209
rect 671158 233135 671214 233144
rect 671160 233028 671212 233034
rect 671160 232970 671212 232976
rect 670884 232824 670936 232830
rect 670884 232766 670936 232772
rect 670896 224346 670924 232766
rect 671172 228426 671200 232970
rect 671172 228398 671292 228426
rect 671068 228268 671120 228274
rect 671068 228210 671120 228216
rect 671080 225729 671108 228210
rect 671066 225720 671122 225729
rect 671066 225655 671122 225664
rect 671066 225312 671122 225321
rect 671066 225247 671068 225256
rect 671120 225247 671122 225256
rect 671068 225218 671120 225224
rect 671068 224936 671120 224942
rect 671066 224904 671068 224913
rect 671120 224904 671122 224913
rect 671066 224839 671122 224848
rect 671020 224496 671076 224505
rect 671020 224431 671022 224440
rect 671074 224431 671076 224440
rect 671022 224402 671074 224408
rect 670896 224318 671016 224346
rect 670712 215266 670832 215294
rect 670606 211168 670662 211177
rect 670606 211103 670662 211112
rect 670606 210896 670662 210905
rect 670606 210831 670662 210840
rect 670620 190369 670648 210831
rect 670804 199374 670832 215266
rect 670792 199368 670844 199374
rect 670792 199310 670844 199316
rect 670988 194426 671016 224318
rect 671264 215294 671292 228398
rect 670804 194398 671016 194426
rect 671172 215266 671292 215294
rect 670804 194342 670832 194398
rect 670792 194336 670844 194342
rect 670792 194278 670844 194284
rect 671172 190454 671200 215266
rect 670804 190426 671200 190454
rect 670606 190360 670662 190369
rect 670606 190295 670662 190304
rect 670804 189446 670832 190426
rect 670792 189440 670844 189446
rect 670792 189382 670844 189388
rect 670606 170368 670662 170377
rect 670606 170303 670662 170312
rect 670332 169720 670384 169726
rect 670332 169662 670384 169668
rect 670330 165608 670386 165617
rect 670330 165543 670386 165552
rect 670148 164960 670200 164966
rect 670148 164902 670200 164908
rect 669964 136400 670016 136406
rect 669964 136342 670016 136348
rect 669780 125588 669832 125594
rect 669780 125530 669832 125536
rect 669962 122768 670018 122777
rect 669962 122703 670018 122712
rect 668582 120864 668638 120873
rect 668582 120799 668638 120808
rect 668950 120184 669006 120193
rect 668950 120119 669006 120128
rect 667938 119232 667994 119241
rect 667938 119167 667994 119176
rect 668032 118516 668084 118522
rect 668032 118458 668084 118464
rect 668044 117609 668072 118458
rect 668030 117600 668086 117609
rect 668030 117535 668086 117544
rect 668964 114345 668992 120119
rect 668950 114336 669006 114345
rect 668950 114271 669006 114280
rect 669976 114170 670004 122703
rect 670344 118522 670372 165543
rect 670620 147665 670648 170303
rect 671356 147674 671384 234586
rect 671448 222194 671476 237118
rect 671620 236972 671672 236978
rect 671620 236914 671672 236920
rect 671632 225604 671660 236914
rect 671804 234048 671856 234054
rect 671804 233990 671856 233996
rect 671816 233374 671844 233990
rect 671804 233368 671856 233374
rect 671804 233310 671856 233316
rect 671802 231432 671858 231441
rect 671802 231367 671858 231376
rect 671816 228478 671844 231367
rect 671804 228472 671856 228478
rect 671804 228414 671856 228420
rect 671804 227860 671856 227866
rect 671804 227802 671856 227808
rect 671816 226001 671844 227802
rect 672000 227066 672028 301951
rect 672184 266529 672212 311199
rect 672170 266520 672226 266529
rect 672170 266455 672226 266464
rect 672172 238060 672224 238066
rect 672172 238002 672224 238008
rect 672184 234569 672212 238002
rect 672170 234560 672226 234569
rect 672170 234495 672226 234504
rect 672368 231854 672396 348463
rect 672552 310049 672580 354583
rect 672538 310040 672594 310049
rect 672538 309975 672594 309984
rect 672736 251174 672764 392527
rect 673012 378049 673040 397151
rect 672998 378040 673054 378049
rect 672998 377975 673054 377984
rect 673196 364334 673224 398783
rect 673366 396400 673422 396409
rect 673366 396335 673422 396344
rect 673380 382265 673408 396335
rect 673826 396128 673882 396137
rect 673826 396063 673882 396072
rect 673366 382256 673422 382265
rect 673366 382191 673422 382200
rect 673840 381449 673868 396063
rect 674010 395720 674066 395729
rect 674010 395655 674066 395664
rect 673826 381440 673882 381449
rect 673826 381375 673882 381384
rect 674024 375465 674052 395655
rect 674010 375456 674066 375465
rect 674010 375391 674066 375400
rect 673196 364306 673408 364334
rect 673182 355464 673238 355473
rect 673182 355399 673238 355408
rect 672998 351384 673054 351393
rect 672998 351319 673054 351328
rect 673012 338065 673040 351319
rect 672998 338056 673054 338065
rect 672998 337991 673054 338000
rect 673196 310865 673224 355399
rect 673380 355065 673408 364306
rect 674208 357513 674236 402183
rect 674654 401432 674710 401441
rect 674654 401367 674710 401376
rect 674470 394496 674526 394505
rect 674470 394431 674526 394440
rect 674484 377777 674512 394431
rect 674470 377768 674526 377777
rect 674470 377703 674526 377712
rect 674668 364334 674696 401367
rect 676034 399392 676090 399401
rect 676034 399327 676090 399336
rect 675852 395752 675904 395758
rect 675036 395700 675852 395706
rect 675036 395694 675904 395700
rect 675036 395678 675892 395694
rect 675036 382582 675064 395678
rect 676048 395570 676076 399327
rect 676218 398440 676274 398449
rect 676218 398375 676274 398384
rect 675128 395542 676076 395570
rect 675128 384449 675156 395542
rect 676232 393314 676260 398375
rect 676402 398032 676458 398041
rect 676402 397967 676458 397976
rect 676416 395758 676444 397967
rect 681002 397624 681058 397633
rect 681002 397559 681058 397568
rect 676404 395752 676456 395758
rect 676404 395694 676456 395700
rect 675312 393286 676260 393314
rect 675312 386186 675340 393286
rect 681016 387705 681044 397559
rect 681002 387696 681058 387705
rect 681002 387631 681058 387640
rect 675312 386158 675432 386186
rect 675404 385696 675432 386158
rect 675772 384985 675800 385084
rect 675758 384976 675814 384985
rect 675758 384911 675814 384920
rect 675128 384421 675418 384449
rect 675312 382622 675432 382650
rect 675312 382582 675340 382622
rect 675036 382554 675340 382582
rect 675404 382568 675432 382622
rect 675390 382256 675446 382265
rect 675390 382191 675446 382200
rect 675404 382024 675432 382191
rect 675114 381440 675170 381449
rect 675170 381398 675418 381426
rect 675114 381375 675170 381384
rect 675772 380633 675800 380732
rect 675758 380624 675814 380633
rect 675758 380559 675814 380568
rect 675758 378720 675814 378729
rect 675758 378655 675814 378664
rect 675772 378284 675800 378655
rect 675114 377768 675170 377777
rect 675170 377726 675340 377754
rect 675114 377703 675170 377712
rect 675312 377618 675340 377726
rect 675404 377618 675432 377740
rect 675312 377590 675432 377618
rect 675758 377360 675814 377369
rect 675758 377295 675814 377304
rect 675772 377060 675800 377295
rect 675206 376952 675262 376961
rect 675206 376887 675262 376896
rect 675220 373994 675248 376887
rect 675404 376281 675432 376448
rect 675390 376272 675446 376281
rect 675390 376207 675446 376216
rect 675390 375456 675446 375465
rect 675390 375391 675446 375400
rect 675404 375224 675432 375391
rect 675220 373966 675340 373994
rect 675312 373402 675340 373966
rect 675312 373374 675418 373402
rect 675758 373008 675814 373017
rect 675758 372943 675814 372952
rect 675772 372776 675800 372943
rect 675114 372600 675170 372609
rect 675114 372535 675170 372544
rect 675128 371566 675156 372535
rect 675128 371538 675418 371566
rect 674484 364306 674696 364334
rect 674194 357504 674250 357513
rect 674194 357439 674250 357448
rect 674484 356697 674512 364306
rect 675850 360904 675906 360913
rect 675850 360839 675906 360848
rect 675864 357921 675892 360839
rect 676034 360088 676090 360097
rect 676034 360023 676090 360032
rect 676048 358329 676076 360023
rect 703694 359380 703722 359516
rect 704154 359380 704182 359516
rect 704614 359380 704642 359516
rect 705074 359380 705102 359516
rect 705534 359380 705562 359516
rect 705994 359380 706022 359516
rect 706454 359380 706482 359516
rect 706914 359380 706942 359516
rect 707374 359380 707402 359516
rect 707834 359380 707862 359516
rect 708294 359380 708322 359516
rect 708754 359380 708782 359516
rect 709214 359380 709242 359516
rect 676034 358320 676090 358329
rect 676034 358255 676090 358264
rect 675850 357912 675906 357921
rect 675850 357847 675906 357856
rect 674654 357096 674710 357105
rect 674654 357031 674710 357040
rect 674470 356688 674526 356697
rect 674470 356623 674526 356632
rect 674102 356280 674158 356289
rect 674102 356215 674158 356224
rect 673366 355056 673422 355065
rect 673366 354991 673422 355000
rect 673918 352608 673974 352617
rect 673918 352543 673974 352552
rect 673550 352200 673606 352209
rect 673550 352135 673606 352144
rect 673366 349752 673422 349761
rect 673366 349687 673422 349696
rect 673380 335889 673408 349687
rect 673366 335880 673422 335889
rect 673366 335815 673422 335824
rect 673564 325689 673592 352135
rect 673734 350568 673790 350577
rect 673734 350503 673790 350512
rect 673748 331129 673776 350503
rect 673932 336705 673960 352543
rect 673918 336696 673974 336705
rect 673918 336631 673974 336640
rect 673734 331120 673790 331129
rect 673734 331055 673790 331064
rect 673550 325680 673606 325689
rect 673550 325615 673606 325624
rect 673918 312080 673974 312089
rect 673918 312015 673974 312024
rect 673182 310856 673238 310865
rect 673182 310791 673238 310800
rect 673366 304736 673422 304745
rect 673366 304671 673422 304680
rect 672998 304328 673054 304337
rect 672998 304263 673054 304272
rect 673012 287881 673040 304263
rect 673380 290601 673408 304671
rect 673734 303920 673790 303929
rect 673734 303855 673790 303864
rect 673366 290592 673422 290601
rect 673366 290527 673422 290536
rect 672998 287872 673054 287881
rect 672998 287807 673054 287816
rect 673748 286521 673776 303855
rect 673734 286512 673790 286521
rect 673734 286447 673790 286456
rect 673932 267481 673960 312015
rect 674116 311681 674144 356215
rect 674470 349480 674526 349489
rect 674470 349415 674526 349424
rect 674286 347712 674342 347721
rect 674286 347647 674342 347656
rect 674300 327593 674328 347647
rect 674484 332897 674512 349415
rect 674668 340874 674696 357031
rect 676034 353832 676090 353841
rect 676090 353790 676260 353818
rect 676034 353767 676090 353776
rect 675942 349208 675998 349217
rect 676232 349194 676260 353790
rect 675998 349166 676260 349194
rect 675942 349143 675998 349152
rect 674576 340846 674696 340874
rect 674576 338114 674604 340846
rect 675114 340776 675170 340785
rect 675114 340711 675170 340720
rect 675128 340558 675156 340711
rect 675128 340530 675340 340558
rect 675312 340490 675340 340530
rect 675404 340490 675432 340544
rect 675312 340462 675432 340490
rect 675758 340368 675814 340377
rect 675758 340303 675814 340312
rect 675772 339864 675800 340303
rect 675404 339017 675432 339252
rect 675390 339008 675446 339017
rect 675390 338943 675446 338952
rect 674576 338086 674696 338114
rect 674470 332888 674526 332897
rect 674470 332823 674526 332832
rect 674286 327584 674342 327593
rect 674286 327519 674342 327528
rect 674668 312497 674696 338086
rect 675114 338056 675170 338065
rect 675114 337991 675170 338000
rect 675128 336857 675156 337991
rect 675574 337784 675630 337793
rect 675574 337719 675630 337728
rect 675588 337416 675616 337719
rect 675128 336829 675418 336857
rect 675114 336696 675170 336705
rect 675114 336631 675170 336640
rect 675758 336696 675814 336705
rect 675758 336631 675814 336640
rect 675128 333078 675156 336631
rect 675772 336192 675800 336631
rect 675482 335880 675538 335889
rect 675482 335815 675538 335824
rect 675496 335580 675524 335815
rect 675128 333050 675418 333078
rect 675390 332888 675446 332897
rect 675390 332823 675446 332832
rect 675404 332520 675432 332823
rect 675114 332344 675170 332353
rect 675114 332279 675170 332288
rect 675128 331242 675156 332279
rect 675758 332208 675814 332217
rect 675758 332143 675814 332152
rect 675772 331875 675800 332143
rect 675128 331214 675418 331242
rect 675114 331120 675170 331129
rect 675114 331055 675170 331064
rect 675128 330049 675156 331055
rect 675128 330021 675418 330049
rect 675758 328400 675814 328409
rect 675758 328335 675814 328344
rect 675772 328168 675800 328335
rect 675114 327584 675170 327593
rect 675170 327542 675418 327570
rect 675114 327519 675170 327528
rect 675312 326454 675432 326482
rect 675312 326346 675340 326454
rect 675128 326318 675340 326346
rect 675404 326332 675432 326454
rect 675128 325689 675156 326318
rect 675114 325680 675170 325689
rect 675114 325615 675170 325624
rect 676034 315480 676090 315489
rect 676034 315415 676090 315424
rect 676048 313313 676076 315415
rect 703694 314364 703722 314500
rect 704154 314364 704182 314500
rect 704614 314364 704642 314500
rect 705074 314364 705102 314500
rect 705534 314364 705562 314500
rect 705994 314364 706022 314500
rect 706454 314364 706482 314500
rect 706914 314364 706942 314500
rect 707374 314364 707402 314500
rect 707834 314364 707862 314500
rect 708294 314364 708322 314500
rect 708754 314364 708782 314500
rect 709214 314364 709242 314500
rect 676034 313304 676090 313313
rect 676034 313239 676090 313248
rect 674654 312488 674710 312497
rect 674654 312423 674710 312432
rect 674102 311672 674158 311681
rect 674102 311607 674158 311616
rect 674194 310448 674250 310457
rect 674194 310383 674250 310392
rect 673918 267472 673974 267481
rect 673918 267407 673974 267416
rect 674010 266248 674066 266257
rect 674010 266183 674066 266192
rect 673090 263800 673146 263809
rect 673090 263735 673146 263744
rect 672906 259176 672962 259185
rect 672906 259111 672962 259120
rect 672460 251146 672764 251174
rect 672460 241514 672488 251146
rect 672920 243085 672948 259111
rect 673104 258074 673132 263735
rect 673366 260400 673422 260409
rect 673366 260335 673422 260344
rect 672828 243057 672948 243085
rect 673012 258046 673132 258074
rect 672828 242865 672856 243057
rect 672814 242856 672870 242865
rect 672814 242791 672870 242800
rect 672460 241486 672856 241514
rect 672632 236156 672684 236162
rect 672632 236098 672684 236104
rect 672644 234818 672672 236098
rect 672644 234790 672764 234818
rect 672540 234660 672592 234666
rect 672276 231826 672396 231854
rect 672460 234608 672540 234614
rect 672460 234602 672592 234608
rect 672460 234586 672580 234602
rect 672276 228857 672304 231826
rect 672262 228848 672318 228857
rect 672262 228783 672318 228792
rect 672460 227610 672488 234586
rect 671908 227038 672028 227066
rect 672092 227582 672488 227610
rect 672604 227656 672656 227662
rect 672656 227604 672672 227610
rect 672604 227598 672672 227604
rect 672616 227582 672672 227598
rect 671908 226114 671936 227038
rect 672092 226896 672120 227582
rect 672448 227452 672500 227458
rect 672448 227394 672500 227400
rect 672460 227089 672488 227394
rect 672644 227202 672672 227582
rect 672736 227338 672764 234790
rect 672828 231854 672856 241486
rect 673012 237425 673040 258046
rect 673182 257136 673238 257145
rect 673182 257071 673238 257080
rect 672998 237416 673054 237425
rect 672998 237351 673054 237360
rect 673196 236722 673224 257071
rect 673380 245041 673408 260335
rect 673734 259720 673790 259729
rect 673734 259655 673790 259664
rect 673748 245585 673776 259655
rect 674024 258618 674052 266183
rect 674208 265849 674236 310383
rect 674562 309632 674618 309641
rect 674562 309567 674618 309576
rect 674378 305552 674434 305561
rect 674378 305487 674434 305496
rect 674392 292641 674420 305487
rect 674576 302234 674604 309567
rect 674838 309224 674894 309233
rect 674838 309159 674894 309168
rect 674852 303657 674880 309159
rect 676034 308408 676090 308417
rect 676090 308366 676260 308394
rect 676034 308343 676090 308352
rect 676232 304994 676260 308366
rect 681002 307592 681058 307601
rect 681002 307527 681058 307536
rect 678242 307184 678298 307193
rect 678242 307119 678298 307128
rect 676402 305960 676458 305969
rect 676402 305895 676458 305904
rect 675864 304966 676260 304994
rect 674838 303648 674894 303657
rect 674838 303583 674894 303592
rect 675390 303648 675446 303657
rect 675390 303583 675446 303592
rect 674576 302206 674696 302234
rect 674668 294794 674696 302206
rect 675114 301744 675170 301753
rect 675114 301679 675170 301688
rect 675128 298092 675156 301679
rect 675128 298064 675340 298092
rect 674838 296848 674894 296857
rect 674838 296783 674894 296792
rect 674668 294766 674788 294794
rect 674378 292632 674434 292641
rect 674378 292567 674434 292576
rect 674760 292482 674788 294766
rect 674484 292454 674788 292482
rect 674484 287722 674512 292454
rect 674654 292360 674710 292369
rect 674654 292295 674710 292304
rect 674668 289814 674696 292295
rect 674392 287694 674512 287722
rect 674576 289786 674696 289814
rect 674392 277394 674420 287694
rect 674576 285070 674604 289786
rect 674852 288062 674880 296783
rect 675022 296576 675078 296585
rect 675022 296511 675078 296520
rect 675036 292574 675064 296511
rect 675312 296426 675340 298064
rect 675220 296398 675340 296426
rect 675220 294386 675248 296398
rect 675404 296290 675432 303583
rect 675864 302234 675892 304966
rect 676034 303512 676090 303521
rect 676034 303447 676090 303456
rect 675680 302206 675892 302234
rect 675680 299474 675708 302206
rect 676048 302025 676076 303447
rect 676034 302016 676090 302025
rect 676034 301951 676090 301960
rect 676416 301481 676444 305895
rect 676586 305144 676642 305153
rect 676586 305079 676642 305088
rect 676600 301617 676628 305079
rect 676586 301608 676642 301617
rect 676586 301543 676642 301552
rect 676402 301472 676458 301481
rect 676402 301407 676458 301416
rect 675588 299446 675708 299474
rect 675588 296313 675616 299446
rect 675852 298104 675904 298110
rect 675852 298046 675904 298052
rect 675864 296585 675892 298046
rect 676128 297900 676180 297906
rect 676128 297842 676180 297848
rect 676140 296857 676168 297842
rect 678256 297401 678284 307119
rect 678978 306368 679034 306377
rect 678978 306303 679034 306312
rect 678992 298110 679020 306303
rect 678980 298104 679032 298110
rect 678980 298046 679032 298052
rect 681016 297906 681044 307527
rect 681004 297900 681056 297906
rect 681004 297842 681056 297848
rect 678242 297392 678298 297401
rect 678242 297327 678298 297336
rect 676126 296848 676182 296857
rect 676126 296783 676182 296792
rect 675850 296576 675906 296585
rect 675850 296511 675906 296520
rect 675312 296262 675432 296290
rect 675574 296304 675630 296313
rect 675312 294522 675340 296262
rect 675574 296239 675630 296248
rect 675482 295896 675538 295905
rect 675482 295831 675538 295840
rect 675496 295528 675524 295831
rect 675758 295216 675814 295225
rect 675758 295151 675814 295160
rect 675772 294879 675800 295151
rect 675312 294494 675432 294522
rect 675220 294358 675340 294386
rect 675036 292546 675156 292574
rect 675128 291870 675156 292546
rect 675312 292414 675340 294358
rect 675404 294236 675432 294494
rect 675312 292386 675418 292414
rect 675128 291842 675418 291870
rect 675758 291544 675814 291553
rect 675758 291479 675814 291488
rect 675772 291176 675800 291479
rect 675114 290592 675170 290601
rect 675170 290550 675418 290578
rect 675114 290527 675170 290536
rect 675312 288102 675432 288130
rect 675312 288062 675340 288102
rect 674852 288034 675340 288062
rect 675404 288048 675432 288102
rect 675114 287872 675170 287881
rect 675114 287807 675170 287816
rect 675128 287518 675156 287807
rect 675128 287490 675418 287518
rect 675758 287056 675814 287065
rect 675758 286991 675814 287000
rect 675772 286892 675800 286991
rect 675390 286512 675446 286521
rect 675390 286447 675446 286456
rect 675404 286212 675432 286447
rect 674576 285042 675340 285070
rect 675312 285002 675340 285042
rect 675404 285002 675432 285056
rect 675312 284974 675432 285002
rect 675758 283656 675814 283665
rect 675758 283591 675814 283600
rect 675772 283220 675800 283591
rect 675666 282840 675722 282849
rect 675666 282775 675722 282784
rect 675680 282540 675708 282775
rect 675666 281616 675722 281625
rect 675666 281551 675722 281560
rect 675680 281355 675708 281551
rect 674392 277366 674512 277394
rect 674194 265840 674250 265849
rect 674194 265775 674250 265784
rect 674286 265432 674342 265441
rect 674286 265367 674342 265376
rect 674300 261066 674328 265367
rect 674484 265033 674512 277366
rect 683118 271144 683174 271153
rect 683118 271079 683174 271088
rect 676034 269784 676090 269793
rect 676034 269719 676090 269728
rect 676048 268297 676076 269719
rect 676034 268288 676090 268297
rect 676034 268223 676090 268232
rect 683132 268161 683160 271079
rect 703694 269348 703722 269484
rect 704154 269348 704182 269484
rect 704614 269348 704642 269484
rect 705074 269348 705102 269484
rect 705534 269348 705562 269484
rect 705994 269348 706022 269484
rect 706454 269348 706482 269484
rect 706914 269348 706942 269484
rect 707374 269348 707402 269484
rect 707834 269348 707862 269484
rect 708294 269348 708322 269484
rect 708754 269348 708782 269484
rect 709214 269348 709242 269484
rect 683118 268152 683174 268161
rect 683118 268087 683174 268096
rect 674654 267064 674710 267073
rect 674654 266999 674710 267008
rect 674470 265024 674526 265033
rect 674470 264959 674526 264968
rect 674300 261038 674420 261066
rect 674194 260944 674250 260953
rect 674194 260879 674250 260888
rect 674024 258590 674144 258618
rect 673918 258496 673974 258505
rect 673918 258431 673974 258440
rect 673734 245576 673790 245585
rect 673734 245511 673790 245520
rect 673366 245032 673422 245041
rect 673366 244967 673422 244976
rect 673932 244274 673960 258431
rect 674116 258074 674144 258590
rect 674024 258046 674144 258074
rect 674024 253934 674052 258046
rect 674208 253934 674236 260879
rect 674392 253934 674420 261038
rect 674024 253906 674144 253934
rect 674208 253906 674328 253934
rect 674392 253906 674512 253934
rect 674116 244274 674144 253906
rect 674300 246945 674328 253906
rect 674286 246936 674342 246945
rect 674286 246871 674342 246880
rect 673932 244246 674052 244274
rect 674116 244246 674236 244274
rect 673302 237144 673358 237153
rect 673302 237079 673304 237088
rect 673356 237079 673358 237088
rect 673304 237050 673356 237056
rect 673414 236904 673466 236910
rect 673414 236846 673466 236852
rect 673196 236694 673316 236722
rect 673000 235748 673052 235754
rect 673000 235690 673052 235696
rect 673012 231854 673040 235690
rect 673288 235634 673316 236694
rect 673426 236586 673454 236846
rect 673526 236736 673582 236745
rect 673526 236671 673528 236680
rect 673580 236671 673582 236680
rect 673528 236642 673580 236648
rect 673426 236558 673592 236586
rect 673414 236496 673466 236502
rect 673196 235606 673316 235634
rect 673380 236444 673414 236450
rect 673380 236438 673466 236444
rect 673380 236422 673454 236438
rect 672828 231826 672948 231854
rect 673012 231826 673132 231854
rect 672920 228585 672948 231826
rect 672906 228576 672962 228585
rect 672906 228511 672962 228520
rect 673104 228256 673132 231826
rect 672828 228228 673132 228256
rect 672828 227610 672856 228228
rect 673046 227928 673098 227934
rect 673196 227916 673224 235606
rect 673380 233322 673408 236422
rect 673564 234036 673592 236558
rect 673752 236292 673804 236298
rect 673752 236234 673804 236240
rect 673764 236178 673792 236234
rect 673748 236150 673792 236178
rect 673748 234138 673776 236150
rect 674024 234954 674052 244246
rect 674208 235657 674236 244246
rect 674194 235648 674250 235657
rect 674194 235583 674250 235592
rect 674484 234977 674512 253906
rect 674470 234968 674526 234977
rect 674024 234926 674328 234954
rect 673748 234110 673868 234138
rect 673564 234008 673776 234036
rect 673288 233294 673408 233322
rect 673288 228018 673316 233294
rect 673552 231056 673604 231062
rect 673604 231004 673684 231010
rect 673552 230998 673684 231004
rect 673564 230982 673684 230998
rect 673460 230852 673512 230858
rect 673460 230794 673512 230800
rect 673472 229809 673500 230794
rect 673656 230110 673684 230982
rect 673748 230330 673776 234008
rect 673840 233594 673868 234110
rect 673840 233566 673960 233594
rect 673932 233322 673960 233566
rect 673932 233294 673988 233322
rect 673960 233186 673988 233294
rect 673932 233158 673988 233186
rect 673932 232937 673960 233158
rect 673918 232928 673974 232937
rect 673918 232863 673974 232872
rect 673920 232076 673972 232082
rect 673920 232018 673972 232024
rect 673932 230738 673960 232018
rect 674300 231854 674328 234926
rect 674470 234903 674526 234912
rect 674426 234796 674478 234802
rect 674426 234738 674478 234744
rect 674438 234614 674466 234738
rect 673840 230710 673960 230738
rect 674208 231826 674328 231854
rect 674392 234586 674466 234614
rect 673840 230466 673868 230710
rect 674010 230616 674066 230625
rect 674010 230551 674012 230560
rect 674064 230551 674066 230560
rect 674012 230522 674064 230528
rect 673840 230450 673960 230466
rect 673840 230444 673972 230450
rect 673840 230438 673920 230444
rect 673920 230386 673972 230392
rect 673748 230314 673868 230330
rect 673748 230308 673880 230314
rect 673748 230302 673828 230308
rect 673828 230250 673880 230256
rect 674058 230240 674110 230246
rect 674208 230228 674236 231826
rect 674184 230217 674236 230228
rect 674058 230182 674110 230188
rect 674170 230208 674236 230217
rect 673644 230104 673696 230110
rect 673644 230046 673696 230052
rect 673826 230072 673882 230081
rect 673826 230007 673882 230016
rect 673458 229800 673514 229809
rect 673458 229735 673514 229744
rect 673840 229498 673868 230007
rect 673948 229968 674000 229974
rect 673946 229936 673948 229945
rect 674000 229936 674002 229945
rect 673946 229871 674002 229880
rect 674070 229786 674098 230182
rect 674226 230200 674236 230208
rect 674170 230143 674226 230152
rect 674392 230160 674420 234586
rect 674668 234433 674696 266999
rect 674838 264480 674894 264489
rect 674838 264415 674894 264424
rect 674852 263809 674880 264415
rect 676494 264072 676550 264081
rect 676494 264007 676550 264016
rect 674838 263800 674894 263809
rect 674838 263735 674894 263744
rect 676508 263673 676536 264007
rect 676494 263664 676550 263673
rect 676494 263599 676550 263608
rect 678242 263256 678298 263265
rect 678242 263191 678298 263200
rect 676218 262848 676274 262857
rect 676218 262783 676274 262792
rect 676232 260522 676260 262783
rect 675496 260494 676260 260522
rect 675298 257544 675354 257553
rect 675298 257479 675354 257488
rect 675312 256737 675340 257479
rect 675298 256728 675354 256737
rect 675298 256663 675354 256672
rect 675496 252362 675524 260494
rect 675942 258768 675998 258777
rect 675942 258703 675998 258712
rect 675956 258233 675984 258703
rect 675942 258224 675998 258233
rect 675942 258159 675998 258168
rect 675220 252334 675524 252362
rect 674930 251560 674986 251569
rect 674930 251495 674986 251504
rect 674944 251174 674972 251495
rect 674944 251146 675156 251174
rect 674930 249384 674986 249393
rect 674930 249319 674986 249328
rect 674944 245426 674972 249319
rect 675128 247058 675156 251146
rect 675220 247398 675248 252334
rect 678256 252278 678284 263191
rect 678426 261216 678482 261225
rect 678426 261151 678482 261160
rect 675852 252272 675904 252278
rect 675312 252220 675852 252226
rect 675312 252214 675904 252220
rect 678244 252272 678296 252278
rect 678244 252214 678296 252220
rect 675312 252198 675892 252214
rect 675312 250526 675340 252198
rect 678440 251598 678468 261151
rect 675852 251592 675904 251598
rect 675850 251560 675852 251569
rect 678428 251592 678480 251598
rect 675904 251560 675906 251569
rect 678428 251534 678480 251540
rect 675850 251495 675906 251504
rect 675312 250498 675418 250526
rect 675758 250336 675814 250345
rect 675758 250271 675814 250280
rect 675772 249900 675800 250271
rect 675390 249656 675446 249665
rect 675390 249591 675446 249600
rect 675404 249220 675432 249591
rect 675220 247370 675418 247398
rect 675128 247030 675340 247058
rect 675114 246936 675170 246945
rect 675114 246871 675170 246880
rect 675128 246213 675156 246871
rect 675312 246854 675340 247030
rect 675312 246826 675418 246854
rect 675128 246185 675418 246213
rect 675114 245576 675170 245585
rect 675170 245534 675418 245562
rect 675114 245511 675170 245520
rect 674944 245398 675156 245426
rect 674838 245304 674894 245313
rect 674838 245239 674894 245248
rect 674852 241890 674880 245239
rect 675128 243085 675156 245398
rect 675128 243057 675418 243085
rect 675390 242856 675446 242865
rect 675390 242791 675446 242800
rect 675404 242519 675432 242791
rect 674852 241862 675418 241890
rect 675114 241496 675170 241505
rect 675114 241431 675170 241440
rect 675128 241245 675156 241431
rect 675128 241217 675418 241245
rect 675206 240272 675262 240281
rect 675206 240207 675262 240216
rect 675220 240054 675248 240207
rect 675220 240026 675418 240054
rect 675114 238232 675170 238241
rect 675170 238190 675418 238218
rect 675114 238167 675170 238176
rect 675312 237646 675432 237674
rect 675312 237538 675340 237646
rect 675128 237510 675340 237538
rect 675404 237524 675432 237646
rect 674838 237416 674894 237425
rect 674838 237351 674894 237360
rect 674852 235249 674880 237351
rect 675128 235929 675156 237510
rect 675390 236872 675446 236881
rect 675390 236807 675446 236816
rect 675404 236368 675432 236807
rect 675114 235920 675170 235929
rect 675114 235855 675170 235864
rect 675666 235512 675722 235521
rect 675666 235447 675722 235456
rect 674838 235240 674894 235249
rect 674838 235175 674894 235184
rect 674654 234424 674710 234433
rect 674654 234359 674710 234368
rect 674886 234320 674938 234326
rect 674760 234268 674886 234274
rect 674760 234262 674938 234268
rect 675680 234274 675708 235447
rect 676034 235240 676090 235249
rect 676034 235175 676090 235184
rect 675850 234968 675906 234977
rect 675850 234903 675906 234912
rect 675864 234598 675892 234903
rect 675852 234592 675904 234598
rect 675852 234534 675904 234540
rect 675850 234424 675906 234433
rect 675850 234359 675852 234368
rect 675904 234359 675906 234368
rect 675852 234330 675904 234336
rect 674564 234252 674616 234258
rect 674564 234194 674616 234200
rect 674760 234246 674926 234262
rect 675680 234258 675892 234274
rect 675680 234252 675904 234258
rect 675680 234246 675852 234252
rect 674576 232082 674604 234194
rect 674760 233034 674788 234246
rect 675852 234194 675904 234200
rect 674978 234116 675030 234122
rect 674978 234058 675030 234064
rect 674990 234002 675018 234058
rect 674990 233974 675892 234002
rect 675096 233912 675148 233918
rect 675148 233860 675156 233900
rect 675096 233854 675156 233860
rect 675128 233492 675156 233854
rect 675864 233714 675892 233974
rect 675852 233708 675904 233714
rect 675852 233650 675904 233656
rect 675036 233464 675156 233492
rect 674748 233028 674800 233034
rect 674748 232970 674800 232976
rect 675036 232830 675064 233464
rect 676048 233442 676076 235175
rect 679624 234592 679676 234598
rect 679624 234534 679676 234540
rect 677784 233708 677836 233714
rect 677784 233650 677836 233656
rect 676036 233436 676088 233442
rect 676036 233378 676088 233384
rect 675024 232824 675076 232830
rect 675024 232766 675076 232772
rect 675484 232552 675536 232558
rect 675852 232552 675904 232558
rect 675536 232500 675852 232506
rect 675484 232494 675904 232500
rect 675496 232478 675892 232494
rect 675346 232348 675398 232354
rect 675346 232290 675398 232296
rect 675358 232082 675386 232290
rect 674564 232076 674616 232082
rect 674564 232018 674616 232024
rect 675346 232076 675398 232082
rect 675346 232018 675398 232024
rect 675178 231840 675234 231849
rect 675178 231775 675180 231784
rect 675232 231775 675234 231784
rect 675180 231746 675232 231752
rect 675070 231600 675122 231606
rect 675068 231568 675070 231577
rect 675122 231568 675124 231577
rect 675068 231503 675124 231512
rect 674956 231328 675008 231334
rect 675008 231276 675892 231282
rect 674956 231270 675892 231276
rect 674968 231266 675892 231270
rect 674968 231260 675904 231266
rect 674968 231254 675852 231260
rect 675852 231202 675904 231208
rect 677600 231260 677652 231266
rect 677600 231202 677652 231208
rect 674840 231192 674892 231198
rect 674838 231160 674840 231169
rect 674892 231160 674894 231169
rect 674838 231095 674894 231104
rect 674564 231056 674616 231062
rect 674564 230998 674616 231004
rect 674576 230738 674604 230998
rect 674732 230920 674784 230926
rect 674730 230888 674732 230897
rect 674784 230888 674786 230897
rect 674730 230823 674786 230832
rect 674838 230752 674894 230761
rect 674576 230710 674838 230738
rect 674838 230687 674894 230696
rect 675850 230752 675906 230761
rect 675850 230687 675906 230696
rect 674518 230512 674570 230518
rect 674746 230480 674802 230489
rect 674570 230460 674746 230466
rect 674518 230454 674746 230460
rect 674530 230438 674746 230454
rect 674746 230415 674802 230424
rect 674392 230132 674512 230160
rect 674070 229758 674236 229786
rect 674208 229673 674236 229758
rect 674194 229664 674250 229673
rect 674194 229599 674250 229608
rect 673828 229492 673880 229498
rect 673828 229434 673880 229440
rect 673458 229392 673514 229401
rect 673458 229327 673460 229336
rect 673512 229327 673514 229336
rect 673460 229298 673512 229304
rect 673596 229120 673652 229129
rect 673596 229055 673598 229064
rect 673650 229055 673652 229064
rect 673598 229026 673650 229032
rect 673506 228880 673558 228886
rect 673504 228848 673506 228857
rect 673558 228848 673560 228857
rect 673504 228783 673560 228792
rect 673386 228576 673442 228585
rect 673386 228511 673388 228520
rect 673440 228511 673442 228520
rect 673388 228482 673440 228488
rect 673288 227990 673684 228018
rect 673196 227888 673500 227916
rect 673046 227870 673098 227876
rect 673058 227746 673086 227870
rect 673058 227718 673224 227746
rect 672828 227582 673040 227610
rect 673012 227474 673040 227582
rect 673012 227446 673086 227474
rect 673058 227372 673086 227446
rect 673058 227344 673132 227372
rect 672736 227310 672948 227338
rect 672920 227202 672948 227310
rect 672644 227174 672856 227202
rect 672920 227174 673040 227202
rect 672604 227112 672656 227118
rect 672446 227080 672502 227089
rect 672446 227015 672502 227024
rect 672602 227080 672604 227089
rect 672656 227080 672658 227089
rect 672602 227015 672658 227024
rect 672494 226908 672546 226914
rect 672092 226868 672212 226896
rect 672184 226658 672212 226868
rect 672546 226868 672672 226896
rect 672494 226850 672546 226856
rect 672378 226808 672434 226817
rect 672378 226743 672380 226752
rect 672432 226743 672434 226752
rect 672380 226714 672432 226720
rect 672184 226630 672304 226658
rect 672034 226296 672086 226302
rect 672032 226264 672034 226273
rect 672086 226264 672088 226273
rect 672032 226199 672088 226208
rect 671908 226086 672028 226114
rect 671802 225992 671858 226001
rect 671802 225927 671858 225936
rect 671820 225752 671872 225758
rect 671818 225720 671820 225729
rect 671872 225720 671874 225729
rect 671818 225655 671874 225664
rect 671608 225576 671660 225604
rect 671608 225468 671636 225576
rect 671712 225548 671764 225554
rect 671712 225490 671764 225496
rect 671608 225440 671660 225468
rect 671448 222166 671568 222194
rect 671540 150249 671568 222166
rect 671632 215294 671660 225440
rect 671724 222194 671752 225490
rect 672000 225434 672028 226086
rect 671954 225406 672028 225434
rect 671954 225162 671982 225406
rect 671908 225134 671982 225162
rect 671724 222166 671844 222194
rect 671816 221513 671844 222166
rect 671908 221626 671936 225134
rect 672078 223000 672134 223009
rect 672078 222935 672134 222944
rect 672092 222194 672120 222935
rect 672092 222166 672212 222194
rect 671908 221598 672028 221626
rect 671802 221504 671858 221513
rect 671802 221439 671858 221448
rect 672000 220153 672028 221598
rect 671986 220144 672042 220153
rect 671986 220079 672042 220088
rect 671894 219464 671950 219473
rect 671894 219399 671950 219408
rect 671632 215266 671752 215294
rect 671724 158409 671752 215266
rect 671908 174865 671936 219399
rect 672184 214962 672212 222166
rect 672092 214934 672212 214962
rect 672092 214849 672120 214934
rect 672078 214840 672134 214849
rect 672078 214775 672134 214784
rect 672276 214554 672304 226630
rect 672644 226624 672672 226868
rect 672552 226596 672672 226624
rect 672552 225593 672580 226596
rect 672828 226545 672856 227174
rect 672814 226536 672870 226545
rect 672814 226471 672870 226480
rect 673012 226386 673040 227174
rect 672920 226358 673040 226386
rect 672538 225584 672594 225593
rect 672538 225519 672594 225528
rect 672722 224904 672778 224913
rect 672722 224839 672778 224848
rect 672538 224632 672594 224641
rect 672538 224567 672594 224576
rect 672552 214849 672580 224567
rect 672736 216345 672764 224839
rect 672722 216336 672778 216345
rect 672722 216271 672778 216280
rect 672538 214840 672594 214849
rect 672538 214775 672594 214784
rect 672276 214526 672488 214554
rect 672170 213752 672226 213761
rect 672170 213687 672226 213696
rect 672184 200841 672212 213687
rect 672460 209774 672488 214526
rect 672722 210216 672778 210225
rect 672722 210151 672778 210160
rect 672460 209746 672580 209774
rect 672170 200832 672226 200841
rect 672170 200767 672226 200776
rect 672552 198801 672580 209746
rect 672538 198792 672594 198801
rect 672538 198727 672594 198736
rect 672078 183560 672134 183569
rect 672078 183495 672134 183504
rect 671894 174856 671950 174865
rect 671894 174791 671950 174800
rect 671894 166968 671950 166977
rect 671894 166903 671950 166912
rect 671710 158400 671766 158409
rect 671710 158335 671766 158344
rect 671526 150240 671582 150249
rect 671526 150175 671582 150184
rect 670606 147656 670662 147665
rect 670606 147591 670662 147600
rect 670804 147646 671384 147674
rect 670804 145586 670832 147646
rect 670792 145580 670844 145586
rect 670792 145522 670844 145528
rect 671342 131744 671398 131753
rect 671342 131679 671398 131688
rect 670332 118516 670384 118522
rect 670332 118458 670384 118464
rect 668124 114164 668176 114170
rect 668124 114106 668176 114112
rect 669964 114164 670016 114170
rect 669964 114106 670016 114112
rect 668136 112713 668164 114106
rect 671356 113174 671384 131679
rect 671526 130928 671582 130937
rect 671526 130863 671582 130872
rect 670804 113146 671384 113174
rect 668122 112704 668178 112713
rect 668122 112639 668178 112648
rect 668582 111888 668638 111897
rect 668582 111823 668638 111832
rect 589924 111104 589976 111110
rect 589924 111046 589976 111052
rect 590106 110120 590162 110129
rect 590106 110055 590162 110064
rect 589372 109744 589424 109750
rect 589372 109686 589424 109692
rect 589462 108488 589518 108497
rect 589462 108423 589518 108432
rect 589476 107710 589504 108423
rect 589464 107704 589516 107710
rect 589464 107646 589516 107652
rect 589462 106856 589518 106865
rect 589462 106791 589518 106800
rect 589476 106350 589504 106791
rect 589464 106344 589516 106350
rect 589464 106286 589516 106292
rect 589462 105224 589518 105233
rect 589462 105159 589518 105168
rect 589476 104922 589504 105159
rect 589464 104916 589516 104922
rect 589464 104858 589516 104864
rect 589554 103592 589610 103601
rect 589554 103527 589610 103536
rect 589568 100774 589596 103527
rect 589922 101960 589978 101969
rect 589922 101895 589978 101904
rect 589556 100768 589608 100774
rect 589556 100710 589608 100716
rect 588544 91792 588596 91798
rect 588544 91734 588596 91740
rect 589936 79490 589964 101895
rect 590120 100026 590148 110055
rect 666650 109372 666706 109381
rect 666650 109307 666706 109316
rect 666664 103514 666692 109307
rect 668400 106208 668452 106214
rect 668122 106176 668178 106185
rect 668122 106111 668178 106120
rect 668398 106176 668400 106185
rect 668452 106176 668454 106185
rect 668398 106111 668454 106120
rect 666572 103486 666692 103514
rect 624792 100156 624844 100162
rect 624792 100098 624844 100104
rect 590108 100020 590160 100026
rect 590108 99962 590160 99968
rect 595272 100014 595608 100042
rect 596344 100014 596496 100042
rect 595272 99142 595300 100014
rect 595260 99136 595312 99142
rect 595260 99078 595312 99084
rect 595272 93854 595300 99078
rect 596180 96960 596232 96966
rect 596180 96902 596232 96908
rect 595272 93826 595484 93854
rect 595456 80714 595484 93826
rect 595444 80708 595496 80714
rect 595444 80650 595496 80656
rect 589924 79484 589976 79490
rect 589924 79426 589976 79432
rect 589922 77344 589978 77353
rect 589922 77279 589978 77288
rect 588544 75948 588596 75954
rect 588544 75890 588596 75896
rect 587164 73160 587216 73166
rect 587164 73102 587216 73108
rect 585784 71256 585836 71262
rect 585784 71198 585836 71204
rect 585784 68332 585836 68338
rect 585784 68274 585836 68280
rect 584404 54936 584456 54942
rect 584404 54878 584456 54884
rect 585796 54777 585824 68274
rect 588556 56574 588584 75890
rect 588544 56568 588596 56574
rect 588544 56510 588596 56516
rect 589936 54806 589964 77279
rect 596192 56030 596220 96902
rect 596468 56166 596496 100014
rect 596744 100014 597080 100042
rect 597664 100014 597816 100042
rect 597940 100014 598552 100042
rect 598952 100014 599288 100042
rect 599504 100014 600024 100042
rect 600332 100014 600760 100042
rect 600884 100014 601496 100042
rect 601896 100014 602232 100042
rect 602356 100014 602968 100042
rect 603092 100014 603704 100042
rect 596744 96966 596772 100014
rect 596732 96960 596784 96966
rect 596732 96902 596784 96908
rect 596456 56160 596508 56166
rect 596456 56102 596508 56108
rect 596180 56024 596232 56030
rect 596180 55966 596232 55972
rect 589924 54800 589976 54806
rect 585782 54768 585838 54777
rect 589924 54742 589976 54748
rect 585782 54703 585838 54712
rect 597664 54670 597692 100014
rect 597652 54664 597704 54670
rect 597652 54606 597704 54612
rect 597940 54534 597968 100014
rect 598952 79354 598980 100014
rect 599504 84194 599532 100014
rect 600332 89010 600360 100014
rect 600320 89004 600372 89010
rect 600320 88946 600372 88952
rect 600884 84194 600912 100014
rect 601896 95946 601924 100014
rect 601884 95940 601936 95946
rect 601884 95882 601936 95888
rect 602356 84194 602384 100014
rect 599136 84166 599532 84194
rect 600516 84166 600912 84194
rect 601896 84166 602384 84194
rect 598940 79348 598992 79354
rect 598940 79290 598992 79296
rect 599136 55894 599164 84166
rect 600516 58682 600544 84166
rect 601896 68338 601924 84166
rect 601884 68332 601936 68338
rect 601884 68274 601936 68280
rect 600504 58676 600556 58682
rect 600504 58618 600556 58624
rect 603092 57254 603120 100014
rect 604426 99770 604454 100028
rect 605176 100014 605512 100042
rect 605912 100014 606248 100042
rect 606648 100014 607168 100042
rect 607384 100014 607720 100042
rect 608120 100014 608548 100042
rect 608856 100014 609192 100042
rect 609592 100014 609928 100042
rect 610328 100014 610664 100042
rect 611064 100014 611308 100042
rect 611800 100014 612136 100042
rect 612536 100014 612688 100042
rect 613272 100014 613608 100042
rect 604426 99742 604500 99770
rect 603080 57248 603132 57254
rect 603080 57190 603132 57196
rect 599124 55888 599176 55894
rect 599124 55830 599176 55836
rect 597928 54528 597980 54534
rect 604472 54505 604500 99742
rect 605484 97986 605512 100014
rect 605472 97980 605524 97986
rect 605472 97922 605524 97928
rect 606220 96762 606248 100014
rect 606484 97980 606536 97986
rect 606484 97922 606536 97928
rect 606208 96756 606260 96762
rect 606208 96698 606260 96704
rect 606496 76566 606524 97922
rect 607140 92614 607168 100014
rect 607692 95946 607720 100014
rect 607680 95940 607732 95946
rect 607680 95882 607732 95888
rect 607128 92608 607180 92614
rect 607128 92550 607180 92556
rect 608520 84182 608548 100014
rect 609164 94518 609192 100014
rect 609152 94512 609204 94518
rect 609152 94454 609204 94460
rect 609900 85542 609928 100014
rect 610636 96082 610664 100014
rect 610624 96076 610676 96082
rect 610624 96018 610676 96024
rect 611280 93158 611308 100014
rect 612108 96898 612136 100014
rect 612660 97102 612688 100014
rect 613580 97442 613608 100014
rect 613994 99770 614022 100028
rect 614744 100014 615172 100042
rect 615480 100014 615816 100042
rect 616216 100014 616644 100042
rect 616952 100014 617288 100042
rect 617688 100014 618024 100042
rect 618424 100014 618760 100042
rect 619160 100014 619588 100042
rect 619896 100014 620232 100042
rect 620632 100014 620968 100042
rect 621368 100014 621704 100042
rect 622104 100014 622348 100042
rect 622840 100014 623176 100042
rect 623576 100014 623728 100042
rect 624312 100014 624648 100042
rect 614856 99952 614908 99958
rect 614856 99894 614908 99900
rect 613994 99742 614068 99770
rect 613568 97436 613620 97442
rect 613568 97378 613620 97384
rect 612648 97096 612700 97102
rect 612648 97038 612700 97044
rect 612096 96892 612148 96898
rect 612096 96834 612148 96840
rect 612648 96892 612700 96898
rect 612648 96834 612700 96840
rect 612004 96756 612056 96762
rect 612004 96698 612056 96704
rect 611268 93152 611320 93158
rect 611268 93094 611320 93100
rect 610072 92608 610124 92614
rect 610072 92550 610124 92556
rect 610084 88330 610112 92550
rect 610072 88324 610124 88330
rect 610072 88266 610124 88272
rect 609888 85536 609940 85542
rect 609888 85478 609940 85484
rect 608508 84176 608560 84182
rect 608508 84118 608560 84124
rect 606484 76560 606536 76566
rect 606484 76502 606536 76508
rect 612016 75342 612044 96698
rect 612660 75478 612688 96834
rect 613382 95840 613438 95849
rect 613382 95775 613438 95784
rect 612648 75472 612700 75478
rect 612648 75414 612700 75420
rect 612004 75336 612056 75342
rect 612004 75278 612056 75284
rect 613396 62082 613424 95775
rect 614040 80850 614068 99742
rect 614028 80844 614080 80850
rect 614028 80786 614080 80792
rect 614868 64870 614896 99894
rect 615144 93854 615172 100014
rect 615788 96966 615816 100014
rect 615776 96960 615828 96966
rect 615776 96902 615828 96908
rect 615144 93826 615448 93854
rect 615420 79354 615448 93826
rect 616616 91798 616644 100014
rect 616788 96960 616840 96966
rect 616788 96902 616840 96908
rect 616604 91792 616656 91798
rect 616604 91734 616656 91740
rect 615408 79348 615460 79354
rect 615408 79290 615460 79296
rect 616800 76702 616828 96902
rect 617260 96898 617288 100014
rect 617248 96892 617300 96898
rect 617248 96834 617300 96840
rect 617996 92478 618024 100014
rect 618732 97986 618760 100014
rect 618720 97980 618772 97986
rect 618720 97922 618772 97928
rect 618904 97436 618956 97442
rect 618904 97378 618956 97384
rect 618168 96892 618220 96898
rect 618168 96834 618220 96840
rect 617984 92472 618036 92478
rect 617984 92414 618036 92420
rect 618180 91050 618208 96834
rect 618168 91044 618220 91050
rect 618168 90986 618220 90992
rect 618916 80986 618944 97378
rect 619560 93838 619588 100014
rect 620204 97442 620232 100014
rect 620192 97436 620244 97442
rect 620192 97378 620244 97384
rect 620940 95198 620968 100014
rect 621676 97714 621704 100014
rect 622320 99346 622348 100014
rect 622308 99340 622360 99346
rect 622308 99282 622360 99288
rect 621664 97708 621716 97714
rect 621664 97650 621716 97656
rect 623148 97306 623176 100014
rect 623700 99210 623728 100014
rect 623688 99204 623740 99210
rect 623688 99146 623740 99152
rect 623136 97300 623188 97306
rect 623136 97242 623188 97248
rect 621664 97096 621716 97102
rect 621664 97038 621716 97044
rect 620928 95192 620980 95198
rect 620928 95134 620980 95140
rect 620284 94512 620336 94518
rect 620284 94454 620336 94460
rect 619548 93832 619600 93838
rect 619548 93774 619600 93780
rect 619548 93152 619600 93158
rect 619548 93094 619600 93100
rect 619560 88194 619588 93094
rect 619548 88188 619600 88194
rect 619548 88130 619600 88136
rect 620296 85406 620324 94454
rect 620284 85400 620336 85406
rect 620284 85342 620336 85348
rect 618904 80980 618956 80986
rect 618904 80922 618956 80928
rect 621676 77994 621704 97038
rect 624620 97034 624648 100014
rect 624608 97028 624660 97034
rect 624608 96970 624660 96976
rect 623044 96076 623096 96082
rect 623044 96018 623096 96024
rect 622308 95940 622360 95946
rect 622308 95882 622360 95888
rect 622320 89690 622348 95882
rect 622308 89684 622360 89690
rect 622308 89626 622360 89632
rect 623056 86358 623084 96018
rect 623044 86352 623096 86358
rect 623044 86294 623096 86300
rect 624804 84194 624832 100098
rect 625034 99770 625062 100028
rect 625784 100014 626120 100042
rect 626520 100014 626856 100042
rect 627256 100014 627592 100042
rect 627992 100014 628328 100042
rect 628728 100014 629064 100042
rect 629464 100014 629800 100042
rect 630200 100014 630536 100042
rect 630936 100014 631272 100042
rect 631672 100014 632008 100042
rect 632408 100014 632744 100042
rect 633144 100014 633296 100042
rect 633880 100014 634216 100042
rect 634616 100014 634768 100042
rect 635352 100014 635596 100042
rect 625034 99742 625108 99770
rect 625080 99074 625108 99742
rect 625068 99068 625120 99074
rect 625068 99010 625120 99016
rect 625804 97980 625856 97986
rect 625804 97922 625856 97928
rect 625816 92041 625844 97922
rect 626092 97578 626120 100014
rect 626080 97572 626132 97578
rect 626080 97514 626132 97520
rect 625988 97436 626040 97442
rect 625988 97378 626040 97384
rect 626000 93673 626028 97378
rect 626828 97170 626856 100014
rect 627564 97850 627592 100014
rect 628300 97986 628328 100014
rect 629036 98938 629064 100014
rect 629024 98932 629076 98938
rect 629024 98874 629076 98880
rect 629772 98802 629800 100014
rect 629760 98796 629812 98802
rect 629760 98738 629812 98744
rect 630508 98666 630536 100014
rect 630772 99340 630824 99346
rect 630772 99282 630824 99288
rect 630496 98660 630548 98666
rect 630496 98602 630548 98608
rect 628288 97980 628340 97986
rect 628288 97922 628340 97928
rect 627552 97844 627604 97850
rect 627552 97786 627604 97792
rect 629300 97708 629352 97714
rect 629300 97650 629352 97656
rect 626816 97164 626868 97170
rect 626816 97106 626868 97112
rect 629312 95826 629340 97650
rect 630784 95826 630812 99282
rect 631244 97442 631272 100014
rect 631980 97714 632008 100014
rect 631968 97708 632020 97714
rect 631968 97650 632020 97656
rect 631232 97436 631284 97442
rect 631232 97378 631284 97384
rect 632716 97306 632744 100014
rect 632060 97300 632112 97306
rect 632060 97242 632112 97248
rect 632704 97300 632756 97306
rect 632704 97242 632756 97248
rect 629280 95798 629340 95826
rect 630752 95798 630812 95826
rect 632072 95826 632100 97242
rect 633268 96898 633296 100014
rect 633440 99204 633492 99210
rect 633440 99146 633492 99152
rect 633256 96892 633308 96898
rect 633256 96834 633308 96840
rect 633452 95826 633480 99146
rect 634188 97850 634216 100014
rect 634176 97844 634228 97850
rect 634176 97786 634228 97792
rect 634740 96762 634768 100014
rect 635568 97034 635596 100014
rect 635752 100014 636088 100042
rect 636824 100014 637068 100042
rect 635004 97028 635056 97034
rect 635004 96970 635056 96976
rect 635556 97028 635608 97034
rect 635556 96970 635608 96976
rect 634728 96756 634780 96762
rect 634728 96698 634780 96704
rect 635016 95826 635044 96970
rect 635752 96121 635780 100014
rect 636292 99068 636344 99074
rect 636292 99010 636344 99016
rect 635738 96112 635794 96121
rect 635738 96047 635794 96056
rect 636304 95826 636332 99010
rect 637040 96937 637068 100014
rect 637546 99770 637574 100028
rect 638296 100014 638632 100042
rect 639032 100014 639644 100042
rect 639768 100014 640104 100042
rect 637546 99742 637620 99770
rect 637026 96928 637082 96937
rect 637026 96863 637082 96872
rect 637592 96218 637620 99742
rect 637764 97572 637816 97578
rect 637764 97514 637816 97520
rect 637580 96212 637632 96218
rect 637580 96154 637632 96160
rect 637776 95826 637804 97514
rect 638604 96626 638632 100014
rect 639052 97572 639104 97578
rect 639052 97514 639104 97520
rect 639064 97034 639092 97514
rect 639236 97164 639288 97170
rect 639236 97106 639288 97112
rect 639052 97028 639104 97034
rect 639052 96970 639104 96976
rect 638592 96620 638644 96626
rect 638592 96562 638644 96568
rect 639248 95826 639276 97106
rect 639420 97028 639472 97034
rect 639420 96970 639472 96976
rect 639432 96762 639460 96970
rect 639420 96756 639472 96762
rect 639420 96698 639472 96704
rect 639616 96490 639644 100014
rect 639788 97436 639840 97442
rect 639788 97378 639840 97384
rect 639800 96898 639828 97378
rect 639788 96892 639840 96898
rect 639788 96834 639840 96840
rect 639604 96484 639656 96490
rect 639604 96426 639656 96432
rect 640076 96354 640104 100014
rect 640490 99770 640518 100028
rect 641240 100014 641576 100042
rect 640490 99742 640564 99770
rect 640064 96348 640116 96354
rect 640064 96290 640116 96296
rect 632072 95798 632224 95826
rect 633452 95798 633696 95826
rect 635016 95798 635168 95826
rect 636304 95798 636640 95826
rect 637776 95798 638112 95826
rect 639248 95798 639584 95826
rect 640536 95470 640564 99742
rect 640708 98048 640760 98054
rect 640708 97990 640760 97996
rect 640720 95826 640748 97990
rect 641548 96082 641576 100014
rect 641962 99770 641990 100028
rect 642712 100014 643048 100042
rect 641962 99742 642036 99770
rect 641536 96076 641588 96082
rect 641536 96018 641588 96024
rect 640720 95798 641056 95826
rect 642008 95606 642036 99742
rect 642180 98184 642232 98190
rect 642180 98126 642232 98132
rect 642192 95826 642220 98126
rect 643020 97578 643048 100014
rect 643434 99770 643462 100028
rect 644184 100014 644336 100042
rect 644920 100014 645348 100042
rect 645656 100014 645808 100042
rect 643434 99742 643508 99770
rect 643008 97572 643060 97578
rect 643008 97514 643060 97520
rect 642640 96484 642692 96490
rect 642640 96426 642692 96432
rect 642192 95798 642528 95826
rect 642652 95742 642680 96426
rect 642640 95736 642692 95742
rect 642640 95678 642692 95684
rect 641996 95600 642048 95606
rect 641996 95542 642048 95548
rect 643480 95470 643508 99742
rect 643652 98932 643704 98938
rect 643652 98874 643704 98880
rect 643664 95826 643692 98874
rect 644308 97170 644336 100014
rect 645124 98796 645176 98802
rect 645124 98738 645176 98744
rect 644296 97164 644348 97170
rect 644296 97106 644348 97112
rect 645136 95826 645164 98738
rect 645320 95946 645348 100014
rect 645780 96626 645808 100014
rect 646378 99770 646406 100028
rect 647114 99770 647142 100028
rect 647864 100014 648200 100042
rect 648600 100014 648936 100042
rect 649336 100014 649764 100042
rect 650072 100014 650408 100042
rect 650808 100014 651144 100042
rect 651544 100014 651880 100042
rect 652280 100014 652616 100042
rect 653016 100014 653352 100042
rect 653752 100014 653996 100042
rect 654488 100014 654824 100042
rect 655224 100014 655468 100042
rect 646378 99742 646452 99770
rect 647114 99742 647188 99770
rect 645768 96620 645820 96626
rect 645768 96562 645820 96568
rect 645308 95940 645360 95946
rect 645308 95882 645360 95888
rect 643664 95798 644000 95826
rect 645136 95798 645472 95826
rect 646424 95606 646452 99742
rect 646596 98660 646648 98666
rect 646596 98602 646648 98608
rect 646608 95826 646636 98602
rect 647160 97850 647188 99742
rect 647148 97844 647200 97850
rect 647148 97786 647200 97792
rect 647056 97436 647108 97442
rect 647056 97378 647108 97384
rect 646608 95798 646944 95826
rect 646228 95600 646280 95606
rect 646226 95568 646228 95577
rect 646412 95600 646464 95606
rect 646280 95568 646282 95577
rect 646412 95542 646464 95548
rect 646226 95503 646282 95512
rect 640524 95464 640576 95470
rect 640524 95406 640576 95412
rect 643468 95464 643520 95470
rect 643468 95406 643520 95412
rect 647068 95198 647096 97378
rect 647516 97028 647568 97034
rect 647516 96970 647568 96976
rect 647332 96892 647384 96898
rect 647332 96834 647384 96840
rect 626448 95192 626500 95198
rect 626448 95134 626500 95140
rect 647056 95192 647108 95198
rect 647056 95134 647108 95140
rect 626460 94489 626488 95134
rect 647344 95033 647372 96834
rect 647330 95024 647386 95033
rect 647330 94959 647386 94968
rect 626446 94480 626502 94489
rect 626446 94415 626502 94424
rect 626448 93832 626500 93838
rect 626448 93774 626500 93780
rect 625986 93664 626042 93673
rect 625986 93599 626042 93608
rect 626460 92857 626488 93774
rect 626446 92848 626502 92857
rect 626446 92783 626502 92792
rect 626448 92472 626500 92478
rect 626448 92414 626500 92420
rect 625802 92032 625858 92041
rect 625802 91967 625858 91976
rect 626264 91792 626316 91798
rect 626264 91734 626316 91740
rect 626276 89593 626304 91734
rect 626460 91225 626488 92414
rect 626446 91216 626502 91225
rect 626446 91151 626502 91160
rect 626448 91044 626500 91050
rect 626448 90986 626500 90992
rect 626460 90409 626488 90986
rect 626446 90400 626502 90409
rect 626446 90335 626502 90344
rect 626448 89684 626500 89690
rect 626448 89626 626500 89632
rect 626262 89584 626318 89593
rect 626262 89519 626318 89528
rect 626460 88777 626488 89626
rect 626446 88768 626502 88777
rect 626446 88703 626502 88712
rect 626448 88324 626500 88330
rect 626448 88266 626500 88272
rect 626264 88188 626316 88194
rect 626264 88130 626316 88136
rect 626276 87145 626304 88130
rect 626460 87961 626488 88266
rect 626446 87952 626502 87961
rect 626446 87887 626502 87896
rect 626262 87136 626318 87145
rect 626262 87071 626318 87080
rect 626448 86352 626500 86358
rect 626446 86320 626448 86329
rect 626500 86320 626502 86329
rect 626446 86255 626502 86264
rect 626448 85536 626500 85542
rect 626446 85504 626448 85513
rect 626500 85504 626502 85513
rect 626446 85439 626502 85448
rect 625252 85400 625304 85406
rect 625252 85342 625304 85348
rect 625264 84697 625292 85342
rect 625250 84688 625306 84697
rect 625250 84623 625306 84632
rect 624436 84166 624832 84194
rect 625804 84176 625856 84182
rect 621664 77988 621716 77994
rect 621664 77930 621716 77936
rect 616788 76696 616840 76702
rect 616788 76638 616840 76644
rect 623044 66292 623096 66298
rect 623044 66234 623096 66240
rect 614856 64864 614908 64870
rect 614856 64806 614908 64812
rect 613384 62076 613436 62082
rect 613384 62018 613436 62024
rect 597928 54470 597980 54476
rect 604458 54496 604514 54505
rect 604458 54431 604514 54440
rect 583024 54392 583076 54398
rect 583024 54334 583076 54340
rect 580264 54256 580316 54262
rect 576858 54224 576914 54233
rect 580264 54198 580316 54204
rect 576858 54159 576914 54168
rect 574928 53848 574980 53854
rect 574928 53790 574980 53796
rect 459834 53680 459890 53689
rect 459834 53615 459890 53624
rect 460754 53680 460810 53689
rect 460754 53615 460810 53624
rect 461674 53680 461730 53689
rect 462594 53680 462650 53689
rect 461674 53615 461730 53624
rect 462228 53644 462280 53650
rect 459468 53508 459520 53514
rect 459468 53450 459520 53456
rect 130384 53372 130436 53378
rect 130384 53314 130436 53320
rect 129004 53100 129056 53106
rect 129004 53042 129056 53048
rect 126428 52012 126480 52018
rect 126428 51954 126480 51960
rect 126440 50794 126468 51954
rect 126428 50788 126480 50794
rect 126428 50730 126480 50736
rect 129016 50674 129044 53042
rect 129464 51876 129516 51882
rect 129464 51818 129516 51824
rect 129280 50788 129332 50794
rect 129280 50730 129332 50736
rect 129016 50646 129228 50674
rect 128636 50516 128688 50522
rect 128636 50458 128688 50464
rect 51724 49156 51776 49162
rect 51724 49098 51776 49104
rect 128452 49156 128504 49162
rect 128452 49098 128504 49104
rect 47584 49020 47636 49026
rect 47584 48962 47636 48968
rect 128464 44674 128492 49098
rect 128648 48142 128676 50458
rect 129004 50380 129056 50386
rect 129004 50322 129056 50328
rect 128636 48136 128688 48142
rect 128636 48078 128688 48084
rect 128452 44668 128504 44674
rect 128452 44610 128504 44616
rect 129016 44198 129044 50322
rect 129200 47734 129228 50646
rect 129292 48314 129320 50730
rect 129292 48286 129412 48314
rect 129188 47728 129240 47734
rect 129188 47670 129240 47676
rect 129384 44538 129412 48286
rect 129476 47682 129504 51818
rect 129648 49020 129700 49026
rect 129648 48962 129700 48968
rect 129660 48314 129688 48962
rect 129660 48286 129780 48314
rect 129476 47654 129596 47682
rect 129568 45082 129596 47654
rect 129556 45076 129608 45082
rect 129556 45018 129608 45024
rect 129752 44946 129780 48286
rect 129740 44940 129792 44946
rect 129740 44882 129792 44888
rect 129372 44532 129424 44538
rect 129372 44474 129424 44480
rect 129004 44192 129056 44198
rect 129004 44134 129056 44140
rect 130396 44062 130424 53314
rect 130568 53236 130620 53242
rect 130568 53178 130620 53184
rect 130384 44056 130436 44062
rect 130384 43998 130436 44004
rect 130580 43926 130608 53178
rect 312360 53168 312412 53174
rect 312018 53116 312360 53122
rect 312018 53110 312412 53116
rect 313740 53168 313792 53174
rect 316316 53168 316368 53174
rect 313792 53116 314042 53122
rect 313740 53110 314042 53116
rect 306024 52494 306052 53108
rect 145380 52488 145432 52494
rect 145380 52430 145432 52436
rect 306012 52488 306064 52494
rect 306012 52430 306064 52436
rect 130752 51740 130804 51746
rect 130752 51682 130804 51688
rect 130764 44334 130792 51682
rect 145392 50810 145420 52430
rect 145084 50782 145420 50810
rect 308048 50289 308076 53108
rect 312018 53094 312400 53110
rect 313752 53108 314042 53110
rect 316020 53116 316316 53122
rect 316020 53110 316368 53116
rect 317696 53168 317748 53174
rect 317748 53116 318380 53122
rect 317696 53110 318380 53116
rect 313752 53094 314056 53108
rect 316020 53094 316356 53110
rect 317708 53094 318380 53110
rect 314028 50386 314056 53094
rect 318352 50522 318380 53094
rect 459480 52578 459508 53450
rect 459848 52578 459876 53615
rect 460388 53372 460440 53378
rect 460388 53314 460440 53320
rect 460400 52578 460428 53314
rect 460768 52578 460796 53615
rect 460986 52760 461038 52766
rect 460986 52702 461038 52708
rect 459172 52550 459508 52578
rect 459632 52550 459876 52578
rect 460092 52550 460428 52578
rect 460552 52550 460796 52578
rect 460998 52564 461026 52702
rect 461688 52578 461716 53615
rect 464342 53680 464398 53689
rect 462594 53615 462650 53624
rect 462780 53644 462832 53650
rect 462228 53586 462280 53592
rect 462240 52578 462268 53586
rect 462608 52578 462636 53615
rect 462780 53586 462832 53592
rect 463608 53644 463660 53650
rect 482282 53680 482338 53689
rect 464342 53615 464344 53624
rect 463608 53586 463660 53592
rect 464396 53615 464398 53624
rect 472716 53644 472768 53650
rect 464344 53586 464396 53592
rect 472716 53586 472768 53592
rect 473176 53644 473228 53650
rect 473176 53586 473228 53592
rect 476764 53644 476816 53650
rect 476764 53586 476816 53592
rect 477868 53644 477920 53650
rect 477868 53586 477920 53592
rect 481732 53644 481784 53650
rect 482282 53615 482284 53624
rect 481732 53586 481784 53592
rect 482336 53615 482338 53624
rect 485228 53644 485280 53650
rect 482284 53586 482336 53592
rect 485228 53586 485280 53592
rect 462792 53378 462820 53586
rect 463148 53508 463200 53514
rect 463148 53450 463200 53456
rect 462780 53372 462832 53378
rect 462780 53314 462832 53320
rect 463160 52578 463188 53450
rect 463424 53236 463476 53242
rect 463424 53178 463476 53184
rect 463436 52578 463464 53178
rect 463620 52766 463648 53586
rect 472532 53576 472584 53582
rect 472532 53518 472584 53524
rect 472544 53417 472572 53518
rect 472530 53408 472586 53417
rect 465448 53372 465500 53378
rect 472530 53343 472586 53352
rect 465448 53314 465500 53320
rect 464528 53100 464580 53106
rect 464528 53042 464580 53048
rect 464068 52964 464120 52970
rect 464068 52906 464120 52912
rect 463608 52760 463660 52766
rect 463608 52702 463660 52708
rect 464080 52578 464108 52906
rect 464540 52578 464568 53042
rect 464666 52828 464718 52834
rect 464666 52770 464718 52776
rect 461472 52550 461716 52578
rect 461932 52550 462268 52578
rect 462392 52550 462636 52578
rect 462852 52550 463188 52578
rect 463312 52550 463464 52578
rect 463772 52550 464108 52578
rect 464232 52550 464568 52578
rect 464678 52564 464706 52770
rect 465460 52578 465488 53314
rect 472728 52698 472756 53586
rect 473188 53106 473216 53586
rect 476776 53242 476804 53586
rect 477132 53508 477184 53514
rect 477132 53450 477184 53456
rect 476764 53236 476816 53242
rect 476764 53178 476816 53184
rect 473176 53100 473228 53106
rect 473176 53042 473228 53048
rect 477144 52970 477172 53450
rect 477880 53378 477908 53586
rect 481744 53417 481772 53586
rect 482112 53514 482508 53530
rect 482100 53508 482520 53514
rect 482152 53502 482468 53508
rect 482100 53450 482152 53456
rect 482468 53450 482520 53456
rect 481730 53408 481786 53417
rect 477868 53372 477920 53378
rect 481730 53343 481786 53352
rect 477868 53314 477920 53320
rect 477132 52964 477184 52970
rect 477132 52906 477184 52912
rect 485240 52834 485268 53586
rect 485228 52828 485280 52834
rect 485228 52770 485280 52776
rect 465908 52692 465960 52698
rect 465908 52634 465960 52640
rect 472716 52692 472768 52698
rect 472716 52634 472768 52640
rect 465920 52578 465948 52634
rect 465152 52550 465488 52578
rect 465612 52550 465948 52578
rect 318340 50516 318392 50522
rect 318340 50458 318392 50464
rect 458364 50516 458416 50522
rect 458364 50458 458416 50464
rect 314016 50380 314068 50386
rect 314016 50322 314068 50328
rect 458180 50380 458232 50386
rect 458180 50322 458232 50328
rect 308034 50280 308090 50289
rect 308034 50215 308090 50224
rect 132132 48136 132184 48142
rect 132132 48078 132184 48084
rect 131856 47728 131908 47734
rect 131856 47670 131908 47676
rect 131868 44606 131896 47670
rect 131856 44600 131908 44606
rect 131856 44542 131908 44548
rect 132144 44506 132172 48078
rect 458192 47025 458220 50322
rect 458178 47016 458234 47025
rect 458178 46951 458234 46960
rect 458376 46753 458404 50458
rect 459172 47654 459232 47682
rect 459632 47654 459968 47682
rect 460092 47654 460152 47682
rect 460552 47654 460888 47682
rect 461012 47654 461164 47682
rect 461472 47654 461808 47682
rect 461932 47654 461992 47682
rect 458362 46744 458418 46753
rect 142370 46702 142660 46730
rect 132132 44500 132184 44506
rect 132132 44442 132184 44448
rect 132408 44464 132460 44470
rect 132236 44412 132408 44418
rect 132236 44406 132460 44412
rect 132236 44390 132448 44406
rect 130752 44328 130804 44334
rect 130752 44270 130804 44276
rect 132236 44198 132264 44390
rect 142632 44305 142660 46702
rect 458362 46679 458418 46688
rect 431222 44840 431278 44849
rect 431222 44775 431278 44784
rect 142618 44296 142674 44305
rect 142618 44231 142674 44240
rect 132224 44192 132276 44198
rect 132224 44134 132276 44140
rect 307298 44160 307354 44169
rect 307298 44095 307354 44104
rect 130568 43920 130620 43926
rect 130568 43862 130620 43868
rect 187332 43580 187384 43586
rect 187332 43522 187384 43528
rect 43444 42832 43496 42838
rect 43444 42774 43496 42780
rect 187344 42092 187372 43522
rect 194322 42120 194378 42129
rect 194074 42078 194322 42106
rect 307312 42106 307340 44095
rect 431236 43654 431264 44775
rect 431224 43648 431276 43654
rect 361762 43616 361818 43625
rect 431224 43590 431276 43596
rect 361762 43551 361818 43560
rect 310428 42764 310480 42770
rect 310428 42706 310480 42712
rect 310440 42106 310468 42706
rect 307004 42078 307340 42106
rect 310132 42078 310468 42106
rect 361776 42092 361804 43551
rect 364892 42764 364944 42770
rect 364892 42706 364944 42712
rect 431224 42764 431276 42770
rect 431224 42706 431276 42712
rect 456064 42764 456116 42770
rect 456064 42706 456116 42712
rect 364904 42092 364932 42706
rect 427084 42628 427136 42634
rect 427084 42570 427136 42576
rect 416594 42392 416650 42401
rect 404452 42356 404504 42362
rect 404452 42298 404504 42304
rect 405188 42356 405240 42362
rect 416594 42327 416650 42336
rect 420736 42356 420788 42362
rect 405188 42298 405240 42304
rect 194322 42055 194378 42064
rect 404464 41478 404492 42298
rect 405200 42106 405228 42298
rect 415766 42120 415822 42129
rect 405200 42078 405582 42106
rect 415426 42078 415766 42106
rect 416608 42092 416636 42327
rect 420736 42298 420788 42304
rect 426900 42356 426952 42362
rect 426900 42298 426952 42304
rect 415766 42055 415822 42064
rect 419906 41848 419962 41857
rect 419750 41806 419906 41834
rect 419906 41783 419962 41792
rect 420748 41478 420776 42298
rect 426912 41478 426940 42298
rect 427096 42090 427124 42570
rect 431236 42090 431264 42706
rect 455420 42492 455472 42498
rect 455420 42434 455472 42440
rect 446402 42256 446458 42265
rect 446402 42191 446458 42200
rect 427084 42084 427136 42090
rect 427084 42026 427136 42032
rect 431224 42084 431276 42090
rect 431224 42026 431276 42032
rect 446416 41585 446444 42191
rect 455432 41954 455460 42434
rect 456076 42090 456104 42706
rect 456064 42084 456116 42090
rect 456064 42026 456116 42032
rect 455420 41948 455472 41954
rect 455420 41890 455472 41896
rect 446402 41576 446458 41585
rect 446402 41511 446458 41520
rect 459204 41478 459232 47654
rect 459940 42106 459968 47654
rect 460124 44849 460152 47654
rect 460110 44840 460166 44849
rect 460110 44775 460166 44784
rect 460860 43897 460888 47654
rect 460846 43888 460902 43897
rect 460846 43823 460902 43832
rect 461136 42265 461164 47654
rect 461780 42945 461808 47654
rect 461964 44441 461992 47654
rect 462378 47410 462406 47668
rect 462332 47382 462406 47410
rect 462516 47654 462852 47682
rect 462976 47654 463312 47682
rect 461950 44432 462006 44441
rect 461950 44367 462006 44376
rect 462332 43217 462360 47382
rect 462516 44441 462544 47654
rect 462502 44432 462558 44441
rect 462502 44367 462558 44376
rect 462318 43208 462374 43217
rect 462318 43143 462374 43152
rect 461766 42936 461822 42945
rect 461766 42871 461822 42880
rect 462976 42498 463004 47654
rect 463758 47410 463786 47668
rect 463712 47382 463786 47410
rect 463896 47654 464232 47682
rect 464356 47654 464692 47682
rect 463712 43058 463740 47382
rect 463896 44169 463924 47654
rect 463882 44160 463938 44169
rect 463882 44095 463938 44104
rect 464356 43625 464384 47654
rect 465138 47410 465166 47668
rect 465092 47382 465166 47410
rect 465276 47654 465612 47682
rect 465092 46753 465120 47382
rect 465276 47025 465304 47654
rect 544028 47569 544056 53108
rect 545684 53094 546020 53122
rect 547892 53094 548044 53122
rect 544014 47560 544070 47569
rect 544014 47495 544070 47504
rect 545684 47297 545712 53094
rect 547892 47841 547920 53094
rect 550008 48929 550036 53108
rect 549994 48920 550050 48929
rect 549994 48855 550050 48864
rect 552032 48113 552060 53108
rect 553688 53094 554024 53122
rect 553688 50289 553716 53094
rect 553674 50280 553730 50289
rect 553674 50215 553730 50224
rect 552018 48104 552074 48113
rect 552018 48039 552074 48048
rect 547878 47832 547934 47841
rect 547878 47767 547934 47776
rect 545670 47288 545726 47297
rect 545670 47223 545726 47232
rect 465262 47016 465318 47025
rect 465262 46951 465318 46960
rect 465078 46744 465134 46753
rect 465078 46679 465134 46688
rect 623056 46510 623084 66234
rect 624436 57934 624464 84166
rect 625804 84118 625856 84124
rect 625816 83881 625844 84118
rect 625802 83872 625858 83881
rect 625802 83807 625858 83816
rect 628746 83328 628802 83337
rect 628746 83263 628802 83272
rect 628760 81122 628788 83263
rect 647528 82793 647556 96970
rect 647884 96348 647936 96354
rect 647884 96290 647936 96296
rect 647698 95568 647754 95577
rect 647698 95503 647754 95512
rect 647712 92818 647740 95503
rect 647700 92812 647752 92818
rect 647700 92754 647752 92760
rect 647896 86630 647924 96290
rect 648172 93906 648200 100014
rect 648620 97708 648672 97714
rect 648620 97650 648672 97656
rect 648160 93900 648212 93906
rect 648160 93842 648212 93848
rect 648632 92041 648660 97650
rect 648908 96354 648936 100014
rect 648896 96348 648948 96354
rect 648896 96290 648948 96296
rect 649448 95940 649500 95946
rect 649448 95882 649500 95888
rect 649264 95464 649316 95470
rect 649264 95406 649316 95412
rect 648896 95192 648948 95198
rect 648896 95134 648948 95140
rect 648618 92032 648674 92041
rect 648618 91967 648674 91976
rect 647884 86624 647936 86630
rect 647884 86566 647936 86572
rect 647514 82784 647570 82793
rect 647514 82719 647570 82728
rect 629206 81696 629262 81705
rect 629206 81631 629262 81640
rect 628748 81116 628800 81122
rect 628748 81058 628800 81064
rect 629220 79490 629248 81631
rect 642456 81116 642508 81122
rect 642456 81058 642508 81064
rect 632808 80974 633144 81002
rect 629208 79484 629260 79490
rect 629208 79426 629260 79432
rect 631048 78124 631100 78130
rect 631048 78066 631100 78072
rect 631060 77450 631088 78066
rect 631048 77444 631100 77450
rect 631048 77386 631100 77392
rect 628472 77308 628524 77314
rect 628472 77250 628524 77256
rect 628484 75954 628512 77250
rect 628472 75948 628524 75954
rect 628472 75890 628524 75896
rect 628484 75290 628512 75890
rect 631060 75290 631088 77386
rect 632808 77314 632836 80974
rect 636108 80708 636160 80714
rect 636108 80650 636160 80656
rect 633898 78568 633954 78577
rect 633898 78503 633954 78512
rect 633912 77353 633940 78503
rect 633898 77344 633954 77353
rect 632796 77308 632848 77314
rect 633898 77279 633954 77288
rect 636120 77294 636148 80650
rect 639602 77888 639658 77897
rect 639602 77823 639658 77832
rect 632796 77250 632848 77256
rect 633912 75290 633940 77279
rect 636120 77266 636332 77294
rect 628176 75262 628512 75290
rect 631028 75262 631088 75290
rect 633880 75262 633940 75290
rect 636304 75154 636332 77266
rect 639616 75290 639644 77823
rect 642468 75290 642496 81058
rect 643080 80974 643140 81002
rect 643112 78130 643140 80974
rect 646044 80844 646096 80850
rect 646044 80786 646096 80792
rect 645308 79484 645360 79490
rect 645308 79426 645360 79432
rect 643100 78124 643152 78130
rect 643100 78066 643152 78072
rect 645320 75290 645348 79426
rect 639584 75262 639644 75290
rect 642436 75262 642496 75290
rect 645288 75262 645348 75290
rect 636304 75126 636732 75154
rect 646056 69034 646084 80786
rect 646228 79348 646280 79354
rect 646228 79290 646280 79296
rect 646240 69193 646268 79290
rect 648712 77988 648764 77994
rect 648712 77930 648764 77936
rect 646780 76696 646832 76702
rect 646780 76638 646832 76644
rect 646596 75472 646648 75478
rect 646596 75414 646648 75420
rect 646412 75336 646464 75342
rect 646412 75278 646464 75284
rect 646424 74497 646452 75278
rect 646410 74488 646466 74497
rect 646410 74423 646466 74432
rect 646226 69184 646282 69193
rect 646226 69119 646282 69128
rect 646056 69006 646268 69034
rect 646240 67153 646268 69006
rect 646226 67144 646282 67153
rect 646226 67079 646282 67088
rect 646608 64874 646636 75414
rect 646792 74534 646820 76638
rect 646792 74506 647280 74534
rect 647252 71777 647280 74506
rect 647238 71768 647294 71777
rect 647238 71703 647294 71712
rect 646424 64846 646636 64874
rect 646424 59401 646452 64846
rect 648724 62121 648752 77930
rect 648710 62112 648766 62121
rect 648710 62047 648766 62056
rect 646410 59392 646466 59401
rect 646410 59327 646466 59336
rect 624424 57928 624476 57934
rect 624424 57870 624476 57876
rect 648908 57361 648936 95134
rect 649276 86766 649304 95406
rect 649460 94858 649488 95882
rect 649448 94852 649500 94858
rect 649448 94794 649500 94800
rect 649736 88806 649764 100014
rect 650380 97034 650408 100014
rect 650736 97980 650788 97986
rect 650736 97922 650788 97928
rect 650552 97300 650604 97306
rect 650552 97242 650604 97248
rect 650368 97028 650420 97034
rect 650368 96970 650420 96976
rect 650184 96756 650236 96762
rect 650184 96698 650236 96704
rect 649954 95940 650006 95946
rect 649954 95882 650006 95888
rect 649966 95826 649994 95882
rect 649920 95798 649994 95826
rect 649920 95198 649948 95798
rect 649908 95192 649960 95198
rect 649908 95134 649960 95140
rect 649724 88800 649776 88806
rect 649724 88742 649776 88748
rect 650196 87145 650224 96698
rect 650564 95826 650592 97242
rect 650472 95798 650592 95826
rect 650472 89593 650500 95798
rect 650458 89584 650514 89593
rect 650458 89519 650514 89528
rect 650182 87136 650238 87145
rect 650182 87071 650238 87080
rect 649264 86760 649316 86766
rect 649264 86702 649316 86708
rect 650748 84697 650776 97922
rect 651116 97442 651144 100014
rect 651104 97436 651156 97442
rect 651104 97378 651156 97384
rect 651852 97306 651880 100014
rect 651840 97300 651892 97306
rect 651840 97242 651892 97248
rect 652588 96626 652616 100014
rect 652024 96620 652076 96626
rect 652024 96562 652076 96568
rect 652576 96620 652628 96626
rect 652576 96562 652628 96568
rect 651840 95736 651892 95742
rect 651840 95678 651892 95684
rect 651852 90681 651880 95678
rect 651838 90672 651894 90681
rect 651838 90607 651894 90616
rect 652036 86902 652064 96562
rect 653324 96490 653352 100014
rect 653968 97714 653996 100014
rect 653956 97708 654008 97714
rect 653956 97650 654008 97656
rect 654600 97436 654652 97442
rect 654600 97378 654652 97384
rect 654324 97300 654376 97306
rect 654324 97242 654376 97248
rect 654336 96830 654364 97242
rect 654324 96824 654376 96830
rect 654324 96766 654376 96772
rect 652208 96484 652260 96490
rect 652208 96426 652260 96432
rect 653312 96484 653364 96490
rect 653312 96426 653364 96432
rect 652220 92478 652248 96426
rect 653404 95328 653456 95334
rect 653404 95270 653456 95276
rect 652208 92472 652260 92478
rect 652208 92414 652260 92420
rect 652024 86896 652076 86902
rect 652024 86838 652076 86844
rect 653416 86222 653444 95270
rect 654416 93900 654468 93906
rect 654416 93842 654468 93848
rect 654428 86358 654456 93842
rect 654612 93401 654640 97378
rect 654796 96966 654824 100014
rect 655440 97986 655468 100014
rect 655808 100014 655960 100042
rect 656696 100014 656848 100042
rect 657432 100014 657768 100042
rect 655428 97980 655480 97986
rect 655428 97922 655480 97928
rect 655060 97708 655112 97714
rect 655060 97650 655112 97656
rect 654784 96960 654836 96966
rect 654784 96902 654836 96908
rect 655072 94217 655100 97650
rect 655428 96960 655480 96966
rect 655428 96902 655480 96908
rect 655058 94208 655114 94217
rect 655058 94143 655114 94152
rect 655440 93854 655468 96902
rect 655072 93826 655468 93854
rect 654598 93392 654654 93401
rect 654598 93327 654654 93336
rect 655072 88330 655100 93826
rect 655428 92812 655480 92818
rect 655428 92754 655480 92760
rect 655440 92585 655468 92754
rect 655426 92576 655482 92585
rect 655426 92511 655482 92520
rect 655244 92472 655296 92478
rect 655244 92414 655296 92420
rect 655256 91497 655284 92414
rect 655242 91488 655298 91497
rect 655242 91423 655298 91432
rect 655808 89865 655836 100014
rect 656820 97374 656848 100014
rect 656808 97368 656860 97374
rect 656808 97310 656860 97316
rect 657740 95132 657768 100014
rect 658154 99770 658182 100028
rect 658904 100014 659240 100042
rect 659640 100014 659976 100042
rect 660376 100014 660712 100042
rect 658154 99742 658228 99770
rect 658200 97510 658228 99742
rect 659212 97850 659240 100014
rect 659016 97844 659068 97850
rect 659016 97786 659068 97792
rect 659200 97844 659252 97850
rect 659200 97786 659252 97792
rect 658188 97504 658240 97510
rect 658188 97446 658240 97452
rect 659028 97238 659056 97786
rect 659948 97714 659976 100014
rect 659936 97708 659988 97714
rect 659936 97650 659988 97656
rect 659752 97640 659804 97646
rect 659752 97582 659804 97588
rect 658832 97232 658884 97238
rect 658832 97174 658884 97180
rect 659016 97232 659068 97238
rect 659016 97174 659068 97180
rect 658280 97096 658332 97102
rect 658280 97038 658332 97044
rect 658292 95132 658320 97038
rect 658844 95132 658872 97174
rect 659568 96824 659620 96830
rect 659568 96766 659620 96772
rect 659580 95132 659608 96766
rect 659764 95146 659792 97582
rect 660684 96966 660712 100014
rect 662512 97980 662564 97986
rect 662512 97922 662564 97928
rect 661408 97368 661460 97374
rect 661408 97310 661460 97316
rect 660672 96960 660724 96966
rect 660672 96902 660724 96908
rect 660672 96212 660724 96218
rect 660672 96154 660724 96160
rect 659764 95118 660146 95146
rect 660684 95132 660712 96154
rect 661420 95132 661448 97310
rect 661960 97232 662012 97238
rect 661960 97174 662012 97180
rect 661972 95132 662000 97174
rect 662524 95132 662552 97922
rect 663892 97844 663944 97850
rect 663892 97786 663944 97792
rect 663064 97504 663116 97510
rect 663064 97446 663116 97452
rect 663076 95132 663104 97446
rect 663248 96960 663300 96966
rect 663248 96902 663300 96908
rect 656164 94852 656216 94858
rect 656164 94794 656216 94800
rect 655794 89856 655850 89865
rect 655794 89791 655850 89800
rect 655060 88324 655112 88330
rect 655060 88266 655112 88272
rect 656176 86494 656204 94794
rect 658556 88800 658608 88806
rect 662328 88800 662380 88806
rect 658608 88748 658858 88754
rect 658556 88742 658858 88748
rect 658568 88726 658858 88742
rect 661986 88748 662328 88754
rect 661986 88742 662380 88748
rect 661986 88726 662368 88742
rect 658306 88330 658504 88346
rect 658306 88324 658516 88330
rect 658306 88318 658464 88324
rect 658464 88266 658516 88272
rect 656164 86488 656216 86494
rect 656164 86430 656216 86436
rect 654416 86352 654468 86358
rect 654416 86294 654468 86300
rect 657188 86222 657216 88196
rect 657740 86902 657768 88196
rect 659580 86970 659608 88196
rect 659568 86964 659620 86970
rect 659568 86906 659620 86912
rect 657728 86896 657780 86902
rect 657728 86838 657780 86844
rect 660132 86630 660160 88196
rect 660120 86624 660172 86630
rect 660120 86566 660172 86572
rect 660684 86494 660712 88196
rect 661420 86766 661448 88196
rect 661408 86760 661460 86766
rect 661408 86702 661460 86708
rect 660672 86488 660724 86494
rect 660672 86430 660724 86436
rect 662524 86358 662552 88196
rect 663260 86970 663288 96902
rect 663708 96076 663760 96082
rect 663708 96018 663760 96024
rect 663720 95962 663748 96018
rect 663720 95934 663840 95962
rect 663812 92970 663840 95934
rect 663720 92942 663840 92970
rect 663720 92857 663748 92942
rect 663706 92848 663762 92857
rect 663706 92783 663762 92792
rect 663904 88806 663932 97786
rect 665364 97708 665416 97714
rect 665364 97650 665416 97656
rect 664352 96620 664404 96626
rect 664352 96562 664404 96568
rect 664168 96348 664220 96354
rect 664168 96290 664220 96296
rect 664180 89865 664208 96290
rect 664364 90681 664392 96562
rect 665180 96484 665232 96490
rect 665180 96426 665232 96432
rect 664536 95940 664588 95946
rect 664536 95882 664588 95888
rect 664548 91769 664576 95882
rect 664534 91760 664590 91769
rect 664534 91695 664590 91704
rect 664350 90672 664406 90681
rect 664350 90607 664406 90616
rect 664166 89856 664222 89865
rect 664166 89791 664222 89800
rect 665192 89049 665220 96426
rect 665376 93401 665404 97650
rect 665362 93392 665418 93401
rect 665362 93327 665418 93336
rect 665178 89040 665234 89049
rect 665178 88975 665234 88984
rect 663892 88800 663944 88806
rect 663892 88742 663944 88748
rect 663248 86964 663300 86970
rect 663248 86906 663300 86912
rect 662512 86352 662564 86358
rect 662512 86294 662564 86300
rect 653404 86216 653456 86222
rect 653404 86158 653456 86164
rect 657176 86216 657228 86222
rect 657176 86158 657228 86164
rect 650734 84688 650790 84697
rect 650734 84623 650790 84632
rect 649080 80980 649132 80986
rect 649080 80922 649132 80928
rect 649092 64433 649120 80922
rect 662420 76560 662472 76566
rect 662420 76502 662472 76508
rect 649078 64424 649134 64433
rect 649078 64359 649134 64368
rect 648894 57352 648950 57361
rect 648894 57287 648950 57296
rect 661590 47789 661646 47798
rect 661590 47724 661646 47733
rect 661604 46510 661632 47724
rect 662432 47433 662460 76502
rect 666572 75206 666600 103486
rect 667938 102776 667994 102785
rect 667938 102711 667994 102720
rect 667952 100026 667980 102711
rect 668136 100162 668164 106111
rect 668596 104553 668624 111823
rect 670804 106214 670832 113146
rect 671540 107817 671568 130863
rect 671908 115841 671936 166903
rect 672092 140457 672120 183495
rect 672262 182064 672318 182073
rect 672262 181999 672318 182008
rect 672276 164257 672304 181999
rect 672538 175264 672594 175273
rect 672538 175199 672594 175208
rect 672262 164248 672318 164257
rect 672262 164183 672318 164192
rect 672078 140448 672134 140457
rect 672078 140383 672134 140392
rect 672552 130529 672580 175199
rect 672538 130520 672594 130529
rect 672538 130455 672594 130464
rect 672736 124137 672764 210151
rect 672920 180794 672948 226358
rect 673104 222194 673132 227344
rect 673196 227202 673224 227718
rect 673472 227372 673500 227888
rect 673656 227508 673684 227990
rect 673656 227480 673776 227508
rect 673472 227344 673684 227372
rect 673196 227174 673500 227202
rect 673472 227089 673500 227174
rect 673458 227080 673514 227089
rect 673458 227015 673514 227024
rect 673656 226930 673684 227344
rect 672828 180766 672948 180794
rect 673012 222166 673132 222194
rect 673196 226902 673684 226930
rect 673196 222194 673224 226902
rect 673550 225312 673606 225321
rect 673550 225247 673606 225256
rect 673564 224954 673592 225247
rect 673564 224926 673684 224954
rect 673196 222166 673316 222194
rect 672828 176654 672856 180766
rect 673012 177993 673040 222166
rect 673288 215294 673316 222166
rect 673656 220810 673684 224926
rect 673564 220782 673684 220810
rect 673564 220697 673592 220782
rect 673550 220688 673606 220697
rect 673550 220623 673606 220632
rect 673550 220280 673606 220289
rect 673550 220215 673606 220224
rect 673564 218657 673592 220215
rect 673550 218648 673606 218657
rect 673550 218583 673606 218592
rect 673458 216200 673514 216209
rect 673458 216135 673514 216144
rect 673472 216050 673500 216135
rect 673196 215266 673316 215294
rect 673380 216022 673500 216050
rect 673196 201770 673224 215266
rect 673380 201929 673408 216022
rect 673550 206952 673606 206961
rect 673550 206887 673606 206896
rect 673366 201920 673422 201929
rect 673366 201855 673422 201864
rect 673196 201742 673316 201770
rect 673288 201657 673316 201742
rect 673274 201648 673330 201657
rect 673274 201583 673330 201592
rect 673564 197713 673592 206887
rect 673550 197704 673606 197713
rect 673550 197639 673606 197648
rect 672998 177984 673054 177993
rect 672998 177919 673054 177928
rect 672828 176626 672948 176654
rect 672920 173097 672948 176626
rect 673366 174448 673422 174457
rect 673366 174383 673422 174392
rect 672906 173088 672962 173097
rect 672906 173023 672962 173032
rect 673182 169960 673238 169969
rect 673182 169895 673238 169904
rect 672998 169144 673054 169153
rect 672998 169079 673054 169088
rect 673012 153105 673040 169079
rect 672998 153096 673054 153105
rect 672998 153031 673054 153040
rect 673196 151745 673224 169895
rect 673182 151736 673238 151745
rect 673182 151671 673238 151680
rect 673380 129713 673408 174383
rect 673748 168473 673776 227480
rect 673918 227080 673974 227089
rect 673918 227015 673974 227024
rect 673932 212945 673960 227015
rect 674102 226264 674158 226273
rect 674102 226199 674158 226208
rect 674116 220289 674144 226199
rect 674102 220280 674158 220289
rect 674102 220215 674158 220224
rect 674484 220130 674512 230132
rect 675864 229906 675892 230687
rect 676770 230480 676826 230489
rect 676770 230415 676826 230424
rect 676586 230208 676642 230217
rect 676586 230143 676642 230152
rect 675852 229900 675904 229906
rect 675852 229842 675904 229848
rect 675114 229664 675170 229673
rect 675170 229634 675892 229650
rect 675170 229628 675904 229634
rect 675170 229622 675852 229628
rect 675114 229599 675170 229608
rect 675852 229570 675904 229576
rect 675114 229392 675170 229401
rect 675852 229356 675904 229362
rect 675170 229336 675852 229344
rect 675114 229327 675852 229336
rect 675128 229316 675852 229327
rect 675852 229298 675904 229304
rect 675114 229120 675170 229129
rect 675170 229090 675892 229106
rect 675170 229084 675904 229090
rect 675170 229078 675852 229084
rect 675114 229055 675170 229064
rect 675852 229026 675904 229032
rect 676404 229084 676456 229090
rect 676404 229026 676456 229032
rect 675114 228848 675170 228857
rect 675170 228818 675892 228834
rect 675170 228812 675904 228818
rect 675170 228806 675852 228812
rect 675114 228783 675170 228792
rect 675852 228754 675904 228760
rect 676220 228812 676272 228818
rect 676220 228754 676272 228760
rect 675390 226808 675446 226817
rect 675390 226743 675446 226752
rect 675022 226536 675078 226545
rect 675022 226471 675078 226480
rect 674838 224360 674894 224369
rect 674838 224295 674894 224304
rect 674852 222193 674880 224295
rect 674838 222184 674894 222193
rect 674838 222119 674894 222128
rect 674654 221912 674710 221921
rect 674654 221847 674710 221856
rect 674392 220102 674512 220130
rect 674392 219994 674420 220102
rect 674116 219966 674420 219994
rect 673918 212936 673974 212945
rect 673918 212871 673974 212880
rect 673918 209672 673974 209681
rect 673918 209607 673974 209616
rect 673932 203561 673960 209607
rect 673918 203552 673974 203561
rect 673918 203487 673974 203496
rect 674116 179489 674144 219966
rect 674668 217274 674696 221847
rect 675036 219745 675064 226471
rect 675206 225584 675262 225593
rect 675206 225519 675262 225528
rect 675022 219736 675078 219745
rect 675022 219671 675078 219680
rect 674838 219056 674894 219065
rect 674838 218991 674894 219000
rect 674392 217246 674696 217274
rect 674102 179480 674158 179489
rect 674102 179415 674158 179424
rect 674392 177313 674420 217246
rect 674852 216730 674880 218991
rect 675022 217832 675078 217841
rect 675022 217767 675078 217776
rect 674852 216702 674972 216730
rect 674746 216608 674802 216617
rect 674746 216543 674802 216552
rect 674562 215384 674618 215393
rect 674562 215319 674618 215328
rect 674378 177304 674434 177313
rect 674378 177239 674434 177248
rect 674286 176896 674342 176905
rect 674286 176831 674342 176840
rect 673918 176080 673974 176089
rect 673918 176015 673974 176024
rect 673734 168464 673790 168473
rect 673734 168399 673790 168408
rect 673932 131345 673960 176015
rect 674102 169552 674158 169561
rect 674102 169487 674158 169496
rect 674116 155417 674144 169487
rect 674102 155408 674158 155417
rect 674102 155343 674158 155352
rect 674300 132161 674328 176831
rect 674576 175681 674604 215319
rect 674760 205057 674788 216543
rect 674746 205048 674802 205057
rect 674746 204983 674802 204992
rect 674944 204513 674972 216702
rect 675036 212534 675064 217767
rect 675220 216889 675248 225519
rect 675206 216880 675262 216889
rect 675206 216815 675262 216824
rect 675206 215384 675262 215393
rect 675206 215319 675262 215328
rect 675036 212506 675156 212534
rect 674930 204504 674986 204513
rect 674930 204439 674986 204448
rect 674838 204232 674894 204241
rect 674838 204167 674894 204176
rect 674852 204049 674880 204167
rect 675128 204082 675156 212506
rect 675220 210474 675248 215319
rect 675404 215294 675432 226743
rect 676036 220720 676088 220726
rect 676034 220688 676036 220697
rect 676088 220688 676090 220697
rect 676034 220623 676090 220632
rect 676034 220416 676090 220425
rect 676232 220402 676260 228754
rect 676416 227390 676444 229026
rect 676404 227384 676456 227390
rect 676404 227326 676456 227332
rect 676090 220374 676260 220402
rect 676034 220351 676090 220360
rect 675852 218680 675904 218686
rect 675680 218628 675852 218634
rect 675680 218622 675904 218628
rect 675680 218606 675892 218622
rect 675680 218385 675708 218606
rect 675666 218376 675722 218385
rect 675666 218311 675722 218320
rect 676404 218136 676456 218142
rect 676404 218078 676456 218084
rect 675404 215266 675708 215294
rect 675680 214577 675708 215266
rect 675944 215144 675996 215150
rect 675942 215112 675944 215121
rect 675996 215112 675998 215121
rect 675942 215047 675998 215056
rect 675666 214568 675722 214577
rect 675666 214503 675722 214512
rect 676416 214146 676444 218078
rect 676600 215294 676628 230143
rect 676784 215294 676812 230415
rect 676956 229900 677008 229906
rect 676956 229842 677008 229848
rect 676968 229242 676996 229842
rect 677140 229628 677192 229634
rect 677140 229570 677192 229576
rect 676232 214118 676444 214146
rect 676508 215266 676628 215294
rect 676692 215266 676812 215294
rect 676876 229214 676996 229242
rect 677152 229242 677180 229570
rect 677324 229356 677376 229362
rect 677324 229298 677376 229304
rect 677152 229214 677272 229242
rect 675852 213988 675904 213994
rect 675852 213930 675904 213936
rect 675220 210446 675340 210474
rect 675312 204241 675340 210446
rect 675864 208321 675892 213930
rect 676034 213480 676090 213489
rect 676232 213466 676260 214118
rect 676508 213994 676536 215266
rect 676496 213988 676548 213994
rect 676496 213930 676548 213936
rect 676090 213438 676260 213466
rect 676034 213415 676090 213424
rect 676034 213208 676090 213217
rect 676692 213194 676720 215266
rect 676090 213166 676720 213194
rect 676034 213143 676090 213152
rect 676876 209681 676904 229214
rect 677048 227384 677100 227390
rect 677048 227326 677100 227332
rect 677060 218686 677088 227326
rect 677048 218680 677100 218686
rect 677048 218622 677100 218628
rect 677244 215150 677272 229214
rect 677336 224954 677364 229298
rect 677336 224926 677456 224954
rect 677428 220726 677456 224926
rect 677416 220720 677468 220726
rect 677416 220662 677468 220668
rect 677612 218142 677640 231202
rect 677600 218136 677652 218142
rect 677600 218078 677652 218084
rect 677232 215144 677284 215150
rect 677232 215086 677284 215092
rect 676862 209672 676918 209681
rect 676862 209607 676918 209616
rect 675850 208312 675906 208321
rect 675850 208247 675906 208256
rect 677796 206961 677824 233650
rect 679254 223816 679310 223825
rect 679254 223751 679310 223760
rect 679268 223582 679296 223751
rect 679256 223576 679308 223582
rect 679256 223518 679308 223524
rect 679636 220697 679664 234534
rect 679992 234388 680044 234394
rect 679992 234330 680044 234336
rect 679808 234252 679860 234258
rect 679808 234194 679860 234200
rect 679820 221513 679848 234194
rect 680004 222329 680032 234330
rect 683854 234152 683910 234161
rect 683854 234087 683910 234096
rect 683302 233880 683358 233889
rect 683302 233815 683358 233824
rect 680176 232552 680228 232558
rect 680176 232494 680228 232500
rect 680188 223582 680216 232494
rect 680176 223576 680228 223582
rect 680176 223518 680228 223524
rect 683316 223145 683344 233815
rect 683488 233436 683540 233442
rect 683488 233378 683540 233384
rect 683302 223136 683358 223145
rect 683302 223071 683358 223080
rect 679990 222320 680046 222329
rect 679990 222255 680046 222264
rect 679806 221504 679862 221513
rect 679806 221439 679862 221448
rect 679622 220688 679678 220697
rect 679622 220623 679678 220632
rect 683500 219881 683528 233378
rect 683868 222737 683896 234087
rect 703694 224196 703722 224264
rect 704154 224196 704182 224264
rect 704614 224196 704642 224264
rect 705074 224196 705102 224264
rect 705534 224196 705562 224264
rect 705994 224196 706022 224264
rect 706454 224196 706482 224264
rect 706914 224196 706942 224264
rect 707374 224196 707402 224264
rect 707834 224196 707862 224264
rect 708294 224196 708322 224264
rect 708754 224196 708782 224264
rect 709214 224196 709242 224264
rect 683854 222728 683910 222737
rect 683854 222663 683910 222672
rect 683486 219872 683542 219881
rect 683486 219807 683542 219816
rect 683302 213344 683358 213353
rect 683302 213279 683358 213288
rect 683118 212528 683174 212537
rect 683118 212463 683174 212472
rect 683132 211177 683160 212463
rect 683118 211168 683174 211177
rect 683118 211103 683174 211112
rect 683316 210361 683344 213279
rect 683302 210352 683358 210361
rect 683302 210287 683358 210296
rect 677782 206952 677838 206961
rect 677782 206887 677838 206896
rect 675758 205592 675814 205601
rect 675758 205527 675814 205536
rect 675772 205323 675800 205527
rect 675482 205048 675538 205057
rect 675482 204983 675538 204992
rect 675496 204680 675524 204983
rect 675482 204504 675538 204513
rect 675482 204439 675538 204448
rect 675298 204232 675354 204241
rect 675298 204167 675354 204176
rect 675128 204054 675248 204082
rect 674852 204021 674972 204049
rect 674944 195974 674972 204021
rect 675220 202874 675248 204054
rect 675496 204035 675524 204439
rect 675128 202846 675248 202874
rect 675128 202209 675156 202846
rect 675128 202181 675418 202209
rect 675482 201920 675538 201929
rect 675482 201855 675538 201864
rect 675496 201620 675524 201855
rect 675128 200994 675418 201022
rect 675128 197985 675156 200994
rect 675298 200832 675354 200841
rect 675298 200767 675354 200776
rect 675114 197976 675170 197985
rect 675114 197911 675170 197920
rect 675312 196466 675340 200767
rect 675758 200696 675814 200705
rect 675758 200631 675814 200640
rect 675772 200328 675800 200631
rect 675574 198248 675630 198257
rect 675574 198183 675630 198192
rect 675588 197880 675616 198183
rect 675496 197169 675524 197336
rect 675482 197160 675538 197169
rect 675482 197095 675538 197104
rect 675758 197160 675814 197169
rect 675758 197095 675814 197104
rect 675772 196656 675800 197095
rect 675312 196438 675432 196466
rect 675404 196044 675432 196438
rect 674852 195946 674972 195974
rect 674852 194834 674880 195946
rect 674852 194806 675418 194834
rect 675666 193216 675722 193225
rect 675666 193151 675722 193160
rect 675680 192984 675708 193151
rect 675404 191978 675432 192372
rect 675312 191950 675432 191978
rect 675312 190369 675340 191950
rect 675758 191584 675814 191593
rect 675758 191519 675814 191528
rect 675772 191148 675800 191519
rect 675298 190360 675354 190369
rect 675298 190295 675354 190304
rect 683118 186960 683174 186969
rect 683118 186895 683174 186904
rect 676494 181384 676550 181393
rect 676494 181319 676550 181328
rect 676034 178120 676090 178129
rect 676508 178106 676536 181319
rect 683132 178809 683160 186895
rect 703694 179180 703722 179316
rect 704154 179180 704182 179316
rect 704614 179180 704642 179316
rect 705074 179180 705102 179316
rect 705534 179180 705562 179316
rect 705994 179180 706022 179316
rect 706454 179180 706482 179316
rect 706914 179180 706942 179316
rect 707374 179180 707402 179316
rect 707834 179180 707862 179316
rect 708294 179180 708322 179316
rect 708754 179180 708782 179316
rect 709214 179180 709242 179316
rect 683118 178800 683174 178809
rect 683118 178735 683174 178744
rect 676090 178078 676536 178106
rect 676034 178055 676090 178064
rect 674562 175672 674618 175681
rect 674562 175607 674618 175616
rect 678242 173224 678298 173233
rect 678242 173159 678298 173168
rect 674838 172816 674894 172825
rect 674838 172751 674894 172760
rect 674470 168736 674526 168745
rect 674470 168671 674526 168680
rect 674484 151042 674512 168671
rect 674852 157593 674880 172751
rect 676586 170776 676642 170785
rect 676586 170711 676642 170720
rect 676034 167920 676090 167929
rect 676034 167855 676090 167864
rect 676048 165617 676076 167855
rect 676600 166433 676628 170711
rect 676586 166424 676642 166433
rect 676586 166359 676642 166368
rect 676034 165608 676090 165617
rect 676034 165543 676090 165552
rect 678256 162858 678284 173159
rect 681002 171592 681058 171601
rect 681002 171527 681058 171536
rect 679622 171184 679678 171193
rect 679622 171119 679678 171128
rect 676128 162852 676180 162858
rect 676128 162794 676180 162800
rect 678244 162852 678296 162858
rect 678244 162794 678296 162800
rect 675944 162648 675996 162654
rect 675944 162590 675996 162596
rect 675956 161945 675984 162590
rect 675942 161936 675998 161945
rect 675942 161871 675998 161880
rect 675852 161764 675904 161770
rect 675852 161706 675904 161712
rect 675864 161242 675892 161706
rect 676140 161401 676168 162794
rect 679636 162654 679664 171119
rect 679624 162648 679676 162654
rect 679624 162590 679676 162596
rect 681016 161770 681044 171527
rect 681004 161764 681056 161770
rect 681004 161706 681056 161712
rect 676126 161392 676182 161401
rect 676126 161327 676182 161336
rect 675312 161214 675892 161242
rect 675312 159678 675340 161214
rect 675758 160712 675814 160721
rect 675758 160647 675814 160656
rect 675772 160344 675800 160647
rect 675312 159650 675418 159678
rect 675758 159352 675814 159361
rect 675758 159287 675814 159296
rect 675772 159052 675800 159287
rect 674838 157584 674894 157593
rect 674838 157519 674894 157528
rect 675482 157584 675538 157593
rect 675482 157519 675538 157528
rect 675496 157216 675524 157519
rect 675390 157040 675446 157049
rect 675390 156975 675446 156984
rect 675404 156643 675432 156975
rect 675758 156360 675814 156369
rect 675758 156295 675814 156304
rect 675772 155992 675800 156295
rect 675114 155408 675170 155417
rect 675170 155366 675340 155394
rect 675114 155343 675170 155352
rect 675312 155258 675340 155366
rect 675404 155258 675432 155380
rect 675312 155230 675432 155258
rect 675114 153096 675170 153105
rect 675114 153031 675170 153040
rect 675758 153096 675814 153105
rect 675758 153031 675814 153040
rect 675128 152334 675156 153031
rect 675772 152864 675800 153031
rect 675128 152306 675418 152334
rect 675114 151736 675170 151745
rect 675170 151680 675418 151689
rect 675114 151671 675418 151680
rect 675128 151661 675418 151671
rect 674484 151014 675418 151042
rect 675128 149821 675418 149849
rect 675128 147665 675156 149821
rect 675666 148472 675722 148481
rect 675666 148407 675722 148416
rect 675680 147968 675708 148407
rect 675114 147656 675170 147665
rect 675114 147591 675170 147600
rect 675666 147656 675722 147665
rect 675666 147591 675722 147600
rect 675680 147356 675708 147591
rect 675772 146033 675800 146132
rect 675758 146024 675814 146033
rect 675758 145959 675814 145968
rect 683118 135960 683174 135969
rect 683118 135895 683174 135904
rect 675850 134600 675906 134609
rect 675850 134535 675906 134544
rect 675864 133958 675892 134535
rect 675852 133952 675904 133958
rect 675852 133894 675904 133900
rect 676496 133952 676548 133958
rect 676496 133894 676548 133900
rect 676508 133113 676536 133894
rect 676494 133104 676550 133113
rect 676494 133039 676550 133048
rect 683132 132705 683160 135895
rect 703694 133892 703722 134028
rect 704154 133892 704182 134028
rect 704614 133892 704642 134028
rect 705074 133892 705102 134028
rect 705534 133892 705562 134028
rect 705994 133892 706022 134028
rect 706454 133892 706482 134028
rect 706914 133892 706942 134028
rect 707374 133892 707402 134028
rect 707834 133892 707862 134028
rect 708294 133892 708322 134028
rect 708754 133892 708782 134028
rect 709214 133892 709242 134028
rect 683118 132696 683174 132705
rect 683118 132631 683174 132640
rect 674286 132152 674342 132161
rect 674286 132087 674342 132096
rect 673918 131336 673974 131345
rect 673918 131271 673974 131280
rect 675942 130112 675998 130121
rect 675942 130047 675998 130056
rect 673366 129704 673422 129713
rect 673366 129639 673422 129648
rect 674102 129296 674158 129305
rect 674102 129231 674158 129240
rect 673090 126032 673146 126041
rect 673090 125967 673146 125976
rect 672906 124400 672962 124409
rect 672906 124335 672962 124344
rect 672722 124128 672778 124137
rect 672722 124063 672778 124072
rect 672538 123856 672594 123865
rect 672538 123791 672594 123800
rect 672354 123176 672410 123185
rect 672354 123111 672410 123120
rect 672368 120193 672396 123111
rect 672354 120184 672410 120193
rect 672354 120119 672410 120128
rect 672552 120034 672580 123791
rect 672368 120006 672580 120034
rect 671894 115832 671950 115841
rect 671894 115767 671950 115776
rect 671526 107808 671582 107817
rect 671526 107743 671582 107752
rect 672368 106457 672396 120006
rect 672920 119898 672948 124335
rect 672552 119870 672948 119898
rect 672552 110265 672580 119870
rect 672722 117872 672778 117881
rect 672722 117807 672778 117816
rect 672736 111081 672764 117807
rect 673104 111489 673132 125967
rect 673366 123584 673422 123593
rect 673366 123519 673422 123528
rect 673090 111480 673146 111489
rect 673090 111415 673146 111424
rect 672722 111072 672778 111081
rect 672722 111007 672778 111016
rect 672538 110256 672594 110265
rect 672538 110191 672594 110200
rect 672354 106448 672410 106457
rect 672354 106383 672410 106392
rect 670792 106208 670844 106214
rect 670792 106150 670844 106156
rect 673380 105641 673408 123519
rect 673918 121680 673974 121689
rect 673918 121615 673974 121624
rect 673932 117881 673960 121615
rect 673918 117872 673974 117881
rect 673918 117807 673974 117816
rect 674116 111897 674144 129231
rect 675956 128353 675984 130047
rect 674286 128344 674342 128353
rect 674286 128279 674342 128288
rect 675942 128344 675998 128353
rect 675942 128279 675998 128288
rect 674102 111888 674158 111897
rect 674102 111823 674158 111832
rect 673366 105632 673422 105641
rect 673366 105567 673422 105576
rect 668582 104544 668638 104553
rect 668582 104479 668638 104488
rect 668596 103514 668624 104479
rect 668320 103486 668624 103514
rect 668124 100156 668176 100162
rect 668124 100098 668176 100104
rect 667940 100020 667992 100026
rect 667940 99962 667992 99968
rect 668320 95849 668348 103486
rect 674300 102377 674328 128279
rect 682382 127800 682438 127809
rect 682382 127735 682438 127744
rect 674838 127664 674894 127673
rect 674838 127599 674894 127608
rect 674654 125624 674710 125633
rect 674654 125559 674710 125568
rect 674470 125216 674526 125225
rect 674470 125151 674526 125160
rect 674484 104666 674512 125151
rect 674668 110786 674696 125559
rect 674852 112010 674880 127599
rect 675022 126440 675078 126449
rect 675022 126375 675078 126384
rect 675036 114493 675064 126375
rect 682396 117298 682424 127735
rect 675852 117292 675904 117298
rect 675852 117234 675904 117240
rect 682384 117292 682436 117298
rect 682384 117234 682436 117240
rect 675864 117178 675892 117234
rect 675312 117150 675892 117178
rect 675312 115138 675340 117150
rect 675312 115110 675418 115138
rect 675036 114465 675418 114493
rect 675312 113818 675418 113846
rect 675312 113121 675340 113818
rect 675298 113112 675354 113121
rect 675298 113047 675354 113056
rect 674852 111982 675418 112010
rect 675114 111480 675170 111489
rect 675170 111438 675418 111466
rect 675114 111415 675170 111424
rect 675312 110894 675432 110922
rect 675312 110786 675340 110894
rect 674668 110758 675340 110786
rect 675404 110772 675432 110894
rect 674654 110256 674710 110265
rect 674710 110214 674880 110242
rect 674654 110191 674710 110200
rect 674852 110174 674880 110214
rect 674852 110146 675418 110174
rect 675666 108080 675722 108089
rect 675666 108015 675722 108024
rect 675680 107644 675708 108015
rect 675312 107222 675432 107250
rect 675312 107114 675340 107222
rect 675128 107086 675340 107114
rect 675404 107100 675432 107222
rect 675128 106457 675156 107086
rect 675114 106448 675170 106457
rect 675114 106383 675170 106392
rect 675772 106185 675800 106488
rect 675758 106176 675814 106185
rect 675758 106111 675814 106120
rect 675312 105862 675432 105890
rect 675312 105822 675340 105862
rect 675128 105794 675340 105822
rect 675404 105808 675432 105862
rect 675128 105641 675156 105794
rect 675114 105632 675170 105641
rect 675114 105567 675170 105576
rect 674484 104638 675340 104666
rect 675312 104530 675340 104638
rect 675404 104530 675432 104652
rect 675312 104502 675432 104530
rect 675758 103184 675814 103193
rect 675758 103119 675814 103128
rect 675772 102816 675800 103119
rect 675666 102640 675722 102649
rect 675666 102575 675722 102584
rect 674286 102368 674342 102377
rect 674286 102303 674342 102312
rect 675680 102136 675708 102575
rect 675758 101416 675814 101425
rect 675758 101351 675814 101360
rect 675772 100980 675800 101351
rect 668306 95840 668362 95849
rect 668306 95775 668362 95784
rect 666560 75200 666612 75206
rect 666560 75142 666612 75148
rect 663798 48512 663854 48521
rect 663798 48447 663854 48456
rect 662418 47424 662474 47433
rect 662418 47359 662474 47368
rect 623044 46504 623096 46510
rect 623044 46446 623096 46452
rect 661592 46504 661644 46510
rect 661592 46446 661644 46452
rect 471058 43888 471114 43897
rect 471058 43823 471114 43832
rect 464342 43616 464398 43625
rect 464342 43551 464398 43560
rect 465814 43208 465870 43217
rect 465814 43143 465870 43152
rect 463712 43030 463924 43058
rect 463698 42936 463754 42945
rect 463698 42871 463754 42880
rect 462964 42492 463016 42498
rect 462964 42434 463016 42440
rect 463712 42378 463740 42871
rect 463896 42770 463924 43030
rect 463884 42764 463936 42770
rect 463884 42706 463936 42712
rect 465828 42500 465856 43143
rect 463712 42350 464036 42378
rect 461122 42256 461178 42265
rect 461122 42191 461178 42200
rect 471072 42106 471100 43823
rect 518806 42800 518862 42809
rect 518806 42735 518862 42744
rect 518820 42364 518848 42735
rect 663812 42231 663840 48447
rect 663800 42225 663852 42231
rect 663800 42167 663852 42173
rect 515402 42120 515458 42129
rect 459940 42078 460368 42106
rect 471072 42078 471408 42106
rect 515154 42078 515402 42106
rect 520922 42120 520978 42129
rect 520674 42078 520922 42106
rect 515402 42055 515458 42064
rect 522026 42120 522082 42129
rect 521870 42078 522026 42106
rect 520922 42055 520978 42064
rect 526442 42120 526498 42129
rect 526194 42078 526442 42106
rect 522026 42055 522082 42064
rect 529570 42120 529626 42129
rect 529322 42078 529570 42106
rect 526442 42055 526498 42064
rect 529570 42055 529626 42064
rect 404452 41472 404504 41478
rect 404452 41414 404504 41420
rect 420736 41472 420788 41478
rect 420736 41414 420788 41420
rect 426900 41472 426952 41478
rect 426900 41414 426952 41420
rect 459192 41472 459244 41478
rect 459192 41414 459244 41420
rect 141698 40488 141754 40497
rect 141698 40423 141754 40432
rect 141712 39984 141740 40423
<< via2 >>
rect 426346 1007140 426402 1007176
rect 426346 1007120 426348 1007140
rect 426348 1007120 426400 1007140
rect 426400 1007120 426402 1007140
rect 358542 1007004 358598 1007040
rect 358542 1006984 358544 1007004
rect 358544 1006984 358596 1007004
rect 358596 1006984 358598 1007004
rect 359370 1006868 359426 1006904
rect 359370 1006848 359372 1006868
rect 359372 1006848 359424 1006868
rect 359424 1006848 359426 1006868
rect 360198 1006732 360254 1006768
rect 360198 1006712 360200 1006732
rect 360200 1006712 360252 1006732
rect 360252 1006712 360254 1006732
rect 101954 1006596 102010 1006632
rect 101954 1006576 101956 1006596
rect 101956 1006576 102008 1006596
rect 102008 1006576 102010 1006596
rect 82266 995696 82322 995752
rect 86498 995696 86554 995752
rect 88982 995696 89038 995752
rect 89626 995696 89682 995752
rect 90270 995696 90326 995752
rect 77022 995016 77078 995072
rect 78678 994744 78734 994800
rect 84658 995424 84714 995480
rect 86038 994472 86094 994528
rect 85026 994200 85082 994256
rect 92478 996920 92534 996976
rect 92662 995968 92718 996024
rect 92478 994472 92534 994528
rect 93122 995696 93178 995752
rect 92846 995424 92902 995480
rect 92662 994200 92718 994256
rect 98274 1006460 98330 1006496
rect 98274 1006440 98276 1006460
rect 98276 1006440 98328 1006460
rect 98328 1006440 98330 1006460
rect 103978 1006324 104034 1006360
rect 103978 1006304 103980 1006324
rect 103980 1006304 104032 1006324
rect 104032 1006304 104034 1006324
rect 108486 1006324 108542 1006360
rect 108486 1006304 108488 1006324
rect 108488 1006304 108540 1006324
rect 108540 1006304 108542 1006324
rect 99470 1006052 99526 1006088
rect 99470 1006032 99472 1006052
rect 99472 1006032 99524 1006052
rect 99524 1006032 99526 1006052
rect 100298 1002652 100354 1002688
rect 100298 1002632 100300 1002652
rect 100300 1002632 100352 1002652
rect 100352 1002632 100354 1002652
rect 94686 997192 94742 997248
rect 87878 993928 87934 993984
rect 93306 993928 93362 993984
rect 41786 967136 41842 967192
rect 42338 966728 42394 966784
rect 42430 964688 42486 964744
rect 42430 963328 42486 963384
rect 42246 962920 42302 962976
rect 41786 962104 41842 962160
rect 42246 961968 42302 962024
rect 41786 959792 41842 959848
rect 41786 959112 41842 959168
rect 42430 958704 42486 958760
rect 41786 957752 41842 957808
rect 41786 955440 41842 955496
rect 41786 954624 41842 954680
rect 41786 954352 41842 954408
rect 35162 952856 35218 952912
rect 31758 946600 31814 946656
rect 28722 942656 28778 942712
rect 33782 938168 33838 938224
rect 37922 952448 37978 952504
rect 35806 943064 35862 943120
rect 35806 941840 35862 941896
rect 35806 940208 35862 940264
rect 36542 938984 36598 939040
rect 39302 952176 39358 952232
rect 37922 938576 37978 938632
rect 35162 937760 35218 937816
rect 40038 951632 40094 951688
rect 39762 943744 39818 943800
rect 39302 937352 39358 937408
rect 39762 935720 39818 935776
rect 40038 934496 40094 934552
rect 42062 940616 42118 940672
rect 42062 939800 42118 939856
rect 41970 935584 42026 935640
rect 43442 966728 43498 966784
rect 43258 964688 43314 964744
rect 42982 963328 43038 963384
rect 42798 936944 42854 937000
rect 43442 962920 43498 962976
rect 43258 935312 43314 935368
rect 44270 961968 44326 962024
rect 43442 934904 43498 934960
rect 44454 958704 44510 958760
rect 46202 946600 46258 946656
rect 45558 943472 45614 943528
rect 44822 941432 44878 941488
rect 44638 941024 44694 941080
rect 44454 936128 44510 936184
rect 44270 934088 44326 934144
rect 42982 933680 43038 933736
rect 43350 933272 43406 933328
rect 42338 932864 42394 932920
rect 41602 911920 41658 911976
rect 41418 911648 41474 911704
rect 43074 892744 43130 892800
rect 42844 892492 42900 892528
rect 42844 892472 42846 892492
rect 42846 892472 42898 892492
rect 42898 892472 42900 892492
rect 42936 892254 42992 892256
rect 42936 892202 42938 892254
rect 42938 892202 42990 892254
rect 42990 892202 42992 892254
rect 42936 892200 42992 892202
rect 41602 885400 41658 885456
rect 41418 885128 41474 885184
rect 35806 817264 35862 817320
rect 35806 816448 35862 816504
rect 42062 884584 42118 884640
rect 35806 814816 35862 814872
rect 41326 812776 41382 812832
rect 40958 812368 41014 812424
rect 35162 811552 35218 811608
rect 35898 811144 35954 811200
rect 40774 808288 40830 808344
rect 40590 805160 40646 805216
rect 40774 805024 40830 805080
rect 41142 811960 41198 812016
rect 40958 804752 41014 804808
rect 41786 808696 41842 808752
rect 43166 810736 43222 810792
rect 42798 809920 42854 809976
rect 42338 806656 42394 806712
rect 41142 804480 41198 804536
rect 41694 802460 41750 802496
rect 41694 802440 41696 802460
rect 41696 802440 41748 802460
rect 41748 802440 41750 802460
rect 41786 800264 41842 800320
rect 41786 799856 41842 799912
rect 42614 802440 42670 802496
rect 42246 798904 42302 798960
rect 42430 798088 42486 798144
rect 42154 797816 42210 797872
rect 42338 797136 42394 797192
rect 42430 796728 42486 796784
rect 42430 794824 42486 794880
rect 41786 794144 41842 794200
rect 42246 792512 42302 792568
rect 42982 807472 43038 807528
rect 42154 789248 42210 789304
rect 41786 788568 41842 788624
rect 42246 788160 42302 788216
rect 41786 786800 41842 786856
rect 42706 788976 42762 789032
rect 42798 788568 42854 788624
rect 35806 773472 35862 773528
rect 35622 769392 35678 769448
rect 35438 768984 35494 769040
rect 35806 769004 35862 769040
rect 35806 768984 35808 769004
rect 35808 768984 35860 769004
rect 35860 768984 35862 769004
rect 31022 768168 31078 768224
rect 35806 767760 35862 767816
rect 35806 767372 35862 767408
rect 35806 767352 35808 767372
rect 35808 767352 35860 767372
rect 35860 767352 35862 767372
rect 35162 766944 35218 767000
rect 37094 763292 37150 763328
rect 37094 763272 37096 763292
rect 37096 763272 37148 763292
rect 37148 763272 37150 763292
rect 41326 765720 41382 765776
rect 40038 764496 40094 764552
rect 39302 759056 39358 759112
rect 36542 757696 36598 757752
rect 40590 758276 40592 758296
rect 40592 758276 40644 758296
rect 40644 758276 40646 758296
rect 40590 758240 40646 758276
rect 42246 765720 42302 765776
rect 42338 759056 42394 759112
rect 42062 758648 42118 758704
rect 42522 758240 42578 758296
rect 40314 757288 40370 757344
rect 40866 757288 40922 757344
rect 41786 756608 41842 756664
rect 42338 754840 42394 754896
rect 42062 754024 42118 754080
rect 42338 753616 42394 753672
rect 42062 752936 42118 752992
rect 41970 751032 42026 751088
rect 41786 750352 41842 750408
rect 41786 747360 41842 747416
rect 42154 746680 42210 746736
rect 42798 754568 42854 754624
rect 42154 746000 42210 746056
rect 42706 746000 42762 746056
rect 42246 745320 42302 745376
rect 41786 743688 41842 743744
rect 42614 744368 42670 744424
rect 42614 743008 42670 743064
rect 42430 741648 42486 741704
rect 35622 731312 35678 731368
rect 35806 730904 35862 730960
rect 41326 726416 41382 726472
rect 41142 726008 41198 726064
rect 31022 725192 31078 725248
rect 36542 724784 36598 724840
rect 33046 723968 33102 724024
rect 33782 723152 33838 723208
rect 40682 724376 40738 724432
rect 40038 720296 40094 720352
rect 39854 715128 39910 715184
rect 40222 715556 40278 715592
rect 40222 715536 40224 715556
rect 40224 715536 40276 715556
rect 40276 715536 40278 715556
rect 41326 725600 41382 725656
rect 41142 721712 41198 721768
rect 41878 722336 41934 722392
rect 41694 719208 41750 719264
rect 41878 718528 41934 718584
rect 42522 719208 42578 719264
rect 42154 718256 42210 718312
rect 40682 714720 40738 714776
rect 40038 714448 40094 714504
rect 42338 715128 42394 715184
rect 42062 714720 42118 714776
rect 42062 714448 42118 714504
rect 41510 714176 41566 714232
rect 41970 713360 42026 713416
rect 42154 711592 42210 711648
rect 42154 710776 42210 710832
rect 42246 709144 42302 709200
rect 42154 708464 42210 708520
rect 42062 707648 42118 707704
rect 41786 707376 41842 707432
rect 42062 706560 42118 706616
rect 42246 705200 42302 705256
rect 42246 703976 42302 704032
rect 42246 703568 42302 703624
rect 42062 703024 42118 703080
rect 42706 715536 42762 715592
rect 42798 703024 42854 703080
rect 42614 702072 42670 702128
rect 42246 701800 42302 701856
rect 42430 701528 42486 701584
rect 41694 697856 41750 697912
rect 35622 691328 35678 691384
rect 35806 687656 35862 687712
rect 35622 687248 35678 687304
rect 35806 683188 35862 683224
rect 35806 683168 35808 683188
rect 35808 683168 35860 683188
rect 35860 683168 35862 683188
rect 35438 682760 35494 682816
rect 35622 682352 35678 682408
rect 35806 681944 35862 682000
rect 35622 681536 35678 681592
rect 35162 680720 35218 680776
rect 35806 681128 35862 681184
rect 41786 680992 41842 681048
rect 42798 679904 42854 679960
rect 39946 677048 40002 677104
rect 39946 672424 40002 672480
rect 38934 672152 38990 672208
rect 42614 674192 42670 674248
rect 42246 672424 42302 672480
rect 42430 672424 42486 672480
rect 39578 671200 39634 671256
rect 41510 671200 41566 671256
rect 37922 670928 37978 670984
rect 41786 670248 41842 670304
rect 41970 668480 42026 668536
rect 41878 667664 41934 667720
rect 42522 672152 42578 672208
rect 42798 672152 42854 672208
rect 42154 665352 42210 665408
rect 42154 664808 42210 664864
rect 41786 664128 41842 664184
rect 42246 663992 42302 664048
rect 42062 662768 42118 662824
rect 42062 661000 42118 661056
rect 42798 667256 42854 667312
rect 42798 663992 42854 664048
rect 42706 663720 42762 663776
rect 42706 661000 42762 661056
rect 42706 660728 42762 660784
rect 42430 658552 42486 658608
rect 42246 658280 42302 658336
rect 42062 657328 42118 657384
rect 42614 657328 42670 657384
rect 35806 646720 35862 646776
rect 35806 644680 35862 644736
rect 41786 641620 41842 641676
rect 41786 641144 41842 641200
rect 35806 639784 35862 639840
rect 35806 638988 35862 639024
rect 35806 638968 35808 638988
rect 35808 638968 35860 638988
rect 35860 638968 35862 638988
rect 35806 638560 35862 638616
rect 32402 638152 32458 638208
rect 41970 638016 42026 638072
rect 40038 637336 40094 637392
rect 41970 637540 42026 637596
rect 42338 633800 42394 633856
rect 41418 627680 41474 627736
rect 42706 627272 42762 627328
rect 42430 624552 42486 624608
rect 42246 623736 42302 623792
rect 42062 623328 42118 623384
rect 42062 620880 42118 620936
rect 42246 620608 42302 620664
rect 41786 620200 41842 620256
rect 42430 620336 42486 620392
rect 42706 619928 42762 619984
rect 42430 618976 42486 619032
rect 42062 615848 42118 615904
rect 42430 615440 42486 615496
rect 42062 615168 42118 615224
rect 41878 614080 41934 614136
rect 43166 788160 43222 788216
rect 43166 766264 43222 766320
rect 43166 752936 43222 752992
rect 43166 723560 43222 723616
rect 43166 705200 43222 705256
rect 43166 679088 43222 679144
rect 43166 663720 43222 663776
rect 43166 636248 43222 636304
rect 43166 624552 43222 624608
rect 43534 932048 43590 932104
rect 44086 891948 44142 891984
rect 44086 891928 44088 891948
rect 44088 891928 44140 891948
rect 44140 891928 44142 891948
rect 44362 816040 44418 816096
rect 44178 814408 44234 814464
rect 43902 809512 43958 809568
rect 43718 806248 43774 806304
rect 43902 797680 43958 797736
rect 48962 940072 49018 940128
rect 51722 942248 51778 942304
rect 50342 939800 50398 939856
rect 47582 891928 47638 891984
rect 44638 815632 44694 815688
rect 44822 815224 44878 815280
rect 44546 810328 44602 810384
rect 44546 789248 44602 789304
rect 44362 773200 44418 773256
rect 44178 771976 44234 772032
rect 44638 772792 44694 772848
rect 44362 771568 44418 771624
rect 44362 771160 44418 771216
rect 44178 729272 44234 729328
rect 45006 813592 45062 813648
rect 44822 772384 44878 772440
rect 45190 807880 45246 807936
rect 45190 796728 45246 796784
rect 45006 770752 45062 770808
rect 45098 770344 45154 770400
rect 44822 766672 44878 766728
rect 44822 746680 44878 746736
rect 44638 730088 44694 730144
rect 44546 729680 44602 729736
rect 44362 728456 44418 728512
rect 44270 727232 44326 727288
rect 43902 721520 43958 721576
rect 43902 708464 43958 708520
rect 44914 728864 44970 728920
rect 44730 721112 44786 721168
rect 44546 686840 44602 686896
rect 44546 686432 44602 686488
rect 44270 684392 44326 684448
rect 44362 683984 44418 684040
rect 44178 680312 44234 680368
rect 44178 662768 44234 662824
rect 45282 764768 45338 764824
rect 45558 764224 45614 764280
rect 45282 753616 45338 753672
rect 45282 728048 45338 728104
rect 45098 727640 45154 727696
rect 45098 722744 45154 722800
rect 45098 707648 45154 707704
rect 44914 686024 44970 686080
rect 45098 685616 45154 685672
rect 44914 684800 44970 684856
rect 45282 685208 45338 685264
rect 45190 679496 45246 679552
rect 45190 664808 45246 664864
rect 44730 653112 44786 653168
rect 44546 643320 44602 643376
rect 44362 641416 44418 641472
rect 44178 636520 44234 636576
rect 43902 635296 43958 635352
rect 43902 620880 43958 620936
rect 44730 642504 44786 642560
rect 44270 623328 44326 623384
rect 44086 620608 44142 620664
rect 45374 643592 45430 643648
rect 45098 643048 45154 643104
rect 44914 642232 44970 642288
rect 45282 641144 45338 641200
rect 44914 640872 44970 640928
rect 44914 635704 44970 635760
rect 44178 614080 44234 614136
rect 42982 612312 43038 612368
rect 43580 612332 43636 612368
rect 43580 612312 43582 612332
rect 43582 612312 43634 612332
rect 43634 612312 43636 612332
rect 42706 610952 42762 611008
rect 44270 610952 44326 611008
rect 44546 600480 44602 600536
rect 44638 600072 44694 600128
rect 40314 597216 40370 597272
rect 42982 596944 43038 597000
rect 42614 596808 42670 596864
rect 40866 596162 40922 596218
rect 41142 596162 41198 596218
rect 32402 595584 32458 595640
rect 36542 595176 36598 595232
rect 35162 594360 35218 594416
rect 37922 594768 37978 594824
rect 41786 595992 41842 596048
rect 41694 594904 41750 594960
rect 39946 590688 40002 590744
rect 39946 585928 40002 585984
rect 37922 585112 37978 585168
rect 40498 585656 40554 585712
rect 39486 584840 39542 584896
rect 40958 589600 41014 589656
rect 41786 593544 41842 593600
rect 42798 593952 42854 594008
rect 41786 593136 41842 593192
rect 41786 592728 41842 592784
rect 41786 589328 41842 589384
rect 42706 586064 42762 586120
rect 42246 585928 42302 585984
rect 41418 585384 41474 585440
rect 42614 585656 42670 585712
rect 42430 585384 42486 585440
rect 40682 584568 40738 584624
rect 42338 581848 42394 581904
rect 42246 581440 42302 581496
rect 42062 581168 42118 581224
rect 42246 580760 42302 580816
rect 41786 580216 41842 580272
rect 41786 578176 41842 578232
rect 41786 577496 41842 577552
rect 42246 576816 42302 576872
rect 42522 576136 42578 576192
rect 42062 573280 42118 573336
rect 42706 573280 42762 573336
rect 41970 572600 42026 572656
rect 42246 572192 42302 572248
rect 42062 570968 42118 571024
rect 42614 571920 42670 571976
rect 42338 569200 42394 569256
rect 35806 558048 35862 558104
rect 42062 558456 42118 558512
rect 42062 557504 42118 557560
rect 44454 591912 44510 591968
rect 43442 590280 43498 590336
rect 35806 554804 35862 554840
rect 35806 554784 35808 554804
rect 35808 554784 35860 554804
rect 35860 554784 35862 554804
rect 35622 553968 35678 554024
rect 35806 553580 35862 553616
rect 35806 553560 35808 553580
rect 35808 553560 35860 553580
rect 35860 553560 35862 553580
rect 40866 553152 40922 553208
rect 33782 551928 33838 551984
rect 31758 547460 31814 547496
rect 31758 547440 31760 547460
rect 31760 547440 31812 547460
rect 31812 547440 31814 547460
rect 41050 552744 41106 552800
rect 41234 551112 41290 551168
rect 41326 548256 41382 548312
rect 41326 546352 41382 546408
rect 41786 553152 41842 553208
rect 42982 552336 43038 552392
rect 41878 551928 41934 551984
rect 42062 550296 42118 550352
rect 41694 547712 41750 547768
rect 42062 545672 42118 545728
rect 41786 541048 41842 541104
rect 41786 540640 41842 540696
rect 42614 540232 42670 540288
rect 42338 538600 42394 538656
rect 42246 538192 42302 538248
rect 42062 537920 42118 537976
rect 42614 537920 42670 537976
rect 42246 536288 42302 536344
rect 42614 537104 42670 537160
rect 42154 533840 42210 533896
rect 42246 533160 42302 533216
rect 42522 532752 42578 532808
rect 43166 549480 43222 549536
rect 42982 533840 43038 533896
rect 43166 533160 43222 533216
rect 42154 530032 42210 530088
rect 41878 529352 41934 529408
rect 42522 530576 42578 530632
rect 42706 530032 42762 530088
rect 42614 529624 42670 529680
rect 42890 529080 42946 529136
rect 41326 425992 41382 426048
rect 40958 425584 41014 425640
rect 36542 424360 36598 424416
rect 41326 423952 41382 424008
rect 41142 418784 41198 418840
rect 41878 422728 41934 422784
rect 41510 418512 41566 418568
rect 42062 421912 42118 421968
rect 41878 417832 41934 417888
rect 42430 419872 42486 419928
rect 42246 418512 42302 418568
rect 42062 417560 42118 417616
rect 42062 411848 42118 411904
rect 42522 411848 42578 411904
rect 41786 409400 41842 409456
rect 42430 408448 42486 408504
rect 42430 407768 42486 407824
rect 42430 406952 42486 407008
rect 41786 406272 41842 406328
rect 42614 405592 42670 405648
rect 41786 403824 41842 403880
rect 42338 402872 42394 402928
rect 41786 401784 41842 401840
rect 42430 400152 42486 400208
rect 42430 399744 42486 399800
rect 43074 423136 43130 423192
rect 43258 421096 43314 421152
rect 43258 407768 43314 407824
rect 43074 402872 43130 402928
rect 41786 398792 41842 398848
rect 41142 387116 41198 387152
rect 41142 387096 41144 387116
rect 41144 387096 41196 387116
rect 41196 387096 41198 387116
rect 41878 386960 41934 387016
rect 41326 386688 41382 386744
rect 41510 386688 41566 386744
rect 41326 382608 41382 382664
rect 40038 382200 40094 382256
rect 37922 381384 37978 381440
rect 33782 380160 33838 380216
rect 28538 376488 28594 376544
rect 28538 373224 28594 373280
rect 35806 379344 35862 379400
rect 35806 376080 35862 376136
rect 40222 380976 40278 381032
rect 40038 376896 40094 376952
rect 41694 375420 41750 375456
rect 41694 375400 41696 375420
rect 41696 375400 41748 375420
rect 41748 375400 41750 375420
rect 41694 372580 41696 372600
rect 41696 372580 41748 372600
rect 41748 372580 41750 372600
rect 41694 372544 41750 372580
rect 33782 371864 33838 371920
rect 42614 372544 42670 372600
rect 41786 368464 41842 368520
rect 42430 366968 42486 367024
rect 42338 365744 42394 365800
rect 42154 364928 42210 364984
rect 44454 581032 44510 581088
rect 44822 599664 44878 599720
rect 44822 599256 44878 599312
rect 44638 557232 44694 557288
rect 45374 633392 45430 633448
rect 46386 763000 46442 763056
rect 46202 754024 46258 754080
rect 45742 676640 45798 676696
rect 46018 637744 46074 637800
rect 46202 636928 46258 636984
rect 46202 618976 46258 619032
rect 46018 615576 46074 615632
rect 46938 719888 46994 719944
rect 47766 817672 47822 817728
rect 50342 816856 50398 816912
rect 47582 710776 47638 710832
rect 47214 677864 47270 677920
rect 53286 892744 53342 892800
rect 97262 996104 97318 996160
rect 98274 1001972 98330 1002008
rect 98274 1001952 98276 1001972
rect 98276 1001952 98328 1001972
rect 98328 1001952 98330 1001972
rect 100298 1002380 100354 1002416
rect 100298 1002360 100300 1002380
rect 100300 1002360 100352 1002380
rect 100352 1002360 100354 1002380
rect 99102 1002108 99158 1002144
rect 99102 1002088 99104 1002108
rect 99104 1002088 99156 1002108
rect 99156 1002088 99158 1002108
rect 101126 1002244 101182 1002280
rect 101126 1002224 101128 1002244
rect 101128 1002224 101180 1002244
rect 101180 1002224 101182 1002244
rect 101126 1001972 101182 1002008
rect 101126 1001952 101128 1001972
rect 101128 1001952 101180 1001972
rect 101180 1001952 101182 1001972
rect 104806 1006188 104862 1006224
rect 104806 1006168 104808 1006188
rect 104808 1006168 104860 1006188
rect 104860 1006168 104862 1006188
rect 106830 1006188 106886 1006224
rect 106830 1006168 106832 1006188
rect 106832 1006168 106884 1006188
rect 106884 1006168 106886 1006188
rect 103150 1006052 103206 1006088
rect 103150 1006032 103152 1006052
rect 103152 1006032 103204 1006052
rect 103204 1006032 103206 1006052
rect 106002 1006052 106058 1006088
rect 106002 1006032 106004 1006052
rect 106004 1006032 106056 1006052
rect 106056 1006032 106058 1006052
rect 108854 1005252 108856 1005272
rect 108856 1005252 108908 1005272
rect 108908 1005252 108910 1005272
rect 101954 1002516 102010 1002552
rect 101954 1002496 101956 1002516
rect 101956 1002496 102008 1002516
rect 102008 1002496 102010 1002516
rect 102322 1002108 102378 1002144
rect 102322 1002088 102324 1002108
rect 102324 1002088 102376 1002108
rect 102376 1002088 102378 1002108
rect 101402 995016 101458 995072
rect 108854 1005216 108910 1005252
rect 108486 1004692 108542 1004728
rect 108486 1004672 108488 1004692
rect 108488 1004672 108540 1004692
rect 108540 1004672 108542 1004692
rect 103150 1002380 103206 1002416
rect 103150 1002360 103152 1002380
rect 103152 1002360 103204 1002380
rect 103204 1002360 103206 1002380
rect 105634 1002244 105690 1002280
rect 105634 1002224 105636 1002244
rect 105636 1002224 105688 1002244
rect 105688 1002224 105690 1002244
rect 103978 1002108 104034 1002144
rect 103978 1002088 103980 1002108
rect 103980 1002088 104032 1002108
rect 104032 1002088 104034 1002108
rect 104806 1001952 104862 1002008
rect 106002 1001972 106058 1002008
rect 106002 1001952 106004 1001972
rect 106004 1001952 106056 1001972
rect 106056 1001952 106058 1001972
rect 104162 994744 104218 994800
rect 107658 1002380 107714 1002416
rect 107658 1002360 107660 1002380
rect 107660 1002360 107712 1002380
rect 107712 1002360 107714 1002380
rect 108026 1002244 108082 1002280
rect 108026 1002224 108028 1002244
rect 108028 1002224 108080 1002244
rect 108080 1002224 108082 1002244
rect 106830 1002108 106886 1002144
rect 106830 1002088 106832 1002108
rect 106832 1002088 106884 1002108
rect 106884 1002088 106886 1002108
rect 109682 1002108 109738 1002144
rect 109682 1002088 109684 1002108
rect 109684 1002088 109736 1002108
rect 109736 1002088 109738 1002108
rect 117226 997192 117282 997248
rect 116950 996920 117006 996976
rect 143814 997192 143870 997248
rect 126242 996240 126298 996296
rect 131854 995696 131910 995752
rect 132958 995696 133014 995752
rect 136730 995696 136786 995752
rect 137374 995696 137430 995752
rect 140410 995696 140466 995752
rect 144366 996376 144422 996432
rect 144182 996104 144238 996160
rect 141790 995560 141846 995616
rect 124862 995016 124918 995072
rect 132406 995288 132462 995344
rect 132130 994744 132186 994800
rect 135902 994744 135958 994800
rect 133142 994472 133198 994528
rect 141882 994744 141938 994800
rect 142066 994744 142122 994800
rect 144826 996920 144882 996976
rect 143722 994200 143778 994256
rect 143906 994200 143962 994256
rect 139214 993928 139270 993984
rect 139398 993928 139454 993984
rect 137742 993656 137798 993712
rect 153750 1006596 153806 1006632
rect 153750 1006576 153752 1006596
rect 153752 1006576 153804 1006596
rect 153804 1006576 153806 1006596
rect 157430 1006596 157486 1006632
rect 157430 1006576 157432 1006596
rect 157432 1006576 157484 1006596
rect 157484 1006576 157486 1006596
rect 152922 1006460 152978 1006496
rect 152922 1006440 152924 1006460
rect 152924 1006440 152976 1006460
rect 152976 1006440 152978 1006460
rect 160282 1006460 160338 1006496
rect 160282 1006440 160284 1006460
rect 160284 1006440 160336 1006460
rect 160336 1006440 160338 1006460
rect 152094 1006324 152150 1006360
rect 152094 1006304 152096 1006324
rect 152096 1006304 152148 1006324
rect 152148 1006304 152150 1006324
rect 158258 1006324 158314 1006360
rect 158258 1006304 158260 1006324
rect 158260 1006304 158312 1006324
rect 158312 1006304 158314 1006324
rect 151266 1006204 151268 1006224
rect 151268 1006204 151320 1006224
rect 151320 1006204 151322 1006224
rect 151266 1006168 151322 1006204
rect 158626 1006188 158682 1006224
rect 158626 1006168 158628 1006188
rect 158628 1006168 158680 1006188
rect 158680 1006168 158682 1006188
rect 147126 1006032 147182 1006088
rect 148874 1006068 148876 1006088
rect 148876 1006068 148928 1006088
rect 148928 1006068 148930 1006088
rect 148874 1006032 148930 1006068
rect 150070 1006068 150072 1006088
rect 150072 1006068 150124 1006088
rect 150124 1006068 150126 1006088
rect 150070 1006032 150126 1006068
rect 145562 993928 145618 993984
rect 142158 993692 142160 993712
rect 142160 993692 142212 993712
rect 142212 993692 142214 993712
rect 142158 993656 142214 993692
rect 142342 993656 142398 993712
rect 158258 1006052 158314 1006088
rect 158258 1006032 158260 1006052
rect 158260 1006032 158312 1006052
rect 158312 1006032 158314 1006052
rect 159454 1006052 159510 1006088
rect 159454 1006032 159456 1006052
rect 159456 1006032 159508 1006052
rect 159508 1006032 159510 1006052
rect 153750 1005100 153806 1005136
rect 153750 1005080 153752 1005100
rect 153752 1005080 153804 1005100
rect 153804 1005080 153806 1005100
rect 147126 995560 147182 995616
rect 149242 1001972 149298 1002008
rect 149242 1001952 149244 1001972
rect 149244 1001952 149296 1001972
rect 149296 1001952 149298 1001972
rect 150898 1002380 150954 1002416
rect 150898 1002360 150900 1002380
rect 150900 1002360 150952 1002380
rect 150952 1002360 150954 1002380
rect 150898 1002108 150954 1002144
rect 150898 1002088 150900 1002108
rect 150900 1002088 150952 1002108
rect 150952 1002088 150954 1002108
rect 152922 1004964 152978 1005000
rect 152922 1004944 152924 1004964
rect 152924 1004944 152976 1004964
rect 152976 1004944 152978 1004964
rect 151726 1004692 151782 1004728
rect 151726 1004672 151728 1004692
rect 151728 1004672 151780 1004692
rect 151780 1004672 151782 1004692
rect 149702 994472 149758 994528
rect 148506 994200 148562 994256
rect 154118 1004828 154174 1004864
rect 154118 1004808 154120 1004828
rect 154120 1004808 154172 1004828
rect 154172 1004808 154174 1004828
rect 160650 1004828 160706 1004864
rect 160650 1004808 160652 1004828
rect 160652 1004808 160704 1004828
rect 160704 1004808 160706 1004828
rect 161110 1004692 161166 1004728
rect 161110 1004672 161112 1004692
rect 161112 1004672 161164 1004692
rect 161164 1004672 161166 1004692
rect 155774 1002244 155830 1002280
rect 155774 1002224 155776 1002244
rect 155776 1002224 155828 1002244
rect 155828 1002224 155830 1002244
rect 154578 1002108 154634 1002144
rect 154578 1002088 154580 1002108
rect 154580 1002088 154632 1002108
rect 154632 1002088 154634 1002108
rect 154302 995696 154358 995752
rect 154302 995016 154358 995072
rect 154946 1001952 155002 1002008
rect 155774 1001952 155830 1002008
rect 156602 1001972 156658 1002008
rect 156602 1001952 156604 1001972
rect 156604 1001952 156656 1001972
rect 156656 1001952 156658 1001972
rect 157798 1002108 157854 1002144
rect 157798 1002088 157800 1002108
rect 157800 1002088 157852 1002108
rect 157852 1002088 157854 1002108
rect 154578 994472 154634 994528
rect 152462 993656 152518 993712
rect 170862 995288 170918 995344
rect 171690 995329 171746 995344
rect 171690 995288 171692 995329
rect 171692 995288 171744 995329
rect 171744 995288 171746 995329
rect 256146 1006460 256202 1006496
rect 256146 1006440 256148 1006460
rect 256148 1006440 256200 1006460
rect 256200 1006440 256202 1006460
rect 354862 1006460 354918 1006496
rect 354862 1006440 354864 1006460
rect 354864 1006440 354916 1006460
rect 354916 1006440 354918 1006460
rect 210422 1006188 210478 1006224
rect 210422 1006168 210424 1006188
rect 210424 1006168 210476 1006188
rect 210476 1006168 210478 1006188
rect 201038 1006052 201094 1006088
rect 201038 1006032 201040 1006052
rect 201040 1006032 201092 1006052
rect 201092 1006032 201094 1006052
rect 208398 1006052 208454 1006088
rect 208398 1006032 208400 1006052
rect 208400 1006032 208452 1006052
rect 208452 1006032 208454 1006052
rect 175922 995832 175978 995888
rect 212078 1005252 212080 1005272
rect 212080 1005252 212132 1005272
rect 212132 1005252 212134 1005272
rect 195058 995832 195114 995888
rect 192482 995730 192538 995786
rect 177302 995560 177358 995616
rect 173162 995016 173218 995072
rect 183834 995288 183890 995344
rect 187606 994744 187662 994800
rect 184846 994200 184902 994256
rect 188802 994472 188858 994528
rect 190366 994472 190422 994528
rect 189446 993928 189502 993984
rect 195058 995288 195114 995344
rect 195242 994744 195298 994800
rect 196070 997736 196126 997792
rect 193126 993656 193182 993712
rect 195334 993656 195390 993712
rect 196070 994472 196126 994528
rect 196622 994200 196678 994256
rect 200210 997736 200266 997792
rect 200210 997228 200212 997248
rect 200212 997228 200264 997248
rect 200264 997228 200266 997248
rect 200210 997192 200266 997228
rect 201866 997908 201868 997928
rect 201868 997908 201920 997928
rect 201920 997908 201922 997928
rect 201866 997872 201922 997908
rect 200210 996648 200266 996704
rect 200670 996260 200726 996296
rect 200670 996240 200672 996260
rect 200672 996240 200724 996260
rect 200724 996240 200726 996260
rect 202694 1001136 202750 1001192
rect 203890 998844 203946 998880
rect 203890 998824 203892 998844
rect 203892 998824 203944 998844
rect 203944 998824 203946 998844
rect 203522 998572 203578 998608
rect 203522 998552 203524 998572
rect 203524 998552 203576 998572
rect 203576 998552 203578 998572
rect 204350 998708 204406 998744
rect 204350 998688 204352 998708
rect 204352 998688 204404 998708
rect 204404 998688 204406 998708
rect 203522 998180 203524 998200
rect 203524 998180 203576 998200
rect 203576 998180 203578 998200
rect 203522 998144 203578 998180
rect 202694 998044 202696 998064
rect 202696 998044 202748 998064
rect 202748 998044 202750 998064
rect 202694 998008 202750 998044
rect 204718 997772 204720 997792
rect 204720 997772 204772 997792
rect 204772 997772 204774 997792
rect 204718 997736 204774 997772
rect 202326 995832 202382 995888
rect 203614 995832 203670 995888
rect 203614 995288 203670 995344
rect 199382 993928 199438 993984
rect 186502 992840 186558 992896
rect 212078 1005216 212134 1005252
rect 209226 1004964 209282 1005000
rect 209226 1004944 209228 1004964
rect 209228 1004944 209280 1004964
rect 209280 1004944 209282 1004964
rect 211250 1004828 211306 1004864
rect 211250 1004808 211252 1004828
rect 211252 1004808 211304 1004828
rect 211304 1004808 211306 1004828
rect 209226 1004692 209282 1004728
rect 209226 1004672 209228 1004692
rect 209228 1004672 209280 1004692
rect 209280 1004672 209282 1004692
rect 206374 1002516 206430 1002552
rect 206374 1002496 206376 1002516
rect 206376 1002496 206428 1002516
rect 206428 1002496 206430 1002516
rect 207202 1002244 207258 1002280
rect 207202 1002224 207204 1002244
rect 207204 1002224 207256 1002244
rect 207256 1002224 207258 1002244
rect 206742 1002108 206798 1002144
rect 206742 1002088 206744 1002108
rect 206744 1002088 206796 1002108
rect 206796 1002088 206798 1002108
rect 210882 1002108 210938 1002144
rect 210882 1002088 210884 1002108
rect 210884 1002088 210936 1002108
rect 210936 1002088 210938 1002108
rect 205546 1001972 205602 1002008
rect 205546 1001952 205548 1001972
rect 205548 1001952 205600 1001972
rect 205600 1001952 205602 1001972
rect 205546 997908 205548 997928
rect 205548 997908 205600 997928
rect 205600 997908 205602 997928
rect 205546 997872 205602 997908
rect 207202 1001952 207258 1002008
rect 207570 1001972 207626 1002008
rect 207570 1001952 207572 1001972
rect 207572 1001952 207624 1001972
rect 207624 1001952 207626 1001972
rect 208398 995832 208454 995888
rect 212538 1001972 212594 1002008
rect 212538 1001952 212540 1001972
rect 212540 1001952 212592 1001972
rect 212592 1001952 212594 1001972
rect 208398 995016 208454 995072
rect 246578 998008 246634 998064
rect 246670 996376 246726 996432
rect 246670 995968 246726 996024
rect 247130 996648 247186 996704
rect 238574 995696 238630 995752
rect 239586 995696 239642 995752
rect 240230 995696 240286 995752
rect 240874 995696 240930 995752
rect 243818 995696 243874 995752
rect 244094 995696 244150 995752
rect 245566 995696 245622 995752
rect 246946 995696 247002 995752
rect 247130 995696 247186 995752
rect 228362 995016 228418 995072
rect 235262 994472 235318 994528
rect 242070 995288 242126 995344
rect 245014 995288 245070 995344
rect 243266 994744 243322 994800
rect 247314 994744 247370 994800
rect 258998 1006324 259054 1006360
rect 258998 1006304 259000 1006324
rect 259000 1006304 259052 1006324
rect 259052 1006304 259054 1006324
rect 307758 1006324 307814 1006360
rect 307758 1006304 307760 1006324
rect 307760 1006304 307812 1006324
rect 307812 1006304 307814 1006324
rect 314658 1006324 314714 1006360
rect 314658 1006304 314660 1006324
rect 314660 1006304 314712 1006324
rect 314712 1006304 314714 1006324
rect 361394 1006324 361450 1006360
rect 361394 1006304 361396 1006324
rect 361396 1006304 361448 1006324
rect 361448 1006304 361450 1006324
rect 235906 994200 235962 994256
rect 247682 994200 247738 994256
rect 252466 1006032 252522 1006088
rect 249062 997192 249118 997248
rect 251178 995424 251234 995480
rect 255318 1003892 255320 1003912
rect 255320 1003892 255372 1003912
rect 255372 1003892 255374 1003912
rect 255318 1003856 255374 1003892
rect 252466 997772 252468 997792
rect 252468 997772 252520 997792
rect 252520 997772 252522 997792
rect 252466 997736 252522 997772
rect 254122 1002532 254124 1002552
rect 254124 1002532 254176 1002552
rect 254176 1002532 254178 1002552
rect 254122 1002496 254178 1002532
rect 254490 1002380 254546 1002416
rect 254490 1002360 254492 1002380
rect 254492 1002360 254544 1002380
rect 254544 1002360 254546 1002380
rect 253662 998164 253718 998200
rect 253662 998144 253664 998164
rect 253664 998144 253716 998164
rect 253716 998144 253718 998164
rect 253662 997908 253664 997928
rect 253664 997908 253716 997928
rect 253716 997908 253718 997928
rect 253662 997872 253718 997908
rect 253386 995696 253442 995752
rect 253110 994472 253166 994528
rect 255318 1002108 255374 1002144
rect 255318 1002088 255320 1002108
rect 255320 1002088 255372 1002108
rect 255372 1002088 255374 1002108
rect 257342 1006188 257398 1006224
rect 257342 1006168 257344 1006188
rect 257344 1006168 257396 1006188
rect 257396 1006168 257398 1006188
rect 262678 1006188 262734 1006224
rect 262678 1006168 262680 1006188
rect 262680 1006168 262732 1006188
rect 262732 1006168 262734 1006188
rect 258170 1006052 258226 1006088
rect 258170 1006032 258172 1006052
rect 258172 1006032 258224 1006052
rect 258224 1006032 258226 1006052
rect 261850 1006052 261906 1006088
rect 261850 1006032 261852 1006052
rect 261852 1006032 261904 1006052
rect 261904 1006032 261906 1006052
rect 256146 1002668 256148 1002688
rect 256148 1002668 256200 1002688
rect 256200 1002668 256202 1002688
rect 256146 1002632 256202 1002668
rect 256514 1002244 256570 1002280
rect 256514 1002224 256516 1002244
rect 256516 1002224 256568 1002244
rect 256568 1002224 256570 1002244
rect 256974 1001972 257030 1002008
rect 256974 1001952 256976 1001972
rect 256976 1001952 257028 1001972
rect 257028 1001952 257030 1001972
rect 263046 1004964 263102 1005000
rect 263046 1004944 263048 1004964
rect 263048 1004944 263100 1004964
rect 263100 1004944 263102 1004964
rect 258170 1004828 258226 1004864
rect 258170 1004808 258172 1004828
rect 258172 1004808 258224 1004828
rect 258224 1004808 258226 1004828
rect 258998 1001952 259054 1002008
rect 261022 1002380 261078 1002416
rect 261022 1002360 261024 1002380
rect 261024 1002360 261076 1002380
rect 261076 1002360 261078 1002380
rect 260194 1002244 260250 1002280
rect 260194 1002224 260196 1002244
rect 260196 1002224 260248 1002244
rect 260248 1002224 260250 1002244
rect 259826 1002108 259882 1002144
rect 259826 1002088 259828 1002108
rect 259828 1002088 259880 1002108
rect 259880 1002088 259882 1002108
rect 260194 1001972 260250 1002008
rect 260194 1001952 260196 1001972
rect 260196 1001952 260248 1001972
rect 260248 1001952 260250 1001972
rect 261850 1001952 261906 1002008
rect 263874 1002108 263930 1002144
rect 263874 1002088 263876 1002108
rect 263876 1002088 263928 1002108
rect 263928 1002088 263930 1002108
rect 263506 1001972 263562 1002008
rect 263506 1001952 263508 1001972
rect 263508 1001952 263560 1001972
rect 263560 1001952 263562 1001972
rect 270406 995016 270462 995072
rect 298282 1002224 298338 1002280
rect 298098 997736 298154 997792
rect 282734 995696 282790 995752
rect 288070 995696 288126 995752
rect 291106 995696 291162 995752
rect 279422 995288 279478 995344
rect 290738 994744 290794 994800
rect 286506 994472 286562 994528
rect 298834 996648 298890 996704
rect 298650 996396 298706 996432
rect 298650 996376 298652 996396
rect 298652 996376 298704 996396
rect 298704 996376 298706 996396
rect 294786 994744 294842 994800
rect 295246 994744 295302 994800
rect 292118 994200 292174 994256
rect 299478 997192 299534 997248
rect 299294 996920 299350 996976
rect 304906 1006188 304962 1006224
rect 304906 1006168 304908 1006188
rect 304908 1006168 304960 1006188
rect 304960 1006168 304962 1006188
rect 301686 1006032 301742 1006088
rect 303250 1006052 303306 1006088
rect 303250 1006032 303252 1006052
rect 303252 1006032 303304 1006052
rect 303304 1006032 303306 1006052
rect 304078 1006052 304134 1006088
rect 304078 1006032 304080 1006052
rect 304080 1006032 304132 1006052
rect 304132 1006032 304134 1006052
rect 311806 1006052 311862 1006088
rect 311806 1006032 311808 1006052
rect 311808 1006032 311860 1006052
rect 311860 1006032 311862 1006052
rect 314658 1006052 314714 1006088
rect 314658 1006032 314660 1006052
rect 314660 1006032 314712 1006052
rect 314712 1006032 314714 1006052
rect 307298 1005236 307354 1005272
rect 307298 1005216 307300 1005236
rect 307300 1005216 307352 1005236
rect 307352 1005216 307354 1005236
rect 303250 1002224 303306 1002280
rect 301686 997736 301742 997792
rect 302882 996104 302938 996160
rect 304078 1002108 304134 1002144
rect 304078 1002088 304080 1002108
rect 304080 1002088 304132 1002108
rect 304132 1002088 304134 1002108
rect 303066 995832 303122 995888
rect 306930 1004964 306986 1005000
rect 306930 1004944 306932 1004964
rect 306932 1004944 306984 1004964
rect 306984 1004944 306986 1004964
rect 308954 1004828 309010 1004864
rect 308954 1004808 308956 1004828
rect 308956 1004808 309008 1004828
rect 309008 1004808 309010 1004828
rect 313830 1004828 313886 1004864
rect 313830 1004808 313832 1004828
rect 313832 1004808 313884 1004828
rect 313884 1004808 313886 1004828
rect 305274 1003332 305330 1003368
rect 305274 1003312 305276 1003332
rect 305276 1003312 305328 1003332
rect 305328 1003312 305330 1003332
rect 308126 1004692 308182 1004728
rect 308126 1004672 308128 1004692
rect 308128 1004672 308180 1004692
rect 308180 1004672 308182 1004692
rect 315486 1004692 315542 1004728
rect 315486 1004672 315488 1004692
rect 315488 1004672 315540 1004692
rect 315540 1004672 315542 1004692
rect 308954 1003196 309010 1003232
rect 308954 1003176 308956 1003196
rect 308956 1003176 309008 1003196
rect 309008 1003176 309010 1003196
rect 310610 1002496 310666 1002552
rect 306102 1002244 306158 1002280
rect 306102 1002224 306104 1002244
rect 306104 1002224 306156 1002244
rect 306156 1002224 306158 1002244
rect 306102 1001972 306158 1002008
rect 306102 1001952 306104 1001972
rect 306104 1001952 306156 1001972
rect 306156 1001952 306158 1001972
rect 301502 994472 301558 994528
rect 306930 1001952 306986 1002008
rect 308770 995560 308826 995616
rect 309782 1001952 309838 1002008
rect 310150 1001972 310206 1002008
rect 310150 1001952 310152 1001972
rect 310152 1001952 310204 1001972
rect 310204 1001952 310206 1001972
rect 310610 1002244 310666 1002280
rect 310610 1002224 310612 1002244
rect 310612 1002224 310664 1002244
rect 310664 1002224 310666 1002244
rect 308770 995016 308826 995072
rect 300306 994200 300362 994256
rect 306378 994200 306434 994256
rect 291750 993928 291806 993984
rect 360566 1006188 360622 1006224
rect 360566 1006168 360568 1006188
rect 360568 1006168 360620 1006188
rect 360620 1006168 360622 1006188
rect 363418 1006188 363474 1006224
rect 363418 1006168 363420 1006188
rect 363420 1006168 363472 1006188
rect 363472 1006168 363474 1006188
rect 358542 1006052 358598 1006088
rect 358542 1006032 358544 1006052
rect 358544 1006032 358596 1006052
rect 358596 1006032 358598 1006052
rect 360566 1005388 360568 1005408
rect 360568 1005388 360620 1005408
rect 360620 1005388 360622 1005408
rect 360566 1005352 360622 1005388
rect 355690 1005252 355692 1005272
rect 355692 1005252 355744 1005272
rect 355744 1005252 355746 1005272
rect 355690 1005216 355746 1005252
rect 356518 1004964 356574 1005000
rect 356518 1004944 356520 1004964
rect 356520 1004944 356572 1004964
rect 356572 1004944 356574 1004964
rect 361394 1004964 361450 1005000
rect 361394 1004944 361396 1004964
rect 361396 1004944 361448 1004964
rect 361448 1004944 361450 1004964
rect 354034 1001972 354090 1002008
rect 354034 1001952 354036 1001972
rect 354036 1001952 354088 1001972
rect 354088 1001952 354090 1001972
rect 355690 1004828 355746 1004864
rect 355690 1004808 355692 1004828
rect 355692 1004808 355744 1004828
rect 355744 1004808 355746 1004828
rect 357714 1002380 357770 1002416
rect 357714 1002360 357716 1002380
rect 357716 1002360 357768 1002380
rect 357768 1002360 357770 1002380
rect 357714 1002108 357770 1002144
rect 357714 1002088 357716 1002108
rect 357716 1002088 357768 1002108
rect 357768 1002088 357770 1002108
rect 356518 1001952 356574 1002008
rect 357346 1001952 357402 1002008
rect 359370 1001952 359426 1002008
rect 362590 1004828 362646 1004864
rect 362590 1004808 362592 1004828
rect 362592 1004808 362644 1004828
rect 362644 1004808 362646 1004828
rect 365074 1006052 365130 1006088
rect 365074 1006032 365076 1006052
rect 365076 1006032 365128 1006052
rect 365128 1006032 365130 1006052
rect 365074 1005100 365130 1005136
rect 365074 1005080 365076 1005100
rect 365076 1005080 365128 1005100
rect 365128 1005080 365130 1005100
rect 364246 1004692 364302 1004728
rect 364246 1004672 364248 1004692
rect 364248 1004672 364300 1004692
rect 364300 1004672 364302 1004692
rect 365902 1001972 365958 1002008
rect 365902 1001952 365904 1001972
rect 365904 1001952 365956 1001972
rect 365956 1001952 365958 1001972
rect 372526 996920 372582 996976
rect 372342 996376 372398 996432
rect 372342 995968 372398 996024
rect 374642 997736 374698 997792
rect 429198 1006748 429200 1006768
rect 429200 1006748 429252 1006768
rect 429252 1006748 429254 1006768
rect 429198 1006712 429254 1006748
rect 431682 1006612 431684 1006632
rect 431684 1006612 431736 1006632
rect 431736 1006612 431738 1006632
rect 431682 1006576 431738 1006612
rect 428370 1006476 428372 1006496
rect 428372 1006476 428424 1006496
rect 428424 1006476 428426 1006496
rect 428370 1006440 428426 1006476
rect 427542 1006324 427598 1006360
rect 427542 1006304 427544 1006324
rect 427544 1006304 427596 1006324
rect 427596 1006304 427598 1006324
rect 380898 995832 380954 995888
rect 382186 995832 382242 995888
rect 382646 995696 382702 995752
rect 382462 995288 382518 995344
rect 382830 995016 382886 995072
rect 383106 994744 383162 994800
rect 399942 996920 399998 996976
rect 400494 996648 400550 996704
rect 400034 996376 400090 996432
rect 385038 995696 385094 995752
rect 389362 995696 389418 995752
rect 389730 995696 389786 995752
rect 392214 995696 392270 995752
rect 396630 995696 396686 995752
rect 386326 995560 386382 995616
rect 388902 995288 388958 995344
rect 386510 994744 386566 994800
rect 387798 994744 387854 994800
rect 400034 995696 400090 995752
rect 429198 1006188 429254 1006224
rect 429198 1006168 429200 1006188
rect 429200 1006168 429252 1006188
rect 429252 1006168 429254 1006188
rect 421838 1006032 421894 1006088
rect 425150 1006052 425206 1006088
rect 425150 1006032 425152 1006052
rect 425152 1006032 425204 1006052
rect 425204 1006032 425206 1006052
rect 431682 1006052 431738 1006088
rect 431682 1006032 431684 1006052
rect 431684 1006032 431736 1006052
rect 431736 1006032 431738 1006052
rect 428370 1005796 428372 1005816
rect 428372 1005796 428424 1005816
rect 428424 1005796 428426 1005816
rect 428370 1005760 428426 1005796
rect 423494 1005660 423496 1005680
rect 423496 1005660 423548 1005680
rect 423548 1005660 423550 1005680
rect 423494 1005624 423550 1005660
rect 423494 1005388 423496 1005408
rect 423496 1005388 423548 1005408
rect 423548 1005388 423550 1005408
rect 423494 1005352 423550 1005388
rect 425518 1005100 425574 1005136
rect 425518 1005080 425520 1005100
rect 425520 1005080 425572 1005100
rect 425572 1005080 425574 1005100
rect 422666 1004828 422722 1004864
rect 422666 1004808 422668 1004828
rect 422668 1004808 422720 1004828
rect 422720 1004808 422722 1004828
rect 414478 996376 414534 996432
rect 400494 995424 400550 995480
rect 383474 994472 383530 994528
rect 392674 994472 392730 994528
rect 416134 995696 416190 995752
rect 415398 995444 415454 995480
rect 415398 995424 415400 995444
rect 415400 995424 415452 995444
rect 415452 995424 415454 995444
rect 424322 1003892 424324 1003912
rect 424324 1003892 424376 1003912
rect 424376 1003892 424378 1003912
rect 424322 1003856 424378 1003892
rect 424690 1002668 424692 1002688
rect 424692 1002668 424744 1002688
rect 424744 1002668 424746 1002688
rect 424690 1002632 424746 1002668
rect 421470 1001972 421526 1002008
rect 421470 1001952 421472 1001972
rect 421472 1001952 421524 1001972
rect 421524 1001952 421526 1001972
rect 425518 1001972 425574 1002008
rect 425518 1001952 425520 1001972
rect 425520 1001952 425572 1001972
rect 425572 1001952 425574 1001972
rect 427174 1005372 427230 1005408
rect 427174 1005352 427176 1005372
rect 427176 1005352 427228 1005372
rect 427228 1005352 427230 1005372
rect 428002 1004964 428058 1005000
rect 428002 1004944 428004 1004964
rect 428004 1004944 428056 1004964
rect 428056 1004944 428058 1004964
rect 553950 1007004 554006 1007040
rect 553950 1006984 553952 1007004
rect 553952 1006984 554004 1007004
rect 554004 1006984 554006 1007004
rect 505006 1006884 505008 1006904
rect 505008 1006884 505060 1006904
rect 505060 1006884 505062 1006904
rect 505006 1006848 505062 1006884
rect 507858 1006732 507914 1006768
rect 507858 1006712 507860 1006732
rect 507860 1006712 507912 1006732
rect 507912 1006712 507914 1006732
rect 505374 1006596 505430 1006632
rect 505374 1006576 505376 1006596
rect 505376 1006576 505428 1006596
rect 505428 1006576 505430 1006596
rect 426346 1002108 426402 1002144
rect 426346 1002088 426348 1002108
rect 426348 1002088 426400 1002108
rect 426400 1002088 426402 1002108
rect 430854 998300 430910 998336
rect 430854 998280 430856 998300
rect 430856 998280 430908 998300
rect 430908 998280 430910 998300
rect 430026 998164 430082 998200
rect 430026 998144 430028 998164
rect 430028 998144 430080 998164
rect 430080 998144 430082 998164
rect 430026 997892 430082 997928
rect 430026 997872 430028 997892
rect 430028 997872 430080 997892
rect 430080 997872 430082 997892
rect 432878 1004692 432934 1004728
rect 432878 1004672 432880 1004692
rect 432880 1004672 432932 1004692
rect 432932 1004672 432934 1004692
rect 432050 998028 432106 998064
rect 432050 998008 432052 998028
rect 432052 998008 432104 998028
rect 432104 998008 432106 998028
rect 435362 997736 435418 997792
rect 440054 997192 440110 997248
rect 439870 996920 439926 996976
rect 439686 996376 439742 996432
rect 451922 996104 451978 996160
rect 448518 995560 448574 995616
rect 458362 995288 458418 995344
rect 464986 995016 465042 995072
rect 457442 994472 457498 994528
rect 443642 994200 443698 994256
rect 506202 1006460 506258 1006496
rect 506202 1006440 506204 1006460
rect 506204 1006440 506256 1006460
rect 506256 1006440 506258 1006460
rect 498842 1006052 498898 1006088
rect 498842 1006032 498844 1006052
rect 498844 1006032 498896 1006052
rect 498896 1006032 498898 1006052
rect 469862 995832 469918 995888
rect 471058 996104 471114 996160
rect 471242 996104 471298 996160
rect 471242 995016 471298 995072
rect 471058 994744 471114 994800
rect 488906 997192 488962 997248
rect 489090 996920 489146 996976
rect 472622 996648 472678 996704
rect 489826 996648 489882 996704
rect 490010 996648 490066 996704
rect 474738 995560 474794 995616
rect 472254 995016 472310 995072
rect 474002 995016 474058 995072
rect 476394 995016 476450 995072
rect 477038 995016 477094 995072
rect 474462 994744 474518 994800
rect 480810 995016 480866 995072
rect 484122 995016 484178 995072
rect 484582 995016 484638 995072
rect 481638 994472 481694 994528
rect 486330 995288 486386 995344
rect 487802 994744 487858 994800
rect 500498 1005388 500500 1005408
rect 500500 1005388 500552 1005408
rect 500552 1005388 500554 1005408
rect 498842 1005252 498844 1005272
rect 498844 1005252 498896 1005272
rect 498896 1005252 498898 1005272
rect 498842 1005216 498898 1005252
rect 500498 1005352 500554 1005388
rect 500498 1004964 500554 1005000
rect 500498 1004944 500500 1004964
rect 500500 1004944 500552 1004964
rect 500552 1004944 500554 1004964
rect 499670 1004828 499726 1004864
rect 499670 1004808 499672 1004828
rect 499672 1004808 499724 1004828
rect 499724 1004808 499726 1004828
rect 555974 1006868 556030 1006904
rect 555974 1006848 555976 1006868
rect 555976 1006848 556028 1006868
rect 556028 1006848 556030 1006868
rect 556802 1006732 556858 1006768
rect 556802 1006712 556804 1006732
rect 556804 1006712 556856 1006732
rect 556856 1006712 556858 1006732
rect 509882 1002516 509938 1002552
rect 509882 1002496 509884 1002516
rect 509884 1002496 509936 1002516
rect 509936 1002496 509938 1002516
rect 501694 1002380 501750 1002416
rect 501694 1002360 501696 1002380
rect 501696 1002360 501748 1002380
rect 501748 1002360 501750 1002380
rect 503350 1002244 503406 1002280
rect 503350 1002224 503352 1002244
rect 503352 1002224 503404 1002244
rect 503404 1002224 503406 1002244
rect 501694 1002088 501750 1002144
rect 502522 1002108 502578 1002144
rect 502522 1002088 502524 1002108
rect 502524 1002088 502576 1002108
rect 502576 1002088 502578 1002108
rect 501326 1001972 501382 1002008
rect 501326 1001952 501328 1001972
rect 501328 1001952 501380 1001972
rect 501380 1001952 501382 1001972
rect 502154 1001952 502210 1002008
rect 503350 1001952 503406 1002008
rect 504178 1002244 504234 1002280
rect 504178 1002224 504180 1002244
rect 504180 1002224 504232 1002244
rect 504232 1002224 504234 1002244
rect 504546 1001972 504602 1002008
rect 504546 1001952 504548 1001972
rect 504548 1001952 504600 1001972
rect 504600 1001952 504602 1001972
rect 505374 998980 505430 999016
rect 505374 998960 505376 998980
rect 505376 998960 505428 998980
rect 505428 998960 505430 998980
rect 507398 999116 507454 999152
rect 507398 999096 507400 999116
rect 507400 999096 507452 999116
rect 507452 999096 507454 999116
rect 507030 998708 507086 998744
rect 507030 998688 507032 998708
rect 507032 998688 507084 998708
rect 507084 998688 507086 998708
rect 509054 998300 509110 998336
rect 509054 998280 509056 998300
rect 509056 998280 509108 998300
rect 509108 998280 509110 998300
rect 508226 998164 508282 998200
rect 508226 998144 508228 998164
rect 508228 998144 508280 998164
rect 508280 998144 508282 998164
rect 508226 997908 508228 997928
rect 508228 997908 508280 997928
rect 508280 997908 508282 997928
rect 508226 997872 508282 997908
rect 512642 997736 512698 997792
rect 511446 997192 511502 997248
rect 478602 994200 478658 994256
rect 485318 994200 485374 994256
rect 511078 994200 511134 994256
rect 467102 993928 467158 993984
rect 474462 993928 474518 993984
rect 516690 998572 516746 998608
rect 516690 998552 516692 998572
rect 516692 998552 516744 998572
rect 516744 998552 516746 998572
rect 516874 996920 516930 996976
rect 516690 996648 516746 996704
rect 518898 998552 518954 998608
rect 519082 996376 519138 996432
rect 518898 995560 518954 995616
rect 518162 995288 518218 995344
rect 555146 1006460 555202 1006496
rect 555146 1006440 555148 1006460
rect 555148 1006440 555200 1006460
rect 555200 1006440 555202 1006460
rect 551466 1006324 551522 1006360
rect 551466 1006304 551468 1006324
rect 551468 1006304 551520 1006324
rect 551520 1006304 551522 1006324
rect 550270 1006052 550326 1006088
rect 550270 1006032 550272 1006052
rect 550272 1006032 550324 1006052
rect 550324 1006032 550326 1006052
rect 554778 1006052 554834 1006088
rect 554778 1006032 554780 1006052
rect 554780 1006032 554832 1006052
rect 554832 1006032 554834 1006052
rect 520922 995016 520978 995072
rect 523498 996648 523554 996704
rect 523866 997600 523922 997656
rect 551466 1005252 551468 1005272
rect 551468 1005252 551520 1005272
rect 551520 1005252 551522 1005272
rect 551466 1005216 551522 1005252
rect 554778 1003312 554834 1003368
rect 553122 1002652 553178 1002688
rect 553122 1002632 553124 1002652
rect 553124 1002632 553176 1002652
rect 553176 1002632 553178 1002652
rect 550270 1001172 550272 1001192
rect 550272 1001172 550324 1001192
rect 550324 1001172 550326 1001192
rect 550270 1001136 550326 1001172
rect 524050 997192 524106 997248
rect 540334 996920 540390 996976
rect 524050 996376 524106 996432
rect 523682 996104 523738 996160
rect 529754 995696 529810 995752
rect 532146 995696 532202 995752
rect 532882 995696 532938 995752
rect 535274 995696 535330 995752
rect 536562 995696 536618 995752
rect 529018 995560 529074 995616
rect 533526 995560 533582 995616
rect 523314 994200 523370 994256
rect 526074 994472 526130 994528
rect 537114 995288 537170 995344
rect 552294 997736 552350 997792
rect 552294 997228 552296 997248
rect 552296 997228 552348 997248
rect 552348 997228 552350 997248
rect 552294 997192 552350 997228
rect 553950 1002124 553952 1002144
rect 553952 1002124 554004 1002144
rect 554004 1002124 554006 1002144
rect 553950 1002088 554006 1002124
rect 555974 1004828 556030 1004864
rect 555974 1004808 555976 1004828
rect 555976 1004808 556028 1004828
rect 556028 1004808 556030 1004828
rect 553122 996512 553178 996568
rect 558826 1006188 558882 1006224
rect 558826 1006168 558828 1006188
rect 558828 1006168 558880 1006188
rect 558880 1006168 558882 1006188
rect 557170 1004964 557226 1005000
rect 557170 1004944 557172 1004964
rect 557172 1004944 557224 1004964
rect 557224 1004944 557226 1004964
rect 557630 1004692 557686 1004728
rect 557630 1004672 557632 1004692
rect 557632 1004672 557684 1004692
rect 557684 1004672 557686 1004692
rect 557998 1002244 558054 1002280
rect 557998 1002224 558000 1002244
rect 558000 1002224 558052 1002244
rect 558052 1002224 558054 1002244
rect 557998 1001972 558054 1002008
rect 557998 1001952 558000 1001972
rect 558000 1001952 558052 1001972
rect 558052 1001952 558054 1001972
rect 560850 1004692 560906 1004728
rect 560850 1004672 560852 1004692
rect 560852 1004672 560904 1004692
rect 560904 1004672 560906 1004692
rect 558826 1002652 558882 1002688
rect 558826 1002632 558828 1002652
rect 558828 1002632 558880 1002652
rect 558880 1002632 558882 1002652
rect 528926 994200 528982 994256
rect 560850 1002516 560906 1002552
rect 560850 1002496 560852 1002516
rect 560852 1002496 560904 1002516
rect 560904 1002496 560906 1002516
rect 560482 1002380 560538 1002416
rect 560482 1002360 560484 1002380
rect 560484 1002360 560536 1002380
rect 560536 1002360 560538 1002380
rect 560022 1002108 560078 1002144
rect 560022 1002088 560024 1002108
rect 560024 1002088 560076 1002108
rect 560076 1002088 560078 1002108
rect 561678 1001972 561734 1002008
rect 561678 1001952 561680 1001972
rect 561680 1001952 561732 1001972
rect 561732 1001952 561734 1001972
rect 572810 994880 572866 994936
rect 570786 994608 570842 994664
rect 590566 996940 590622 996976
rect 590566 996920 590568 996940
rect 590568 996920 590620 996940
rect 590620 996920 590622 996940
rect 590566 996684 590568 996704
rect 590568 996684 590620 996704
rect 590620 996684 590622 996704
rect 590566 996648 590622 996684
rect 590566 996376 590622 996432
rect 590566 995288 590622 995344
rect 590566 995016 590622 995072
rect 625066 997192 625122 997248
rect 625250 997192 625306 997248
rect 625158 994472 625214 994528
rect 625618 995968 625674 996024
rect 625802 995696 625858 995752
rect 627182 995696 627238 995752
rect 629206 995696 629262 995752
rect 629850 995696 629906 995752
rect 630310 995730 630366 995786
rect 635646 995696 635702 995752
rect 637026 995696 637082 995752
rect 635186 995560 635242 995616
rect 627918 994744 627974 994800
rect 635830 995288 635886 995344
rect 635646 994744 635702 994800
rect 640982 995016 641038 995072
rect 62118 975976 62174 976032
rect 651654 975840 651710 975896
rect 62118 962920 62174 962976
rect 651470 962512 651526 962568
rect 62118 949864 62174 949920
rect 652206 949320 652262 949376
rect 651470 936128 651526 936184
rect 661682 957752 661738 957808
rect 660302 937216 660358 937272
rect 664442 947280 664498 947336
rect 663062 941704 663118 941760
rect 665822 939800 665878 939856
rect 674378 966048 674434 966104
rect 673366 962784 673422 962840
rect 673090 962512 673146 962568
rect 672906 958704 672962 958760
rect 668582 938440 668638 938496
rect 672170 938032 672226 938088
rect 667202 937760 667258 937816
rect 672814 937760 672870 937816
rect 672630 937488 672686 937544
rect 672170 937216 672226 937272
rect 671802 936672 671858 936728
rect 658922 935992 658978 936048
rect 671618 935720 671674 935776
rect 62118 923752 62174 923808
rect 651470 922664 651526 922720
rect 62118 910696 62174 910752
rect 652390 909492 652446 909528
rect 652390 909472 652392 909492
rect 652392 909472 652444 909492
rect 652444 909472 652446 909492
rect 62118 897776 62174 897832
rect 651470 896144 651526 896200
rect 54482 892200 54538 892256
rect 55862 892200 55918 892256
rect 651654 882816 651710 882872
rect 62118 871664 62174 871720
rect 651470 869624 651526 869680
rect 62762 858608 62818 858664
rect 62118 845552 62174 845608
rect 53102 799176 53158 799232
rect 62118 832496 62174 832552
rect 54482 774288 54538 774344
rect 62118 819440 62174 819496
rect 62118 806520 62174 806576
rect 652390 856296 652446 856352
rect 652022 842968 652078 843024
rect 651470 829776 651526 829832
rect 651470 816448 651526 816504
rect 651470 803276 651526 803312
rect 651470 803256 651472 803276
rect 651472 803256 651524 803276
rect 651524 803256 651526 803276
rect 62946 793600 63002 793656
rect 62762 788568 62818 788624
rect 62762 780408 62818 780464
rect 55862 772792 55918 772848
rect 62118 767372 62174 767408
rect 62118 767352 62120 767372
rect 62120 767352 62172 767372
rect 62172 767352 62174 767372
rect 62118 754296 62174 754352
rect 50342 730496 50398 730552
rect 48962 669296 49018 669352
rect 47398 638016 47454 638072
rect 47398 620336 47454 620392
rect 45190 598848 45246 598904
rect 45190 598440 45246 598496
rect 45006 598032 45062 598088
rect 62762 743008 62818 743064
rect 651470 789928 651526 789984
rect 651470 776600 651526 776656
rect 651470 763292 651526 763328
rect 651470 763272 651472 763292
rect 651472 763272 651524 763292
rect 651524 763272 651526 763292
rect 651470 750080 651526 750136
rect 62946 741648 63002 741704
rect 62118 741240 62174 741296
rect 51722 691328 51778 691384
rect 51722 646584 51778 646640
rect 62762 728184 62818 728240
rect 62118 715264 62174 715320
rect 62118 702208 62174 702264
rect 54482 688064 54538 688120
rect 53102 644680 53158 644736
rect 50342 627272 50398 627328
rect 51722 601704 51778 601760
rect 48962 601296 49018 601352
rect 651470 723424 651526 723480
rect 652574 736752 652630 736808
rect 652022 718256 652078 718312
rect 660302 778912 660358 778968
rect 658922 715944 658978 716000
rect 652574 710232 652630 710288
rect 62762 697856 62818 697912
rect 652390 696940 652392 696960
rect 652392 696940 652444 696960
rect 652444 696940 652446 696960
rect 652390 696904 652446 696940
rect 62118 689152 62174 689208
rect 652022 683576 652078 683632
rect 62118 676096 62174 676152
rect 651470 670384 651526 670440
rect 62118 663040 62174 663096
rect 651470 657056 651526 657112
rect 62118 649984 62174 650040
rect 651470 643728 651526 643784
rect 55862 643184 55918 643240
rect 62118 637064 62174 637120
rect 651470 630536 651526 630592
rect 62118 624008 62174 624064
rect 651470 617208 651526 617264
rect 62118 610952 62174 611008
rect 54482 600888 54538 600944
rect 47582 582392 47638 582448
rect 44822 556416 44878 556472
rect 44362 556008 44418 556064
rect 44178 548664 44234 548720
rect 43626 547712 43682 547768
rect 43810 547032 43866 547088
rect 43350 375400 43406 375456
rect 42798 365744 42854 365800
rect 42430 364248 42486 364304
rect 41786 363568 41842 363624
rect 41786 360032 41842 360088
rect 42154 359896 42210 359952
rect 41786 359352 41842 359408
rect 41786 358672 41842 358728
rect 42430 356904 42486 356960
rect 42154 356360 42210 356416
rect 43350 355816 43406 355872
rect 41878 355680 41934 355736
rect 44178 536832 44234 536888
rect 48962 557776 49018 557832
rect 51722 557504 51778 557560
rect 45558 556824 45614 556880
rect 45006 555600 45062 555656
rect 44822 555192 44878 555248
rect 44638 554376 44694 554432
rect 44362 428848 44418 428904
rect 44178 428440 44234 428496
rect 43994 419464 44050 419520
rect 44454 427624 44510 427680
rect 44178 385600 44234 385656
rect 45006 551520 45062 551576
rect 45190 550704 45246 550760
rect 45374 549072 45430 549128
rect 45374 537104 45430 537160
rect 45190 532752 45246 532808
rect 45006 529624 45062 529680
rect 45558 429664 45614 429720
rect 45006 429256 45062 429312
rect 44822 428032 44878 428088
rect 44638 427216 44694 427272
rect 44638 421504 44694 421560
rect 44822 420688 44878 420744
rect 44638 406952 44694 407008
rect 44638 385192 44694 385248
rect 44454 384784 44510 384840
rect 45190 426808 45246 426864
rect 45006 386688 45062 386744
rect 45006 384376 45062 384432
rect 44454 377848 44510 377904
rect 44270 377440 44326 377496
rect 44454 364928 44510 364984
rect 44270 356632 44326 356688
rect 45558 426400 45614 426456
rect 45374 422320 45430 422376
rect 45374 405592 45430 405648
rect 45558 399744 45614 399800
rect 45374 386008 45430 386064
rect 45190 383968 45246 384024
rect 45190 383560 45246 383616
rect 43902 354184 43958 354240
rect 44730 353776 44786 353832
rect 28538 351192 28594 351248
rect 40222 345344 40278 345400
rect 28906 344256 28962 344312
rect 28538 343848 28594 343904
rect 45006 341672 45062 341728
rect 45558 380704 45614 380760
rect 45742 379888 45798 379944
rect 47582 430072 47638 430128
rect 46938 423544 46994 423600
rect 46938 400152 46994 400208
rect 46938 383152 46994 383208
rect 46202 366968 46258 367024
rect 45742 359896 45798 359952
rect 45558 356904 45614 356960
rect 45650 356632 45706 356688
rect 45926 355816 45982 355872
rect 45374 343304 45430 343360
rect 45190 340856 45246 340912
rect 45558 340040 45614 340096
rect 35806 339768 35862 339824
rect 35806 338952 35862 339008
rect 31022 338544 31078 338600
rect 31022 329024 31078 329080
rect 45374 337184 45430 337240
rect 42890 334600 42946 334656
rect 43258 334600 43314 334656
rect 44178 334600 44234 334656
rect 37922 334464 37978 334520
rect 42614 334328 42670 334384
rect 36542 328344 36598 328400
rect 41786 326712 41842 326768
rect 42614 326440 42670 326496
rect 41786 325352 41842 325408
rect 41878 324672 41934 324728
rect 42062 322768 42118 322824
rect 42430 321408 42486 321464
rect 41786 321000 41842 321056
rect 42982 326440 43038 326496
rect 43258 322768 43314 322824
rect 42430 318960 42486 319016
rect 42430 317328 42486 317384
rect 44178 317328 44234 317384
rect 42430 316376 42486 316432
rect 42154 315968 42210 316024
rect 45466 315968 45522 316024
rect 41786 315560 41842 315616
rect 42154 313656 42210 313712
rect 45650 313656 45706 313712
rect 42430 312704 42486 312760
rect 41786 312568 41842 312624
rect 44730 311752 44786 311808
rect 44178 311480 44234 311536
rect 41786 303048 41842 303104
rect 41786 300872 41842 300928
rect 44546 311208 44602 311264
rect 44178 299240 44234 299296
rect 44270 298832 44326 298888
rect 43258 298016 43314 298072
rect 42890 297200 42946 297256
rect 41786 296792 41842 296848
rect 32402 294752 32458 294808
rect 42062 295976 42118 296032
rect 41786 292712 41842 292768
rect 42062 292304 42118 292360
rect 42246 291080 42302 291136
rect 42062 290400 42118 290456
rect 41326 290264 41382 290320
rect 42062 289856 42118 289912
rect 42246 289856 42302 289912
rect 41970 281424 42026 281480
rect 42154 279792 42210 279848
rect 42430 278704 42486 278760
rect 42430 278160 42486 278216
rect 41786 277888 41842 277944
rect 42338 277616 42394 277672
rect 42062 277072 42118 277128
rect 42062 276528 42118 276584
rect 41786 274216 41842 274272
rect 42062 273400 42118 273456
rect 42062 272856 42118 272912
rect 41786 270408 41842 270464
rect 42430 270408 42486 270464
rect 41786 269048 41842 269104
rect 43074 293528 43130 293584
rect 43074 273400 43130 273456
rect 40682 267008 40738 267064
rect 35806 257080 35862 257136
rect 42890 254768 42946 254824
rect 35622 253408 35678 253464
rect 35438 253000 35494 253056
rect 35806 253000 35862 253056
rect 35806 252184 35862 252240
rect 41694 242836 41696 242856
rect 41696 242836 41748 242856
rect 41748 242836 41750 242856
rect 41694 242800 41750 242836
rect 40682 242528 40738 242584
rect 41786 240080 41842 240136
rect 42062 238448 42118 238504
rect 42706 242800 42762 242856
rect 42522 237360 42578 237416
rect 41786 235864 41842 235920
rect 42430 235864 42486 235920
rect 42246 234504 42302 234560
rect 42338 234096 42394 234152
rect 42338 233144 42394 233200
rect 42338 231784 42394 231840
rect 42154 230288 42210 230344
rect 42338 229336 42394 229392
rect 42430 227568 42486 227624
rect 41970 227296 42026 227352
rect 43442 294344 43498 294400
rect 43626 293120 43682 293176
rect 43810 291896 43866 291952
rect 43626 279792 43682 279848
rect 43810 277072 43866 277128
rect 43442 270408 43498 270464
rect 43718 256400 43774 256456
rect 43442 255584 43498 255640
rect 43258 255176 43314 255232
rect 43074 254360 43130 254416
rect 43074 249056 43130 249112
rect 43534 251096 43590 251152
rect 43258 242528 43314 242584
rect 43074 231784 43130 231840
rect 42430 225664 42486 225720
rect 43166 225664 43222 225720
rect 43534 227568 43590 227624
rect 40682 222808 40738 222864
rect 35530 217912 35586 217968
rect 35530 214240 35586 214296
rect 35806 214240 35862 214296
rect 44730 300056 44786 300112
rect 44730 299648 44786 299704
rect 44546 298424 44602 298480
rect 44454 291488 44510 291544
rect 44454 278160 44510 278216
rect 44638 256808 44694 256864
rect 44270 255992 44326 256048
rect 44178 253952 44234 254008
rect 43718 213696 43774 213752
rect 43442 212880 43498 212936
rect 43442 212472 43498 212528
rect 42890 212064 42946 212120
rect 35806 211384 35862 211440
rect 42798 209344 42854 209400
rect 35806 208936 35862 208992
rect 41694 208936 41750 208992
rect 40038 207712 40094 207768
rect 35622 204040 35678 204096
rect 35806 203632 35862 203688
rect 35622 202136 35678 202192
rect 37922 197784 37978 197840
rect 41786 197104 41842 197160
rect 41878 195744 41934 195800
rect 41786 195200 41842 195256
rect 42246 194928 42302 194984
rect 42246 193160 42302 193216
rect 42338 192888 42394 192944
rect 42338 191664 42394 191720
rect 42430 191120 42486 191176
rect 42430 190440 42486 190496
rect 42430 189896 42486 189952
rect 42430 187584 42486 187640
rect 41786 187176 41842 187232
rect 42338 186224 42394 186280
rect 42154 185952 42210 186008
rect 42430 184864 42486 184920
rect 42430 183096 42486 183152
rect 43258 207984 43314 208040
rect 42982 206352 43038 206408
rect 42982 191120 43038 191176
rect 44638 251912 44694 251968
rect 44546 248648 44602 248704
rect 44362 248240 44418 248296
rect 44362 235864 44418 235920
rect 44546 234096 44602 234152
rect 44546 233144 44602 233200
rect 45006 295160 45062 295216
rect 45190 293936 45246 293992
rect 45006 276528 45062 276584
rect 45190 272856 45246 272912
rect 47122 379072 47178 379128
rect 47122 364248 47178 364304
rect 46938 356360 46994 356416
rect 47582 345344 47638 345400
rect 46938 338408 46994 338464
rect 47582 333104 47638 333160
rect 46938 318960 46994 319016
rect 46386 303048 46442 303104
rect 46202 257896 46258 257952
rect 45834 250688 45890 250744
rect 45558 250280 45614 250336
rect 45558 230288 45614 230344
rect 46018 249464 46074 249520
rect 46202 247832 46258 247888
rect 46018 234504 46074 234560
rect 45834 229336 45890 229392
rect 44822 214920 44878 214976
rect 44178 211248 44234 211304
rect 44178 210432 44234 210488
rect 43810 206760 43866 206816
rect 43442 206216 43498 206272
rect 43626 205536 43682 205592
rect 43442 202136 43498 202192
rect 43258 183096 43314 183152
rect 43994 205128 44050 205184
rect 43810 192888 43866 192944
rect 43994 191664 44050 191720
rect 43626 190440 43682 190496
rect 44546 208528 44602 208584
rect 44362 205944 44418 206000
rect 44822 204720 44878 204776
rect 44546 189896 44602 189952
rect 44362 187584 44418 187640
rect 44178 184864 44234 184920
rect 46938 247016 46994 247072
rect 46938 238448 46994 238504
rect 46386 203496 46442 203552
rect 50342 430888 50398 430944
rect 48962 386960 49018 387016
rect 51722 386688 51778 386744
rect 51906 386416 51962 386472
rect 50526 351192 50582 351248
rect 48962 334056 49018 334112
rect 47766 300464 47822 300520
rect 47766 247424 47822 247480
rect 47950 213288 48006 213344
rect 48134 210840 48190 210896
rect 48778 206216 48834 206272
rect 48134 194384 48190 194440
rect 48778 192344 48834 192400
rect 47950 190440 48006 190496
rect 54482 430480 54538 430536
rect 651470 603880 651526 603936
rect 62118 597896 62174 597952
rect 651470 590708 651526 590744
rect 651470 590688 651472 590708
rect 651472 590688 651524 590708
rect 651524 590688 651526 590708
rect 62118 584840 62174 584896
rect 669226 879144 669282 879200
rect 664442 868672 664498 868728
rect 668214 868128 668270 868184
rect 663062 760824 663118 760880
rect 661682 760416 661738 760472
rect 660302 625232 660358 625288
rect 660302 599528 660358 599584
rect 652022 582936 652078 582992
rect 666282 777008 666338 777064
rect 664442 716488 664498 716544
rect 663062 689288 663118 689344
rect 661866 643728 661922 643784
rect 661682 581032 661738 581088
rect 651470 577360 651526 577416
rect 62118 571784 62174 571840
rect 62118 569200 62174 569256
rect 651654 564032 651710 564088
rect 62118 558728 62174 558784
rect 658922 553968 658978 554024
rect 651470 550840 651526 550896
rect 62118 545808 62174 545864
rect 56046 540232 56102 540288
rect 651470 537512 651526 537568
rect 62118 532772 62174 532808
rect 62118 532752 62120 532772
rect 62120 532752 62172 532772
rect 62172 532752 62174 532772
rect 651838 524184 651894 524240
rect 62118 519696 62174 519752
rect 651470 510992 651526 511048
rect 62118 506640 62174 506696
rect 651470 497664 651526 497720
rect 62118 493584 62174 493640
rect 651470 484492 651526 484528
rect 651470 484472 651472 484492
rect 651472 484472 651524 484492
rect 651524 484472 651526 484492
rect 62118 480528 62174 480584
rect 651470 471144 651526 471200
rect 62118 467472 62174 467528
rect 652390 457816 652446 457872
rect 62118 454552 62174 454608
rect 651470 444508 651526 444544
rect 651470 444488 651472 444508
rect 651472 444488 651524 444508
rect 651524 444488 651526 444508
rect 62118 441496 62174 441552
rect 651470 431296 651526 431352
rect 62118 428440 62174 428496
rect 651838 417968 651894 418024
rect 62118 415420 62120 415440
rect 62120 415420 62172 415440
rect 62172 415420 62174 415440
rect 62118 415384 62174 415420
rect 55862 408448 55918 408504
rect 651470 404640 651526 404696
rect 62118 402328 62174 402384
rect 54482 344256 54538 344312
rect 53102 321408 53158 321464
rect 51722 301280 51778 301336
rect 49146 290400 49202 290456
rect 50342 290128 50398 290184
rect 49514 208936 49570 208992
rect 49514 196424 49570 196480
rect 51722 289856 51778 289912
rect 50526 246472 50582 246528
rect 53286 257488 53342 257544
rect 652574 391448 652630 391504
rect 62118 389292 62174 389328
rect 62118 389272 62120 389292
rect 62120 389272 62172 389292
rect 62172 389272 62174 389292
rect 652022 378120 652078 378176
rect 62118 376216 62174 376272
rect 651654 364792 651710 364848
rect 62118 363296 62174 363352
rect 651470 351600 651526 351656
rect 62762 350240 62818 350296
rect 62118 337184 62174 337240
rect 62118 324128 62174 324184
rect 62118 311072 62174 311128
rect 62118 298172 62174 298208
rect 62118 298152 62120 298172
rect 62120 298152 62172 298172
rect 62172 298152 62174 298172
rect 55862 278704 55918 278760
rect 651470 338272 651526 338328
rect 651470 324944 651526 325000
rect 651470 311752 651526 311808
rect 651470 285232 651526 285288
rect 62946 285096 63002 285152
rect 62762 267008 62818 267064
rect 54482 217912 54538 217968
rect 136546 269728 136602 269784
rect 139950 269764 139952 269784
rect 139952 269764 140004 269784
rect 140004 269764 140006 269784
rect 139950 269728 140006 269764
rect 473266 266620 473322 266656
rect 473266 266600 473268 266620
rect 473268 266600 473320 266620
rect 473320 266600 473322 266620
rect 474830 266620 474886 266656
rect 474830 266600 474832 266620
rect 474832 266600 474884 266620
rect 474884 266600 474886 266620
rect 494334 270308 494336 270328
rect 494336 270308 494388 270328
rect 494388 270308 494390 270328
rect 494334 270272 494390 270308
rect 494150 270000 494206 270056
rect 494886 270272 494942 270328
rect 499762 267164 499818 267200
rect 499762 267144 499764 267164
rect 499764 267144 499816 267164
rect 499816 267144 499818 267164
rect 501050 267164 501106 267200
rect 501050 267144 501052 267164
rect 501052 267144 501104 267164
rect 501104 267144 501106 267164
rect 502338 269592 502394 269648
rect 504178 270544 504234 270600
rect 504546 269628 504548 269648
rect 504548 269628 504600 269648
rect 504600 269628 504602 269648
rect 504546 269592 504602 269628
rect 506202 267144 506258 267200
rect 507858 270544 507914 270600
rect 507858 267164 507914 267200
rect 507858 267144 507860 267164
rect 507860 267144 507912 267164
rect 507912 267144 507914 267164
rect 511722 271396 511724 271416
rect 511724 271396 511776 271416
rect 511776 271396 511778 271416
rect 511722 271360 511778 271396
rect 509882 269728 509938 269784
rect 513194 272312 513250 272368
rect 515310 271396 515312 271416
rect 515312 271396 515364 271416
rect 515364 271396 515366 271416
rect 515310 271360 515366 271396
rect 516598 274100 516654 274136
rect 516598 274080 516600 274100
rect 516600 274080 516652 274100
rect 516652 274080 516654 274100
rect 518438 272312 518494 272368
rect 519726 274080 519782 274136
rect 518438 268504 518494 268560
rect 518990 268504 519046 268560
rect 519174 268368 519230 268424
rect 518898 267300 518954 267336
rect 518898 267280 518900 267300
rect 518900 267280 518952 267300
rect 518952 267280 518954 267300
rect 518714 266756 518770 266792
rect 518714 266736 518716 266756
rect 518716 266736 518768 266756
rect 518768 266736 518770 266756
rect 518898 266736 518954 266792
rect 521106 273672 521162 273728
rect 520462 268388 520518 268424
rect 520462 268368 520464 268388
rect 520464 268368 520516 268388
rect 520516 268368 520518 268388
rect 521474 272448 521530 272504
rect 524234 273672 524290 273728
rect 523958 271632 524014 271688
rect 523958 270852 523960 270872
rect 523960 270852 524012 270872
rect 524012 270852 524014 270872
rect 523958 270816 524014 270852
rect 523314 269728 523370 269784
rect 521658 269456 521714 269512
rect 524878 272448 524934 272504
rect 524602 272176 524658 272232
rect 525798 275712 525854 275768
rect 524786 271632 524842 271688
rect 524878 270852 524880 270872
rect 524880 270852 524932 270872
rect 524932 270852 524934 270872
rect 524878 270816 524934 270852
rect 526258 271088 526314 271144
rect 525522 268640 525578 268696
rect 524510 267008 524566 267064
rect 525890 267028 525946 267064
rect 525890 267008 525892 267028
rect 525892 267008 525944 267028
rect 525944 267008 525946 267028
rect 527822 274624 527878 274680
rect 527178 267280 527234 267336
rect 527638 267280 527694 267336
rect 530858 275732 530914 275768
rect 530858 275712 530860 275732
rect 530860 275712 530912 275732
rect 530912 275712 530914 275732
rect 528650 270716 528652 270736
rect 528652 270716 528704 270736
rect 528704 270716 528706 270736
rect 528650 270680 528706 270716
rect 529570 271124 529572 271144
rect 529572 271124 529624 271144
rect 529624 271124 529626 271144
rect 529570 271088 529626 271124
rect 529754 271088 529810 271144
rect 531502 272176 531558 272232
rect 535090 275304 535146 275360
rect 534078 272720 534134 272776
rect 533526 272448 533582 272504
rect 534170 272484 534172 272504
rect 534172 272484 534224 272504
rect 534224 272484 534226 272504
rect 534170 272448 534226 272484
rect 533158 270680 533214 270736
rect 531410 270000 531466 270056
rect 532882 269728 532938 269784
rect 532698 269456 532754 269512
rect 532238 266872 532294 266928
rect 533894 270816 533950 270872
rect 534354 270816 534410 270872
rect 533894 269728 533950 269784
rect 533894 268640 533950 268696
rect 533894 267688 533950 267744
rect 533710 267280 533766 267336
rect 533894 267144 533950 267200
rect 534170 267144 534226 267200
rect 534078 266600 534134 266656
rect 536838 275596 536894 275632
rect 536838 275576 536840 275596
rect 536840 275576 536892 275596
rect 536892 275576 536894 275596
rect 536746 273808 536802 273864
rect 535918 269456 535974 269512
rect 535458 267688 535514 267744
rect 537942 275596 537998 275632
rect 537942 275576 537944 275596
rect 537944 275576 537996 275596
rect 537996 275576 537998 275596
rect 538678 275324 538734 275360
rect 538678 275304 538680 275324
rect 538680 275304 538732 275324
rect 538732 275304 538734 275324
rect 538678 274896 538734 274952
rect 537022 269220 537024 269240
rect 537024 269220 537076 269240
rect 537076 269220 537078 269240
rect 537022 269184 537078 269220
rect 538126 269728 538182 269784
rect 537574 267552 537630 267608
rect 537390 266600 537446 266656
rect 541162 274896 541218 274952
rect 539506 270544 539562 270600
rect 538678 269184 538734 269240
rect 539230 268096 539286 268152
rect 543186 274624 543242 274680
rect 544842 272720 544898 272776
rect 543002 272448 543058 272504
rect 541990 269456 542046 269512
rect 542174 267280 542230 267336
rect 543554 271496 543610 271552
rect 546222 271496 546278 271552
rect 543554 270544 543610 270600
rect 543554 267552 543610 267608
rect 547510 268388 547566 268424
rect 547510 268368 547512 268388
rect 547512 268368 547564 268388
rect 547564 268368 547566 268388
rect 547694 268096 547750 268152
rect 552202 270680 552258 270736
rect 549258 268368 549314 268424
rect 553398 270680 553454 270736
rect 574466 270272 574522 270328
rect 607862 267280 607918 267336
rect 625066 271088 625122 271144
rect 627918 270000 627974 270056
rect 635646 273808 635702 273864
rect 637578 269728 637634 269784
rect 645122 272448 645178 272504
rect 629298 267008 629354 267064
rect 554410 262112 554466 262168
rect 554318 259936 554374 259992
rect 553950 257760 554006 257816
rect 553674 255584 553730 255640
rect 553490 251252 553546 251288
rect 553490 251232 553492 251252
rect 553492 251232 553544 251252
rect 553544 251232 553546 251252
rect 554502 253428 554558 253464
rect 554502 253408 554504 253428
rect 554504 253408 554556 253428
rect 554556 253408 554558 253428
rect 553858 249056 553914 249112
rect 554410 246880 554466 246936
rect 554502 244704 554558 244760
rect 553950 242528 554006 242584
rect 553858 240352 553914 240408
rect 554318 238176 554374 238232
rect 554502 236036 554504 236056
rect 554504 236036 554556 236056
rect 554556 236036 554558 236056
rect 554502 236000 554558 236036
rect 554410 233824 554466 233880
rect 62946 222808 63002 222864
rect 73066 226888 73122 226944
rect 68926 224168 68982 224224
rect 69754 220088 69810 220144
rect 72882 220360 72938 220416
rect 79966 228248 80022 228304
rect 103610 229744 103666 229800
rect 101862 221448 101918 221504
rect 123482 222808 123538 222864
rect 135166 227976 135222 228032
rect 134982 226616 135038 226672
rect 135626 226636 135682 226672
rect 135626 226616 135628 226636
rect 135628 226616 135680 226636
rect 135680 226616 135682 226636
rect 139306 226480 139362 226536
rect 136546 226072 136602 226128
rect 138478 221176 138534 221232
rect 141146 227976 141202 228032
rect 142158 227160 142214 227216
rect 142250 226500 142306 226536
rect 142250 226480 142252 226500
rect 142252 226480 142304 226500
rect 142304 226480 142306 226500
rect 143078 227160 143134 227216
rect 141698 226108 141700 226128
rect 141700 226108 141752 226128
rect 141752 226108 141754 226128
rect 141698 226072 141754 226108
rect 142158 224576 142214 224632
rect 141790 223896 141846 223952
rect 140778 219564 140834 219600
rect 140778 219544 140780 219564
rect 140780 219544 140832 219564
rect 140832 219544 140834 219564
rect 143170 225528 143226 225584
rect 142618 223896 142674 223952
rect 142986 222436 142988 222456
rect 142988 222436 143040 222456
rect 143040 222436 143042 222456
rect 142986 222400 143042 222436
rect 142158 221856 142214 221912
rect 142250 221196 142306 221232
rect 142250 221176 142252 221196
rect 142252 221176 142304 221196
rect 142304 221176 142306 221196
rect 142158 220768 142214 220824
rect 141974 219816 142030 219872
rect 142250 219816 142306 219872
rect 142158 219564 142214 219600
rect 142158 219544 142160 219564
rect 142160 219544 142212 219564
rect 142212 219544 142214 219564
rect 142250 218748 142306 218784
rect 142250 218728 142252 218748
rect 142252 218728 142304 218748
rect 142304 218728 142306 218748
rect 145654 229744 145710 229800
rect 146298 229220 146354 229256
rect 146298 229200 146300 229220
rect 146300 229200 146352 229220
rect 146352 229200 146354 229220
rect 145930 225256 145986 225312
rect 145562 224032 145618 224088
rect 145010 222436 145012 222456
rect 145012 222436 145064 222456
rect 145064 222436 145066 222456
rect 145010 222400 145066 222436
rect 147954 229200 148010 229256
rect 146942 225936 146998 225992
rect 147126 225564 147128 225584
rect 147128 225564 147180 225584
rect 147180 225564 147182 225584
rect 147126 225528 147182 225564
rect 147678 228520 147734 228576
rect 147310 224576 147366 224632
rect 147678 223932 147680 223952
rect 147680 223932 147732 223952
rect 147732 223932 147734 223952
rect 147678 223896 147734 223932
rect 148414 220768 148470 220824
rect 148414 219292 148470 219328
rect 148414 219272 148422 219292
rect 148422 219272 148470 219292
rect 149794 228520 149850 228576
rect 150162 227180 150218 227216
rect 150162 227160 150164 227180
rect 150164 227160 150216 227180
rect 150216 227160 150218 227180
rect 149058 221856 149114 221912
rect 150714 220768 150770 220824
rect 148598 218728 148654 218784
rect 151910 227432 151966 227488
rect 151726 223760 151782 223816
rect 151082 220088 151138 220144
rect 152922 227432 152978 227488
rect 153106 226072 153162 226128
rect 152830 225936 152886 225992
rect 152554 224304 152610 224360
rect 152922 219272 152978 219328
rect 153290 225256 153346 225312
rect 153658 220496 153714 220552
rect 152094 218884 152150 218920
rect 152094 218864 152096 218884
rect 152096 218864 152148 218884
rect 152148 218864 152150 218884
rect 154578 227160 154634 227216
rect 155866 227976 155922 228032
rect 155314 226888 155370 226944
rect 154578 224168 154634 224224
rect 155038 222536 155094 222592
rect 153842 218864 153898 218920
rect 156142 220768 156198 220824
rect 157430 228520 157486 228576
rect 157982 228928 158038 228984
rect 157798 227976 157854 228032
rect 157614 226108 157616 226128
rect 157616 226108 157668 226128
rect 157668 226108 157670 226128
rect 157614 226072 157670 226108
rect 156878 223760 156934 223816
rect 156878 223252 156880 223272
rect 156880 223252 156932 223272
rect 156932 223252 156934 223272
rect 156878 223216 156934 223252
rect 157338 224576 157394 224632
rect 157430 224168 157486 224224
rect 157430 223252 157432 223272
rect 157432 223252 157484 223272
rect 157484 223252 157486 223272
rect 157430 223216 157486 223252
rect 157246 222536 157302 222592
rect 157338 220516 157394 220552
rect 157338 220496 157340 220516
rect 157340 220496 157392 220516
rect 157392 220496 157394 220516
rect 157246 218592 157302 218648
rect 158810 228520 158866 228576
rect 159638 227452 159694 227488
rect 159638 227432 159640 227452
rect 159640 227432 159692 227452
rect 159692 227432 159694 227452
rect 160466 228248 160522 228304
rect 158350 223080 158406 223136
rect 157706 218476 157762 218512
rect 157706 218456 157708 218476
rect 157708 218456 157760 218476
rect 157760 218456 157762 218476
rect 161202 226072 161258 226128
rect 162306 226072 162362 226128
rect 162306 225528 162362 225584
rect 161754 220496 161810 220552
rect 161938 220496 161994 220552
rect 159638 218204 159694 218240
rect 159638 218184 159640 218204
rect 159640 218184 159692 218204
rect 159692 218184 159694 218204
rect 163870 228928 163926 228984
rect 162950 224576 163006 224632
rect 163962 224440 164018 224496
rect 162858 220516 162914 220552
rect 162858 220496 162860 220516
rect 162860 220496 162912 220516
rect 162912 220496 162914 220516
rect 165066 223116 165068 223136
rect 165068 223116 165120 223136
rect 165120 223116 165122 223136
rect 162858 218184 162914 218240
rect 165066 223080 165122 223116
rect 166446 228812 166502 228848
rect 166446 228792 166448 228812
rect 166448 228792 166500 228812
rect 166500 228792 166502 228812
rect 166446 228384 166502 228440
rect 166630 227432 166686 227488
rect 166814 225972 166816 225992
rect 166816 225972 166868 225992
rect 166868 225972 166870 225992
rect 166814 225936 166870 225972
rect 166906 225528 166962 225584
rect 166446 225020 166448 225040
rect 166448 225020 166500 225040
rect 166500 225020 166502 225040
rect 166446 224984 166502 225020
rect 166446 223080 166502 223136
rect 165618 222808 165674 222864
rect 166262 219272 166318 219328
rect 166998 225256 167054 225312
rect 166078 218884 166134 218920
rect 166078 218864 166080 218884
rect 166080 218864 166132 218884
rect 166132 218864 166134 218884
rect 167642 229200 167698 229256
rect 167366 225020 167368 225040
rect 167368 225020 167420 225040
rect 167420 225020 167422 225040
rect 167366 224984 167422 225020
rect 168194 228792 168250 228848
rect 168010 228384 168066 228440
rect 169206 226072 169262 226128
rect 169022 225936 169078 225992
rect 167090 218864 167146 218920
rect 169114 219292 169170 219328
rect 169114 219272 169116 219292
rect 169116 219272 169168 219292
rect 169168 219272 169170 219292
rect 169850 225256 169906 225312
rect 170770 224440 170826 224496
rect 172426 229220 172482 229256
rect 172426 229200 172428 229220
rect 172428 229200 172480 229220
rect 172480 229200 172482 229220
rect 172426 228928 172482 228984
rect 170954 224168 171010 224224
rect 171414 224168 171470 224224
rect 170402 223080 170458 223136
rect 171230 222264 171286 222320
rect 171046 221856 171102 221912
rect 171506 221876 171562 221912
rect 171506 221856 171508 221876
rect 171508 221856 171560 221876
rect 171560 221856 171562 221876
rect 175646 228948 175702 228984
rect 175646 228928 175648 228948
rect 175648 228928 175700 228948
rect 175700 228928 175702 228948
rect 176474 225528 176530 225584
rect 177026 225528 177082 225584
rect 176474 225256 176530 225312
rect 177210 225256 177266 225312
rect 176106 222028 176108 222048
rect 176108 222028 176160 222048
rect 176160 222028 176162 222048
rect 176106 221992 176162 222028
rect 177026 221992 177082 222048
rect 178682 225972 178684 225992
rect 178684 225972 178736 225992
rect 178736 225972 178738 225992
rect 178682 225936 178738 225972
rect 178038 221448 178094 221504
rect 180614 228928 180670 228984
rect 179970 222264 180026 222320
rect 181258 228692 181260 228712
rect 181260 228692 181312 228712
rect 181312 228692 181314 228712
rect 181258 228656 181314 228692
rect 181074 227996 181130 228032
rect 181074 227976 181076 227996
rect 181076 227976 181128 227996
rect 181128 227976 181130 227996
rect 180614 221176 180670 221232
rect 180890 221176 180946 221232
rect 180798 220768 180854 220824
rect 181902 228948 181958 228984
rect 181902 228928 181904 228948
rect 181904 228928 181956 228948
rect 181956 228928 181958 228948
rect 181902 228656 181958 228712
rect 181718 227976 181774 228032
rect 183282 225120 183338 225176
rect 184846 225664 184902 225720
rect 185674 225936 185730 225992
rect 185674 225392 185730 225448
rect 185674 224848 185730 224904
rect 185950 220768 186006 220824
rect 187330 225664 187386 225720
rect 187054 224848 187110 224904
rect 187514 225120 187570 225176
rect 190550 228812 190606 228848
rect 190550 228792 190552 228812
rect 190552 228792 190604 228812
rect 190604 228792 190606 228812
rect 192850 228792 192906 228848
rect 195426 225936 195482 225992
rect 194874 225392 194930 225448
rect 194782 220788 194838 220824
rect 194782 220768 194784 220788
rect 194784 220768 194836 220788
rect 194836 220768 194838 220788
rect 195058 219272 195114 219328
rect 196070 220788 196126 220824
rect 196070 220768 196072 220788
rect 196072 220768 196124 220788
rect 196124 220768 196126 220788
rect 196070 219292 196126 219328
rect 196070 219272 196072 219292
rect 196072 219272 196124 219292
rect 196124 219272 196126 219292
rect 484582 219408 484638 219464
rect 486606 220904 486662 220960
rect 487802 218048 487858 218104
rect 490562 219136 490618 219192
rect 491114 219136 491170 219192
rect 490286 218864 490342 218920
rect 491114 218592 491170 218648
rect 492126 217096 492182 217152
rect 492954 219136 493010 219192
rect 493598 219136 493654 219192
rect 494794 219680 494850 219736
rect 493598 217232 493654 217288
rect 497738 219136 497794 219192
rect 496910 218320 496966 218376
rect 497554 217232 497610 217288
rect 498658 217504 498714 217560
rect 500038 218340 500094 218376
rect 500038 218320 500040 218340
rect 500040 218320 500092 218340
rect 500092 218320 500094 218340
rect 500222 218320 500278 218376
rect 502522 219136 502578 219192
rect 502706 219136 502762 219192
rect 503534 217504 503590 217560
rect 505098 219136 505154 219192
rect 505282 219136 505338 219192
rect 504822 218592 504878 218648
rect 505282 218626 505338 218682
rect 504638 218320 504694 218376
rect 504822 217776 504878 217832
rect 505466 217812 505468 217832
rect 505468 217812 505520 217832
rect 505520 217812 505522 217832
rect 505466 217776 505522 217812
rect 506018 217504 506074 217560
rect 507306 218320 507362 218376
rect 508502 217776 508558 217832
rect 510986 219952 511042 220008
rect 513378 221876 513434 221912
rect 513378 221856 513380 221876
rect 513380 221856 513432 221876
rect 513432 221856 513434 221876
rect 512642 219952 512698 220008
rect 515954 221176 516010 221232
rect 514482 219136 514538 219192
rect 514758 219136 514814 219192
rect 514666 218286 514722 218342
rect 516598 219136 516654 219192
rect 517794 221448 517850 221504
rect 519542 220224 519598 220280
rect 519542 219680 519598 219736
rect 519818 219680 519874 219736
rect 522578 219680 522634 219736
rect 524418 219156 524474 219192
rect 524418 219136 524420 219156
rect 524420 219136 524472 219156
rect 524472 219136 524474 219156
rect 524602 219136 524658 219192
rect 524142 218320 524198 218376
rect 524602 218320 524658 218376
rect 524418 217776 524474 217832
rect 524602 217776 524658 217832
rect 530030 219952 530086 220008
rect 530306 219952 530362 220008
rect 534170 219136 534226 219192
rect 533710 218320 533766 218376
rect 533894 218320 533950 218376
rect 534078 218048 534134 218104
rect 534262 218048 534318 218104
rect 534630 219136 534686 219192
rect 542542 220224 542598 220280
rect 542358 219136 542414 219192
rect 541990 217232 542046 217288
rect 545026 220496 545082 220552
rect 545302 220496 545358 220552
rect 543370 220224 543426 220280
rect 543370 219136 543426 219192
rect 544014 218320 544070 218376
rect 543462 218048 543518 218104
rect 543646 218048 543702 218104
rect 543830 217232 543886 217288
rect 553030 220224 553086 220280
rect 555790 222012 555846 222048
rect 555790 221992 555792 222012
rect 555792 221992 555844 222012
rect 555844 221992 555846 222012
rect 556710 220224 556766 220280
rect 558366 218320 558422 218376
rect 558550 218320 558606 218376
rect 560666 222264 560722 222320
rect 561954 222264 562010 222320
rect 562690 222264 562746 222320
rect 563426 222012 563482 222048
rect 563426 221992 563428 222012
rect 563428 221992 563480 222012
rect 563480 221992 563482 222012
rect 562506 220224 562562 220280
rect 562874 220224 562930 220280
rect 563058 217776 563114 217832
rect 563242 217776 563298 217832
rect 564346 217776 564402 217832
rect 564530 217776 564586 217832
rect 565634 222536 565690 222592
rect 566830 220496 566886 220552
rect 567014 220496 567070 220552
rect 567658 219136 567714 219192
rect 568118 218320 568174 218376
rect 572304 221992 572360 222048
rect 572994 220224 573050 220280
rect 571614 218320 571670 218376
rect 571154 217776 571210 217832
rect 575846 220224 575902 220280
rect 574374 217776 574430 217832
rect 574558 217776 574614 217832
rect 576582 221992 576638 222048
rect 577318 216416 577374 216472
rect 577318 215872 577374 215928
rect 577042 215056 577098 215112
rect 575662 213560 575718 213616
rect 582194 222264 582250 222320
rect 577686 220496 577742 220552
rect 582378 220632 582434 220688
rect 591854 220632 591910 220688
rect 582194 220380 582250 220416
rect 582194 220360 582196 220380
rect 582196 220360 582248 220380
rect 582248 220360 582250 220380
rect 582378 220380 582434 220416
rect 582378 220360 582380 220380
rect 582380 220360 582432 220380
rect 582432 220360 582434 220380
rect 591854 220380 591910 220416
rect 592314 220632 592370 220688
rect 591854 220360 591856 220380
rect 591856 220360 591908 220380
rect 591908 220360 591910 220380
rect 592130 220360 592186 220416
rect 592130 219156 592186 219192
rect 592130 219136 592132 219156
rect 592132 219136 592184 219156
rect 592184 219136 592186 219156
rect 592314 219136 592370 219192
rect 582102 218320 582158 218376
rect 582286 218320 582342 218376
rect 582746 218320 582802 218376
rect 582930 218320 582986 218376
rect 591946 218320 592002 218376
rect 592130 218320 592186 218376
rect 582930 218048 582986 218104
rect 591854 218048 591910 218104
rect 582378 217776 582434 217832
rect 591670 217776 591726 217832
rect 592130 217912 592186 217968
rect 590106 217504 590162 217560
rect 582332 216960 582388 217016
rect 582378 216416 582434 216472
rect 582562 216416 582618 216472
rect 582746 216144 582802 216200
rect 591762 217232 591818 217288
rect 592222 217232 592278 217288
rect 591762 216416 591818 216472
rect 592038 216452 592040 216472
rect 592040 216452 592092 216472
rect 592092 216452 592094 216472
rect 592038 216416 592094 216452
rect 592222 216300 592278 216336
rect 592222 216280 592224 216300
rect 592224 216280 592276 216300
rect 592276 216280 592278 216300
rect 578882 213968 578938 214024
rect 578514 211676 578570 211712
rect 578514 211656 578516 211676
rect 578516 211656 578568 211676
rect 578568 211656 578570 211676
rect 579250 209788 579252 209808
rect 579252 209788 579304 209808
rect 579304 209788 579306 209808
rect 579250 209752 579306 209788
rect 599490 221720 599546 221776
rect 601514 221720 601570 221776
rect 602250 221720 602306 221776
rect 596546 219136 596602 219192
rect 597006 218864 597062 218920
rect 594798 217232 594854 217288
rect 595166 216688 595222 216744
rect 597558 216552 597614 216608
rect 595718 216280 595774 216336
rect 595902 216280 595958 216336
rect 599030 216280 599086 216336
rect 600594 221176 600650 221232
rect 600410 220632 600466 220688
rect 603078 219136 603134 219192
rect 616878 221448 616934 221504
rect 611634 220904 611690 220960
rect 610806 220224 610862 220280
rect 610806 219680 610862 219736
rect 611358 215872 611414 215928
rect 614486 218592 614542 218648
rect 617062 219952 617118 220008
rect 618902 215600 618958 215656
rect 620558 215328 620614 215384
rect 626446 218048 626502 218104
rect 630954 219680 631010 219736
rect 630770 219408 630826 219464
rect 629942 218320 629998 218376
rect 631138 218592 631194 218648
rect 652206 298424 652262 298480
rect 640246 231376 640302 231432
rect 639602 230016 639658 230072
rect 638866 219136 638922 219192
rect 640062 218864 640118 218920
rect 650642 223080 650698 223136
rect 643190 220360 643246 220416
rect 641442 220088 641498 220144
rect 642086 217232 642142 217288
rect 643006 215872 643062 215928
rect 642178 213152 642234 213208
rect 644938 217504 644994 217560
rect 646594 216144 646650 216200
rect 649906 218592 649962 218648
rect 647146 214512 647202 214568
rect 652022 222808 652078 222864
rect 651286 214784 651342 214840
rect 579526 207440 579582 207496
rect 579526 205828 579582 205864
rect 579526 205808 579528 205828
rect 579528 205808 579580 205828
rect 579580 205808 579582 205828
rect 578330 203224 578386 203280
rect 578790 200776 578846 200832
rect 660302 405592 660358 405648
rect 659106 360032 659162 360088
rect 666466 742736 666522 742792
rect 666282 705472 666338 705528
rect 667754 786664 667810 786720
rect 667570 743144 667626 743200
rect 667202 671064 667258 671120
rect 668398 783808 668454 783864
rect 668214 752256 668270 752312
rect 668214 733352 668270 733408
rect 667754 710776 667810 710832
rect 667754 688880 667810 688936
rect 667570 665896 667626 665952
rect 666466 665352 666522 665408
rect 665822 626048 665878 626104
rect 664442 579672 664498 579728
rect 662050 491952 662106 492008
rect 661866 406272 661922 406328
rect 661682 313520 661738 313576
rect 666466 603064 666522 603120
rect 668398 708736 668454 708792
rect 668398 693232 668454 693288
rect 668214 662496 668270 662552
rect 668214 654200 668270 654256
rect 667754 621152 667810 621208
rect 668950 773744 669006 773800
rect 668766 734304 668822 734360
rect 668766 731448 668822 731504
rect 668582 670520 668638 670576
rect 671158 872208 671214 872264
rect 670606 867856 670662 867912
rect 669778 864184 669834 864240
rect 669594 789384 669650 789440
rect 669226 755112 669282 755168
rect 669410 741104 669466 741160
rect 668950 709960 669006 710016
rect 669226 705064 669282 705120
rect 668766 664536 668822 664592
rect 669042 648624 669098 648680
rect 668398 620200 668454 620256
rect 668398 601704 668454 601760
rect 668214 574096 668270 574152
rect 668214 564440 668270 564496
rect 667202 534112 667258 534168
rect 666466 529896 666522 529952
rect 665822 494672 665878 494728
rect 664626 493992 664682 494048
rect 668858 593680 668914 593736
rect 668582 535880 668638 535936
rect 669042 573144 669098 573200
rect 669042 559136 669098 559192
rect 668858 528536 668914 528592
rect 668398 526496 668454 526552
rect 668214 485152 668270 485208
rect 663246 358536 663302 358592
rect 669042 483112 669098 483168
rect 669778 750896 669834 750952
rect 669778 738520 669834 738576
rect 669594 709552 669650 709608
rect 669594 695136 669650 695192
rect 669410 663584 669466 663640
rect 670330 782992 670386 783048
rect 670146 780680 670202 780736
rect 670146 710368 670202 710424
rect 670974 778640 671030 778696
rect 670606 751712 670662 751768
rect 670790 750080 670846 750136
rect 671342 763000 671398 763056
rect 673090 934632 673146 934688
rect 674194 957072 674250 957128
rect 673366 932592 673422 932648
rect 673090 930552 673146 930608
rect 675206 966048 675262 966104
rect 675758 965096 675814 965152
rect 675206 963600 675262 963656
rect 675390 963328 675446 963384
rect 674930 962512 674986 962568
rect 674654 962104 674710 962160
rect 674378 933000 674434 933056
rect 675482 962784 675538 962840
rect 675390 962104 675446 962160
rect 675206 959248 675262 959304
rect 675114 958704 675170 958760
rect 675298 957752 675354 957808
rect 675758 957752 675814 957808
rect 675482 957072 675538 957128
rect 675758 956392 675814 956448
rect 675022 954488 675078 954544
rect 674838 953400 674894 953456
rect 674654 932184 674710 932240
rect 674194 930144 674250 930200
rect 671986 928240 672042 928296
rect 671802 758648 671858 758704
rect 671526 758240 671582 758296
rect 671158 752528 671214 752584
rect 671158 737024 671214 737080
rect 671066 730496 671122 730552
rect 670790 727912 670846 727968
rect 670790 712408 670846 712464
rect 670330 707512 670386 707568
rect 670606 699760 670662 699816
rect 670330 687384 670386 687440
rect 669962 673104 670018 673160
rect 669778 666168 669834 666224
rect 669962 648080 670018 648136
rect 669778 645360 669834 645416
rect 669594 620608 669650 620664
rect 669778 574912 669834 574968
rect 669962 571648 670018 571704
rect 669410 570832 669466 570888
rect 669594 556144 669650 556200
rect 669410 500928 669466 500984
rect 669778 553832 669834 553888
rect 670974 706696 671030 706752
rect 670974 685480 671030 685536
rect 670790 667664 670846 667720
rect 671158 662360 671214 662416
rect 671158 640464 671214 640520
rect 670790 623872 670846 623928
rect 670606 619384 670662 619440
rect 670330 618160 670386 618216
rect 670606 607960 670662 608016
rect 670330 598032 670386 598088
rect 670146 537784 670202 537840
rect 669778 483520 669834 483576
rect 669594 482296 669650 482352
rect 669226 456456 669282 456512
rect 667202 360848 667258 360904
rect 665822 315424 665878 315480
rect 664442 271088 664498 271144
rect 663062 268096 663118 268152
rect 661866 234096 661922 234152
rect 658922 233824 658978 233880
rect 661682 230288 661738 230344
rect 660946 229744 661002 229800
rect 652758 226344 652814 226400
rect 658922 225528 658978 225584
rect 655518 225256 655574 225312
rect 654782 224984 654838 225040
rect 653034 220632 653090 220688
rect 654046 216416 654102 216472
rect 656622 223896 656678 223952
rect 658186 223624 658242 223680
rect 658002 221448 658058 221504
rect 659290 224440 659346 224496
rect 659474 221720 659530 221776
rect 659658 215056 659714 215112
rect 663062 231648 663118 231704
rect 664442 230832 664498 230888
rect 663706 230560 663762 230616
rect 661498 213424 661554 213480
rect 664258 220360 664314 220416
rect 664258 219680 664314 219736
rect 664258 216688 664314 216744
rect 664258 216144 664314 216200
rect 664810 213696 664866 213752
rect 665822 231104 665878 231160
rect 666650 223216 666706 223272
rect 666834 222808 666890 222864
rect 666650 221040 666706 221096
rect 589462 207984 589518 208040
rect 589462 206352 589518 206408
rect 589646 204720 589702 204776
rect 589462 203088 589518 203144
rect 589462 201456 589518 201512
rect 579526 198872 579582 198928
rect 578514 196424 578570 196480
rect 579526 194928 579582 194984
rect 579526 192208 579582 192264
rect 579526 190712 579582 190768
rect 579526 187992 579582 188048
rect 579526 186260 579528 186280
rect 579528 186260 579580 186280
rect 579580 186260 579582 186280
rect 579526 186224 579582 186260
rect 579526 184320 579582 184376
rect 579526 181872 579582 181928
rect 578790 180104 578846 180160
rect 579526 177656 579582 177712
rect 578790 175072 578846 175128
rect 578422 173440 578478 173496
rect 578238 170992 578294 171048
rect 578698 169224 578754 169280
rect 579526 166912 579582 166968
rect 578882 164464 578938 164520
rect 579526 162696 579582 162752
rect 578238 159840 578294 159896
rect 578422 158344 578478 158400
rect 578882 155896 578938 155952
rect 578330 153992 578386 154048
rect 578238 151680 578294 151736
rect 578330 149640 578386 149696
rect 578698 147228 578700 147248
rect 578700 147228 578752 147248
rect 578752 147228 578754 147248
rect 578698 147192 578754 147228
rect 578606 140528 578662 140584
rect 578606 138760 578662 138816
rect 579250 144644 579252 144664
rect 579252 144644 579304 144664
rect 579304 144644 579306 144664
rect 579250 144608 579306 144644
rect 579526 142976 579582 143032
rect 578882 136584 578938 136640
rect 578698 134408 578754 134464
rect 579066 132232 579122 132288
rect 578330 123528 578386 123584
rect 578698 118360 578754 118416
rect 578698 116864 578754 116920
rect 579066 129648 579122 129704
rect 579158 127744 579214 127800
rect 579526 125332 579528 125352
rect 579528 125332 579580 125352
rect 579580 125332 579582 125352
rect 579526 125296 579582 125332
rect 579526 121080 579582 121136
rect 579250 114452 579252 114472
rect 579252 114452 579304 114472
rect 579304 114452 579306 114472
rect 579250 114416 579306 114452
rect 579158 112512 579214 112568
rect 578882 110336 578938 110392
rect 578882 108296 578938 108352
rect 578330 103300 578332 103320
rect 578332 103300 578384 103320
rect 578384 103300 578386 103320
rect 578330 103264 578386 103300
rect 578514 101632 578570 101688
rect 578330 97416 578386 97472
rect 578330 86400 578386 86456
rect 579066 105848 579122 105904
rect 579250 99220 579252 99240
rect 579252 99220 579304 99240
rect 579304 99220 579306 99240
rect 579250 99184 579306 99220
rect 579434 95004 579436 95024
rect 579436 95004 579488 95024
rect 579488 95004 579490 95024
rect 579434 94968 579490 95004
rect 579526 93064 579582 93120
rect 579342 90888 579398 90944
rect 579526 88032 579582 88088
rect 579526 83988 579528 84008
rect 579528 83988 579580 84008
rect 579580 83988 579582 84008
rect 579526 83952 579582 83988
rect 579434 82184 579490 82240
rect 578882 80008 578938 80064
rect 578422 77832 578478 77888
rect 578330 75656 578386 75712
rect 578514 61784 578570 61840
rect 578882 60424 578938 60480
rect 589462 199824 589518 199880
rect 590382 198192 590438 198248
rect 589462 196560 589518 196616
rect 589278 194928 589334 194984
rect 589462 193296 589518 193352
rect 589462 191664 589518 191720
rect 590566 190032 590622 190088
rect 589646 188400 589702 188456
rect 589462 186768 589518 186824
rect 589462 185136 589518 185192
rect 589462 183504 589518 183560
rect 590566 181872 590622 181928
rect 589646 180240 589702 180296
rect 589462 178608 589518 178664
rect 589646 176976 589702 177032
rect 589462 175364 589518 175400
rect 589462 175344 589464 175364
rect 589464 175344 589516 175364
rect 589516 175344 589518 175364
rect 666650 176432 666706 176488
rect 589462 173712 589518 173768
rect 589462 172080 589518 172136
rect 589462 170448 589518 170504
rect 589462 168816 589518 168872
rect 589462 167184 589518 167240
rect 589462 165552 589518 165608
rect 589462 163920 589518 163976
rect 589462 162288 589518 162344
rect 589462 160656 589518 160712
rect 589830 159024 589886 159080
rect 589462 157412 589518 157448
rect 589462 157392 589464 157412
rect 589464 157392 589516 157412
rect 589516 157392 589518 157412
rect 589462 155760 589518 155816
rect 589462 154128 589518 154184
rect 589462 152496 589518 152552
rect 590014 150864 590070 150920
rect 589462 149232 589518 149288
rect 588542 147600 588598 147656
rect 579526 73108 579528 73128
rect 579528 73108 579580 73128
rect 579580 73108 579582 73128
rect 579526 73072 579582 73108
rect 579526 71204 579528 71224
rect 579528 71204 579580 71224
rect 579580 71204 579582 71224
rect 579526 71168 579582 71204
rect 579526 66292 579582 66328
rect 579526 66272 579528 66292
rect 579528 66272 579580 66292
rect 579580 66272 579582 66292
rect 579526 64504 579582 64560
rect 579526 57876 579528 57896
rect 579528 57876 579580 57896
rect 579580 57876 579582 57896
rect 579526 57840 579582 57876
rect 579526 56072 579582 56128
rect 577502 54984 577558 55040
rect 589462 145968 589518 146024
rect 589462 144336 589518 144392
rect 589830 142704 589886 142760
rect 589462 141072 589518 141128
rect 589462 139460 589518 139496
rect 589462 139440 589464 139460
rect 589464 139440 589516 139460
rect 589516 139440 589518 139460
rect 589462 137808 589518 137864
rect 589462 136176 589518 136232
rect 590290 134544 590346 134600
rect 588726 132912 588782 132968
rect 583022 77832 583078 77888
rect 588542 114960 588598 115016
rect 667018 178744 667074 178800
rect 671710 757832 671766 757888
rect 671710 757424 671766 757480
rect 671526 713632 671582 713688
rect 671526 713224 671582 713280
rect 672538 873568 672594 873624
rect 672354 784352 672410 784408
rect 672170 770616 672226 770672
rect 672170 733624 672226 733680
rect 671986 732808 672042 732864
rect 671710 712816 671766 712872
rect 671986 688608 672042 688664
rect 671618 668480 671674 668536
rect 671802 668072 671858 668128
rect 671526 667256 671582 667312
rect 671526 627816 671582 627872
rect 671802 624416 671858 624472
rect 671618 623464 671674 623520
rect 671710 623056 671766 623112
rect 671526 622648 671582 622704
rect 670790 578992 670846 579048
rect 670790 578584 670846 578640
rect 670882 577768 670938 577824
rect 671250 594768 671306 594824
rect 671066 576136 671122 576192
rect 671434 579808 671490 579864
rect 671434 579400 671490 579456
rect 673366 929464 673422 929520
rect 672998 870032 673054 870088
rect 672722 760280 672778 760336
rect 672722 759872 672778 759928
rect 672538 754160 672594 754216
rect 672538 738248 672594 738304
rect 673182 759056 673238 759112
rect 672998 755384 673054 755440
rect 672906 751304 672962 751360
rect 672354 709144 672410 709200
rect 672446 670248 672502 670304
rect 672446 668888 672502 668944
rect 672170 661544 672226 661600
rect 672814 715264 672870 715320
rect 672814 714856 672870 714912
rect 675390 953400 675446 953456
rect 675206 951360 675262 951416
rect 675850 951360 675906 951416
rect 675206 951088 675262 951144
rect 675022 934224 675078 934280
rect 677506 951496 677562 951552
rect 676218 941704 676274 941760
rect 676218 939256 676274 939312
rect 676494 938032 676550 938088
rect 676034 937760 676090 937816
rect 675206 933816 675262 933872
rect 678242 950680 678298 950736
rect 678242 935584 678298 935640
rect 683118 947280 683174 947336
rect 683118 939664 683174 939720
rect 682382 935176 682438 935232
rect 681002 933544 681058 933600
rect 677506 931096 677562 931152
rect 683118 929056 683174 929112
rect 675298 879144 675354 879200
rect 675758 875880 675814 875936
rect 675390 873976 675446 874032
rect 675390 873568 675446 873624
rect 675114 873160 675170 873216
rect 675390 872208 675446 872264
rect 674930 870848 674986 870904
rect 675114 870032 675170 870088
rect 673918 864864 673974 864920
rect 673734 779320 673790 779376
rect 673550 777416 673606 777472
rect 673366 732808 673422 732864
rect 673918 771976 673974 772032
rect 674470 788024 674526 788080
rect 674286 780000 674342 780056
rect 673918 752120 673974 752176
rect 673366 730088 673422 730144
rect 673366 728476 673422 728512
rect 673366 728456 673368 728476
rect 673368 728456 673420 728476
rect 673420 728456 673422 728476
rect 673182 714448 673238 714504
rect 672998 714040 673054 714096
rect 673182 698264 673238 698320
rect 672998 685752 673054 685808
rect 672814 669840 672870 669896
rect 672814 669432 672870 669488
rect 672630 662360 672686 662416
rect 672630 661136 672686 661192
rect 672354 638696 672410 638752
rect 672170 635432 672226 635488
rect 672170 619792 672226 619848
rect 672170 616664 672226 616720
rect 671986 614896 672042 614952
rect 671710 578176 671766 578232
rect 670790 535064 670846 535120
rect 671158 569608 671214 569664
rect 670882 533024 670938 533080
rect 671710 555192 671766 555248
rect 671434 534656 671490 534712
rect 671434 534384 671490 534440
rect 670606 528944 670662 529000
rect 670330 527720 670386 527776
rect 670882 524864 670938 524920
rect 671526 532752 671582 532808
rect 671342 490864 671398 490920
rect 671526 489232 671582 489288
rect 671710 485968 671766 486024
rect 672170 604696 672226 604752
rect 672538 604288 672594 604344
rect 673826 728184 673882 728240
rect 673826 727640 673882 727696
rect 673550 724104 673606 724160
rect 673550 689560 673606 689616
rect 673366 666440 673422 666496
rect 673366 660728 673422 660784
rect 673366 659912 673422 659968
rect 673182 622240 673238 622296
rect 672998 621560 673054 621616
rect 672906 615712 672962 615768
rect 672446 576952 672502 577008
rect 673182 577360 673238 577416
rect 672998 574504 673054 574560
rect 672906 559000 672962 559056
rect 672630 546216 672686 546272
rect 672538 533432 672594 533488
rect 672262 531392 672318 531448
rect 672170 530168 672226 530224
rect 672354 529352 672410 529408
rect 672722 531800 672778 531856
rect 673182 548392 673238 548448
rect 672722 490048 672778 490104
rect 672446 489640 672502 489696
rect 671986 455368 672042 455424
rect 672262 453736 672318 453792
rect 669962 403688 670018 403744
rect 670606 393488 670662 393544
rect 669962 347248 670018 347304
rect 668582 312840 668638 312896
rect 668306 302232 668362 302288
rect 667570 186904 667626 186960
rect 667386 181328 667442 181384
rect 667938 223896 667994 223952
rect 667938 192616 667994 192672
rect 667938 189388 667940 189408
rect 667940 189388 667992 189408
rect 667992 189388 667994 189408
rect 667938 189352 667994 189388
rect 668490 234504 668546 234560
rect 668306 229472 668362 229528
rect 668306 226344 668362 226400
rect 668306 225256 668362 225312
rect 668122 182824 668178 182880
rect 667938 174700 667940 174720
rect 667940 174700 667992 174720
rect 667992 174700 667994 174720
rect 667938 174664 667994 174700
rect 668030 169668 668032 169688
rect 668032 169668 668084 169688
rect 668084 169668 668086 169688
rect 668030 169632 668086 169668
rect 667938 164908 667940 164928
rect 667940 164908 667992 164928
rect 667992 164908 667994 164928
rect 667938 164872 667994 164908
rect 668306 163240 668362 163296
rect 668950 236680 669006 236736
rect 669410 224984 669466 225040
rect 669410 223624 669466 223680
rect 669410 214104 669466 214160
rect 669226 208256 669282 208312
rect 669226 207304 669282 207360
rect 669226 202408 669282 202464
rect 669134 199316 669136 199336
rect 669136 199316 669188 199336
rect 669188 199316 669190 199336
rect 669134 199280 669190 199316
rect 669226 198736 669282 198792
rect 669410 197104 669466 197160
rect 669134 194284 669136 194304
rect 669136 194284 669188 194304
rect 669188 194284 669190 194304
rect 669134 194248 669190 194284
rect 669134 187584 669190 187640
rect 669226 184456 669282 184512
rect 669778 168136 669834 168192
rect 669134 164192 669190 164248
rect 668950 159976 669006 160032
rect 668766 153448 668822 153504
rect 668766 149096 668822 149152
rect 668490 148552 668546 148608
rect 668582 145288 668638 145344
rect 667754 135904 667810 135960
rect 667938 135496 667994 135552
rect 667202 134544 667258 134600
rect 666834 133048 666890 133104
rect 589462 131300 589518 131336
rect 589462 131280 589464 131300
rect 589464 131280 589516 131300
rect 589516 131280 589518 131300
rect 589646 129648 589702 129704
rect 589462 128016 589518 128072
rect 668582 128288 668638 128344
rect 590106 126384 590162 126440
rect 589922 124752 589978 124808
rect 589462 123120 589518 123176
rect 589278 121508 589334 121544
rect 589278 121488 589280 121508
rect 589280 121488 589332 121508
rect 589332 121488 589334 121508
rect 589462 119856 589518 119912
rect 589462 118224 589518 118280
rect 589462 116592 589518 116648
rect 589462 113328 589518 113384
rect 589370 111696 589426 111752
rect 669134 138760 669190 138816
rect 668766 125704 668822 125760
rect 670422 256672 670478 256728
rect 670422 235864 670478 235920
rect 670330 233144 670386 233200
rect 670146 232872 670202 232928
rect 672906 488416 672962 488472
rect 672630 488008 672686 488064
rect 672446 401648 672502 401704
rect 672446 400424 672502 400480
rect 672262 393896 672318 393952
rect 672262 376216 672318 376272
rect 673182 485560 673238 485616
rect 672998 484744 673054 484800
rect 674148 727912 674204 727968
rect 675298 868400 675354 868456
rect 674838 868128 674894 868184
rect 674838 867448 674894 867504
rect 675482 867856 675538 867912
rect 675482 867448 675538 867504
rect 675390 864864 675446 864920
rect 675482 864184 675538 864240
rect 675298 863096 675354 863152
rect 674838 796864 674894 796920
rect 675206 796864 675262 796920
rect 675206 789384 675262 789440
rect 675390 788024 675446 788080
rect 674838 784080 674894 784136
rect 674838 778912 674894 778968
rect 674838 776464 674894 776520
rect 674838 775784 674894 775840
rect 675298 786664 675354 786720
rect 675390 784352 675446 784408
rect 675298 784080 675354 784136
rect 675022 774832 675078 774888
rect 674838 768168 674894 768224
rect 675482 783808 675538 783864
rect 675482 782992 675538 783048
rect 675482 780680 675538 780736
rect 675482 780000 675538 780056
rect 675482 779320 675538 779376
rect 675482 778640 675538 778696
rect 675482 777416 675538 777472
rect 675482 776464 675538 776520
rect 675482 775784 675538 775840
rect 675666 775648 675722 775704
rect 675482 773744 675538 773800
rect 682382 772656 682438 772712
rect 675206 766536 675262 766592
rect 674654 757152 674710 757208
rect 676126 768168 676182 768224
rect 676126 766536 676182 766592
rect 676034 763000 676090 763056
rect 677046 761912 677102 761968
rect 676770 761776 676826 761832
rect 676034 760688 676090 760744
rect 676034 757172 676090 757208
rect 676034 757152 676036 757172
rect 676036 757152 676088 757172
rect 676088 757152 676090 757172
rect 675850 755792 675906 755848
rect 676770 754976 676826 755032
rect 683210 771976 683266 772032
rect 683394 770888 683450 770944
rect 682382 757016 682438 757072
rect 677046 754568 677102 754624
rect 683578 770616 683634 770672
rect 683578 759464 683634 759520
rect 683302 756608 683358 756664
rect 683486 753752 683542 753808
rect 683118 752936 683174 752992
rect 675114 743144 675170 743200
rect 674930 742736 674986 742792
rect 675390 742464 675446 742520
rect 675114 741512 675170 741568
rect 674930 741104 674986 741160
rect 675114 739608 675170 739664
rect 675022 738520 675078 738576
rect 675206 738316 675262 738372
rect 675114 737024 675170 737080
rect 674286 726824 674342 726880
rect 674930 734304 674986 734360
rect 675114 733624 675170 733680
rect 675114 733352 675170 733408
rect 675114 731448 675170 731504
rect 675482 730496 675538 730552
rect 675298 730088 675354 730144
rect 674746 727640 674802 727696
rect 683486 726824 683542 726880
rect 674010 726552 674066 726608
rect 674562 726552 674618 726608
rect 682382 725736 682438 725792
rect 677322 724260 677378 724296
rect 677322 724240 677324 724260
rect 677324 724240 677376 724260
rect 677376 724240 677378 724260
rect 676034 718256 676090 718312
rect 676034 715672 676090 715728
rect 683118 725464 683174 725520
rect 682382 711592 682438 711648
rect 683118 708328 683174 708384
rect 683302 707920 683358 707976
rect 683670 726416 683726 726472
rect 683670 711184 683726 711240
rect 683486 707104 683542 707160
rect 674378 706288 674434 706344
rect 674010 692960 674066 693016
rect 673734 680992 673790 681048
rect 673734 647808 673790 647864
rect 673550 636792 673606 636848
rect 673550 625096 673606 625152
rect 673550 603472 673606 603528
rect 674194 690104 674250 690160
rect 674930 699760 674986 699816
rect 675114 698264 675170 698320
rect 675390 696768 675446 696824
rect 675114 695136 675170 695192
rect 675666 694320 675722 694376
rect 674930 693232 674986 693288
rect 675114 692960 675170 693016
rect 675390 690104 675446 690160
rect 675298 689560 675354 689616
rect 674930 688880 674986 688936
rect 675298 688880 675354 688936
rect 675114 688608 675170 688664
rect 674838 686432 674894 686488
rect 675482 687384 675538 687440
rect 675482 685752 675538 685808
rect 675206 685480 675262 685536
rect 674562 648896 674618 648952
rect 675022 651480 675078 651536
rect 674838 647536 674894 647592
rect 674470 645088 674526 645144
rect 674194 641688 674250 641744
rect 673918 617344 673974 617400
rect 674010 599528 674066 599584
rect 673642 595584 673698 595640
rect 674010 599256 674066 599312
rect 674378 624824 674434 624880
rect 674378 606464 674434 606520
rect 674010 595312 674066 595368
rect 674286 592864 674342 592920
rect 673918 591640 673974 591696
rect 683210 682624 683266 682680
rect 676494 673104 676550 673160
rect 676494 671064 676550 671120
rect 676494 670248 676550 670304
rect 676494 669432 676550 669488
rect 676494 666168 676550 666224
rect 676494 665352 676550 665408
rect 683670 682352 683726 682408
rect 683486 680992 683542 681048
rect 683210 664536 683266 664592
rect 683670 666984 683726 667040
rect 683486 662904 683542 662960
rect 675390 654200 675446 654256
rect 675574 652840 675630 652896
rect 675390 651480 675446 651536
rect 675206 650120 675262 650176
rect 675390 648896 675446 648952
rect 675482 648624 675538 648680
rect 675482 647808 675538 647864
rect 675298 647192 675354 647248
rect 675298 646040 675354 646096
rect 675482 645768 675538 645824
rect 675758 645496 675814 645552
rect 675482 645360 675538 645416
rect 675298 644272 675354 644328
rect 675758 644272 675814 644328
rect 674930 644000 674986 644056
rect 675114 643728 675170 643784
rect 675482 643456 675538 643512
rect 675298 641688 675354 641744
rect 674930 640736 674986 640792
rect 675390 640464 675446 640520
rect 674930 631352 674986 631408
rect 674746 618568 674802 618624
rect 674838 603064 674894 603120
rect 675022 601704 675078 601760
rect 674838 601024 674894 601080
rect 675022 600480 675078 600536
rect 675022 598984 675078 599040
rect 675022 596808 675078 596864
rect 675482 638696 675538 638752
rect 675390 638016 675446 638072
rect 677506 637880 677562 637936
rect 675758 637608 675814 637664
rect 674930 595448 674986 595504
rect 674654 592592 674710 592648
rect 675758 631352 675814 631408
rect 675850 627816 675906 627872
rect 676494 625640 676550 625696
rect 683394 636792 683450 636848
rect 683210 635432 683266 635488
rect 683394 624824 683450 624880
rect 683210 624416 683266 624472
rect 677506 621968 677562 622024
rect 676494 621560 676550 621616
rect 676494 621152 676550 621208
rect 683578 617888 683634 617944
rect 683394 617072 683450 617128
rect 675482 608232 675538 608288
rect 675482 607960 675538 608016
rect 675482 606464 675538 606520
rect 675482 604696 675538 604752
rect 675482 604288 675538 604344
rect 675482 603472 675538 603528
rect 675482 602792 675538 602848
rect 675482 601024 675538 601080
rect 675482 600480 675538 600536
rect 675482 599256 675538 599312
rect 675666 599120 675722 599176
rect 675482 598032 675538 598088
rect 675482 596808 675538 596864
rect 675390 595448 675446 595504
rect 675482 594768 675538 594824
rect 675390 593680 675446 593736
rect 683302 592864 683358 592920
rect 675758 592320 675814 592376
rect 675574 592048 675630 592104
rect 674194 552064 674250 552120
rect 674010 545672 674066 545728
rect 674010 535336 674066 535392
rect 674010 534112 674066 534168
rect 673826 532480 673882 532536
rect 673642 528264 673698 528320
rect 675574 586200 675630 586256
rect 676034 582936 676090 582992
rect 676034 580216 676090 580272
rect 675758 576544 675814 576600
rect 682382 575592 682438 575648
rect 683486 592592 683542 592648
rect 683762 591368 683818 591424
rect 683486 573960 683542 574016
rect 683302 573144 683358 573200
rect 683762 572328 683818 572384
rect 683118 570696 683174 570752
rect 675206 564440 675262 564496
rect 674654 558320 674710 558376
rect 674378 547032 674434 547088
rect 674470 535064 674526 535120
rect 674470 534112 674526 534168
rect 674470 532208 674526 532264
rect 674470 531392 674526 531448
rect 675390 563080 675446 563136
rect 675482 561176 675538 561232
rect 675298 559000 675354 559056
rect 675206 558728 675262 558784
rect 675390 558320 675446 558376
rect 675206 556144 675262 556200
rect 675390 555192 675446 555248
rect 675758 554648 675814 554704
rect 675390 553832 675446 553888
rect 675206 553424 675262 553480
rect 675390 552064 675446 552120
rect 675758 550704 675814 550760
rect 675390 549616 675446 549672
rect 675482 548392 675538 548448
rect 675114 547848 675170 547904
rect 674838 547304 674894 547360
rect 674838 543768 674894 543824
rect 675206 547576 675262 547632
rect 674930 503784 674986 503840
rect 675850 547304 675906 547360
rect 676402 546216 676458 546272
rect 676034 537784 676090 537840
rect 676034 535676 676090 535732
rect 675850 532480 675906 532536
rect 675758 529352 675814 529408
rect 675942 529352 675998 529408
rect 675758 528740 675814 528796
rect 675942 528536 675998 528592
rect 675022 503512 675078 503568
rect 675022 503240 675078 503296
rect 675850 503784 675906 503840
rect 676034 503532 676090 503568
rect 676034 503512 676036 503532
rect 676036 503512 676088 503532
rect 676088 503512 676090 503532
rect 676034 503240 676090 503296
rect 674930 500928 674986 500984
rect 674654 484336 674710 484392
rect 674194 483928 674250 483984
rect 674746 464752 674802 464808
rect 673826 456864 673882 456920
rect 674746 456864 674802 456920
rect 673946 456476 674002 456512
rect 673946 456456 673948 456476
rect 673948 456456 674000 456476
rect 674000 456456 674002 456476
rect 673596 455660 673652 455696
rect 673596 455640 673598 455660
rect 673598 455640 673650 455660
rect 673650 455640 673652 455660
rect 673504 455388 673560 455424
rect 673504 455368 673506 455388
rect 673506 455368 673558 455388
rect 673558 455368 673560 455388
rect 673386 455132 673388 455152
rect 673388 455132 673440 455152
rect 673440 455132 673442 455152
rect 673386 455096 673442 455132
rect 675298 486376 675354 486432
rect 673162 454844 673218 454880
rect 673162 454824 673164 454844
rect 673164 454824 673216 454844
rect 673216 454824 673218 454844
rect 674930 454824 674986 454880
rect 676586 532244 676588 532264
rect 676588 532244 676640 532264
rect 676640 532244 676642 532264
rect 676586 532208 676642 532244
rect 683210 547032 683266 547088
rect 679622 546488 679678 546544
rect 678242 531392 678298 531448
rect 683394 545672 683450 545728
rect 683210 531800 683266 531856
rect 679622 530984 679678 531040
rect 683578 532208 683634 532264
rect 683394 527720 683450 527776
rect 683578 526496 683634 526552
rect 676862 525680 676918 525736
rect 677874 524456 677930 524512
rect 683210 503648 683266 503704
rect 676034 493992 676090 494048
rect 673044 454588 673046 454608
rect 673046 454588 673098 454608
rect 673098 454588 673100 454608
rect 673044 454552 673100 454588
rect 675482 454552 675538 454608
rect 675850 481888 675906 481944
rect 672952 454316 672954 454336
rect 672954 454316 673006 454336
rect 673006 454316 673008 454336
rect 672952 454280 673008 454316
rect 675666 454280 675722 454336
rect 672814 454044 672816 454064
rect 672816 454044 672868 454064
rect 672868 454044 672870 454064
rect 672814 454008 672870 454044
rect 676034 480664 676090 480720
rect 677322 492360 677378 492416
rect 676954 488824 677010 488880
rect 677322 487192 677378 487248
rect 681002 487600 681058 487656
rect 679622 486784 679678 486840
rect 676954 485732 677010 485788
rect 683578 494672 683634 494728
rect 683394 491680 683450 491736
rect 683578 491272 683634 491328
rect 683210 482704 683266 482760
rect 682382 481480 682438 481536
rect 676770 455640 676826 455696
rect 676034 454008 676090 454064
rect 675850 453736 675906 453792
rect 683118 406272 683174 406328
rect 676034 405592 676090 405648
rect 676034 403416 676090 403472
rect 683118 403280 683174 403336
rect 674194 402192 674250 402248
rect 672630 400016 672686 400072
rect 673182 398792 673238 398848
rect 672998 397160 673054 397216
rect 672722 392536 672778 392592
rect 672446 355816 672502 355872
rect 672538 354592 672594 354648
rect 672170 353368 672226 353424
rect 671986 348880 672042 348936
rect 672354 348472 672410 348528
rect 672170 340720 672226 340776
rect 671986 332288 672042 332344
rect 672170 311208 672226 311264
rect 671986 301960 672042 302016
rect 671342 269728 671398 269784
rect 671342 264016 671398 264072
rect 671710 261976 671766 262032
rect 671526 257896 671582 257952
rect 671710 244704 671766 244760
rect 671526 241440 671582 241496
rect 671342 238176 671398 238232
rect 671158 233144 671214 233200
rect 671066 225664 671122 225720
rect 671066 225276 671122 225312
rect 671066 225256 671068 225276
rect 671068 225256 671120 225276
rect 671120 225256 671122 225276
rect 671066 224884 671068 224904
rect 671068 224884 671120 224904
rect 671120 224884 671122 224904
rect 671066 224848 671122 224884
rect 671020 224460 671076 224496
rect 671020 224440 671022 224460
rect 671022 224440 671074 224460
rect 671074 224440 671076 224460
rect 670606 211112 670662 211168
rect 670606 210840 670662 210896
rect 670606 190304 670662 190360
rect 670606 170312 670662 170368
rect 670330 165552 670386 165608
rect 669962 122712 670018 122768
rect 668582 120808 668638 120864
rect 668950 120128 669006 120184
rect 667938 119176 667994 119232
rect 668030 117544 668086 117600
rect 668950 114280 669006 114336
rect 671802 231376 671858 231432
rect 672170 266464 672226 266520
rect 672170 234504 672226 234560
rect 672538 309984 672594 310040
rect 672998 377984 673054 378040
rect 673366 396344 673422 396400
rect 673826 396072 673882 396128
rect 673366 382200 673422 382256
rect 674010 395664 674066 395720
rect 673826 381384 673882 381440
rect 674010 375400 674066 375456
rect 673182 355408 673238 355464
rect 672998 351328 673054 351384
rect 672998 338000 673054 338056
rect 674654 401376 674710 401432
rect 674470 394440 674526 394496
rect 674470 377712 674526 377768
rect 676034 399336 676090 399392
rect 676218 398384 676274 398440
rect 676402 397976 676458 398032
rect 681002 397568 681058 397624
rect 681002 387640 681058 387696
rect 675758 384920 675814 384976
rect 675390 382200 675446 382256
rect 675114 381384 675170 381440
rect 675758 380568 675814 380624
rect 675758 378664 675814 378720
rect 675114 377712 675170 377768
rect 675758 377304 675814 377360
rect 675206 376896 675262 376952
rect 675390 376216 675446 376272
rect 675390 375400 675446 375456
rect 675758 372952 675814 373008
rect 675114 372544 675170 372600
rect 674194 357448 674250 357504
rect 675850 360848 675906 360904
rect 676034 360032 676090 360088
rect 676034 358264 676090 358320
rect 675850 357856 675906 357912
rect 674654 357040 674710 357096
rect 674470 356632 674526 356688
rect 674102 356224 674158 356280
rect 673366 355000 673422 355056
rect 673918 352552 673974 352608
rect 673550 352144 673606 352200
rect 673366 349696 673422 349752
rect 673366 335824 673422 335880
rect 673734 350512 673790 350568
rect 673918 336640 673974 336696
rect 673734 331064 673790 331120
rect 673550 325624 673606 325680
rect 673918 312024 673974 312080
rect 673182 310800 673238 310856
rect 673366 304680 673422 304736
rect 672998 304272 673054 304328
rect 673734 303864 673790 303920
rect 673366 290536 673422 290592
rect 672998 287816 673054 287872
rect 673734 286456 673790 286512
rect 674470 349424 674526 349480
rect 674286 347656 674342 347712
rect 676034 353776 676090 353832
rect 675942 349152 675998 349208
rect 675114 340720 675170 340776
rect 675758 340312 675814 340368
rect 675390 338952 675446 339008
rect 674470 332832 674526 332888
rect 674286 327528 674342 327584
rect 675114 338000 675170 338056
rect 675574 337728 675630 337784
rect 675114 336640 675170 336696
rect 675758 336640 675814 336696
rect 675482 335824 675538 335880
rect 675390 332832 675446 332888
rect 675114 332288 675170 332344
rect 675758 332152 675814 332208
rect 675114 331064 675170 331120
rect 675758 328344 675814 328400
rect 675114 327528 675170 327584
rect 675114 325624 675170 325680
rect 676034 315424 676090 315480
rect 676034 313248 676090 313304
rect 674654 312432 674710 312488
rect 674102 311616 674158 311672
rect 674194 310392 674250 310448
rect 673918 267416 673974 267472
rect 674010 266192 674066 266248
rect 673090 263744 673146 263800
rect 672906 259120 672962 259176
rect 673366 260344 673422 260400
rect 672814 242800 672870 242856
rect 672262 228792 672318 228848
rect 673182 257080 673238 257136
rect 672998 237360 673054 237416
rect 673734 259664 673790 259720
rect 674562 309576 674618 309632
rect 674378 305496 674434 305552
rect 674838 309168 674894 309224
rect 676034 308352 676090 308408
rect 681002 307536 681058 307592
rect 678242 307128 678298 307184
rect 676402 305904 676458 305960
rect 674838 303592 674894 303648
rect 675390 303592 675446 303648
rect 675114 301688 675170 301744
rect 674838 296792 674894 296848
rect 674378 292576 674434 292632
rect 674654 292304 674710 292360
rect 675022 296520 675078 296576
rect 676034 303456 676090 303512
rect 676034 301960 676090 302016
rect 676586 305088 676642 305144
rect 676586 301552 676642 301608
rect 676402 301416 676458 301472
rect 678978 306312 679034 306368
rect 678242 297336 678298 297392
rect 676126 296792 676182 296848
rect 675850 296520 675906 296576
rect 675574 296248 675630 296304
rect 675482 295840 675538 295896
rect 675758 295160 675814 295216
rect 675758 291488 675814 291544
rect 675114 290536 675170 290592
rect 675114 287816 675170 287872
rect 675758 287000 675814 287056
rect 675390 286456 675446 286512
rect 675758 283600 675814 283656
rect 675666 282784 675722 282840
rect 675666 281560 675722 281616
rect 674194 265784 674250 265840
rect 674286 265376 674342 265432
rect 683118 271088 683174 271144
rect 676034 269728 676090 269784
rect 676034 268232 676090 268288
rect 683118 268096 683174 268152
rect 674654 267008 674710 267064
rect 674470 264968 674526 265024
rect 674194 260888 674250 260944
rect 673918 258440 673974 258496
rect 673734 245520 673790 245576
rect 673366 244976 673422 245032
rect 674286 246880 674342 246936
rect 673302 237108 673358 237144
rect 673302 237088 673304 237108
rect 673304 237088 673356 237108
rect 673356 237088 673358 237108
rect 673526 236700 673582 236736
rect 673526 236680 673528 236700
rect 673528 236680 673580 236700
rect 673580 236680 673582 236700
rect 672906 228520 672962 228576
rect 674194 235592 674250 235648
rect 673918 232872 673974 232928
rect 674470 234912 674526 234968
rect 674010 230580 674066 230616
rect 674010 230560 674012 230580
rect 674012 230560 674064 230580
rect 674064 230560 674066 230580
rect 673826 230016 673882 230072
rect 673458 229744 673514 229800
rect 673946 229916 673948 229936
rect 673948 229916 674000 229936
rect 674000 229916 674002 229936
rect 673946 229880 674002 229916
rect 674170 230152 674226 230208
rect 674838 264424 674894 264480
rect 676494 264016 676550 264072
rect 674838 263744 674894 263800
rect 676494 263608 676550 263664
rect 678242 263200 678298 263256
rect 676218 262792 676274 262848
rect 675298 257488 675354 257544
rect 675298 256672 675354 256728
rect 675942 258712 675998 258768
rect 675942 258168 675998 258224
rect 674930 251504 674986 251560
rect 674930 249328 674986 249384
rect 678426 261160 678482 261216
rect 675850 251540 675852 251560
rect 675852 251540 675904 251560
rect 675904 251540 675906 251560
rect 675850 251504 675906 251540
rect 675758 250280 675814 250336
rect 675390 249600 675446 249656
rect 675114 246880 675170 246936
rect 675114 245520 675170 245576
rect 674838 245248 674894 245304
rect 675390 242800 675446 242856
rect 675114 241440 675170 241496
rect 675206 240216 675262 240272
rect 675114 238176 675170 238232
rect 674838 237360 674894 237416
rect 675390 236816 675446 236872
rect 675114 235864 675170 235920
rect 675666 235456 675722 235512
rect 674838 235184 674894 235240
rect 674654 234368 674710 234424
rect 676034 235184 676090 235240
rect 675850 234912 675906 234968
rect 675850 234388 675906 234424
rect 675850 234368 675852 234388
rect 675852 234368 675904 234388
rect 675904 234368 675906 234388
rect 675178 231804 675234 231840
rect 675178 231784 675180 231804
rect 675180 231784 675232 231804
rect 675232 231784 675234 231804
rect 675068 231548 675070 231568
rect 675070 231548 675122 231568
rect 675122 231548 675124 231568
rect 675068 231512 675124 231548
rect 674838 231140 674840 231160
rect 674840 231140 674892 231160
rect 674892 231140 674894 231160
rect 674838 231104 674894 231140
rect 674730 230868 674732 230888
rect 674732 230868 674784 230888
rect 674784 230868 674786 230888
rect 674730 230832 674786 230868
rect 674838 230696 674894 230752
rect 675850 230696 675906 230752
rect 674746 230424 674802 230480
rect 674194 229608 674250 229664
rect 673458 229356 673514 229392
rect 673458 229336 673460 229356
rect 673460 229336 673512 229356
rect 673512 229336 673514 229356
rect 673596 229084 673652 229120
rect 673596 229064 673598 229084
rect 673598 229064 673650 229084
rect 673650 229064 673652 229084
rect 673504 228828 673506 228848
rect 673506 228828 673558 228848
rect 673558 228828 673560 228848
rect 673504 228792 673560 228828
rect 673386 228540 673442 228576
rect 673386 228520 673388 228540
rect 673388 228520 673440 228540
rect 673440 228520 673442 228540
rect 672446 227024 672502 227080
rect 672602 227060 672604 227080
rect 672604 227060 672656 227080
rect 672656 227060 672658 227080
rect 672602 227024 672658 227060
rect 672378 226772 672434 226808
rect 672378 226752 672380 226772
rect 672380 226752 672432 226772
rect 672432 226752 672434 226772
rect 672032 226244 672034 226264
rect 672034 226244 672086 226264
rect 672086 226244 672088 226264
rect 672032 226208 672088 226244
rect 671802 225936 671858 225992
rect 671818 225700 671820 225720
rect 671820 225700 671872 225720
rect 671872 225700 671874 225720
rect 671818 225664 671874 225700
rect 672078 222944 672134 223000
rect 671802 221448 671858 221504
rect 671986 220088 672042 220144
rect 671894 219408 671950 219464
rect 672078 214784 672134 214840
rect 672814 226480 672870 226536
rect 672538 225528 672594 225584
rect 672722 224848 672778 224904
rect 672538 224576 672594 224632
rect 672722 216280 672778 216336
rect 672538 214784 672594 214840
rect 672170 213696 672226 213752
rect 672722 210160 672778 210216
rect 672170 200776 672226 200832
rect 672538 198736 672594 198792
rect 672078 183504 672134 183560
rect 671894 174800 671950 174856
rect 671894 166912 671950 166968
rect 671710 158344 671766 158400
rect 671526 150184 671582 150240
rect 670606 147600 670662 147656
rect 671342 131688 671398 131744
rect 671526 130872 671582 130928
rect 668122 112648 668178 112704
rect 668582 111832 668638 111888
rect 590106 110064 590162 110120
rect 589462 108432 589518 108488
rect 589462 106800 589518 106856
rect 589462 105168 589518 105224
rect 589554 103536 589610 103592
rect 589922 101904 589978 101960
rect 666650 109316 666706 109372
rect 668122 106120 668178 106176
rect 668398 106156 668400 106176
rect 668400 106156 668452 106176
rect 668452 106156 668454 106176
rect 668398 106120 668454 106156
rect 589922 77288 589978 77344
rect 585782 54712 585838 54768
rect 613382 95784 613438 95840
rect 635738 96056 635794 96112
rect 637026 96872 637082 96928
rect 646226 95548 646228 95568
rect 646228 95548 646280 95568
rect 646280 95548 646282 95568
rect 646226 95512 646282 95548
rect 647330 94968 647386 95024
rect 626446 94424 626502 94480
rect 625986 93608 626042 93664
rect 626446 92792 626502 92848
rect 625802 91976 625858 92032
rect 626446 91160 626502 91216
rect 626446 90344 626502 90400
rect 626262 89528 626318 89584
rect 626446 88712 626502 88768
rect 626446 87896 626502 87952
rect 626262 87080 626318 87136
rect 626446 86300 626448 86320
rect 626448 86300 626500 86320
rect 626500 86300 626502 86320
rect 626446 86264 626502 86300
rect 626446 85484 626448 85504
rect 626448 85484 626500 85504
rect 626500 85484 626502 85504
rect 626446 85448 626502 85484
rect 625250 84632 625306 84688
rect 604458 54440 604514 54496
rect 576858 54168 576914 54224
rect 459834 53624 459890 53680
rect 460754 53624 460810 53680
rect 461674 53624 461730 53680
rect 462594 53624 462650 53680
rect 464342 53644 464398 53680
rect 464342 53624 464344 53644
rect 464344 53624 464396 53644
rect 464396 53624 464398 53644
rect 482282 53644 482338 53680
rect 482282 53624 482284 53644
rect 482284 53624 482336 53644
rect 482336 53624 482338 53644
rect 472530 53352 472586 53408
rect 481730 53352 481786 53408
rect 308034 50224 308090 50280
rect 458178 46960 458234 47016
rect 458362 46688 458418 46744
rect 431222 44784 431278 44840
rect 142618 44240 142674 44296
rect 307298 44104 307354 44160
rect 194322 42064 194378 42120
rect 361762 43560 361818 43616
rect 416594 42336 416650 42392
rect 415766 42064 415822 42120
rect 419906 41792 419962 41848
rect 446402 42200 446458 42256
rect 446402 41520 446458 41576
rect 460110 44784 460166 44840
rect 460846 43832 460902 43888
rect 461950 44376 462006 44432
rect 462502 44376 462558 44432
rect 462318 43152 462374 43208
rect 461766 42880 461822 42936
rect 463882 44104 463938 44160
rect 544014 47504 544070 47560
rect 549994 48864 550050 48920
rect 553674 50224 553730 50280
rect 552018 48048 552074 48104
rect 547878 47776 547934 47832
rect 545670 47232 545726 47288
rect 465262 46960 465318 47016
rect 465078 46688 465134 46744
rect 625802 83816 625858 83872
rect 628746 83272 628802 83328
rect 647698 95512 647754 95568
rect 648618 91976 648674 92032
rect 647514 82728 647570 82784
rect 629206 81640 629262 81696
rect 633898 78512 633954 78568
rect 633898 77288 633954 77344
rect 639602 77832 639658 77888
rect 646410 74432 646466 74488
rect 646226 69128 646282 69184
rect 646226 67088 646282 67144
rect 647238 71712 647294 71768
rect 648710 62056 648766 62112
rect 646410 59336 646466 59392
rect 650458 89528 650514 89584
rect 650182 87080 650238 87136
rect 651838 90616 651894 90672
rect 655058 94152 655114 94208
rect 654598 93336 654654 93392
rect 655426 92520 655482 92576
rect 655242 91432 655298 91488
rect 655794 89800 655850 89856
rect 663706 92792 663762 92848
rect 664534 91704 664590 91760
rect 664350 90616 664406 90672
rect 664166 89800 664222 89856
rect 665362 93336 665418 93392
rect 665178 88984 665234 89040
rect 650734 84632 650790 84688
rect 649078 64368 649134 64424
rect 648894 57296 648950 57352
rect 661590 47733 661646 47789
rect 667938 102720 667994 102776
rect 672262 182008 672318 182064
rect 672538 175208 672594 175264
rect 672262 164192 672318 164248
rect 672078 140392 672134 140448
rect 672538 130464 672594 130520
rect 673458 227024 673514 227080
rect 673550 225256 673606 225312
rect 673550 220632 673606 220688
rect 673550 220224 673606 220280
rect 673550 218592 673606 218648
rect 673458 216144 673514 216200
rect 673550 206896 673606 206952
rect 673366 201864 673422 201920
rect 673274 201592 673330 201648
rect 673550 197648 673606 197704
rect 672998 177928 673054 177984
rect 673366 174392 673422 174448
rect 672906 173032 672962 173088
rect 673182 169904 673238 169960
rect 672998 169088 673054 169144
rect 672998 153040 673054 153096
rect 673182 151680 673238 151736
rect 673918 227024 673974 227080
rect 674102 226208 674158 226264
rect 674102 220224 674158 220280
rect 676770 230424 676826 230480
rect 676586 230152 676642 230208
rect 675114 229608 675170 229664
rect 675114 229336 675170 229392
rect 675114 229064 675170 229120
rect 675114 228792 675170 228848
rect 675390 226752 675446 226808
rect 675022 226480 675078 226536
rect 674838 224304 674894 224360
rect 674838 222128 674894 222184
rect 674654 221856 674710 221912
rect 673918 212880 673974 212936
rect 673918 209616 673974 209672
rect 673918 203496 673974 203552
rect 675206 225528 675262 225584
rect 675022 219680 675078 219736
rect 674838 219000 674894 219056
rect 674102 179424 674158 179480
rect 675022 217776 675078 217832
rect 674746 216552 674802 216608
rect 674562 215328 674618 215384
rect 674378 177248 674434 177304
rect 674286 176840 674342 176896
rect 673918 176024 673974 176080
rect 673734 168408 673790 168464
rect 674102 169496 674158 169552
rect 674102 155352 674158 155408
rect 674746 204992 674802 205048
rect 675206 216824 675262 216880
rect 675206 215328 675262 215384
rect 674930 204448 674986 204504
rect 674838 204176 674894 204232
rect 676034 220668 676036 220688
rect 676036 220668 676088 220688
rect 676088 220668 676090 220688
rect 676034 220632 676090 220668
rect 676034 220360 676090 220416
rect 675666 218320 675722 218376
rect 675942 215092 675944 215112
rect 675944 215092 675996 215112
rect 675996 215092 675998 215112
rect 675942 215056 675998 215092
rect 675666 214512 675722 214568
rect 676034 213424 676090 213480
rect 676034 213152 676090 213208
rect 676862 209616 676918 209672
rect 675850 208256 675906 208312
rect 679254 223760 679310 223816
rect 683854 234096 683910 234152
rect 683302 233824 683358 233880
rect 683302 223080 683358 223136
rect 679990 222264 680046 222320
rect 679806 221448 679862 221504
rect 679622 220632 679678 220688
rect 683854 222672 683910 222728
rect 683486 219816 683542 219872
rect 683302 213288 683358 213344
rect 683118 212472 683174 212528
rect 683118 211112 683174 211168
rect 683302 210296 683358 210352
rect 677782 206896 677838 206952
rect 675758 205536 675814 205592
rect 675482 204992 675538 205048
rect 675482 204448 675538 204504
rect 675298 204176 675354 204232
rect 675482 201864 675538 201920
rect 675298 200776 675354 200832
rect 675114 197920 675170 197976
rect 675758 200640 675814 200696
rect 675574 198192 675630 198248
rect 675482 197104 675538 197160
rect 675758 197104 675814 197160
rect 675666 193160 675722 193216
rect 675758 191528 675814 191584
rect 675298 190304 675354 190360
rect 683118 186904 683174 186960
rect 676494 181328 676550 181384
rect 676034 178064 676090 178120
rect 683118 178744 683174 178800
rect 674562 175616 674618 175672
rect 678242 173168 678298 173224
rect 674838 172760 674894 172816
rect 674470 168680 674526 168736
rect 676586 170720 676642 170776
rect 676034 167864 676090 167920
rect 676586 166368 676642 166424
rect 676034 165552 676090 165608
rect 681002 171536 681058 171592
rect 679622 171128 679678 171184
rect 675942 161880 675998 161936
rect 676126 161336 676182 161392
rect 675758 160656 675814 160712
rect 675758 159296 675814 159352
rect 674838 157528 674894 157584
rect 675482 157528 675538 157584
rect 675390 156984 675446 157040
rect 675758 156304 675814 156360
rect 675114 155352 675170 155408
rect 675114 153040 675170 153096
rect 675758 153040 675814 153096
rect 675114 151680 675170 151736
rect 675666 148416 675722 148472
rect 675114 147600 675170 147656
rect 675666 147600 675722 147656
rect 675758 145968 675814 146024
rect 683118 135904 683174 135960
rect 675850 134544 675906 134600
rect 676494 133048 676550 133104
rect 683118 132640 683174 132696
rect 674286 132096 674342 132152
rect 673918 131280 673974 131336
rect 675942 130056 675998 130112
rect 673366 129648 673422 129704
rect 674102 129240 674158 129296
rect 673090 125976 673146 126032
rect 672906 124344 672962 124400
rect 672722 124072 672778 124128
rect 672538 123800 672594 123856
rect 672354 123120 672410 123176
rect 672354 120128 672410 120184
rect 671894 115776 671950 115832
rect 671526 107752 671582 107808
rect 672722 117816 672778 117872
rect 673366 123528 673422 123584
rect 673090 111424 673146 111480
rect 672722 111016 672778 111072
rect 672538 110200 672594 110256
rect 672354 106392 672410 106448
rect 673918 121624 673974 121680
rect 673918 117816 673974 117872
rect 674286 128288 674342 128344
rect 675942 128288 675998 128344
rect 674102 111832 674158 111888
rect 673366 105576 673422 105632
rect 668582 104488 668638 104544
rect 682382 127744 682438 127800
rect 674838 127608 674894 127664
rect 674654 125568 674710 125624
rect 674470 125160 674526 125216
rect 675022 126384 675078 126440
rect 675298 113056 675354 113112
rect 675114 111424 675170 111480
rect 674654 110200 674710 110256
rect 675666 108024 675722 108080
rect 675114 106392 675170 106448
rect 675758 106120 675814 106176
rect 675114 105576 675170 105632
rect 675758 103128 675814 103184
rect 675666 102584 675722 102640
rect 674286 102312 674342 102368
rect 675758 101360 675814 101416
rect 668306 95784 668362 95840
rect 663798 48456 663854 48512
rect 662418 47368 662474 47424
rect 471058 43832 471114 43888
rect 464342 43560 464398 43616
rect 465814 43152 465870 43208
rect 463698 42880 463754 42936
rect 461122 42200 461178 42256
rect 518806 42744 518862 42800
rect 515402 42064 515458 42120
rect 520922 42064 520978 42120
rect 522026 42064 522082 42120
rect 526442 42064 526498 42120
rect 529570 42064 529626 42120
rect 141698 40432 141754 40488
<< metal3 >>
rect 426341 1007178 426407 1007181
rect 426341 1007176 426604 1007178
rect 426341 1007120 426346 1007176
rect 426402 1007120 426604 1007176
rect 426341 1007118 426604 1007120
rect 426341 1007115 426407 1007118
rect 358537 1007042 358603 1007045
rect 553945 1007042 554011 1007045
rect 358537 1007040 358800 1007042
rect 358537 1006984 358542 1007040
rect 358598 1006984 358800 1007040
rect 358537 1006982 358800 1006984
rect 553748 1007040 554011 1007042
rect 553748 1006984 553950 1007040
rect 554006 1006984 554011 1007040
rect 553748 1006982 554011 1006984
rect 358537 1006979 358603 1006982
rect 553945 1006979 554011 1006982
rect 359365 1006906 359431 1006909
rect 505001 1006906 505067 1006909
rect 359168 1006904 359431 1006906
rect 359168 1006848 359370 1006904
rect 359426 1006848 359431 1006904
rect 359168 1006846 359431 1006848
rect 504804 1006904 505067 1006906
rect 504804 1006848 505006 1006904
rect 505062 1006848 505067 1006904
rect 504804 1006846 505067 1006848
rect 359365 1006843 359431 1006846
rect 505001 1006843 505067 1006846
rect 555969 1006906 556035 1006909
rect 555969 1006904 556232 1006906
rect 555969 1006848 555974 1006904
rect 556030 1006848 556232 1006904
rect 555969 1006846 556232 1006848
rect 555969 1006843 556035 1006846
rect 360193 1006770 360259 1006773
rect 429193 1006770 429259 1006773
rect 507853 1006770 507919 1006773
rect 556797 1006770 556863 1006773
rect 359996 1006768 360259 1006770
rect 359996 1006712 360198 1006768
rect 360254 1006712 360259 1006768
rect 359996 1006710 360259 1006712
rect 428996 1006768 429259 1006770
rect 428996 1006712 429198 1006768
rect 429254 1006712 429259 1006768
rect 428996 1006710 429259 1006712
rect 507656 1006768 507919 1006770
rect 507656 1006712 507858 1006768
rect 507914 1006712 507919 1006768
rect 507656 1006710 507919 1006712
rect 556600 1006768 556863 1006770
rect 556600 1006712 556802 1006768
rect 556858 1006712 556863 1006768
rect 556600 1006710 556863 1006712
rect 360193 1006707 360259 1006710
rect 429193 1006707 429259 1006710
rect 507853 1006707 507919 1006710
rect 556797 1006707 556863 1006710
rect 101949 1006634 102015 1006637
rect 153745 1006634 153811 1006637
rect 157425 1006634 157491 1006637
rect 101949 1006632 102212 1006634
rect 101949 1006576 101954 1006632
rect 102010 1006576 102212 1006632
rect 101949 1006574 102212 1006576
rect 153548 1006632 153811 1006634
rect 153548 1006576 153750 1006632
rect 153806 1006576 153811 1006632
rect 153548 1006574 153811 1006576
rect 157228 1006632 157491 1006634
rect 157228 1006576 157430 1006632
rect 157486 1006576 157491 1006632
rect 157228 1006574 157491 1006576
rect 101949 1006571 102015 1006574
rect 153745 1006571 153811 1006574
rect 157425 1006571 157491 1006574
rect 431677 1006634 431743 1006637
rect 505369 1006634 505435 1006637
rect 431677 1006632 431940 1006634
rect 431677 1006576 431682 1006632
rect 431738 1006576 431940 1006632
rect 431677 1006574 431940 1006576
rect 505172 1006632 505435 1006634
rect 505172 1006576 505374 1006632
rect 505430 1006576 505435 1006632
rect 505172 1006574 505435 1006576
rect 431677 1006571 431743 1006574
rect 505369 1006571 505435 1006574
rect 98269 1006498 98335 1006501
rect 152917 1006498 152983 1006501
rect 160277 1006498 160343 1006501
rect 256141 1006498 256207 1006501
rect 98269 1006496 98532 1006498
rect 98269 1006440 98274 1006496
rect 98330 1006468 98532 1006496
rect 152720 1006496 152983 1006498
rect 98330 1006440 98562 1006468
rect 98269 1006438 98562 1006440
rect 152720 1006440 152922 1006496
rect 152978 1006440 152983 1006496
rect 152720 1006438 152983 1006440
rect 160080 1006496 160343 1006498
rect 160080 1006440 160282 1006496
rect 160338 1006440 160343 1006496
rect 160080 1006438 160343 1006440
rect 255944 1006496 256207 1006498
rect 255944 1006440 256146 1006496
rect 256202 1006440 256207 1006496
rect 255944 1006438 256207 1006440
rect 98269 1006435 98335 1006438
rect 98502 1006090 98562 1006438
rect 152917 1006435 152983 1006438
rect 160277 1006435 160343 1006438
rect 256141 1006435 256207 1006438
rect 354857 1006498 354923 1006501
rect 428365 1006498 428431 1006501
rect 506197 1006498 506263 1006501
rect 354857 1006496 355120 1006498
rect 354857 1006440 354862 1006496
rect 354918 1006468 355120 1006496
rect 428365 1006496 428628 1006498
rect 354918 1006440 355150 1006468
rect 354857 1006438 355150 1006440
rect 354857 1006435 354923 1006438
rect 103973 1006362 104039 1006365
rect 108481 1006362 108547 1006365
rect 103973 1006360 104236 1006362
rect 103973 1006304 103978 1006360
rect 104034 1006304 104236 1006360
rect 103973 1006302 104236 1006304
rect 108284 1006360 108547 1006362
rect 108284 1006304 108486 1006360
rect 108542 1006304 108547 1006360
rect 108284 1006302 108547 1006304
rect 103973 1006299 104039 1006302
rect 108481 1006299 108547 1006302
rect 152089 1006362 152155 1006365
rect 158253 1006362 158319 1006365
rect 152089 1006360 152352 1006362
rect 152089 1006304 152094 1006360
rect 152150 1006304 152352 1006360
rect 152089 1006302 152352 1006304
rect 158056 1006360 158319 1006362
rect 158056 1006304 158258 1006360
rect 158314 1006304 158319 1006360
rect 158056 1006302 158319 1006304
rect 152089 1006299 152155 1006302
rect 158253 1006299 158319 1006302
rect 258993 1006362 259059 1006365
rect 307753 1006362 307819 1006365
rect 314653 1006362 314719 1006365
rect 258993 1006360 259164 1006362
rect 258993 1006304 258998 1006360
rect 259054 1006304 259164 1006360
rect 258993 1006302 259164 1006304
rect 307753 1006360 307924 1006362
rect 307753 1006304 307758 1006360
rect 307814 1006304 307924 1006360
rect 307753 1006302 307924 1006304
rect 314653 1006360 314916 1006362
rect 314653 1006304 314658 1006360
rect 314714 1006304 314916 1006360
rect 314653 1006302 314916 1006304
rect 258993 1006299 259059 1006302
rect 307753 1006299 307819 1006302
rect 314653 1006299 314719 1006302
rect 104801 1006226 104867 1006229
rect 106825 1006226 106891 1006229
rect 104604 1006224 104867 1006226
rect 104604 1006168 104806 1006224
rect 104862 1006168 104867 1006224
rect 104604 1006166 104867 1006168
rect 106628 1006224 106891 1006226
rect 106628 1006168 106830 1006224
rect 106886 1006168 106891 1006224
rect 106628 1006166 106891 1006168
rect 104801 1006163 104867 1006166
rect 106825 1006163 106891 1006166
rect 151261 1006226 151327 1006229
rect 158621 1006226 158687 1006229
rect 210417 1006226 210483 1006229
rect 151261 1006224 151524 1006226
rect 151261 1006168 151266 1006224
rect 151322 1006168 151524 1006224
rect 151261 1006166 151524 1006168
rect 158621 1006224 158884 1006226
rect 158621 1006168 158626 1006224
rect 158682 1006168 158884 1006224
rect 158621 1006166 158884 1006168
rect 210220 1006224 210483 1006226
rect 210220 1006168 210422 1006224
rect 210478 1006168 210483 1006224
rect 210220 1006166 210483 1006168
rect 151261 1006163 151327 1006166
rect 158621 1006163 158687 1006166
rect 210417 1006163 210483 1006166
rect 257337 1006226 257403 1006229
rect 262673 1006226 262739 1006229
rect 257337 1006224 257600 1006226
rect 257337 1006168 257342 1006224
rect 257398 1006168 257600 1006224
rect 257337 1006166 257600 1006168
rect 262476 1006224 262739 1006226
rect 262476 1006168 262678 1006224
rect 262734 1006168 262739 1006224
rect 262476 1006166 262739 1006168
rect 257337 1006163 257403 1006166
rect 262673 1006163 262739 1006166
rect 304901 1006226 304967 1006229
rect 304901 1006224 305164 1006226
rect 304901 1006168 304906 1006224
rect 304962 1006168 305164 1006224
rect 304901 1006166 305164 1006168
rect 304901 1006163 304967 1006166
rect 99465 1006090 99531 1006093
rect 103145 1006090 103211 1006093
rect 105997 1006090 106063 1006093
rect 98502 1006060 98900 1006090
rect 98532 1006030 98900 1006060
rect 99465 1006088 99728 1006090
rect 99465 1006032 99470 1006088
rect 99526 1006032 99728 1006088
rect 99465 1006030 99728 1006032
rect 103145 1006088 103408 1006090
rect 103145 1006032 103150 1006088
rect 103206 1006032 103408 1006088
rect 103145 1006030 103408 1006032
rect 105892 1006088 106063 1006090
rect 105892 1006032 106002 1006088
rect 106058 1006032 106063 1006088
rect 105892 1006030 106063 1006032
rect 99465 1006027 99531 1006030
rect 103145 1006027 103211 1006030
rect 105997 1006027 106063 1006030
rect 147121 1006090 147187 1006093
rect 148869 1006090 148935 1006093
rect 150065 1006090 150131 1006093
rect 158253 1006090 158319 1006093
rect 159449 1006090 159515 1006093
rect 201033 1006090 201099 1006093
rect 208393 1006090 208459 1006093
rect 252461 1006090 252527 1006093
rect 258165 1006090 258231 1006093
rect 261845 1006090 261911 1006093
rect 147121 1006088 148935 1006090
rect 147121 1006032 147126 1006088
rect 147182 1006032 148874 1006088
rect 148930 1006032 148935 1006088
rect 147121 1006030 148935 1006032
rect 149868 1006088 150328 1006090
rect 149868 1006032 150070 1006088
rect 150126 1006032 150328 1006088
rect 149868 1006030 150328 1006032
rect 158253 1006088 158516 1006090
rect 158253 1006032 158258 1006088
rect 158314 1006032 158516 1006088
rect 158253 1006030 158516 1006032
rect 159449 1006088 159712 1006090
rect 159449 1006032 159454 1006088
rect 159510 1006032 159712 1006088
rect 159449 1006030 159712 1006032
rect 201033 1006088 201756 1006090
rect 201033 1006032 201038 1006088
rect 201094 1006032 201756 1006088
rect 201033 1006030 201756 1006032
rect 208393 1006088 208656 1006090
rect 208393 1006032 208398 1006088
rect 208454 1006032 208656 1006088
rect 208393 1006030 208656 1006032
rect 252461 1006088 253092 1006090
rect 252461 1006032 252466 1006088
rect 252522 1006032 253092 1006088
rect 252461 1006030 253092 1006032
rect 258165 1006088 258428 1006090
rect 258165 1006032 258170 1006088
rect 258226 1006032 258428 1006088
rect 258165 1006030 258428 1006032
rect 261648 1006088 261911 1006090
rect 261648 1006032 261850 1006088
rect 261906 1006032 261911 1006088
rect 261648 1006030 261911 1006032
rect 147121 1006027 147187 1006030
rect 148869 1006027 148935 1006030
rect 150065 1006027 150131 1006030
rect 158253 1006027 158319 1006030
rect 159449 1006027 159515 1006030
rect 201033 1006027 201099 1006030
rect 208393 1006027 208459 1006030
rect 252461 1006027 252527 1006030
rect 258165 1006027 258231 1006030
rect 261845 1006027 261911 1006030
rect 301681 1006090 301747 1006093
rect 303245 1006090 303311 1006093
rect 301681 1006088 303311 1006090
rect 301681 1006032 301686 1006088
rect 301742 1006032 303250 1006088
rect 303306 1006032 303311 1006088
rect 301681 1006030 303311 1006032
rect 301681 1006027 301747 1006030
rect 303245 1006027 303311 1006030
rect 304073 1006090 304139 1006093
rect 311801 1006090 311867 1006093
rect 314653 1006090 314719 1006093
rect 355090 1006090 355150 1006438
rect 428365 1006440 428370 1006496
rect 428426 1006440 428628 1006496
rect 428365 1006438 428628 1006440
rect 506000 1006496 506263 1006498
rect 506000 1006440 506202 1006496
rect 506258 1006440 506263 1006496
rect 506000 1006438 506263 1006440
rect 428365 1006435 428431 1006438
rect 506197 1006435 506263 1006438
rect 555141 1006498 555207 1006501
rect 555141 1006496 555404 1006498
rect 555141 1006440 555146 1006496
rect 555202 1006440 555404 1006496
rect 555141 1006438 555404 1006440
rect 555141 1006435 555207 1006438
rect 361389 1006362 361455 1006365
rect 427537 1006362 427603 1006365
rect 361192 1006360 361455 1006362
rect 361192 1006304 361394 1006360
rect 361450 1006304 361455 1006360
rect 361192 1006302 361455 1006304
rect 427340 1006360 427603 1006362
rect 427340 1006304 427542 1006360
rect 427598 1006304 427603 1006360
rect 427340 1006302 427603 1006304
rect 361389 1006299 361455 1006302
rect 427537 1006299 427603 1006302
rect 551461 1006362 551527 1006365
rect 551461 1006360 551724 1006362
rect 551461 1006304 551466 1006360
rect 551522 1006304 551724 1006360
rect 551461 1006302 551724 1006304
rect 551461 1006299 551527 1006302
rect 360561 1006226 360627 1006229
rect 363413 1006226 363479 1006229
rect 360561 1006224 360824 1006226
rect 360561 1006168 360566 1006224
rect 360622 1006168 360824 1006224
rect 360561 1006166 360824 1006168
rect 363308 1006224 363479 1006226
rect 363308 1006168 363418 1006224
rect 363474 1006168 363479 1006224
rect 363308 1006166 363479 1006168
rect 360561 1006163 360627 1006166
rect 363413 1006163 363479 1006166
rect 429193 1006226 429259 1006229
rect 558821 1006226 558887 1006229
rect 429193 1006224 429456 1006226
rect 429193 1006168 429198 1006224
rect 429254 1006168 429456 1006224
rect 429193 1006166 429456 1006168
rect 558624 1006224 558887 1006226
rect 558624 1006168 558826 1006224
rect 558882 1006168 558887 1006224
rect 558624 1006166 558887 1006168
rect 429193 1006163 429259 1006166
rect 558821 1006163 558887 1006166
rect 358537 1006090 358603 1006093
rect 365069 1006090 365135 1006093
rect 304073 1006088 304704 1006090
rect 304073 1006032 304078 1006088
rect 304134 1006032 304704 1006088
rect 304073 1006030 304704 1006032
rect 311801 1006088 312064 1006090
rect 311801 1006032 311806 1006088
rect 311862 1006032 312064 1006088
rect 311801 1006030 312064 1006032
rect 314548 1006088 314719 1006090
rect 314548 1006032 314658 1006088
rect 314714 1006032 314719 1006088
rect 314548 1006030 314719 1006032
rect 354660 1006060 355150 1006090
rect 358340 1006088 358603 1006090
rect 354660 1006030 355120 1006060
rect 358340 1006032 358542 1006088
rect 358598 1006032 358603 1006088
rect 358340 1006030 358603 1006032
rect 364872 1006088 365135 1006090
rect 364872 1006032 365074 1006088
rect 365130 1006032 365135 1006088
rect 364872 1006030 365135 1006032
rect 304073 1006027 304139 1006030
rect 311801 1006027 311867 1006030
rect 314653 1006027 314719 1006030
rect 358537 1006027 358603 1006030
rect 365069 1006027 365135 1006030
rect 421833 1006090 421899 1006093
rect 425145 1006090 425211 1006093
rect 431677 1006090 431743 1006093
rect 421833 1006088 422556 1006090
rect 421833 1006032 421838 1006088
rect 421894 1006032 422556 1006088
rect 421833 1006030 422556 1006032
rect 424948 1006088 425211 1006090
rect 424948 1006032 425150 1006088
rect 425206 1006032 425211 1006088
rect 424948 1006030 425211 1006032
rect 431480 1006088 431743 1006090
rect 431480 1006032 431682 1006088
rect 431738 1006032 431743 1006088
rect 431480 1006030 431743 1006032
rect 421833 1006027 421899 1006030
rect 425145 1006027 425211 1006030
rect 431677 1006027 431743 1006030
rect 498837 1006090 498903 1006093
rect 550265 1006090 550331 1006093
rect 554773 1006090 554839 1006093
rect 498837 1006088 499468 1006090
rect 498837 1006032 498842 1006088
rect 498898 1006032 499468 1006088
rect 498837 1006030 499468 1006032
rect 550265 1006088 550896 1006090
rect 550265 1006032 550270 1006088
rect 550326 1006032 550896 1006088
rect 550265 1006030 550896 1006032
rect 554576 1006088 554839 1006090
rect 554576 1006032 554778 1006088
rect 554834 1006032 554839 1006088
rect 554576 1006030 554839 1006032
rect 498837 1006027 498903 1006030
rect 550265 1006027 550331 1006030
rect 554773 1006027 554839 1006030
rect 428365 1005818 428431 1005821
rect 428260 1005816 428431 1005818
rect 428260 1005760 428370 1005816
rect 428426 1005760 428431 1005816
rect 428260 1005758 428431 1005760
rect 428365 1005755 428431 1005758
rect 423489 1005682 423555 1005685
rect 423489 1005680 423752 1005682
rect 423489 1005624 423494 1005680
rect 423550 1005624 423752 1005680
rect 423489 1005622 423752 1005624
rect 423489 1005619 423555 1005622
rect 360561 1005410 360627 1005413
rect 423489 1005410 423555 1005413
rect 427169 1005410 427235 1005413
rect 360364 1005408 360627 1005410
rect 360364 1005352 360566 1005408
rect 360622 1005352 360627 1005408
rect 360364 1005350 360627 1005352
rect 423292 1005408 423555 1005410
rect 423292 1005352 423494 1005408
rect 423550 1005352 423555 1005408
rect 423292 1005350 423555 1005352
rect 426972 1005408 427235 1005410
rect 426972 1005352 427174 1005408
rect 427230 1005352 427235 1005408
rect 426972 1005350 427235 1005352
rect 360561 1005347 360627 1005350
rect 423489 1005347 423555 1005350
rect 427169 1005347 427235 1005350
rect 500493 1005410 500559 1005413
rect 500493 1005408 500756 1005410
rect 500493 1005352 500498 1005408
rect 500554 1005352 500756 1005408
rect 500493 1005350 500756 1005352
rect 500493 1005347 500559 1005350
rect 108849 1005274 108915 1005277
rect 212073 1005274 212139 1005277
rect 108849 1005272 109112 1005274
rect 108849 1005216 108854 1005272
rect 108910 1005216 109112 1005272
rect 108849 1005214 109112 1005216
rect 211876 1005272 212139 1005274
rect 211876 1005216 212078 1005272
rect 212134 1005216 212139 1005272
rect 211876 1005214 212139 1005216
rect 108849 1005211 108915 1005214
rect 212073 1005211 212139 1005214
rect 307293 1005274 307359 1005277
rect 355685 1005274 355751 1005277
rect 498837 1005274 498903 1005277
rect 551461 1005274 551527 1005277
rect 307293 1005272 307556 1005274
rect 307293 1005216 307298 1005272
rect 307354 1005216 307556 1005272
rect 307293 1005214 307556 1005216
rect 355685 1005272 355948 1005274
rect 355685 1005216 355690 1005272
rect 355746 1005216 355948 1005272
rect 355685 1005214 355948 1005216
rect 498732 1005272 498903 1005274
rect 498732 1005216 498842 1005272
rect 498898 1005216 498903 1005272
rect 498732 1005214 498903 1005216
rect 551356 1005272 551527 1005274
rect 551356 1005216 551466 1005272
rect 551522 1005216 551527 1005272
rect 551356 1005214 551527 1005216
rect 307293 1005211 307359 1005214
rect 355685 1005211 355751 1005214
rect 498837 1005211 498903 1005214
rect 551461 1005211 551527 1005214
rect 153745 1005138 153811 1005141
rect 365069 1005138 365135 1005141
rect 425513 1005138 425579 1005141
rect 153745 1005136 153916 1005138
rect 153745 1005080 153750 1005136
rect 153806 1005080 153916 1005136
rect 153745 1005078 153916 1005080
rect 365069 1005136 365332 1005138
rect 365069 1005080 365074 1005136
rect 365130 1005080 365332 1005136
rect 365069 1005078 365332 1005080
rect 425513 1005136 425776 1005138
rect 425513 1005080 425518 1005136
rect 425574 1005080 425776 1005136
rect 425513 1005078 425776 1005080
rect 153745 1005075 153811 1005078
rect 365069 1005075 365135 1005078
rect 425513 1005075 425579 1005078
rect 152917 1005002 152983 1005005
rect 209221 1005002 209287 1005005
rect 263041 1005002 263107 1005005
rect 152917 1005000 153180 1005002
rect 152917 1004944 152922 1005000
rect 152978 1004944 153180 1005000
rect 152917 1004942 153180 1004944
rect 209221 1005000 209484 1005002
rect 209221 1004944 209226 1005000
rect 209282 1004944 209484 1005000
rect 209221 1004942 209484 1004944
rect 262844 1005000 263107 1005002
rect 262844 1004944 263046 1005000
rect 263102 1004944 263107 1005000
rect 262844 1004942 263107 1004944
rect 152917 1004939 152983 1004942
rect 209221 1004939 209287 1004942
rect 263041 1004939 263107 1004942
rect 306925 1005002 306991 1005005
rect 356513 1005002 356579 1005005
rect 306925 1005000 307188 1005002
rect 306925 1004944 306930 1005000
rect 306986 1004944 307188 1005000
rect 306925 1004942 307188 1004944
rect 356316 1005000 356579 1005002
rect 356316 1004944 356518 1005000
rect 356574 1004944 356579 1005000
rect 356316 1004942 356579 1004944
rect 306925 1004939 306991 1004942
rect 356513 1004939 356579 1004942
rect 361389 1005002 361455 1005005
rect 427997 1005002 428063 1005005
rect 500493 1005002 500559 1005005
rect 557165 1005002 557231 1005005
rect 361389 1005000 361652 1005002
rect 361389 1004944 361394 1005000
rect 361450 1004944 361652 1005000
rect 361389 1004942 361652 1004944
rect 427800 1005000 428063 1005002
rect 427800 1004944 428002 1005000
rect 428058 1004944 428063 1005000
rect 427800 1004942 428063 1004944
rect 500296 1005000 500559 1005002
rect 500296 1004944 500498 1005000
rect 500554 1004944 500559 1005000
rect 500296 1004942 500559 1004944
rect 557060 1005000 557231 1005002
rect 557060 1004944 557170 1005000
rect 557226 1004944 557231 1005000
rect 557060 1004942 557231 1004944
rect 361389 1004939 361455 1004942
rect 427997 1004939 428063 1004942
rect 500493 1004939 500559 1004942
rect 557165 1004939 557231 1004942
rect 154113 1004866 154179 1004869
rect 160645 1004866 160711 1004869
rect 154113 1004864 154376 1004866
rect 154113 1004808 154118 1004864
rect 154174 1004808 154376 1004864
rect 154113 1004806 154376 1004808
rect 160540 1004864 160711 1004866
rect 160540 1004808 160650 1004864
rect 160706 1004808 160711 1004864
rect 160540 1004806 160711 1004808
rect 154113 1004803 154179 1004806
rect 160645 1004803 160711 1004806
rect 211245 1004866 211311 1004869
rect 258165 1004866 258231 1004869
rect 308949 1004866 309015 1004869
rect 313825 1004866 313891 1004869
rect 355685 1004866 355751 1004869
rect 362585 1004866 362651 1004869
rect 211245 1004864 211508 1004866
rect 211245 1004808 211250 1004864
rect 211306 1004808 211508 1004864
rect 211245 1004806 211508 1004808
rect 257968 1004864 258231 1004866
rect 257968 1004808 258170 1004864
rect 258226 1004808 258231 1004864
rect 257968 1004806 258231 1004808
rect 308752 1004864 309015 1004866
rect 308752 1004808 308954 1004864
rect 309010 1004808 309015 1004864
rect 308752 1004806 309015 1004808
rect 313628 1004864 313891 1004866
rect 313628 1004808 313830 1004864
rect 313886 1004808 313891 1004864
rect 313628 1004806 313891 1004808
rect 355488 1004864 355751 1004866
rect 355488 1004808 355690 1004864
rect 355746 1004808 355751 1004864
rect 355488 1004806 355751 1004808
rect 362388 1004864 362651 1004866
rect 362388 1004808 362590 1004864
rect 362646 1004808 362651 1004864
rect 362388 1004806 362651 1004808
rect 211245 1004803 211311 1004806
rect 258165 1004803 258231 1004806
rect 308949 1004803 309015 1004806
rect 313825 1004803 313891 1004806
rect 355685 1004803 355751 1004806
rect 362585 1004803 362651 1004806
rect 422661 1004866 422727 1004869
rect 499665 1004866 499731 1004869
rect 555969 1004866 556035 1004869
rect 422661 1004864 422924 1004866
rect 422661 1004808 422666 1004864
rect 422722 1004808 422924 1004864
rect 422661 1004806 422924 1004808
rect 499665 1004864 499928 1004866
rect 499665 1004808 499670 1004864
rect 499726 1004808 499928 1004864
rect 499665 1004806 499928 1004808
rect 555772 1004864 556035 1004866
rect 555772 1004808 555974 1004864
rect 556030 1004808 556035 1004864
rect 555772 1004806 556035 1004808
rect 422661 1004803 422727 1004806
rect 499665 1004803 499731 1004806
rect 555969 1004803 556035 1004806
rect 108481 1004730 108547 1004733
rect 151721 1004730 151787 1004733
rect 161105 1004730 161171 1004733
rect 209221 1004730 209287 1004733
rect 108481 1004728 108652 1004730
rect 108481 1004672 108486 1004728
rect 108542 1004672 108652 1004728
rect 108481 1004670 108652 1004672
rect 151721 1004728 151892 1004730
rect 151721 1004672 151726 1004728
rect 151782 1004672 151892 1004728
rect 151721 1004670 151892 1004672
rect 160908 1004728 161171 1004730
rect 160908 1004672 161110 1004728
rect 161166 1004672 161171 1004728
rect 160908 1004670 161171 1004672
rect 209024 1004728 209287 1004730
rect 209024 1004672 209226 1004728
rect 209282 1004672 209287 1004728
rect 209024 1004670 209287 1004672
rect 108481 1004667 108547 1004670
rect 151721 1004667 151787 1004670
rect 161105 1004667 161171 1004670
rect 209221 1004667 209287 1004670
rect 308121 1004730 308187 1004733
rect 315481 1004730 315547 1004733
rect 364241 1004730 364307 1004733
rect 432873 1004730 432939 1004733
rect 557625 1004730 557691 1004733
rect 308121 1004728 308384 1004730
rect 308121 1004672 308126 1004728
rect 308182 1004672 308384 1004728
rect 308121 1004670 308384 1004672
rect 315284 1004728 315547 1004730
rect 315284 1004672 315486 1004728
rect 315542 1004672 315547 1004728
rect 315284 1004670 315547 1004672
rect 364044 1004728 364307 1004730
rect 364044 1004672 364246 1004728
rect 364302 1004672 364307 1004728
rect 364044 1004670 364307 1004672
rect 432676 1004728 432939 1004730
rect 432676 1004672 432878 1004728
rect 432934 1004672 432939 1004728
rect 432676 1004670 432939 1004672
rect 557428 1004728 557691 1004730
rect 557428 1004672 557630 1004728
rect 557686 1004672 557691 1004728
rect 557428 1004670 557691 1004672
rect 308121 1004667 308187 1004670
rect 315481 1004667 315547 1004670
rect 364241 1004667 364307 1004670
rect 432873 1004667 432939 1004670
rect 557625 1004667 557691 1004670
rect 560845 1004730 560911 1004733
rect 560845 1004728 561108 1004730
rect 560845 1004672 560850 1004728
rect 560906 1004672 561108 1004728
rect 560845 1004670 561108 1004672
rect 560845 1004667 560911 1004670
rect 255313 1003914 255379 1003917
rect 424317 1003914 424383 1003917
rect 255116 1003912 255379 1003914
rect 255116 1003856 255318 1003912
rect 255374 1003856 255379 1003912
rect 255116 1003854 255379 1003856
rect 424120 1003912 424383 1003914
rect 424120 1003856 424322 1003912
rect 424378 1003856 424383 1003912
rect 424120 1003854 424383 1003856
rect 255313 1003851 255379 1003854
rect 424317 1003851 424383 1003854
rect 305269 1003370 305335 1003373
rect 554773 1003370 554839 1003373
rect 305269 1003368 305532 1003370
rect 305269 1003312 305274 1003368
rect 305330 1003312 305532 1003368
rect 305269 1003310 305532 1003312
rect 554773 1003368 555036 1003370
rect 554773 1003312 554778 1003368
rect 554834 1003312 555036 1003368
rect 554773 1003310 555036 1003312
rect 305269 1003307 305335 1003310
rect 554773 1003307 554839 1003310
rect 308949 1003234 309015 1003237
rect 308949 1003232 309212 1003234
rect 308949 1003176 308954 1003232
rect 309010 1003176 309212 1003232
rect 308949 1003174 309212 1003176
rect 308949 1003171 309015 1003174
rect 100293 1002690 100359 1002693
rect 256141 1002690 256207 1002693
rect 424685 1002690 424751 1002693
rect 100293 1002688 100556 1002690
rect 100293 1002632 100298 1002688
rect 100354 1002632 100556 1002688
rect 100293 1002630 100556 1002632
rect 256141 1002688 256404 1002690
rect 256141 1002632 256146 1002688
rect 256202 1002632 256404 1002688
rect 256141 1002630 256404 1002632
rect 424580 1002688 424751 1002690
rect 424580 1002632 424690 1002688
rect 424746 1002632 424751 1002688
rect 424580 1002630 424751 1002632
rect 100293 1002627 100359 1002630
rect 256141 1002627 256207 1002630
rect 424685 1002627 424751 1002630
rect 553117 1002690 553183 1002693
rect 558821 1002690 558887 1002693
rect 553117 1002688 553380 1002690
rect 553117 1002632 553122 1002688
rect 553178 1002632 553380 1002688
rect 553117 1002630 553380 1002632
rect 558821 1002688 559084 1002690
rect 558821 1002632 558826 1002688
rect 558882 1002632 559084 1002688
rect 558821 1002630 559084 1002632
rect 553117 1002627 553183 1002630
rect 558821 1002627 558887 1002630
rect 101949 1002554 102015 1002557
rect 206369 1002554 206435 1002557
rect 101752 1002552 102015 1002554
rect 101752 1002496 101954 1002552
rect 102010 1002496 102015 1002552
rect 101752 1002494 102015 1002496
rect 206172 1002552 206435 1002554
rect 206172 1002496 206374 1002552
rect 206430 1002496 206435 1002552
rect 206172 1002494 206435 1002496
rect 101949 1002491 102015 1002494
rect 206369 1002491 206435 1002494
rect 254117 1002554 254183 1002557
rect 310605 1002554 310671 1002557
rect 509877 1002554 509943 1002557
rect 560845 1002554 560911 1002557
rect 254117 1002552 254380 1002554
rect 254117 1002496 254122 1002552
rect 254178 1002496 254380 1002552
rect 254117 1002494 254380 1002496
rect 310408 1002552 310671 1002554
rect 310408 1002496 310610 1002552
rect 310666 1002496 310671 1002552
rect 310408 1002494 310671 1002496
rect 509680 1002552 509943 1002554
rect 509680 1002496 509882 1002552
rect 509938 1002496 509943 1002552
rect 509680 1002494 509943 1002496
rect 560740 1002552 560911 1002554
rect 560740 1002496 560850 1002552
rect 560906 1002496 560911 1002552
rect 560740 1002494 560911 1002496
rect 254117 1002491 254183 1002494
rect 310605 1002491 310671 1002494
rect 509877 1002491 509943 1002494
rect 560845 1002491 560911 1002494
rect 100293 1002418 100359 1002421
rect 103145 1002418 103211 1002421
rect 107653 1002418 107719 1002421
rect 100096 1002416 100359 1002418
rect 100096 1002360 100298 1002416
rect 100354 1002360 100359 1002416
rect 100096 1002358 100359 1002360
rect 102948 1002416 103211 1002418
rect 102948 1002360 103150 1002416
rect 103206 1002360 103211 1002416
rect 102948 1002358 103211 1002360
rect 107456 1002416 107719 1002418
rect 107456 1002360 107658 1002416
rect 107714 1002360 107719 1002416
rect 107456 1002358 107719 1002360
rect 100293 1002355 100359 1002358
rect 103145 1002355 103211 1002358
rect 107653 1002355 107719 1002358
rect 150893 1002418 150959 1002421
rect 254485 1002418 254551 1002421
rect 261017 1002418 261083 1002421
rect 357709 1002418 357775 1002421
rect 501689 1002418 501755 1002421
rect 560477 1002418 560543 1002421
rect 150893 1002416 151156 1002418
rect 150893 1002360 150898 1002416
rect 150954 1002360 151156 1002416
rect 150893 1002358 151156 1002360
rect 254485 1002416 254748 1002418
rect 254485 1002360 254490 1002416
rect 254546 1002360 254748 1002416
rect 254485 1002358 254748 1002360
rect 260820 1002416 261083 1002418
rect 260820 1002360 261022 1002416
rect 261078 1002360 261083 1002416
rect 260820 1002358 261083 1002360
rect 357604 1002416 357775 1002418
rect 357604 1002360 357714 1002416
rect 357770 1002360 357775 1002416
rect 357604 1002358 357775 1002360
rect 501492 1002416 501755 1002418
rect 501492 1002360 501694 1002416
rect 501750 1002360 501755 1002416
rect 501492 1002358 501755 1002360
rect 560280 1002416 560543 1002418
rect 560280 1002360 560482 1002416
rect 560538 1002360 560543 1002416
rect 560280 1002358 560543 1002360
rect 150893 1002355 150959 1002358
rect 254485 1002355 254551 1002358
rect 261017 1002355 261083 1002358
rect 357709 1002355 357775 1002358
rect 501689 1002355 501755 1002358
rect 560477 1002355 560543 1002358
rect 101121 1002282 101187 1002285
rect 105629 1002282 105695 1002285
rect 108021 1002282 108087 1002285
rect 155769 1002282 155835 1002285
rect 100924 1002280 101187 1002282
rect 100924 1002224 101126 1002280
rect 101182 1002224 101187 1002280
rect 100924 1002222 101187 1002224
rect 105432 1002280 105695 1002282
rect 105432 1002224 105634 1002280
rect 105690 1002224 105695 1002280
rect 105432 1002222 105695 1002224
rect 107916 1002280 108087 1002282
rect 107916 1002224 108026 1002280
rect 108082 1002224 108087 1002280
rect 107916 1002222 108087 1002224
rect 155572 1002280 155835 1002282
rect 155572 1002224 155774 1002280
rect 155830 1002224 155835 1002280
rect 155572 1002222 155835 1002224
rect 101121 1002219 101187 1002222
rect 105629 1002219 105695 1002222
rect 108021 1002219 108087 1002222
rect 155769 1002219 155835 1002222
rect 207197 1002282 207263 1002285
rect 256509 1002282 256575 1002285
rect 260189 1002282 260255 1002285
rect 207197 1002280 207460 1002282
rect 207197 1002224 207202 1002280
rect 207258 1002224 207460 1002280
rect 207197 1002222 207460 1002224
rect 256509 1002280 256772 1002282
rect 256509 1002224 256514 1002280
rect 256570 1002224 256772 1002280
rect 256509 1002222 256772 1002224
rect 260084 1002280 260255 1002282
rect 260084 1002224 260194 1002280
rect 260250 1002224 260255 1002280
rect 260084 1002222 260255 1002224
rect 207197 1002219 207263 1002222
rect 256509 1002219 256575 1002222
rect 260189 1002219 260255 1002222
rect 298277 1002282 298343 1002285
rect 303245 1002282 303311 1002285
rect 298277 1002280 303311 1002282
rect 298277 1002224 298282 1002280
rect 298338 1002224 303250 1002280
rect 303306 1002224 303311 1002280
rect 298277 1002222 303311 1002224
rect 298277 1002219 298343 1002222
rect 303245 1002219 303311 1002222
rect 306097 1002282 306163 1002285
rect 310605 1002282 310671 1002285
rect 503345 1002282 503411 1002285
rect 504173 1002282 504239 1002285
rect 306097 1002280 306360 1002282
rect 306097 1002224 306102 1002280
rect 306158 1002224 306360 1002280
rect 306097 1002222 306360 1002224
rect 310605 1002280 310868 1002282
rect 310605 1002224 310610 1002280
rect 310666 1002224 310868 1002280
rect 310605 1002222 310868 1002224
rect 503148 1002280 503411 1002282
rect 503148 1002224 503350 1002280
rect 503406 1002224 503411 1002280
rect 503148 1002222 503411 1002224
rect 503976 1002280 504239 1002282
rect 503976 1002224 504178 1002280
rect 504234 1002224 504239 1002280
rect 503976 1002222 504239 1002224
rect 306097 1002219 306163 1002222
rect 310605 1002219 310671 1002222
rect 503345 1002219 503411 1002222
rect 504173 1002219 504239 1002222
rect 557993 1002282 558059 1002285
rect 557993 1002280 558256 1002282
rect 557993 1002224 557998 1002280
rect 558054 1002224 558256 1002280
rect 557993 1002222 558256 1002224
rect 557993 1002219 558059 1002222
rect 99097 1002146 99163 1002149
rect 102317 1002146 102383 1002149
rect 103973 1002146 104039 1002149
rect 99097 1002144 99268 1002146
rect 99097 1002088 99102 1002144
rect 99158 1002088 99268 1002144
rect 99097 1002086 99268 1002088
rect 102317 1002144 102580 1002146
rect 102317 1002088 102322 1002144
rect 102378 1002088 102580 1002144
rect 102317 1002086 102580 1002088
rect 103776 1002144 104039 1002146
rect 103776 1002088 103978 1002144
rect 104034 1002088 104039 1002144
rect 103776 1002086 104039 1002088
rect 99097 1002083 99163 1002086
rect 102317 1002083 102383 1002086
rect 103973 1002083 104039 1002086
rect 106825 1002146 106891 1002149
rect 109677 1002146 109743 1002149
rect 150893 1002146 150959 1002149
rect 106825 1002144 107088 1002146
rect 106825 1002088 106830 1002144
rect 106886 1002088 107088 1002144
rect 106825 1002086 107088 1002088
rect 109480 1002144 109743 1002146
rect 109480 1002088 109682 1002144
rect 109738 1002088 109743 1002144
rect 109480 1002086 109743 1002088
rect 150696 1002144 150959 1002146
rect 150696 1002088 150898 1002144
rect 150954 1002088 150959 1002144
rect 150696 1002086 150959 1002088
rect 106825 1002083 106891 1002086
rect 109677 1002083 109743 1002086
rect 150893 1002083 150959 1002086
rect 154573 1002146 154639 1002149
rect 157793 1002146 157859 1002149
rect 206737 1002146 206803 1002149
rect 154573 1002144 154836 1002146
rect 154573 1002088 154578 1002144
rect 154634 1002088 154836 1002144
rect 154573 1002086 154836 1002088
rect 157596 1002144 157859 1002146
rect 157596 1002088 157798 1002144
rect 157854 1002088 157859 1002144
rect 157596 1002086 157859 1002088
rect 206540 1002144 206803 1002146
rect 206540 1002088 206742 1002144
rect 206798 1002088 206803 1002144
rect 206540 1002086 206803 1002088
rect 154573 1002083 154639 1002086
rect 157793 1002083 157859 1002086
rect 206737 1002083 206803 1002086
rect 210877 1002146 210943 1002149
rect 255313 1002146 255379 1002149
rect 259821 1002146 259887 1002149
rect 263869 1002146 263935 1002149
rect 304073 1002146 304139 1002149
rect 210877 1002144 211140 1002146
rect 210877 1002088 210882 1002144
rect 210938 1002088 211140 1002144
rect 210877 1002086 211140 1002088
rect 255313 1002144 255576 1002146
rect 255313 1002088 255318 1002144
rect 255374 1002088 255576 1002144
rect 255313 1002086 255576 1002088
rect 259624 1002144 259887 1002146
rect 259624 1002088 259826 1002144
rect 259882 1002088 259887 1002144
rect 259624 1002086 259887 1002088
rect 263764 1002144 263935 1002146
rect 263764 1002088 263874 1002144
rect 263930 1002088 263935 1002144
rect 263764 1002086 263935 1002088
rect 303876 1002144 304139 1002146
rect 303876 1002088 304078 1002144
rect 304134 1002088 304139 1002144
rect 303876 1002086 304139 1002088
rect 210877 1002083 210943 1002086
rect 255313 1002083 255379 1002086
rect 259821 1002083 259887 1002086
rect 263869 1002083 263935 1002086
rect 304073 1002083 304139 1002086
rect 357709 1002146 357775 1002149
rect 426341 1002146 426407 1002149
rect 357709 1002144 357972 1002146
rect 357709 1002088 357714 1002144
rect 357770 1002088 357972 1002144
rect 357709 1002086 357972 1002088
rect 426144 1002144 426407 1002146
rect 426144 1002088 426346 1002144
rect 426402 1002088 426407 1002144
rect 426144 1002086 426407 1002088
rect 357709 1002083 357775 1002086
rect 426341 1002083 426407 1002086
rect 501689 1002146 501755 1002149
rect 502517 1002146 502583 1002149
rect 553945 1002146 554011 1002149
rect 560017 1002146 560083 1002149
rect 501689 1002144 501952 1002146
rect 501689 1002088 501694 1002144
rect 501750 1002088 501952 1002144
rect 501689 1002086 501952 1002088
rect 502517 1002144 502780 1002146
rect 502517 1002088 502522 1002144
rect 502578 1002088 502780 1002144
rect 502517 1002086 502780 1002088
rect 553945 1002144 554116 1002146
rect 553945 1002088 553950 1002144
rect 554006 1002088 554116 1002144
rect 553945 1002086 554116 1002088
rect 559820 1002144 560083 1002146
rect 559820 1002088 560022 1002144
rect 560078 1002088 560083 1002144
rect 559820 1002086 560083 1002088
rect 501689 1002083 501755 1002086
rect 502517 1002083 502583 1002086
rect 553945 1002083 554011 1002086
rect 560017 1002083 560083 1002086
rect 98269 1002010 98335 1002013
rect 98072 1002008 98335 1002010
rect 98072 1001952 98274 1002008
rect 98330 1001952 98335 1002008
rect 98072 1001950 98335 1001952
rect 98269 1001947 98335 1001950
rect 101121 1002010 101187 1002013
rect 104801 1002010 104867 1002013
rect 105997 1002010 106063 1002013
rect 149237 1002010 149303 1002013
rect 154941 1002010 155007 1002013
rect 155769 1002010 155835 1002013
rect 156597 1002010 156663 1002013
rect 101121 1002008 101292 1002010
rect 101121 1001952 101126 1002008
rect 101182 1001952 101292 1002008
rect 101121 1001950 101292 1001952
rect 104801 1002008 104972 1002010
rect 104801 1001952 104806 1002008
rect 104862 1001952 104972 1002008
rect 104801 1001950 104972 1001952
rect 105997 1002008 106260 1002010
rect 105997 1001952 106002 1002008
rect 106058 1001952 106260 1002008
rect 105997 1001950 106260 1001952
rect 149237 1002008 149500 1002010
rect 149237 1001952 149242 1002008
rect 149298 1001952 149500 1002008
rect 149237 1001950 149500 1001952
rect 154941 1002008 155204 1002010
rect 154941 1001952 154946 1002008
rect 155002 1001952 155204 1002008
rect 154941 1001950 155204 1001952
rect 155769 1002008 156032 1002010
rect 155769 1001952 155774 1002008
rect 155830 1001952 156032 1002008
rect 155769 1001950 156032 1001952
rect 156400 1002008 156663 1002010
rect 156400 1001952 156602 1002008
rect 156658 1001952 156663 1002008
rect 156400 1001950 156663 1001952
rect 101121 1001947 101187 1001950
rect 104801 1001947 104867 1001950
rect 105997 1001947 106063 1001950
rect 149237 1001947 149303 1001950
rect 154941 1001947 155007 1001950
rect 155769 1001947 155835 1001950
rect 156597 1001947 156663 1001950
rect 205541 1002010 205607 1002013
rect 207197 1002010 207263 1002013
rect 205541 1002008 205804 1002010
rect 205541 1001952 205546 1002008
rect 205602 1001952 205804 1002008
rect 205541 1001950 205804 1001952
rect 207000 1002008 207263 1002010
rect 207000 1001952 207202 1002008
rect 207258 1001952 207263 1002008
rect 207000 1001950 207263 1001952
rect 205541 1001947 205607 1001950
rect 207197 1001947 207263 1001950
rect 207565 1002010 207631 1002013
rect 212533 1002010 212599 1002013
rect 207565 1002008 207828 1002010
rect 207565 1001952 207570 1002008
rect 207626 1001952 207828 1002008
rect 207565 1001950 207828 1001952
rect 212336 1002008 212599 1002010
rect 212336 1001952 212538 1002008
rect 212594 1001952 212599 1002008
rect 212336 1001950 212599 1001952
rect 207565 1001947 207631 1001950
rect 212533 1001947 212599 1001950
rect 256969 1002010 257035 1002013
rect 258993 1002010 259059 1002013
rect 256969 1002008 257140 1002010
rect 256969 1001952 256974 1002008
rect 257030 1001952 257140 1002008
rect 256969 1001950 257140 1001952
rect 258796 1002008 259059 1002010
rect 258796 1001952 258998 1002008
rect 259054 1001952 259059 1002008
rect 258796 1001950 259059 1001952
rect 256969 1001947 257035 1001950
rect 258993 1001947 259059 1001950
rect 260189 1002010 260255 1002013
rect 261845 1002010 261911 1002013
rect 263501 1002010 263567 1002013
rect 306097 1002010 306163 1002013
rect 306925 1002010 306991 1002013
rect 309777 1002010 309843 1002013
rect 310145 1002010 310211 1002013
rect 260189 1002008 260452 1002010
rect 260189 1001952 260194 1002008
rect 260250 1001952 260452 1002008
rect 260189 1001950 260452 1001952
rect 261845 1002008 262108 1002010
rect 261845 1001952 261850 1002008
rect 261906 1001952 262108 1002008
rect 261845 1001950 262108 1001952
rect 263304 1002008 263567 1002010
rect 263304 1001952 263506 1002008
rect 263562 1001952 263567 1002008
rect 263304 1001950 263567 1001952
rect 305900 1002008 306163 1002010
rect 305900 1001952 306102 1002008
rect 306158 1001952 306163 1002008
rect 305900 1001950 306163 1001952
rect 306728 1002008 306991 1002010
rect 306728 1001952 306930 1002008
rect 306986 1001952 306991 1002008
rect 306728 1001950 306991 1001952
rect 309580 1002008 309843 1002010
rect 309580 1001952 309782 1002008
rect 309838 1001952 309843 1002008
rect 309580 1001950 309843 1001952
rect 309948 1002008 310211 1002010
rect 309948 1001952 310150 1002008
rect 310206 1001952 310211 1002008
rect 309948 1001950 310211 1001952
rect 260189 1001947 260255 1001950
rect 261845 1001947 261911 1001950
rect 263501 1001947 263567 1001950
rect 306097 1001947 306163 1001950
rect 306925 1001947 306991 1001950
rect 309777 1001947 309843 1001950
rect 310145 1001947 310211 1001950
rect 354029 1002010 354095 1002013
rect 356513 1002010 356579 1002013
rect 357341 1002010 357407 1002013
rect 354029 1002008 354292 1002010
rect 354029 1001952 354034 1002008
rect 354090 1001952 354292 1002008
rect 354029 1001950 354292 1001952
rect 356513 1002008 356684 1002010
rect 356513 1001952 356518 1002008
rect 356574 1001952 356684 1002008
rect 356513 1001950 356684 1001952
rect 357144 1002008 357407 1002010
rect 357144 1001952 357346 1002008
rect 357402 1001952 357407 1002008
rect 357144 1001950 357407 1001952
rect 354029 1001947 354095 1001950
rect 356513 1001947 356579 1001950
rect 357341 1001947 357407 1001950
rect 359365 1002010 359431 1002013
rect 365897 1002010 365963 1002013
rect 359365 1002008 359628 1002010
rect 359365 1001952 359370 1002008
rect 359426 1001952 359628 1002008
rect 359365 1001950 359628 1001952
rect 365700 1002008 365963 1002010
rect 365700 1001952 365902 1002008
rect 365958 1001952 365963 1002008
rect 365700 1001950 365963 1001952
rect 359365 1001947 359431 1001950
rect 365897 1001947 365963 1001950
rect 421465 1002010 421531 1002013
rect 425513 1002010 425579 1002013
rect 501321 1002010 501387 1002013
rect 421465 1002008 421636 1002010
rect 421465 1001952 421470 1002008
rect 421526 1001952 421636 1002008
rect 421465 1001950 421636 1001952
rect 425316 1002008 425579 1002010
rect 425316 1001952 425518 1002008
rect 425574 1001952 425579 1002008
rect 425316 1001950 425579 1001952
rect 501124 1002008 501387 1002010
rect 501124 1001952 501326 1002008
rect 501382 1001952 501387 1002008
rect 501124 1001950 501387 1001952
rect 421465 1001947 421531 1001950
rect 425513 1001947 425579 1001950
rect 501321 1001947 501387 1001950
rect 502149 1002010 502215 1002013
rect 503345 1002010 503411 1002013
rect 504541 1002010 504607 1002013
rect 557993 1002010 558059 1002013
rect 561673 1002010 561739 1002013
rect 502149 1002008 502412 1002010
rect 502149 1001952 502154 1002008
rect 502210 1001952 502412 1002008
rect 502149 1001950 502412 1001952
rect 503345 1002008 503608 1002010
rect 503345 1001952 503350 1002008
rect 503406 1001952 503608 1002008
rect 503345 1001950 503608 1001952
rect 504436 1002008 504607 1002010
rect 504436 1001952 504546 1002008
rect 504602 1001952 504607 1002008
rect 504436 1001950 504607 1001952
rect 557796 1002008 558059 1002010
rect 557796 1001952 557998 1002008
rect 558054 1001952 558059 1002008
rect 557796 1001950 558059 1001952
rect 561476 1002008 561739 1002010
rect 561476 1001952 561678 1002008
rect 561734 1001952 561739 1002008
rect 561476 1001950 561739 1001952
rect 502149 1001947 502215 1001950
rect 503345 1001947 503411 1001950
rect 504541 1001947 504607 1001950
rect 557993 1001947 558059 1001950
rect 561673 1001947 561739 1001950
rect 202689 1001194 202755 1001197
rect 550265 1001194 550331 1001197
rect 202689 1001192 202952 1001194
rect 202689 1001136 202694 1001192
rect 202750 1001136 202952 1001192
rect 202689 1001134 202952 1001136
rect 550068 1001192 550331 1001194
rect 550068 1001136 550270 1001192
rect 550326 1001136 550331 1001192
rect 550068 1001134 550331 1001136
rect 202689 1001131 202755 1001134
rect 550265 1001131 550331 1001134
rect 507393 999154 507459 999157
rect 507196 999152 507459 999154
rect 507196 999096 507398 999152
rect 507454 999096 507459 999152
rect 507196 999094 507459 999096
rect 507393 999091 507459 999094
rect 505369 999018 505435 999021
rect 505369 999016 505632 999018
rect 505369 998960 505374 999016
rect 505430 998960 505632 999016
rect 505369 998958 505632 998960
rect 505369 998955 505435 998958
rect 203885 998882 203951 998885
rect 203885 998880 204148 998882
rect 203885 998824 203890 998880
rect 203946 998824 204148 998880
rect 203885 998822 204148 998824
rect 203885 998819 203951 998822
rect 204345 998746 204411 998749
rect 507025 998746 507091 998749
rect 204345 998744 204516 998746
rect 204345 998688 204350 998744
rect 204406 998688 204516 998744
rect 204345 998686 204516 998688
rect 506828 998744 507091 998746
rect 506828 998688 507030 998744
rect 507086 998688 507091 998744
rect 506828 998686 507091 998688
rect 204345 998683 204411 998686
rect 507025 998683 507091 998686
rect 203517 998610 203583 998613
rect 203320 998608 203583 998610
rect 203320 998552 203522 998608
rect 203578 998552 203583 998608
rect 203320 998550 203583 998552
rect 203517 998547 203583 998550
rect 516685 998610 516751 998613
rect 518893 998610 518959 998613
rect 516685 998608 518959 998610
rect 516685 998552 516690 998608
rect 516746 998552 518898 998608
rect 518954 998552 518959 998608
rect 516685 998550 518959 998552
rect 516685 998547 516751 998550
rect 518893 998547 518959 998550
rect 430849 998338 430915 998341
rect 430652 998336 430915 998338
rect 430652 998280 430854 998336
rect 430910 998280 430915 998336
rect 430652 998278 430915 998280
rect 430849 998275 430915 998278
rect 509049 998338 509115 998341
rect 509049 998336 509312 998338
rect 509049 998280 509054 998336
rect 509110 998280 509312 998336
rect 509049 998278 509312 998280
rect 509049 998275 509115 998278
rect 203517 998202 203583 998205
rect 253657 998202 253723 998205
rect 430021 998202 430087 998205
rect 203517 998200 203780 998202
rect 203517 998144 203522 998200
rect 203578 998144 203780 998200
rect 203517 998142 203780 998144
rect 253460 998200 253723 998202
rect 253460 998144 253662 998200
rect 253718 998144 253723 998200
rect 253460 998142 253723 998144
rect 429824 998200 430087 998202
rect 429824 998144 430026 998200
rect 430082 998144 430087 998200
rect 429824 998142 430087 998144
rect 203517 998139 203583 998142
rect 253657 998139 253723 998142
rect 430021 998139 430087 998142
rect 508221 998202 508287 998205
rect 508221 998200 508484 998202
rect 508221 998144 508226 998200
rect 508282 998144 508484 998200
rect 508221 998142 508484 998144
rect 508221 998139 508287 998142
rect 202689 998066 202755 998069
rect 202492 998064 202755 998066
rect 202492 998008 202694 998064
rect 202750 998008 202755 998064
rect 202492 998006 202755 998008
rect 202689 998003 202755 998006
rect 246573 998066 246639 998069
rect 432045 998066 432111 998069
rect 246573 998064 246682 998066
rect 246573 998008 246578 998064
rect 246634 998008 246682 998064
rect 246573 998003 246682 998008
rect 432045 998064 432308 998066
rect 432045 998008 432050 998064
rect 432106 998008 432308 998064
rect 432045 998006 432308 998008
rect 432045 998003 432111 998006
rect 201861 997930 201927 997933
rect 205541 997930 205607 997933
rect 201861 997928 202124 997930
rect 201861 997872 201866 997928
rect 201922 997872 202124 997928
rect 201861 997870 202124 997872
rect 205344 997928 205607 997930
rect 205344 997872 205546 997928
rect 205602 997872 205607 997928
rect 205344 997870 205607 997872
rect 201861 997867 201927 997870
rect 205541 997867 205607 997870
rect 196065 997794 196131 997797
rect 200205 997794 200271 997797
rect 196065 997792 200271 997794
rect 196065 997736 196070 997792
rect 196126 997736 200210 997792
rect 200266 997736 200271 997792
rect 196065 997734 200271 997736
rect 196065 997731 196131 997734
rect 200205 997731 200271 997734
rect 204713 997794 204779 997797
rect 204713 997792 204976 997794
rect 204713 997736 204718 997792
rect 204774 997736 204976 997792
rect 204713 997734 204976 997736
rect 204713 997731 204779 997734
rect 246622 997660 246682 998003
rect 253657 997930 253723 997933
rect 430021 997930 430087 997933
rect 508221 997930 508287 997933
rect 253657 997928 253920 997930
rect 253657 997872 253662 997928
rect 253718 997872 253920 997928
rect 253657 997870 253920 997872
rect 430021 997928 430284 997930
rect 430021 997872 430026 997928
rect 430082 997872 430284 997928
rect 430021 997870 430284 997872
rect 508116 997928 508287 997930
rect 508116 997872 508226 997928
rect 508282 997872 508287 997928
rect 508116 997870 508287 997872
rect 253657 997867 253723 997870
rect 430021 997867 430087 997870
rect 508221 997867 508287 997870
rect 252461 997794 252527 997797
rect 252264 997792 252527 997794
rect 252264 997736 252466 997792
rect 252522 997736 252527 997792
rect 252264 997734 252527 997736
rect 252461 997731 252527 997734
rect 298093 997794 298159 997797
rect 301681 997794 301747 997797
rect 298093 997792 301747 997794
rect 298093 997736 298098 997792
rect 298154 997736 301686 997792
rect 301742 997736 301747 997792
rect 298093 997734 301747 997736
rect 298093 997731 298159 997734
rect 301681 997731 301747 997734
rect 374637 997794 374703 997797
rect 435357 997794 435423 997797
rect 512637 997794 512703 997797
rect 552289 997794 552355 997797
rect 374637 997792 383762 997794
rect 374637 997736 374642 997792
rect 374698 997736 383762 997792
rect 374637 997734 383762 997736
rect 433136 997792 435423 997794
rect 433136 997736 435362 997792
rect 435418 997736 435423 997792
rect 433136 997734 435423 997736
rect 510140 997792 512703 997794
rect 510140 997736 512642 997792
rect 512698 997736 512703 997792
rect 510140 997734 512703 997736
rect 552092 997792 552355 997794
rect 552092 997736 552294 997792
rect 552350 997736 552355 997792
rect 552092 997734 552355 997736
rect 374637 997731 374703 997734
rect 246614 997596 246620 997660
rect 246684 997596 246690 997660
rect 86534 997188 86540 997252
rect 86604 997250 86610 997252
rect 94681 997250 94747 997253
rect 86604 997248 94747 997250
rect 86604 997192 94686 997248
rect 94742 997192 94747 997248
rect 86604 997190 94747 997192
rect 86604 997188 86610 997190
rect 94681 997187 94747 997190
rect 117221 997250 117287 997253
rect 143809 997250 143875 997253
rect 117221 997248 143875 997250
rect 117221 997192 117226 997248
rect 117282 997192 143814 997248
rect 143870 997192 143875 997248
rect 117221 997190 143875 997192
rect 117221 997187 117287 997190
rect 143809 997187 143875 997190
rect 192518 997188 192524 997252
rect 192588 997250 192594 997252
rect 200205 997250 200271 997253
rect 249057 997250 249123 997253
rect 192588 997248 200271 997250
rect 192588 997192 200210 997248
rect 200266 997192 200271 997248
rect 192588 997190 200271 997192
rect 192588 997188 192594 997190
rect 200205 997187 200271 997190
rect 238526 997248 249123 997250
rect 238526 997192 249062 997248
rect 249118 997192 249123 997248
rect 238526 997190 249123 997192
rect 89662 996916 89668 996980
rect 89732 996978 89738 996980
rect 92473 996978 92539 996981
rect 89732 996976 92539 996978
rect 89732 996920 92478 996976
rect 92534 996920 92539 996976
rect 89732 996918 92539 996920
rect 89732 996916 89738 996918
rect 92473 996915 92539 996918
rect 116945 996978 117011 996981
rect 144821 996978 144887 996981
rect 116945 996976 144887 996978
rect 116945 996920 116950 996976
rect 117006 996920 144826 996976
rect 144882 996920 144887 996976
rect 116945 996918 144887 996920
rect 116945 996915 117011 996918
rect 144821 996915 144887 996918
rect 200205 996706 200271 996709
rect 195930 996704 200271 996706
rect 195930 996648 200210 996704
rect 200266 996648 200271 996704
rect 195930 996646 200271 996648
rect 188838 996508 188844 996572
rect 188908 996570 188914 996572
rect 195930 996570 195990 996646
rect 200205 996643 200271 996646
rect 188908 996510 195990 996570
rect 188908 996508 188914 996510
rect 144361 996434 144427 996437
rect 82310 996374 86970 996434
rect 82310 995757 82370 996374
rect 86910 996298 86970 996374
rect 138430 996432 144427 996434
rect 138430 996376 144366 996432
rect 144422 996376 144427 996432
rect 138430 996374 144427 996376
rect 126237 996298 126303 996301
rect 86910 996238 93870 996298
rect 93810 996162 93870 996238
rect 126237 996296 136466 996298
rect 126237 996240 126242 996296
rect 126298 996240 136466 996296
rect 126237 996238 136466 996240
rect 126237 996235 126303 996238
rect 97257 996162 97323 996165
rect 93810 996160 97323 996162
rect 93810 996104 97262 996160
rect 97318 996104 97323 996160
rect 93810 996102 97323 996104
rect 97257 996099 97323 996102
rect 92657 996026 92723 996029
rect 89302 996024 92723 996026
rect 89302 995968 92662 996024
rect 92718 995968 92723 996024
rect 89302 995966 92723 995968
rect 82261 995752 82370 995757
rect 86493 995756 86559 995757
rect 86493 995754 86540 995756
rect 82261 995696 82266 995752
rect 82322 995696 82370 995752
rect 82261 995694 82370 995696
rect 86448 995752 86540 995754
rect 86448 995696 86498 995752
rect 86448 995694 86540 995696
rect 82261 995691 82327 995694
rect 86493 995692 86540 995694
rect 86604 995692 86610 995756
rect 88977 995754 89043 995757
rect 89302 995754 89362 995966
rect 92657 995963 92723 995966
rect 132350 995964 132356 996028
rect 132420 996026 132426 996028
rect 132420 995966 132970 996026
rect 132420 995964 132426 995966
rect 132910 995757 132970 995966
rect 89621 995756 89687 995757
rect 89621 995754 89668 995756
rect 88977 995752 89362 995754
rect 88977 995696 88982 995752
rect 89038 995696 89362 995752
rect 88977 995694 89362 995696
rect 89576 995752 89668 995754
rect 89576 995696 89626 995752
rect 89576 995694 89668 995696
rect 86493 995691 86559 995692
rect 88977 995691 89043 995694
rect 89621 995692 89668 995694
rect 89732 995692 89738 995756
rect 90265 995754 90331 995757
rect 93117 995754 93183 995757
rect 90265 995752 93183 995754
rect 90265 995696 90270 995752
rect 90326 995696 93122 995752
rect 93178 995696 93183 995752
rect 90265 995694 93183 995696
rect 89621 995691 89687 995692
rect 90265 995691 90331 995694
rect 93117 995691 93183 995694
rect 131849 995754 131915 995757
rect 132534 995754 132540 995756
rect 131849 995752 132540 995754
rect 131849 995696 131854 995752
rect 131910 995696 132540 995752
rect 131849 995694 132540 995696
rect 131849 995691 131915 995694
rect 132534 995692 132540 995694
rect 132604 995692 132610 995756
rect 132910 995752 133019 995757
rect 132910 995696 132958 995752
rect 133014 995696 133019 995752
rect 132910 995694 133019 995696
rect 132953 995691 133019 995694
rect 84653 995482 84719 995485
rect 92841 995482 92907 995485
rect 84653 995480 92907 995482
rect 84653 995424 84658 995480
rect 84714 995424 92846 995480
rect 92902 995424 92907 995480
rect 84653 995422 92907 995424
rect 84653 995419 84719 995422
rect 92841 995419 92907 995422
rect 132401 995348 132467 995349
rect 132350 995346 132356 995348
rect 132310 995286 132356 995346
rect 132420 995344 132467 995348
rect 132462 995288 132467 995344
rect 132350 995284 132356 995286
rect 132420 995284 132467 995288
rect 136406 995346 136466 996238
rect 138430 996026 138490 996374
rect 144361 996371 144427 996374
rect 200665 996298 200731 996301
rect 200665 996296 200836 996298
rect 200665 996240 200670 996296
rect 200726 996240 200836 996296
rect 200665 996238 200836 996240
rect 200665 996235 200731 996238
rect 144177 996162 144243 996165
rect 195278 996162 195284 996164
rect 137142 995966 138490 996026
rect 139534 996160 144243 996162
rect 139534 996104 144182 996160
rect 144238 996104 144243 996160
rect 139534 996102 144243 996104
rect 136725 995754 136791 995757
rect 137142 995754 137202 995966
rect 136725 995752 137202 995754
rect 136725 995696 136730 995752
rect 136786 995696 137202 995752
rect 136725 995694 137202 995696
rect 137369 995754 137435 995757
rect 139534 995754 139594 996102
rect 144177 996099 144243 996102
rect 142286 995890 142292 995892
rect 141558 995830 142292 995890
rect 137369 995752 139594 995754
rect 137369 995696 137374 995752
rect 137430 995696 139594 995752
rect 137369 995694 139594 995696
rect 140405 995754 140471 995757
rect 141558 995754 141618 995830
rect 142286 995828 142292 995830
rect 142356 995828 142362 995892
rect 140405 995752 141618 995754
rect 140405 995696 140410 995752
rect 140466 995696 141618 995752
rect 140405 995694 141618 995696
rect 154297 995754 154363 995757
rect 156830 995754 156890 996132
rect 154297 995752 156890 995754
rect 154297 995696 154302 995752
rect 154358 995696 156890 995752
rect 154297 995694 156890 995696
rect 136725 995691 136791 995694
rect 137369 995691 137435 995694
rect 140405 995691 140471 995694
rect 154297 995691 154363 995694
rect 141785 995618 141851 995621
rect 147121 995618 147187 995621
rect 141785 995616 147187 995618
rect 141785 995560 141790 995616
rect 141846 995560 147126 995616
rect 147182 995560 147187 995616
rect 141785 995558 147187 995560
rect 141785 995555 141851 995558
rect 147121 995555 147187 995558
rect 159222 995482 159282 996132
rect 192342 996102 195284 996162
rect 192342 996026 192402 996102
rect 195278 996100 195284 996102
rect 195348 996100 195354 996164
rect 176610 995966 192402 996026
rect 175917 995890 175983 995893
rect 176610 995890 176670 995966
rect 175917 995888 176670 995890
rect 175917 995832 175922 995888
rect 175978 995832 176670 995888
rect 175917 995830 176670 995832
rect 195053 995890 195119 995893
rect 202321 995890 202387 995893
rect 195053 995888 202387 995890
rect 195053 995832 195058 995888
rect 195114 995832 202326 995888
rect 202382 995832 202387 995888
rect 195053 995830 202387 995832
rect 175917 995827 175983 995830
rect 195053 995827 195119 995830
rect 202321 995827 202387 995830
rect 203609 995890 203675 995893
rect 208166 995890 208226 996132
rect 203609 995888 208226 995890
rect 203609 995832 203614 995888
rect 203670 995832 208226 995888
rect 203609 995830 208226 995832
rect 208393 995890 208459 995893
rect 209822 995890 209882 996132
rect 208393 995888 209882 995890
rect 208393 995832 208398 995888
rect 208454 995832 209882 995888
rect 208393 995830 209882 995832
rect 203609 995827 203675 995830
rect 208393 995827 208459 995830
rect 192477 995790 192543 995791
rect 192477 995788 192524 995790
rect 192432 995786 192524 995788
rect 192432 995730 192482 995786
rect 192432 995728 192524 995730
rect 192477 995726 192524 995728
rect 192588 995726 192594 995790
rect 192477 995725 192543 995726
rect 177297 995618 177363 995621
rect 210650 995618 210710 996132
rect 238526 995757 238586 997190
rect 249057 997187 249123 997190
rect 295190 997188 295196 997252
rect 295260 997250 295266 997252
rect 299473 997250 299539 997253
rect 295260 997248 299539 997250
rect 295260 997192 299478 997248
rect 299534 997192 299539 997248
rect 295260 997190 299539 997192
rect 383702 997250 383762 997734
rect 435357 997731 435423 997734
rect 512637 997731 512703 997734
rect 552289 997731 552355 997734
rect 523861 997660 523927 997661
rect 523861 997658 523908 997660
rect 523816 997656 523908 997658
rect 523816 997600 523866 997656
rect 523816 997598 523908 997600
rect 523861 997596 523908 997598
rect 523972 997596 523978 997660
rect 523861 997595 523927 997596
rect 387742 997250 387748 997252
rect 383702 997190 387748 997250
rect 295260 997188 295266 997190
rect 299473 997187 299539 997190
rect 387742 997188 387748 997190
rect 387812 997188 387818 997252
rect 440049 997250 440115 997253
rect 488901 997250 488967 997253
rect 440049 997248 488967 997250
rect 440049 997192 440054 997248
rect 440110 997192 488906 997248
rect 488962 997192 488967 997248
rect 440049 997190 488967 997192
rect 440049 997187 440115 997190
rect 488901 997187 488967 997190
rect 511441 997250 511507 997253
rect 511942 997250 511948 997252
rect 511441 997248 511948 997250
rect 511441 997192 511446 997248
rect 511502 997192 511948 997248
rect 511441 997190 511948 997192
rect 511441 997187 511507 997190
rect 511942 997188 511948 997190
rect 512012 997188 512018 997252
rect 524045 997250 524111 997253
rect 533470 997250 533476 997252
rect 524045 997248 533476 997250
rect 524045 997192 524050 997248
rect 524106 997192 533476 997248
rect 524045 997190 533476 997192
rect 524045 997187 524111 997190
rect 533470 997188 533476 997190
rect 533540 997188 533546 997252
rect 552289 997250 552355 997253
rect 625061 997250 625127 997253
rect 625245 997250 625311 997253
rect 552289 997248 552552 997250
rect 552289 997192 552294 997248
rect 552350 997192 552552 997248
rect 552289 997190 552552 997192
rect 625016 997248 625311 997250
rect 625016 997192 625066 997248
rect 625122 997192 625250 997248
rect 625306 997192 625311 997248
rect 625016 997190 625311 997192
rect 552289 997187 552355 997190
rect 625061 997187 625127 997190
rect 625245 997187 625311 997190
rect 246614 996978 246620 996980
rect 241102 996918 246620 996978
rect 241102 996570 241162 996918
rect 246614 996916 246620 996918
rect 246684 996916 246690 996980
rect 290774 996916 290780 996980
rect 290844 996978 290850 996980
rect 299289 996978 299355 996981
rect 290844 996976 299355 996978
rect 290844 996920 299294 996976
rect 299350 996920 299355 996976
rect 290844 996918 299355 996920
rect 290844 996916 290850 996918
rect 299289 996915 299355 996918
rect 372521 996978 372587 996981
rect 399937 996978 400003 996981
rect 372521 996976 400003 996978
rect 372521 996920 372526 996976
rect 372582 996920 399942 996976
rect 399998 996920 400003 996976
rect 372521 996918 400003 996920
rect 372521 996915 372587 996918
rect 399937 996915 400003 996918
rect 439865 996978 439931 996981
rect 489085 996978 489151 996981
rect 439865 996976 489151 996978
rect 439865 996920 439870 996976
rect 439926 996920 489090 996976
rect 489146 996920 489151 996976
rect 439865 996918 489151 996920
rect 439865 996915 439931 996918
rect 489085 996915 489151 996918
rect 516869 996978 516935 996981
rect 540329 996978 540395 996981
rect 516869 996976 540395 996978
rect 516869 996920 516874 996976
rect 516930 996920 540334 996976
rect 540390 996920 540395 996976
rect 516869 996918 540395 996920
rect 516869 996915 516935 996918
rect 540329 996915 540395 996918
rect 590561 996978 590627 996981
rect 629886 996978 629892 996980
rect 590561 996976 629892 996978
rect 590561 996920 590566 996976
rect 590622 996920 629892 996976
rect 590561 996918 629892 996920
rect 590561 996915 590627 996918
rect 629886 996916 629892 996918
rect 629956 996916 629962 996980
rect 247125 996706 247191 996709
rect 298829 996706 298895 996709
rect 240550 996510 241162 996570
rect 242758 996704 247191 996706
rect 242758 996648 247130 996704
rect 247186 996648 247191 996704
rect 242758 996646 247191 996648
rect 240550 996162 240610 996510
rect 242758 996298 242818 996646
rect 247125 996643 247191 996646
rect 282686 996704 298895 996706
rect 282686 996648 298834 996704
rect 298890 996648 298895 996704
rect 282686 996646 298895 996648
rect 243854 996372 243860 996436
rect 243924 996434 243930 996436
rect 246665 996434 246731 996437
rect 243924 996432 246731 996434
rect 243924 996376 246670 996432
rect 246726 996376 246731 996432
rect 243924 996374 246731 996376
rect 243924 996372 243930 996374
rect 246665 996371 246731 996374
rect 239998 996102 240610 996162
rect 240734 996238 242818 996298
rect 238526 995752 238635 995757
rect 238526 995696 238574 995752
rect 238630 995696 238635 995752
rect 238526 995694 238635 995696
rect 238569 995691 238635 995694
rect 239581 995754 239647 995757
rect 239998 995754 240058 996102
rect 240734 995890 240794 996238
rect 245142 996026 245148 996028
rect 240550 995830 240794 995890
rect 242390 995966 245148 996026
rect 239581 995752 240058 995754
rect 239581 995696 239586 995752
rect 239642 995696 240058 995752
rect 239581 995694 240058 995696
rect 240225 995754 240291 995757
rect 240550 995754 240610 995830
rect 240225 995752 240610 995754
rect 240225 995696 240230 995752
rect 240286 995696 240610 995752
rect 240225 995694 240610 995696
rect 240869 995754 240935 995757
rect 242390 995754 242450 995966
rect 245142 995964 245148 995966
rect 245212 995964 245218 996028
rect 246665 996026 246731 996029
rect 245334 996024 246731 996026
rect 245334 995968 246670 996024
rect 246726 995968 246731 996024
rect 245334 995966 246731 995968
rect 243813 995756 243879 995757
rect 243813 995754 243860 995756
rect 240869 995752 242450 995754
rect 240869 995696 240874 995752
rect 240930 995696 242450 995752
rect 240869 995694 242450 995696
rect 243768 995752 243860 995754
rect 243768 995696 243818 995752
rect 243768 995694 243860 995696
rect 239581 995691 239647 995694
rect 240225 995691 240291 995694
rect 240869 995691 240935 995694
rect 243813 995692 243860 995694
rect 243924 995692 243930 995756
rect 244089 995754 244155 995757
rect 245334 995754 245394 995966
rect 246665 995963 246731 995966
rect 244089 995752 245394 995754
rect 244089 995696 244094 995752
rect 244150 995696 245394 995752
rect 244089 995694 245394 995696
rect 245561 995754 245627 995757
rect 246941 995754 247007 995757
rect 245561 995752 247007 995754
rect 245561 995696 245566 995752
rect 245622 995696 246946 995752
rect 247002 995696 247007 995752
rect 245561 995694 247007 995696
rect 243813 995691 243879 995692
rect 244089 995691 244155 995694
rect 245561 995691 245627 995694
rect 246941 995691 247007 995694
rect 247125 995754 247191 995757
rect 253381 995754 253447 995757
rect 247125 995752 253447 995754
rect 247125 995696 247130 995752
rect 247186 995696 253386 995752
rect 253442 995696 253447 995752
rect 247125 995694 253447 995696
rect 247125 995691 247191 995694
rect 253381 995691 253447 995694
rect 177297 995616 210710 995618
rect 177297 995560 177302 995616
rect 177358 995560 210710 995616
rect 177297 995558 210710 995560
rect 177297 995555 177363 995558
rect 151770 995422 159282 995482
rect 151770 995346 151830 995422
rect 245142 995420 245148 995484
rect 245212 995482 245218 995484
rect 251173 995482 251239 995485
rect 245212 995480 251239 995482
rect 245212 995424 251178 995480
rect 251234 995424 251239 995480
rect 245212 995422 251239 995424
rect 245212 995420 245218 995422
rect 251173 995419 251239 995422
rect 136406 995286 151830 995346
rect 170857 995346 170923 995349
rect 171685 995346 171751 995349
rect 170857 995344 171751 995346
rect 170857 995288 170862 995344
rect 170918 995288 171690 995344
rect 171746 995288 171751 995344
rect 170857 995286 171751 995288
rect 132401 995283 132467 995284
rect 170857 995283 170923 995286
rect 171685 995283 171751 995286
rect 183829 995346 183895 995349
rect 195053 995346 195119 995349
rect 183829 995344 195119 995346
rect 183829 995288 183834 995344
rect 183890 995288 195058 995344
rect 195114 995288 195119 995344
rect 183829 995286 195119 995288
rect 183829 995283 183895 995286
rect 195053 995283 195119 995286
rect 195278 995284 195284 995348
rect 195348 995346 195354 995348
rect 203609 995346 203675 995349
rect 195348 995344 203675 995346
rect 195348 995288 203614 995344
rect 203670 995288 203675 995344
rect 195348 995286 203675 995288
rect 195348 995284 195354 995286
rect 203609 995283 203675 995286
rect 242065 995346 242131 995349
rect 245009 995346 245075 995349
rect 242065 995344 245075 995346
rect 242065 995288 242070 995344
rect 242126 995288 245014 995344
rect 245070 995288 245075 995344
rect 242065 995286 245075 995288
rect 242065 995283 242131 995286
rect 245009 995283 245075 995286
rect 77017 995074 77083 995077
rect 101397 995074 101463 995077
rect 77017 995072 101463 995074
rect 77017 995016 77022 995072
rect 77078 995016 101402 995072
rect 101458 995016 101463 995072
rect 77017 995014 101463 995016
rect 77017 995011 77083 995014
rect 101397 995011 101463 995014
rect 124857 995074 124923 995077
rect 154297 995074 154363 995077
rect 124857 995072 154363 995074
rect 124857 995016 124862 995072
rect 124918 995016 154302 995072
rect 154358 995016 154363 995072
rect 124857 995014 154363 995016
rect 124857 995011 124923 995014
rect 154297 995011 154363 995014
rect 173157 995074 173223 995077
rect 208393 995074 208459 995077
rect 173157 995072 208459 995074
rect 173157 995016 173162 995072
rect 173218 995016 208398 995072
rect 208454 995016 208459 995072
rect 173157 995014 208459 995016
rect 173157 995011 173223 995014
rect 208393 995011 208459 995014
rect 228357 995074 228423 995077
rect 261250 995074 261310 996132
rect 282686 995757 282746 996646
rect 298829 996643 298895 996646
rect 391974 996644 391980 996708
rect 392044 996706 392050 996708
rect 400489 996706 400555 996709
rect 392044 996704 400555 996706
rect 392044 996648 400494 996704
rect 400550 996648 400555 996704
rect 392044 996646 400555 996648
rect 392044 996644 392050 996646
rect 400489 996643 400555 996646
rect 472617 996706 472683 996709
rect 480478 996706 480484 996708
rect 472617 996704 480484 996706
rect 472617 996648 472622 996704
rect 472678 996648 480484 996704
rect 472617 996646 480484 996648
rect 472617 996643 472683 996646
rect 480478 996644 480484 996646
rect 480548 996644 480554 996708
rect 489821 996706 489887 996709
rect 490005 996706 490071 996709
rect 489821 996704 490071 996706
rect 489821 996648 489826 996704
rect 489882 996648 490010 996704
rect 490066 996648 490071 996704
rect 489821 996646 490071 996648
rect 489821 996643 489887 996646
rect 490005 996643 490071 996646
rect 516685 996706 516751 996709
rect 523493 996706 523559 996709
rect 516685 996704 523559 996706
rect 516685 996648 516690 996704
rect 516746 996648 523498 996704
rect 523554 996648 523559 996704
rect 516685 996646 523559 996648
rect 516685 996643 516751 996646
rect 523493 996643 523559 996646
rect 590561 996706 590627 996709
rect 630254 996706 630260 996708
rect 590561 996704 630260 996706
rect 590561 996648 590566 996704
rect 590622 996648 630260 996704
rect 590561 996646 630260 996648
rect 590561 996643 590627 996646
rect 630254 996644 630260 996646
rect 630324 996644 630330 996708
rect 553117 996570 553183 996573
rect 552920 996568 553183 996570
rect 552920 996512 553122 996568
rect 553178 996512 553183 996568
rect 552920 996510 553183 996512
rect 553117 996507 553183 996510
rect 294822 996372 294828 996436
rect 294892 996434 294898 996436
rect 298645 996434 298711 996437
rect 294892 996432 298711 996434
rect 294892 996376 298650 996432
rect 298706 996376 298711 996432
rect 294892 996374 298711 996376
rect 294892 996372 294898 996374
rect 298645 996371 298711 996374
rect 372337 996434 372403 996437
rect 400029 996434 400095 996437
rect 414473 996434 414539 996437
rect 372337 996432 392226 996434
rect 372337 996376 372342 996432
rect 372398 996376 392226 996432
rect 372337 996374 392226 996376
rect 372337 996371 372403 996374
rect 291878 996162 291884 996164
rect 290782 996102 291884 996162
rect 282686 995752 282795 995757
rect 282686 995696 282734 995752
rect 282790 995696 282795 995752
rect 282686 995694 282795 995696
rect 282729 995691 282795 995694
rect 288065 995754 288131 995757
rect 290782 995754 290842 996102
rect 291878 996100 291884 996102
rect 291948 996100 291954 996164
rect 302877 996162 302943 996165
rect 391974 996162 391980 996164
rect 292530 996160 302943 996162
rect 292530 996104 302882 996160
rect 302938 996104 302943 996160
rect 292530 996102 302943 996104
rect 292530 995890 292590 996102
rect 302877 996099 302943 996102
rect 303061 995890 303127 995893
rect 291702 995830 292590 995890
rect 302190 995888 303127 995890
rect 302190 995832 303066 995888
rect 303122 995832 303127 995888
rect 302190 995830 303127 995832
rect 288065 995752 290842 995754
rect 288065 995696 288070 995752
rect 288126 995696 290842 995752
rect 288065 995694 290842 995696
rect 291101 995754 291167 995757
rect 291702 995754 291762 995830
rect 291101 995752 291762 995754
rect 291101 995696 291106 995752
rect 291162 995696 291762 995752
rect 291101 995694 291762 995696
rect 288065 995691 288131 995694
rect 291101 995691 291167 995694
rect 291878 995556 291884 995620
rect 291948 995618 291954 995620
rect 302190 995618 302250 995830
rect 303061 995827 303127 995830
rect 291948 995558 302250 995618
rect 308765 995618 308831 995621
rect 311206 995618 311266 996132
rect 308765 995616 311266 995618
rect 308765 995560 308770 995616
rect 308826 995560 311266 995616
rect 308765 995558 311266 995560
rect 291948 995556 291954 995558
rect 308765 995555 308831 995558
rect 279417 995346 279483 995349
rect 312862 995346 312922 996132
rect 373950 996102 389190 996162
rect 372337 996026 372403 996029
rect 373950 996026 374010 996102
rect 372337 996024 374010 996026
rect 372337 995968 372342 996024
rect 372398 995968 374010 996024
rect 372337 995966 374010 995968
rect 372337 995963 372403 995966
rect 380893 995890 380959 995893
rect 382181 995890 382247 995893
rect 380893 995888 382247 995890
rect 380893 995832 380898 995888
rect 380954 995832 382186 995888
rect 382242 995832 382247 995888
rect 380893 995830 382247 995832
rect 380893 995827 380959 995830
rect 382181 995827 382247 995830
rect 382641 995754 382707 995757
rect 385033 995754 385099 995757
rect 382641 995752 385099 995754
rect 382641 995696 382646 995752
rect 382702 995696 385038 995752
rect 385094 995696 385099 995752
rect 382641 995694 385099 995696
rect 389130 995754 389190 996102
rect 389774 996102 391980 996162
rect 389774 995757 389834 996102
rect 391974 996100 391980 996102
rect 392044 996100 392050 996164
rect 389357 995754 389423 995757
rect 389130 995752 389423 995754
rect 389130 995696 389362 995752
rect 389418 995696 389423 995752
rect 389130 995694 389423 995696
rect 382641 995691 382707 995694
rect 385033 995691 385099 995694
rect 389357 995691 389423 995694
rect 389725 995752 389834 995757
rect 389725 995696 389730 995752
rect 389786 995696 389834 995752
rect 389725 995694 389834 995696
rect 392166 995757 392226 996374
rect 400029 996432 414539 996434
rect 400029 996376 400034 996432
rect 400090 996376 414478 996432
rect 414534 996376 414539 996432
rect 400029 996374 414539 996376
rect 400029 996371 400095 996374
rect 414473 996371 414539 996374
rect 439681 996434 439747 996437
rect 476982 996434 476988 996436
rect 439681 996432 476988 996434
rect 439681 996376 439686 996432
rect 439742 996376 476988 996432
rect 439681 996374 476988 996376
rect 439681 996371 439747 996374
rect 476982 996372 476988 996374
rect 477052 996372 477058 996436
rect 519077 996434 519143 996437
rect 524045 996434 524111 996437
rect 519077 996432 524111 996434
rect 519077 996376 519082 996432
rect 519138 996376 524050 996432
rect 524106 996376 524111 996432
rect 519077 996374 524111 996376
rect 519077 996371 519143 996374
rect 524045 996371 524111 996374
rect 590561 996434 590627 996437
rect 629150 996434 629156 996436
rect 590561 996432 629156 996434
rect 590561 996376 590566 996432
rect 590622 996376 629156 996432
rect 590561 996374 629156 996376
rect 590561 996371 590627 996374
rect 629150 996372 629156 996374
rect 629220 996372 629226 996436
rect 451917 996162 451983 996165
rect 471053 996162 471119 996165
rect 451917 996160 471119 996162
rect 392166 995752 392275 995757
rect 392166 995696 392214 995752
rect 392270 995696 392275 995752
rect 392166 995694 392275 995696
rect 389725 995691 389791 995694
rect 392209 995691 392275 995694
rect 396625 995754 396691 995757
rect 400029 995754 400095 995757
rect 416129 995754 416195 995757
rect 396625 995752 400095 995754
rect 396625 995696 396630 995752
rect 396686 995696 400034 995752
rect 400090 995696 400095 995752
rect 396625 995694 400095 995696
rect 396625 995691 396691 995694
rect 400029 995691 400095 995694
rect 400262 995752 416195 995754
rect 400262 995696 416134 995752
rect 416190 995696 416195 995752
rect 400262 995694 416195 995696
rect 386321 995618 386387 995621
rect 386321 995616 389098 995618
rect 386321 995560 386326 995616
rect 386382 995560 389098 995616
rect 386321 995558 389098 995560
rect 386321 995555 386387 995558
rect 389038 995482 389098 995558
rect 400262 995482 400322 995694
rect 416129 995691 416195 995694
rect 389038 995422 400322 995482
rect 400489 995482 400555 995485
rect 415393 995482 415459 995485
rect 400489 995480 415459 995482
rect 400489 995424 400494 995480
rect 400550 995424 415398 995480
rect 415454 995424 415459 995480
rect 400489 995422 415459 995424
rect 400489 995419 400555 995422
rect 415393 995419 415459 995422
rect 279417 995344 312922 995346
rect 279417 995288 279422 995344
rect 279478 995288 312922 995344
rect 279417 995286 312922 995288
rect 382457 995346 382523 995349
rect 388897 995346 388963 995349
rect 382457 995344 388963 995346
rect 382457 995288 382462 995344
rect 382518 995288 388902 995344
rect 388958 995288 388963 995344
rect 382457 995286 388963 995288
rect 279417 995283 279483 995286
rect 382457 995283 382523 995286
rect 388897 995283 388963 995286
rect 228357 995072 261310 995074
rect 228357 995016 228362 995072
rect 228418 995016 261310 995072
rect 228357 995014 261310 995016
rect 270401 995074 270467 995077
rect 308765 995074 308831 995077
rect 270401 995072 308831 995074
rect 270401 995016 270406 995072
rect 270462 995016 308770 995072
rect 308826 995016 308831 995072
rect 270401 995014 308831 995016
rect 228357 995011 228423 995014
rect 270401 995011 270467 995014
rect 308765 995011 308831 995014
rect 382825 995074 382891 995077
rect 430990 995074 431050 996132
rect 451917 996104 451922 996160
rect 451978 996104 471058 996160
rect 471114 996104 471119 996160
rect 451917 996102 471119 996104
rect 451917 996099 451983 996102
rect 471053 996099 471119 996102
rect 471237 996162 471303 996165
rect 523677 996162 523743 996165
rect 471237 996160 476130 996162
rect 471237 996104 471242 996160
rect 471298 996104 476130 996160
rect 523677 996160 524430 996162
rect 471237 996102 476130 996104
rect 471237 996099 471303 996102
rect 469857 995890 469923 995893
rect 476070 995890 476130 996102
rect 484342 995890 484348 995892
rect 469857 995888 475026 995890
rect 469857 995832 469862 995888
rect 469918 995832 475026 995888
rect 469857 995830 475026 995832
rect 476070 995830 484348 995890
rect 469857 995827 469923 995830
rect 448513 995618 448579 995621
rect 474733 995618 474799 995621
rect 448513 995616 474799 995618
rect 448513 995560 448518 995616
rect 448574 995560 474738 995616
rect 474794 995560 474799 995616
rect 448513 995558 474799 995560
rect 474966 995618 475026 995830
rect 484342 995828 484348 995830
rect 484412 995828 484418 995892
rect 474966 995558 489930 995618
rect 448513 995555 448579 995558
rect 474733 995555 474799 995558
rect 458357 995346 458423 995349
rect 486325 995346 486391 995349
rect 458357 995344 486391 995346
rect 458357 995288 458362 995344
rect 458418 995288 486330 995344
rect 486386 995288 486391 995344
rect 458357 995286 486391 995288
rect 489870 995346 489930 995558
rect 506430 995346 506490 996132
rect 489870 995286 506490 995346
rect 458357 995283 458423 995286
rect 486325 995283 486391 995286
rect 382825 995072 431050 995074
rect 382825 995016 382830 995072
rect 382886 995016 431050 995072
rect 382825 995014 431050 995016
rect 464981 995074 465047 995077
rect 471237 995074 471303 995077
rect 464981 995072 471303 995074
rect 464981 995016 464986 995072
rect 465042 995016 471242 995072
rect 471298 995016 471303 995072
rect 464981 995014 471303 995016
rect 382825 995011 382891 995014
rect 464981 995011 465047 995014
rect 471237 995011 471303 995014
rect 472249 995074 472315 995077
rect 473997 995074 474063 995077
rect 476389 995074 476455 995077
rect 477033 995076 477099 995077
rect 472249 995072 474063 995074
rect 472249 995016 472254 995072
rect 472310 995016 474002 995072
rect 474058 995016 474063 995072
rect 472249 995014 474063 995016
rect 472249 995011 472315 995014
rect 473997 995011 474063 995014
rect 474230 995072 476455 995074
rect 474230 995016 476394 995072
rect 476450 995016 476455 995072
rect 474230 995014 476455 995016
rect 78673 994802 78739 994805
rect 104157 994802 104223 994805
rect 78673 994800 104223 994802
rect 78673 994744 78678 994800
rect 78734 994744 104162 994800
rect 104218 994744 104223 994800
rect 78673 994742 104223 994744
rect 78673 994739 78739 994742
rect 104157 994739 104223 994742
rect 132125 994802 132191 994805
rect 135897 994802 135963 994805
rect 141877 994802 141943 994805
rect 132125 994800 132970 994802
rect 132125 994744 132130 994800
rect 132186 994744 132970 994800
rect 132125 994742 132970 994744
rect 132125 994739 132191 994742
rect 86033 994530 86099 994533
rect 92473 994530 92539 994533
rect 86033 994528 92539 994530
rect 86033 994472 86038 994528
rect 86094 994472 92478 994528
rect 92534 994472 92539 994528
rect 86033 994470 92539 994472
rect 86033 994467 86099 994470
rect 92473 994467 92539 994470
rect 85021 994258 85087 994261
rect 92657 994258 92723 994261
rect 85021 994256 92723 994258
rect 85021 994200 85026 994256
rect 85082 994200 92662 994256
rect 92718 994200 92723 994256
rect 85021 994198 92723 994200
rect 132910 994258 132970 994742
rect 135897 994800 141943 994802
rect 135897 994744 135902 994800
rect 135958 994744 141882 994800
rect 141938 994744 141943 994800
rect 135897 994742 141943 994744
rect 135897 994739 135963 994742
rect 141877 994739 141943 994742
rect 142061 994802 142127 994805
rect 187601 994802 187667 994805
rect 195237 994802 195303 994805
rect 142061 994800 151830 994802
rect 142061 994744 142066 994800
rect 142122 994744 151830 994800
rect 142061 994742 151830 994744
rect 142061 994739 142127 994742
rect 133137 994530 133203 994533
rect 149697 994530 149763 994533
rect 133137 994528 149763 994530
rect 133137 994472 133142 994528
rect 133198 994472 149702 994528
rect 149758 994472 149763 994528
rect 133137 994470 149763 994472
rect 151770 994530 151830 994742
rect 187601 994800 195303 994802
rect 187601 994744 187606 994800
rect 187662 994744 195242 994800
rect 195298 994744 195303 994800
rect 187601 994742 195303 994744
rect 187601 994739 187667 994742
rect 195237 994739 195303 994742
rect 243261 994802 243327 994805
rect 247309 994802 247375 994805
rect 290733 994804 290799 994805
rect 294781 994804 294847 994805
rect 295241 994804 295307 994805
rect 290733 994802 290780 994804
rect 243261 994800 247375 994802
rect 243261 994744 243266 994800
rect 243322 994744 247314 994800
rect 247370 994744 247375 994800
rect 243261 994742 247375 994744
rect 290688 994800 290780 994802
rect 290688 994744 290738 994800
rect 290688 994742 290780 994744
rect 243261 994739 243327 994742
rect 247309 994739 247375 994742
rect 290733 994740 290780 994742
rect 290844 994740 290850 994804
rect 294781 994802 294828 994804
rect 294736 994800 294828 994802
rect 294736 994744 294786 994800
rect 294736 994742 294828 994744
rect 294781 994740 294828 994742
rect 294892 994740 294898 994804
rect 295190 994740 295196 994804
rect 295260 994802 295307 994804
rect 383101 994802 383167 994805
rect 386505 994802 386571 994805
rect 387793 994804 387859 994805
rect 295260 994800 295352 994802
rect 295302 994744 295352 994800
rect 295260 994742 295352 994744
rect 383101 994800 386571 994802
rect 383101 994744 383106 994800
rect 383162 994744 386510 994800
rect 386566 994744 386571 994800
rect 383101 994742 386571 994744
rect 295260 994740 295307 994742
rect 290733 994739 290799 994740
rect 294781 994739 294847 994740
rect 295241 994739 295307 994740
rect 383101 994739 383167 994742
rect 386505 994739 386571 994742
rect 387742 994740 387748 994804
rect 387812 994802 387859 994804
rect 471053 994802 471119 994805
rect 474230 994802 474290 995014
rect 476389 995011 476455 995014
rect 476982 995012 476988 995076
rect 477052 995074 477099 995076
rect 477052 995072 477144 995074
rect 477094 995016 477144 995072
rect 477052 995014 477144 995016
rect 477052 995012 477099 995014
rect 480478 995012 480484 995076
rect 480548 995074 480554 995076
rect 480805 995074 480871 995077
rect 480548 995072 480871 995074
rect 480548 995016 480810 995072
rect 480866 995016 480871 995072
rect 480548 995014 480871 995016
rect 480548 995012 480554 995014
rect 477033 995011 477099 995012
rect 480805 995011 480871 995014
rect 484117 995074 484183 995077
rect 484342 995074 484348 995076
rect 484117 995072 484348 995074
rect 484117 995016 484122 995072
rect 484178 995016 484348 995072
rect 484117 995014 484348 995016
rect 484117 995011 484183 995014
rect 484342 995012 484348 995014
rect 484412 995012 484418 995076
rect 484577 995074 484643 995077
rect 508822 995074 508882 996132
rect 523677 996104 523682 996160
rect 523738 996104 524430 996160
rect 523677 996102 524430 996104
rect 523677 996099 523743 996102
rect 524370 995890 524430 996102
rect 524370 995830 529306 995890
rect 529246 995754 529306 995830
rect 532926 995830 533722 995890
rect 532926 995757 532986 995830
rect 529749 995754 529815 995757
rect 529246 995752 529815 995754
rect 529246 995696 529754 995752
rect 529810 995696 529815 995752
rect 529246 995694 529815 995696
rect 529749 995691 529815 995694
rect 531446 995692 531452 995756
rect 531516 995754 531522 995756
rect 532141 995754 532207 995757
rect 531516 995752 532207 995754
rect 531516 995696 532146 995752
rect 532202 995696 532207 995752
rect 531516 995694 532207 995696
rect 531516 995692 531522 995694
rect 532141 995691 532207 995694
rect 532877 995752 532986 995757
rect 532877 995696 532882 995752
rect 532938 995696 532986 995752
rect 532877 995694 532986 995696
rect 533662 995754 533722 995830
rect 535269 995754 535335 995757
rect 536557 995756 536623 995757
rect 536557 995754 536604 995756
rect 533662 995752 535335 995754
rect 533662 995696 535274 995752
rect 535330 995696 535335 995752
rect 533662 995694 535335 995696
rect 536512 995752 536604 995754
rect 536512 995696 536562 995752
rect 536512 995694 536604 995696
rect 532877 995691 532943 995694
rect 535269 995691 535335 995694
rect 536557 995692 536604 995694
rect 536668 995692 536674 995756
rect 536557 995691 536623 995692
rect 518893 995618 518959 995621
rect 529013 995618 529079 995621
rect 533521 995620 533587 995621
rect 518893 995616 529079 995618
rect 518893 995560 518898 995616
rect 518954 995560 529018 995616
rect 529074 995560 529079 995616
rect 518893 995558 529079 995560
rect 518893 995555 518959 995558
rect 529013 995555 529079 995558
rect 533470 995556 533476 995620
rect 533540 995618 533587 995620
rect 533540 995616 533632 995618
rect 533582 995560 533632 995616
rect 533540 995558 533632 995560
rect 533540 995556 533587 995558
rect 533521 995555 533587 995556
rect 518157 995346 518223 995349
rect 537109 995346 537175 995349
rect 518157 995344 537175 995346
rect 518157 995288 518162 995344
rect 518218 995288 537114 995344
rect 537170 995288 537175 995344
rect 518157 995286 537175 995288
rect 518157 995283 518223 995286
rect 537109 995283 537175 995286
rect 484577 995072 508882 995074
rect 484577 995016 484582 995072
rect 484638 995016 508882 995072
rect 484577 995014 508882 995016
rect 520917 995074 520983 995077
rect 520917 995072 522682 995074
rect 520917 995016 520922 995072
rect 520978 995016 522682 995072
rect 520917 995014 522682 995016
rect 484577 995011 484643 995014
rect 520917 995011 520983 995014
rect 387812 994800 387904 994802
rect 387854 994744 387904 994800
rect 387812 994742 387904 994744
rect 471053 994800 474290 994802
rect 471053 994744 471058 994800
rect 471114 994744 474290 994800
rect 471053 994742 474290 994744
rect 474457 994802 474523 994805
rect 487797 994802 487863 994805
rect 474457 994800 487863 994802
rect 474457 994744 474462 994800
rect 474518 994744 487802 994800
rect 487858 994744 487863 994800
rect 474457 994742 487863 994744
rect 522622 994802 522682 995014
rect 522798 995012 522804 995076
rect 522868 995074 522874 995076
rect 524454 995074 524460 995076
rect 522868 995014 524460 995074
rect 522868 995012 522874 995014
rect 524454 995012 524460 995014
rect 524524 995012 524530 995076
rect 559422 995074 559482 996132
rect 625613 996026 625679 996029
rect 625613 996024 630138 996026
rect 625613 995968 625618 996024
rect 625674 995968 630138 996024
rect 625613 995966 630138 995968
rect 625613 995963 625679 995966
rect 625797 995754 625863 995757
rect 627177 995754 627243 995757
rect 629201 995756 629267 995757
rect 625797 995752 627243 995754
rect 625797 995696 625802 995752
rect 625858 995696 627182 995752
rect 627238 995696 627243 995752
rect 625797 995694 627243 995696
rect 625797 995691 625863 995694
rect 627177 995691 627243 995694
rect 629150 995692 629156 995756
rect 629220 995754 629267 995756
rect 629845 995756 629911 995757
rect 629845 995754 629892 995756
rect 629220 995752 629312 995754
rect 629262 995696 629312 995752
rect 629220 995694 629312 995696
rect 629800 995752 629892 995754
rect 629800 995696 629850 995752
rect 629800 995694 629892 995696
rect 629220 995692 629267 995694
rect 629201 995691 629267 995692
rect 629845 995692 629892 995694
rect 629956 995692 629962 995756
rect 629845 995691 629911 995692
rect 630078 995618 630138 995966
rect 630305 995790 630371 995791
rect 630254 995726 630260 995790
rect 630324 995788 630371 995790
rect 630324 995786 630416 995788
rect 630366 995730 630416 995786
rect 630324 995728 630416 995730
rect 635641 995754 635707 995757
rect 637021 995754 637087 995757
rect 635641 995752 637087 995754
rect 630324 995726 630371 995728
rect 630305 995725 630371 995726
rect 635641 995696 635646 995752
rect 635702 995696 637026 995752
rect 637082 995696 637087 995752
rect 635641 995694 637087 995696
rect 635641 995691 635707 995694
rect 637021 995691 637087 995694
rect 635181 995618 635247 995621
rect 630078 995616 635247 995618
rect 630078 995560 635186 995616
rect 635242 995560 635247 995616
rect 630078 995558 635247 995560
rect 635181 995555 635247 995558
rect 590561 995346 590627 995349
rect 635825 995346 635891 995349
rect 590561 995344 635891 995346
rect 590561 995288 590566 995344
rect 590622 995288 635830 995344
rect 635886 995288 635891 995344
rect 590561 995286 635891 995288
rect 590561 995283 590627 995286
rect 635825 995283 635891 995286
rect 524646 995014 559482 995074
rect 590561 995074 590627 995077
rect 640977 995074 641043 995077
rect 590561 995072 641043 995074
rect 590561 995016 590566 995072
rect 590622 995016 640982 995072
rect 641038 995016 641043 995072
rect 590561 995014 641043 995016
rect 524646 994802 524706 995014
rect 590561 995011 590627 995014
rect 640977 995011 641043 995014
rect 569902 994876 569908 994940
rect 569972 994938 569978 994940
rect 572805 994938 572871 994941
rect 569972 994936 572871 994938
rect 569972 994880 572810 994936
rect 572866 994880 572871 994936
rect 569972 994878 572871 994880
rect 569972 994876 569978 994878
rect 572805 994875 572871 994878
rect 627913 994802 627979 994805
rect 635641 994802 635707 994805
rect 522622 994742 524706 994802
rect 576810 994800 627979 994802
rect 576810 994744 627918 994800
rect 627974 994744 627979 994800
rect 576810 994742 627979 994744
rect 387812 994740 387859 994742
rect 387793 994739 387859 994740
rect 471053 994739 471119 994742
rect 474457 994739 474523 994742
rect 487797 994739 487863 994742
rect 570781 994666 570847 994669
rect 576810 994666 576870 994742
rect 627913 994739 627979 994742
rect 634770 994800 635707 994802
rect 634770 994744 635646 994800
rect 635702 994744 635707 994800
rect 634770 994742 635707 994744
rect 570781 994664 576870 994666
rect 570781 994608 570786 994664
rect 570842 994608 576870 994664
rect 570781 994606 576870 994608
rect 570781 994603 570847 994606
rect 154573 994530 154639 994533
rect 188797 994532 188863 994533
rect 188797 994530 188844 994532
rect 151770 994528 154639 994530
rect 151770 994472 154578 994528
rect 154634 994472 154639 994528
rect 151770 994470 154639 994472
rect 188752 994528 188844 994530
rect 188752 994472 188802 994528
rect 188752 994470 188844 994472
rect 133137 994467 133203 994470
rect 149697 994467 149763 994470
rect 154573 994467 154639 994470
rect 188797 994468 188844 994470
rect 188908 994468 188914 994532
rect 190361 994530 190427 994533
rect 196065 994530 196131 994533
rect 190361 994528 196131 994530
rect 190361 994472 190366 994528
rect 190422 994472 196070 994528
rect 196126 994472 196131 994528
rect 190361 994470 196131 994472
rect 188797 994467 188863 994468
rect 190361 994467 190427 994470
rect 196065 994467 196131 994470
rect 235257 994530 235323 994533
rect 253105 994530 253171 994533
rect 235257 994528 253171 994530
rect 235257 994472 235262 994528
rect 235318 994472 253110 994528
rect 253166 994472 253171 994528
rect 235257 994470 253171 994472
rect 235257 994467 235323 994470
rect 253105 994467 253171 994470
rect 286501 994530 286567 994533
rect 301497 994530 301563 994533
rect 286501 994528 301563 994530
rect 286501 994472 286506 994528
rect 286562 994472 301502 994528
rect 301558 994472 301563 994528
rect 286501 994470 301563 994472
rect 286501 994467 286567 994470
rect 301497 994467 301563 994470
rect 383469 994530 383535 994533
rect 392669 994530 392735 994533
rect 383469 994528 392735 994530
rect 383469 994472 383474 994528
rect 383530 994472 392674 994528
rect 392730 994472 392735 994528
rect 383469 994470 392735 994472
rect 383469 994467 383535 994470
rect 392669 994467 392735 994470
rect 457437 994530 457503 994533
rect 481633 994530 481699 994533
rect 457437 994528 481699 994530
rect 457437 994472 457442 994528
rect 457498 994472 481638 994528
rect 481694 994472 481699 994528
rect 457437 994470 481699 994472
rect 457437 994467 457503 994470
rect 481633 994467 481699 994470
rect 524454 994468 524460 994532
rect 524524 994530 524530 994532
rect 526069 994530 526135 994533
rect 524524 994528 526135 994530
rect 524524 994472 526074 994528
rect 526130 994472 526135 994528
rect 524524 994470 526135 994472
rect 524524 994468 524530 994470
rect 526069 994467 526135 994470
rect 625153 994530 625219 994533
rect 634770 994530 634830 994742
rect 635641 994739 635707 994742
rect 625153 994528 634830 994530
rect 625153 994472 625158 994528
rect 625214 994472 634830 994528
rect 625153 994470 634830 994472
rect 625153 994467 625219 994470
rect 143717 994258 143783 994261
rect 132910 994256 143783 994258
rect 132910 994200 143722 994256
rect 143778 994200 143783 994256
rect 132910 994198 143783 994200
rect 85021 994195 85087 994198
rect 92657 994195 92723 994198
rect 143717 994195 143783 994198
rect 143901 994258 143967 994261
rect 148501 994258 148567 994261
rect 143901 994256 148567 994258
rect 143901 994200 143906 994256
rect 143962 994200 148506 994256
rect 148562 994200 148567 994256
rect 143901 994198 148567 994200
rect 143901 994195 143967 994198
rect 148501 994195 148567 994198
rect 184841 994258 184907 994261
rect 196617 994258 196683 994261
rect 184841 994256 196683 994258
rect 184841 994200 184846 994256
rect 184902 994200 196622 994256
rect 196678 994200 196683 994256
rect 184841 994198 196683 994200
rect 184841 994195 184907 994198
rect 196617 994195 196683 994198
rect 235901 994258 235967 994261
rect 247677 994258 247743 994261
rect 235901 994256 247743 994258
rect 235901 994200 235906 994256
rect 235962 994200 247682 994256
rect 247738 994200 247743 994256
rect 235901 994198 247743 994200
rect 235901 994195 235967 994198
rect 247677 994195 247743 994198
rect 292113 994258 292179 994261
rect 300301 994258 300367 994261
rect 306373 994258 306439 994261
rect 292113 994256 300367 994258
rect 292113 994200 292118 994256
rect 292174 994200 300306 994256
rect 300362 994200 300367 994256
rect 292113 994198 300367 994200
rect 292113 994195 292179 994198
rect 300301 994195 300367 994198
rect 302190 994256 306439 994258
rect 302190 994200 306378 994256
rect 306434 994200 306439 994256
rect 302190 994198 306439 994200
rect 87873 993986 87939 993989
rect 93301 993986 93367 993989
rect 87873 993984 93367 993986
rect 87873 993928 87878 993984
rect 87934 993928 93306 993984
rect 93362 993928 93367 993984
rect 87873 993926 93367 993928
rect 87873 993923 87939 993926
rect 93301 993923 93367 993926
rect 132534 993924 132540 993988
rect 132604 993986 132610 993988
rect 139209 993986 139275 993989
rect 132604 993984 139275 993986
rect 132604 993928 139214 993984
rect 139270 993928 139275 993984
rect 132604 993926 139275 993928
rect 132604 993924 132610 993926
rect 139209 993923 139275 993926
rect 139393 993986 139459 993989
rect 145557 993986 145623 993989
rect 139393 993984 145623 993986
rect 139393 993928 139398 993984
rect 139454 993928 145562 993984
rect 145618 993928 145623 993984
rect 139393 993926 145623 993928
rect 139393 993923 139459 993926
rect 145557 993923 145623 993926
rect 189441 993986 189507 993989
rect 199377 993986 199443 993989
rect 189441 993984 199443 993986
rect 189441 993928 189446 993984
rect 189502 993928 199382 993984
rect 199438 993928 199443 993984
rect 189441 993926 199443 993928
rect 189441 993923 189507 993926
rect 199377 993923 199443 993926
rect 291745 993986 291811 993989
rect 302190 993986 302250 994198
rect 306373 994195 306439 994198
rect 443637 994258 443703 994261
rect 478597 994258 478663 994261
rect 443637 994256 478663 994258
rect 443637 994200 443642 994256
rect 443698 994200 478602 994256
rect 478658 994200 478663 994256
rect 443637 994198 478663 994200
rect 443637 994195 443703 994198
rect 478597 994195 478663 994198
rect 485313 994258 485379 994261
rect 511073 994258 511139 994261
rect 485313 994256 511139 994258
rect 485313 994200 485318 994256
rect 485374 994200 511078 994256
rect 511134 994200 511139 994256
rect 485313 994198 511139 994200
rect 485313 994195 485379 994198
rect 511073 994195 511139 994198
rect 523309 994258 523375 994261
rect 528921 994258 528987 994261
rect 523309 994256 528987 994258
rect 523309 994200 523314 994256
rect 523370 994200 528926 994256
rect 528982 994200 528987 994256
rect 523309 994198 528987 994200
rect 523309 994195 523375 994198
rect 528921 994195 528987 994198
rect 291745 993984 302250 993986
rect 291745 993928 291750 993984
rect 291806 993928 302250 993984
rect 291745 993926 302250 993928
rect 467097 993986 467163 993989
rect 474457 993986 474523 993989
rect 467097 993984 474523 993986
rect 467097 993928 467102 993984
rect 467158 993928 474462 993984
rect 474518 993928 474523 993984
rect 467097 993926 474523 993928
rect 291745 993923 291811 993926
rect 467097 993923 467163 993926
rect 474457 993923 474523 993926
rect 137737 993714 137803 993717
rect 142153 993714 142219 993717
rect 137737 993712 142219 993714
rect 137737 993656 137742 993712
rect 137798 993656 142158 993712
rect 142214 993656 142219 993712
rect 137737 993654 142219 993656
rect 137737 993651 137803 993654
rect 142153 993651 142219 993654
rect 142337 993714 142403 993717
rect 152457 993714 152523 993717
rect 142337 993712 152523 993714
rect 142337 993656 142342 993712
rect 142398 993656 152462 993712
rect 152518 993656 152523 993712
rect 142337 993654 152523 993656
rect 142337 993651 142403 993654
rect 152457 993651 152523 993654
rect 193121 993714 193187 993717
rect 195329 993714 195395 993717
rect 193121 993712 195395 993714
rect 193121 993656 193126 993712
rect 193182 993656 195334 993712
rect 195390 993656 195395 993712
rect 193121 993654 195395 993656
rect 193121 993651 193187 993654
rect 195329 993651 195395 993654
rect 142286 992836 142292 992900
rect 142356 992898 142362 992900
rect 186497 992898 186563 992901
rect 142356 992896 186563 992898
rect 142356 992840 186502 992896
rect 186558 992840 186563 992896
rect 142356 992838 186563 992840
rect 142356 992836 142362 992838
rect 186497 992835 186563 992838
rect 62113 976034 62179 976037
rect 62113 976032 64492 976034
rect 62113 975976 62118 976032
rect 62174 975976 64492 976032
rect 62113 975974 64492 975976
rect 62113 975971 62179 975974
rect 651649 975898 651715 975901
rect 650164 975896 651715 975898
rect 650164 975840 651654 975896
rect 651710 975840 651715 975896
rect 650164 975838 651715 975840
rect 651649 975835 651715 975838
rect 41454 967132 41460 967196
rect 41524 967194 41530 967196
rect 41781 967194 41847 967197
rect 41524 967192 41847 967194
rect 41524 967136 41786 967192
rect 41842 967136 41847 967192
rect 41524 967134 41847 967136
rect 41524 967132 41530 967134
rect 41781 967131 41847 967134
rect 42333 966786 42399 966789
rect 43437 966786 43503 966789
rect 42333 966784 43503 966786
rect 42333 966728 42338 966784
rect 42394 966728 43442 966784
rect 43498 966728 43503 966784
rect 42333 966726 43503 966728
rect 42333 966723 42399 966726
rect 43437 966723 43503 966726
rect 674373 966106 674439 966109
rect 675201 966106 675267 966109
rect 674373 966104 675267 966106
rect 674373 966048 674378 966104
rect 674434 966048 675206 966104
rect 675262 966048 675267 966104
rect 674373 966046 675267 966048
rect 674373 966043 674439 966046
rect 675201 966043 675267 966046
rect 675753 965154 675819 965157
rect 676070 965154 676076 965156
rect 675753 965152 676076 965154
rect 675753 965096 675758 965152
rect 675814 965096 676076 965152
rect 675753 965094 676076 965096
rect 675753 965091 675819 965094
rect 676070 965092 676076 965094
rect 676140 965092 676146 965156
rect 42425 964746 42491 964749
rect 43253 964746 43319 964749
rect 42425 964744 43319 964746
rect 42425 964688 42430 964744
rect 42486 964688 43258 964744
rect 43314 964688 43319 964744
rect 42425 964686 43319 964688
rect 42425 964683 42491 964686
rect 43253 964683 43319 964686
rect 675201 963658 675267 963661
rect 676622 963658 676628 963660
rect 675201 963656 676628 963658
rect 675201 963600 675206 963656
rect 675262 963600 676628 963656
rect 675201 963598 676628 963600
rect 675201 963595 675267 963598
rect 676622 963596 676628 963598
rect 676692 963596 676698 963660
rect 42425 963386 42491 963389
rect 42977 963386 43043 963389
rect 675385 963388 675451 963389
rect 675334 963386 675340 963388
rect 42425 963384 43043 963386
rect 42425 963328 42430 963384
rect 42486 963328 42982 963384
rect 43038 963328 43043 963384
rect 42425 963326 43043 963328
rect 675294 963326 675340 963386
rect 675404 963384 675451 963388
rect 675446 963328 675451 963384
rect 42425 963323 42491 963326
rect 42977 963323 43043 963326
rect 675334 963324 675340 963326
rect 675404 963324 675451 963328
rect 675385 963323 675451 963324
rect 42241 962978 42307 962981
rect 43437 962978 43503 962981
rect 42241 962976 43503 962978
rect 42241 962920 42246 962976
rect 42302 962920 43442 962976
rect 43498 962920 43503 962976
rect 42241 962918 43503 962920
rect 42241 962915 42307 962918
rect 43437 962915 43503 962918
rect 62113 962978 62179 962981
rect 62113 962976 64492 962978
rect 62113 962920 62118 962976
rect 62174 962920 64492 962976
rect 62113 962918 64492 962920
rect 62113 962915 62179 962918
rect 673361 962842 673427 962845
rect 675477 962842 675543 962845
rect 673361 962840 675543 962842
rect 673361 962784 673366 962840
rect 673422 962784 675482 962840
rect 675538 962784 675543 962840
rect 673361 962782 675543 962784
rect 673361 962779 673427 962782
rect 675477 962779 675543 962782
rect 651465 962570 651531 962573
rect 650164 962568 651531 962570
rect 650164 962512 651470 962568
rect 651526 962512 651531 962568
rect 650164 962510 651531 962512
rect 651465 962507 651531 962510
rect 673085 962570 673151 962573
rect 674925 962570 674991 962573
rect 673085 962568 674991 962570
rect 673085 962512 673090 962568
rect 673146 962512 674930 962568
rect 674986 962512 674991 962568
rect 673085 962510 674991 962512
rect 673085 962507 673151 962510
rect 674925 962507 674991 962510
rect 41781 962164 41847 962165
rect 41781 962160 41828 962164
rect 41892 962162 41898 962164
rect 674649 962162 674715 962165
rect 675385 962162 675451 962165
rect 41781 962104 41786 962160
rect 41781 962100 41828 962104
rect 41892 962102 41938 962162
rect 674649 962160 675451 962162
rect 674649 962104 674654 962160
rect 674710 962104 675390 962160
rect 675446 962104 675451 962160
rect 674649 962102 675451 962104
rect 41892 962100 41898 962102
rect 41781 962099 41847 962100
rect 674649 962099 674715 962102
rect 675385 962099 675451 962102
rect 42241 962026 42307 962029
rect 44265 962026 44331 962029
rect 42241 962024 44331 962026
rect 42241 961968 42246 962024
rect 42302 961968 44270 962024
rect 44326 961968 44331 962024
rect 42241 961966 44331 961968
rect 42241 961963 42307 961966
rect 44265 961963 44331 961966
rect 41270 959788 41276 959852
rect 41340 959850 41346 959852
rect 41781 959850 41847 959853
rect 41340 959848 41847 959850
rect 41340 959792 41786 959848
rect 41842 959792 41847 959848
rect 41340 959790 41847 959792
rect 41340 959788 41346 959790
rect 41781 959787 41847 959790
rect 675201 959308 675267 959309
rect 675150 959306 675156 959308
rect 675110 959246 675156 959306
rect 675220 959304 675267 959308
rect 675262 959248 675267 959304
rect 675150 959244 675156 959246
rect 675220 959244 675267 959248
rect 675201 959243 675267 959244
rect 40534 959108 40540 959172
rect 40604 959170 40610 959172
rect 41781 959170 41847 959173
rect 40604 959168 41847 959170
rect 40604 959112 41786 959168
rect 41842 959112 41847 959168
rect 40604 959110 41847 959112
rect 40604 959108 40610 959110
rect 41781 959107 41847 959110
rect 42425 958762 42491 958765
rect 44449 958762 44515 958765
rect 42425 958760 44515 958762
rect 42425 958704 42430 958760
rect 42486 958704 44454 958760
rect 44510 958704 44515 958760
rect 42425 958702 44515 958704
rect 42425 958699 42491 958702
rect 44449 958699 44515 958702
rect 672901 958762 672967 958765
rect 675109 958762 675175 958765
rect 672901 958760 675175 958762
rect 672901 958704 672906 958760
rect 672962 958704 675114 958760
rect 675170 958704 675175 958760
rect 672901 958702 675175 958704
rect 672901 958699 672967 958702
rect 675109 958699 675175 958702
rect 41781 957812 41847 957813
rect 41781 957808 41828 957812
rect 41892 957810 41898 957812
rect 661677 957810 661743 957813
rect 675293 957810 675359 957813
rect 41781 957752 41786 957808
rect 41781 957748 41828 957752
rect 41892 957750 41938 957810
rect 661677 957808 675359 957810
rect 661677 957752 661682 957808
rect 661738 957752 675298 957808
rect 675354 957752 675359 957808
rect 661677 957750 675359 957752
rect 41892 957748 41898 957750
rect 41781 957747 41847 957748
rect 661677 957747 661743 957750
rect 675293 957747 675359 957750
rect 675753 957810 675819 957813
rect 676990 957810 676996 957812
rect 675753 957808 676996 957810
rect 675753 957752 675758 957808
rect 675814 957752 676996 957808
rect 675753 957750 676996 957752
rect 675753 957747 675819 957750
rect 676990 957748 676996 957750
rect 677060 957748 677066 957812
rect 674189 957130 674255 957133
rect 675477 957130 675543 957133
rect 674189 957128 675543 957130
rect 674189 957072 674194 957128
rect 674250 957072 675482 957128
rect 675538 957072 675543 957128
rect 674189 957070 675543 957072
rect 674189 957067 674255 957070
rect 675477 957067 675543 957070
rect 675753 956450 675819 956453
rect 676806 956450 676812 956452
rect 675753 956448 676812 956450
rect 675753 956392 675758 956448
rect 675814 956392 676812 956448
rect 675753 956390 676812 956392
rect 675753 956387 675819 956390
rect 676806 956388 676812 956390
rect 676876 956388 676882 956452
rect 40718 955436 40724 955500
rect 40788 955498 40794 955500
rect 41781 955498 41847 955501
rect 40788 955496 41847 955498
rect 40788 955440 41786 955496
rect 41842 955440 41847 955496
rect 40788 955438 41847 955440
rect 40788 955436 40794 955438
rect 41781 955435 41847 955438
rect 41781 954680 41847 954685
rect 41781 954624 41786 954680
rect 41842 954624 41847 954680
rect 41781 954619 41847 954624
rect 41784 954413 41844 954619
rect 675017 954546 675083 954549
rect 675334 954546 675340 954548
rect 675017 954544 675340 954546
rect 675017 954488 675022 954544
rect 675078 954488 675340 954544
rect 675017 954486 675340 954488
rect 675017 954483 675083 954486
rect 675334 954484 675340 954486
rect 675404 954484 675410 954548
rect 41781 954408 41847 954413
rect 41781 954352 41786 954408
rect 41842 954352 41847 954408
rect 41781 954347 41847 954352
rect 674833 953458 674899 953461
rect 675385 953458 675451 953461
rect 674833 953456 675451 953458
rect 674833 953400 674838 953456
rect 674894 953400 675390 953456
rect 675446 953400 675451 953456
rect 674833 953398 675451 953400
rect 674833 953395 674899 953398
rect 675385 953395 675451 953398
rect 35157 952914 35223 952917
rect 41822 952914 41828 952916
rect 35157 952912 41828 952914
rect 35157 952856 35162 952912
rect 35218 952856 41828 952912
rect 35157 952854 41828 952856
rect 35157 952851 35223 952854
rect 41822 952852 41828 952854
rect 41892 952852 41898 952916
rect 37917 952506 37983 952509
rect 41454 952506 41460 952508
rect 37917 952504 41460 952506
rect 37917 952448 37922 952504
rect 37978 952448 41460 952504
rect 37917 952446 41460 952448
rect 37917 952443 37983 952446
rect 41454 952444 41460 952446
rect 41524 952444 41530 952508
rect 39297 952234 39363 952237
rect 41638 952234 41644 952236
rect 39297 952232 41644 952234
rect 39297 952176 39302 952232
rect 39358 952176 41644 952232
rect 39297 952174 41644 952176
rect 39297 952171 39363 952174
rect 41638 952172 41644 952174
rect 41708 952172 41714 952236
rect 40033 951690 40099 951693
rect 41270 951690 41276 951692
rect 40033 951688 41276 951690
rect 40033 951632 40038 951688
rect 40094 951632 41276 951688
rect 40033 951630 41276 951632
rect 40033 951627 40099 951630
rect 41270 951628 41276 951630
rect 41340 951628 41346 951692
rect 676622 951492 676628 951556
rect 676692 951554 676698 951556
rect 677501 951554 677567 951557
rect 676692 951552 677567 951554
rect 676692 951496 677506 951552
rect 677562 951496 677567 951552
rect 676692 951494 677567 951496
rect 676692 951492 676698 951494
rect 677501 951491 677567 951494
rect 675201 951418 675267 951421
rect 675845 951418 675911 951421
rect 675201 951416 675911 951418
rect 675201 951360 675206 951416
rect 675262 951360 675850 951416
rect 675906 951360 675911 951416
rect 675201 951358 675911 951360
rect 675201 951355 675267 951358
rect 675845 951355 675911 951358
rect 675201 951148 675267 951149
rect 675150 951146 675156 951148
rect 675110 951086 675156 951146
rect 675220 951144 675267 951148
rect 675262 951088 675267 951144
rect 675150 951084 675156 951086
rect 675220 951084 675267 951088
rect 675201 951083 675267 951084
rect 676070 950676 676076 950740
rect 676140 950738 676146 950740
rect 678237 950738 678303 950741
rect 676140 950736 678303 950738
rect 676140 950680 678242 950736
rect 678298 950680 678303 950736
rect 676140 950678 678303 950680
rect 676140 950676 676146 950678
rect 678237 950675 678303 950678
rect 62113 949922 62179 949925
rect 62113 949920 64492 949922
rect 62113 949864 62118 949920
rect 62174 949864 64492 949920
rect 62113 949862 64492 949864
rect 62113 949859 62179 949862
rect 652201 949378 652267 949381
rect 650164 949376 652267 949378
rect 650164 949320 652206 949376
rect 652262 949320 652267 949376
rect 650164 949318 652267 949320
rect 652201 949315 652267 949318
rect 664437 947338 664503 947341
rect 683113 947338 683179 947341
rect 664437 947336 683179 947338
rect 664437 947280 664442 947336
rect 664498 947280 683118 947336
rect 683174 947280 683179 947336
rect 664437 947278 683179 947280
rect 664437 947275 664503 947278
rect 683113 947275 683179 947278
rect 31753 946658 31819 946661
rect 46197 946658 46263 946661
rect 31753 946656 46263 946658
rect 31753 946600 31758 946656
rect 31814 946600 46202 946656
rect 46258 946600 46263 946656
rect 31753 946598 46263 946600
rect 31753 946595 31819 946598
rect 46197 946595 46263 946598
rect 39757 943804 39823 943805
rect 39757 943800 39804 943804
rect 39868 943802 39874 943804
rect 39757 943744 39762 943800
rect 39757 943740 39804 943744
rect 39868 943742 39914 943802
rect 39868 943740 39874 943742
rect 40718 943740 40724 943804
rect 40788 943802 40794 943804
rect 42006 943802 42012 943804
rect 40788 943742 42012 943802
rect 40788 943740 40794 943742
rect 42006 943740 42012 943742
rect 42076 943740 42082 943804
rect 39757 943739 39823 943740
rect 45553 943530 45619 943533
rect 41492 943528 45619 943530
rect 41492 943472 45558 943528
rect 45614 943472 45619 943528
rect 41492 943470 45619 943472
rect 45553 943467 45619 943470
rect 35801 943122 35867 943125
rect 35788 943120 35867 943122
rect 35788 943064 35806 943120
rect 35862 943064 35867 943120
rect 35788 943062 35867 943064
rect 35801 943059 35867 943062
rect 28717 942714 28783 942717
rect 28717 942712 28796 942714
rect 28717 942656 28722 942712
rect 28778 942656 28796 942712
rect 28717 942654 28796 942656
rect 28717 942651 28783 942654
rect 51717 942306 51783 942309
rect 41492 942304 51783 942306
rect 41492 942248 51722 942304
rect 51778 942248 51783 942304
rect 41492 942246 51783 942248
rect 51717 942243 51783 942246
rect 35801 941898 35867 941901
rect 35788 941896 35867 941898
rect 35788 941840 35806 941896
rect 35862 941840 35867 941896
rect 35788 941838 35867 941840
rect 35801 941835 35867 941838
rect 663057 941762 663123 941765
rect 676213 941762 676279 941765
rect 663057 941760 676279 941762
rect 663057 941704 663062 941760
rect 663118 941704 676218 941760
rect 676274 941704 676279 941760
rect 663057 941702 676279 941704
rect 663057 941699 663123 941702
rect 676213 941699 676279 941702
rect 44817 941490 44883 941493
rect 41492 941488 44883 941490
rect 41492 941432 44822 941488
rect 44878 941432 44883 941488
rect 41492 941430 44883 941432
rect 44817 941427 44883 941430
rect 44633 941082 44699 941085
rect 41492 941080 44699 941082
rect 41492 941024 44638 941080
rect 44694 941024 44699 941080
rect 41492 941022 44699 941024
rect 44633 941019 44699 941022
rect 42057 940674 42123 940677
rect 41492 940672 42123 940674
rect 41492 940616 42062 940672
rect 42118 940616 42123 940672
rect 41492 940614 42123 940616
rect 42057 940611 42123 940614
rect 35801 940266 35867 940269
rect 35788 940264 35867 940266
rect 35788 940208 35806 940264
rect 35862 940208 35867 940264
rect 35788 940206 35867 940208
rect 35801 940203 35867 940206
rect 48957 940130 49023 940133
rect 41830 940128 49023 940130
rect 41830 940072 48962 940128
rect 49018 940072 49023 940128
rect 41830 940070 49023 940072
rect 41830 939858 41890 940070
rect 48957 940067 49023 940070
rect 41492 939798 41890 939858
rect 42057 939858 42123 939861
rect 50337 939858 50403 939861
rect 42057 939856 50403 939858
rect 42057 939800 42062 939856
rect 42118 939800 50342 939856
rect 50398 939800 50403 939856
rect 42057 939798 50403 939800
rect 42057 939795 42123 939798
rect 50337 939795 50403 939798
rect 665817 939858 665883 939861
rect 676262 939858 676322 939964
rect 665817 939856 676322 939858
rect 665817 939800 665822 939856
rect 665878 939800 676322 939856
rect 665817 939798 676322 939800
rect 665817 939795 665883 939798
rect 683113 939722 683179 939725
rect 683070 939720 683179 939722
rect 683070 939664 683118 939720
rect 683174 939664 683179 939720
rect 683070 939659 683179 939664
rect 683070 939556 683130 939659
rect 41776 939450 41782 939452
rect 41492 939390 41782 939450
rect 41776 939388 41782 939390
rect 41846 939388 41852 939452
rect 676213 939314 676279 939317
rect 676213 939312 676322 939314
rect 676213 939256 676218 939312
rect 676274 939256 676322 939312
rect 676213 939251 676322 939256
rect 676262 939148 676322 939251
rect 36537 939042 36603 939045
rect 36524 939040 36603 939042
rect 36524 938984 36542 939040
rect 36598 938984 36603 939040
rect 36524 938982 36603 938984
rect 36537 938979 36603 938982
rect 37917 938634 37983 938637
rect 37917 938632 37996 938634
rect 37917 938576 37922 938632
rect 37978 938576 37996 938632
rect 37917 938574 37996 938576
rect 37917 938571 37983 938574
rect 668577 938498 668643 938501
rect 676262 938498 676322 938740
rect 668577 938496 676322 938498
rect 668577 938440 668582 938496
rect 668638 938440 676322 938496
rect 668577 938438 676322 938440
rect 668577 938435 668643 938438
rect 33777 938226 33843 938229
rect 33764 938224 33843 938226
rect 33764 938168 33782 938224
rect 33838 938168 33843 938224
rect 33764 938166 33843 938168
rect 33777 938163 33843 938166
rect 676446 938093 676506 938332
rect 672165 938090 672231 938093
rect 672165 938088 676322 938090
rect 672165 938032 672170 938088
rect 672226 938032 676322 938088
rect 672165 938030 676322 938032
rect 676446 938088 676555 938093
rect 676446 938032 676494 938088
rect 676550 938032 676555 938088
rect 676446 938030 676555 938032
rect 672165 938027 672231 938030
rect 676262 937924 676322 938030
rect 676489 938027 676555 938030
rect 35157 937818 35223 937821
rect 667197 937818 667263 937821
rect 672809 937818 672875 937821
rect 676029 937818 676095 937821
rect 35157 937816 35236 937818
rect 35157 937760 35162 937816
rect 35218 937760 35236 937816
rect 35157 937758 35236 937760
rect 667197 937816 672458 937818
rect 667197 937760 667202 937816
rect 667258 937760 672458 937816
rect 667197 937758 672458 937760
rect 35157 937755 35223 937758
rect 667197 937755 667263 937758
rect 39297 937410 39363 937413
rect 39284 937408 39363 937410
rect 39284 937352 39302 937408
rect 39358 937352 39363 937408
rect 39284 937350 39363 937352
rect 39297 937347 39363 937350
rect 660297 937274 660363 937277
rect 672165 937274 672231 937277
rect 660297 937272 672231 937274
rect 660297 937216 660302 937272
rect 660358 937216 672170 937272
rect 672226 937216 672231 937272
rect 660297 937214 672231 937216
rect 672398 937274 672458 937758
rect 672809 937816 676095 937818
rect 672809 937760 672814 937816
rect 672870 937760 676034 937816
rect 676090 937760 676095 937816
rect 672809 937758 676095 937760
rect 672809 937755 672875 937758
rect 676029 937755 676095 937758
rect 672625 937546 672691 937549
rect 672625 937544 676292 937546
rect 672625 937488 672630 937544
rect 672686 937488 676292 937544
rect 672625 937486 676292 937488
rect 672625 937483 672691 937486
rect 672398 937214 676322 937274
rect 660297 937211 660363 937214
rect 672165 937211 672231 937214
rect 676262 937108 676322 937214
rect 42793 937002 42859 937005
rect 41492 937000 42859 937002
rect 41492 936944 42798 937000
rect 42854 936944 42859 937000
rect 41492 936942 42859 936944
rect 42793 936939 42859 936942
rect 41822 936730 41828 936732
rect 41784 936668 41828 936730
rect 41892 936668 41898 936732
rect 41784 936594 41844 936668
rect 41492 936534 41844 936594
rect 44449 936186 44515 936189
rect 41492 936184 44515 936186
rect 41492 936128 44454 936184
rect 44510 936128 44515 936184
rect 41492 936126 44515 936128
rect 44449 936123 44515 936126
rect 39757 935778 39823 935781
rect 64462 935778 64522 936836
rect 671797 936730 671863 936733
rect 671797 936728 676292 936730
rect 671797 936672 671802 936728
rect 671858 936672 676292 936728
rect 671797 936670 676292 936672
rect 671797 936667 671863 936670
rect 651465 936186 651531 936189
rect 650164 936184 651531 936186
rect 650164 936128 651470 936184
rect 651526 936128 651531 936184
rect 650164 936126 651531 936128
rect 651465 936123 651531 936126
rect 658917 936050 658983 936053
rect 676262 936050 676322 936292
rect 658917 936048 676322 936050
rect 658917 935992 658922 936048
rect 658978 935992 676322 936048
rect 658917 935990 676322 935992
rect 658917 935987 658983 935990
rect 39757 935776 39836 935778
rect 39757 935720 39762 935776
rect 39818 935720 39836 935776
rect 39757 935718 39836 935720
rect 48270 935718 64522 935778
rect 671613 935778 671679 935781
rect 676262 935778 676322 935884
rect 671613 935776 676322 935778
rect 671613 935720 671618 935776
rect 671674 935720 676322 935776
rect 671613 935718 676322 935720
rect 39757 935715 39823 935718
rect 41965 935642 42031 935645
rect 48270 935642 48330 935718
rect 671613 935715 671679 935718
rect 41965 935640 48330 935642
rect 41965 935584 41970 935640
rect 42026 935584 48330 935640
rect 41965 935582 48330 935584
rect 678237 935642 678303 935645
rect 678237 935640 678346 935642
rect 678237 935584 678242 935640
rect 678298 935584 678346 935640
rect 41965 935579 42031 935582
rect 678237 935579 678346 935584
rect 678286 935476 678346 935579
rect 43253 935370 43319 935373
rect 41492 935368 43319 935370
rect 41492 935312 43258 935368
rect 43314 935312 43319 935368
rect 41492 935310 43319 935312
rect 43253 935307 43319 935310
rect 682377 935234 682443 935237
rect 682334 935232 682443 935234
rect 682334 935176 682382 935232
rect 682438 935176 682443 935232
rect 682334 935171 682443 935176
rect 682334 935068 682394 935171
rect 43437 934962 43503 934965
rect 41492 934960 43503 934962
rect 41492 934904 43442 934960
rect 43498 934904 43503 934960
rect 41492 934902 43503 934904
rect 43437 934899 43503 934902
rect 673085 934690 673151 934693
rect 673085 934688 676292 934690
rect 673085 934632 673090 934688
rect 673146 934632 676292 934688
rect 673085 934630 676292 934632
rect 673085 934627 673151 934630
rect 40033 934554 40099 934557
rect 40020 934552 40099 934554
rect 40020 934496 40038 934552
rect 40094 934496 40099 934552
rect 40020 934494 40099 934496
rect 40033 934491 40099 934494
rect 675017 934282 675083 934285
rect 675017 934280 676292 934282
rect 675017 934224 675022 934280
rect 675078 934224 676292 934280
rect 675017 934222 676292 934224
rect 675017 934219 675083 934222
rect 44265 934146 44331 934149
rect 41492 934144 44331 934146
rect 41492 934088 44270 934144
rect 44326 934088 44331 934144
rect 41492 934086 44331 934088
rect 44265 934083 44331 934086
rect 675201 933874 675267 933877
rect 675201 933872 676292 933874
rect 675201 933816 675206 933872
rect 675262 933816 676292 933872
rect 675201 933814 676292 933816
rect 675201 933811 675267 933814
rect 42977 933738 43043 933741
rect 41492 933736 43043 933738
rect 41492 933680 42982 933736
rect 43038 933680 43043 933736
rect 41492 933678 43043 933680
rect 42977 933675 43043 933678
rect 680997 933602 681063 933605
rect 680997 933600 681106 933602
rect 680997 933544 681002 933600
rect 681058 933544 681106 933600
rect 680997 933539 681106 933544
rect 681046 933436 681106 933539
rect 43345 933330 43411 933333
rect 41492 933328 43411 933330
rect 41492 933272 43350 933328
rect 43406 933272 43411 933328
rect 41492 933270 43411 933272
rect 43345 933267 43411 933270
rect 674373 933058 674439 933061
rect 674373 933056 676292 933058
rect 674373 933000 674378 933056
rect 674434 933000 676292 933056
rect 674373 932998 676292 933000
rect 674373 932995 674439 932998
rect 42333 932922 42399 932925
rect 41492 932920 42399 932922
rect 41492 932864 42338 932920
rect 42394 932864 42399 932920
rect 41492 932862 42399 932864
rect 42333 932859 42399 932862
rect 673361 932650 673427 932653
rect 673361 932648 676292 932650
rect 673361 932592 673366 932648
rect 673422 932592 676292 932648
rect 673361 932590 676292 932592
rect 673361 932587 673427 932590
rect 674649 932242 674715 932245
rect 674649 932240 676292 932242
rect 674649 932184 674654 932240
rect 674710 932184 676292 932240
rect 674649 932182 676292 932184
rect 674649 932179 674715 932182
rect 43529 932106 43595 932109
rect 41492 932104 43595 932106
rect 41492 932048 43534 932104
rect 43590 932048 43595 932104
rect 41492 932046 43595 932048
rect 43529 932043 43595 932046
rect 676806 931908 676812 931972
rect 676876 931908 676882 931972
rect 676814 931804 676874 931908
rect 676990 931500 676996 931564
rect 677060 931500 677066 931564
rect 676998 931396 677058 931500
rect 677501 931154 677567 931157
rect 677501 931152 677610 931154
rect 677501 931096 677506 931152
rect 677562 931096 677610 931152
rect 677501 931091 677610 931096
rect 677550 930988 677610 931091
rect 673085 930610 673151 930613
rect 673085 930608 676292 930610
rect 673085 930552 673090 930608
rect 673146 930552 676292 930608
rect 673085 930550 676292 930552
rect 673085 930547 673151 930550
rect 674189 930202 674255 930205
rect 674189 930200 676292 930202
rect 674189 930144 674194 930200
rect 674250 930144 676292 930200
rect 674189 930142 676292 930144
rect 674189 930139 674255 930142
rect 673361 929522 673427 929525
rect 676262 929522 676322 929764
rect 673361 929520 676322 929522
rect 673361 929464 673366 929520
rect 673422 929464 676322 929520
rect 673361 929462 676322 929464
rect 673361 929459 673427 929462
rect 682886 929114 682946 929356
rect 683113 929114 683179 929117
rect 682886 929112 683179 929114
rect 682886 929056 683118 929112
rect 683174 929056 683179 929112
rect 682886 929054 683179 929056
rect 682886 928948 682946 929054
rect 683113 929051 683179 929054
rect 671981 928298 672047 928301
rect 676262 928298 676322 928540
rect 671981 928296 676322 928298
rect 671981 928240 671986 928296
rect 672042 928240 676322 928296
rect 671981 928238 676322 928240
rect 671981 928235 672047 928238
rect 62113 923810 62179 923813
rect 62113 923808 64492 923810
rect 62113 923752 62118 923808
rect 62174 923752 64492 923808
rect 62113 923750 64492 923752
rect 62113 923747 62179 923750
rect 651465 922722 651531 922725
rect 650164 922720 651531 922722
rect 650164 922664 651470 922720
rect 651526 922664 651531 922720
rect 650164 922662 651531 922664
rect 651465 922659 651531 922662
rect 41597 911978 41663 911981
rect 42006 911978 42012 911980
rect 41597 911976 42012 911978
rect 41597 911920 41602 911976
rect 41658 911920 42012 911976
rect 41597 911918 42012 911920
rect 41597 911915 41663 911918
rect 42006 911916 42012 911918
rect 42076 911916 42082 911980
rect 41413 911706 41479 911709
rect 42190 911706 42196 911708
rect 41413 911704 42196 911706
rect 41413 911648 41418 911704
rect 41474 911648 42196 911704
rect 41413 911646 42196 911648
rect 41413 911643 41479 911646
rect 42190 911644 42196 911646
rect 42260 911644 42266 911708
rect 62113 910754 62179 910757
rect 62113 910752 64492 910754
rect 62113 910696 62118 910752
rect 62174 910696 64492 910752
rect 62113 910694 64492 910696
rect 62113 910691 62179 910694
rect 652385 909530 652451 909533
rect 650164 909528 652451 909530
rect 650164 909472 652390 909528
rect 652446 909472 652451 909528
rect 650164 909470 652451 909472
rect 652385 909467 652451 909470
rect 62113 897834 62179 897837
rect 62113 897832 64492 897834
rect 62113 897776 62118 897832
rect 62174 897776 64492 897832
rect 62113 897774 64492 897776
rect 62113 897771 62179 897774
rect 651465 896202 651531 896205
rect 650164 896200 651531 896202
rect 650164 896144 651470 896200
rect 651526 896144 651531 896200
rect 650164 896142 651531 896144
rect 651465 896139 651531 896142
rect 43069 892802 43135 892805
rect 53281 892802 53347 892805
rect 43069 892800 53347 892802
rect 43069 892744 43074 892800
rect 43130 892744 53286 892800
rect 53342 892744 53347 892800
rect 43069 892742 53347 892744
rect 43069 892739 43135 892742
rect 53281 892739 53347 892742
rect 42839 892530 42905 892533
rect 42839 892528 55230 892530
rect 42839 892472 42844 892528
rect 42900 892472 55230 892528
rect 42839 892470 55230 892472
rect 42839 892467 42905 892470
rect 42931 892258 42997 892261
rect 54477 892258 54543 892261
rect 42931 892256 54543 892258
rect 42931 892200 42936 892256
rect 42992 892200 54482 892256
rect 54538 892200 54543 892256
rect 42931 892198 54543 892200
rect 55170 892258 55230 892470
rect 55857 892258 55923 892261
rect 55170 892256 55923 892258
rect 55170 892200 55862 892256
rect 55918 892200 55923 892256
rect 55170 892198 55923 892200
rect 42931 892195 42997 892198
rect 54477 892195 54543 892198
rect 55857 892195 55923 892198
rect 44081 891986 44147 891989
rect 47577 891986 47643 891989
rect 44081 891984 47643 891986
rect 44081 891928 44086 891984
rect 44142 891928 47582 891984
rect 47638 891928 47643 891984
rect 44081 891926 47643 891928
rect 44081 891923 44147 891926
rect 47577 891923 47643 891926
rect 41597 885458 41663 885461
rect 42006 885458 42012 885460
rect 41597 885456 42012 885458
rect 41597 885400 41602 885456
rect 41658 885400 42012 885456
rect 41597 885398 42012 885400
rect 41597 885395 41663 885398
rect 42006 885396 42012 885398
rect 42076 885396 42082 885460
rect 41413 885186 41479 885189
rect 42190 885186 42196 885188
rect 41413 885184 42196 885186
rect 41413 885128 41418 885184
rect 41474 885128 42196 885184
rect 41413 885126 42196 885128
rect 41413 885123 41479 885126
rect 42190 885124 42196 885126
rect 42260 885124 42266 885188
rect 45510 884718 64492 884778
rect 42057 884642 42123 884645
rect 45510 884642 45570 884718
rect 42057 884640 45570 884642
rect 42057 884584 42062 884640
rect 42118 884584 45570 884640
rect 42057 884582 45570 884584
rect 42057 884579 42123 884582
rect 651649 882874 651715 882877
rect 650164 882872 651715 882874
rect 650164 882816 651654 882872
rect 651710 882816 651715 882872
rect 650164 882814 651715 882816
rect 651649 882811 651715 882814
rect 669221 879202 669287 879205
rect 675293 879202 675359 879205
rect 669221 879200 675359 879202
rect 669221 879144 669226 879200
rect 669282 879144 675298 879200
rect 675354 879144 675359 879200
rect 669221 879142 675359 879144
rect 669221 879139 669287 879142
rect 675293 879139 675359 879142
rect 675753 875938 675819 875941
rect 676070 875938 676076 875940
rect 675753 875936 676076 875938
rect 675753 875880 675758 875936
rect 675814 875880 676076 875936
rect 675753 875878 676076 875880
rect 675753 875875 675819 875878
rect 676070 875876 676076 875878
rect 676140 875876 676146 875940
rect 675385 874036 675451 874037
rect 675334 874034 675340 874036
rect 675294 873974 675340 874034
rect 675404 874032 675451 874036
rect 675446 873976 675451 874032
rect 675334 873972 675340 873974
rect 675404 873972 675451 873976
rect 675385 873971 675451 873972
rect 672533 873626 672599 873629
rect 675385 873626 675451 873629
rect 672533 873624 675451 873626
rect 672533 873568 672538 873624
rect 672594 873568 675390 873624
rect 675446 873568 675451 873624
rect 672533 873566 675451 873568
rect 672533 873563 672599 873566
rect 675385 873563 675451 873566
rect 673862 873156 673868 873220
rect 673932 873218 673938 873220
rect 675109 873218 675175 873221
rect 673932 873216 675175 873218
rect 673932 873160 675114 873216
rect 675170 873160 675175 873216
rect 673932 873158 675175 873160
rect 673932 873156 673938 873158
rect 675109 873155 675175 873158
rect 671153 872266 671219 872269
rect 675385 872266 675451 872269
rect 671153 872264 675451 872266
rect 671153 872208 671158 872264
rect 671214 872208 675390 872264
rect 675446 872208 675451 872264
rect 671153 872206 675451 872208
rect 671153 872203 671219 872206
rect 675385 872203 675451 872206
rect 62113 871722 62179 871725
rect 62113 871720 64492 871722
rect 62113 871664 62118 871720
rect 62174 871664 64492 871720
rect 62113 871662 64492 871664
rect 62113 871659 62179 871662
rect 674925 870906 674991 870909
rect 676990 870906 676996 870908
rect 674925 870904 676996 870906
rect 674925 870848 674930 870904
rect 674986 870848 676996 870904
rect 674925 870846 676996 870848
rect 674925 870843 674991 870846
rect 676990 870844 676996 870846
rect 677060 870844 677066 870908
rect 672993 870090 673059 870093
rect 675109 870090 675175 870093
rect 672993 870088 675175 870090
rect 672993 870032 672998 870088
rect 673054 870032 675114 870088
rect 675170 870032 675175 870088
rect 672993 870030 675175 870032
rect 672993 870027 673059 870030
rect 675109 870027 675175 870030
rect 651465 869682 651531 869685
rect 650164 869680 651531 869682
rect 650164 869624 651470 869680
rect 651526 869624 651531 869680
rect 650164 869622 651531 869624
rect 651465 869619 651531 869622
rect 664437 868730 664503 868733
rect 664437 868728 669330 868730
rect 664437 868672 664442 868728
rect 664498 868672 669330 868728
rect 664437 868670 669330 868672
rect 664437 868667 664503 868670
rect 669270 868458 669330 868670
rect 675293 868458 675359 868461
rect 669270 868456 675359 868458
rect 669270 868400 675298 868456
rect 675354 868400 675359 868456
rect 669270 868398 675359 868400
rect 675293 868395 675359 868398
rect 668209 868186 668275 868189
rect 674833 868186 674899 868189
rect 668209 868184 674899 868186
rect 668209 868128 668214 868184
rect 668270 868128 674838 868184
rect 674894 868128 674899 868184
rect 668209 868126 674899 868128
rect 668209 868123 668275 868126
rect 674833 868123 674899 868126
rect 670601 867914 670667 867917
rect 675477 867914 675543 867917
rect 670601 867912 675543 867914
rect 670601 867856 670606 867912
rect 670662 867856 675482 867912
rect 675538 867856 675543 867912
rect 670601 867854 675543 867856
rect 670601 867851 670667 867854
rect 675477 867851 675543 867854
rect 674833 867506 674899 867509
rect 675477 867506 675543 867509
rect 674833 867504 675543 867506
rect 674833 867448 674838 867504
rect 674894 867448 675482 867504
rect 675538 867448 675543 867504
rect 674833 867446 675543 867448
rect 674833 867443 674899 867446
rect 675477 867443 675543 867446
rect 673913 864922 673979 864925
rect 675385 864922 675451 864925
rect 673913 864920 675451 864922
rect 673913 864864 673918 864920
rect 673974 864864 675390 864920
rect 675446 864864 675451 864920
rect 673913 864862 675451 864864
rect 673913 864859 673979 864862
rect 675385 864859 675451 864862
rect 669773 864242 669839 864245
rect 675477 864242 675543 864245
rect 669773 864240 675543 864242
rect 669773 864184 669778 864240
rect 669834 864184 675482 864240
rect 675538 864184 675543 864240
rect 669773 864182 675543 864184
rect 669773 864179 669839 864182
rect 675477 864179 675543 864182
rect 675293 863156 675359 863157
rect 675293 863154 675340 863156
rect 675248 863152 675340 863154
rect 675248 863096 675298 863152
rect 675248 863094 675340 863096
rect 675293 863092 675340 863094
rect 675404 863092 675410 863156
rect 675293 863091 675359 863092
rect 62757 858666 62823 858669
rect 62757 858664 64492 858666
rect 62757 858608 62762 858664
rect 62818 858608 64492 858664
rect 62757 858606 64492 858608
rect 62757 858603 62823 858606
rect 652385 856354 652451 856357
rect 650164 856352 652451 856354
rect 650164 856296 652390 856352
rect 652446 856296 652451 856352
rect 650164 856294 652451 856296
rect 652385 856291 652451 856294
rect 62113 845610 62179 845613
rect 62113 845608 64492 845610
rect 62113 845552 62118 845608
rect 62174 845552 64492 845608
rect 62113 845550 64492 845552
rect 62113 845547 62179 845550
rect 652017 843026 652083 843029
rect 650164 843024 652083 843026
rect 650164 842968 652022 843024
rect 652078 842968 652083 843024
rect 650164 842966 652083 842968
rect 652017 842963 652083 842966
rect 62113 832554 62179 832557
rect 62113 832552 64492 832554
rect 62113 832496 62118 832552
rect 62174 832496 64492 832552
rect 62113 832494 64492 832496
rect 62113 832491 62179 832494
rect 651465 829834 651531 829837
rect 650164 829832 651531 829834
rect 650164 829776 651470 829832
rect 651526 829776 651531 829832
rect 650164 829774 651531 829776
rect 651465 829771 651531 829774
rect 62113 819498 62179 819501
rect 62113 819496 64492 819498
rect 62113 819440 62118 819496
rect 62174 819440 64492 819496
rect 62113 819438 64492 819440
rect 62113 819435 62179 819438
rect 47761 817730 47827 817733
rect 41492 817728 47827 817730
rect 41492 817672 47766 817728
rect 47822 817672 47827 817728
rect 41492 817670 47827 817672
rect 47761 817667 47827 817670
rect 35801 817322 35867 817325
rect 35788 817320 35867 817322
rect 35788 817264 35806 817320
rect 35862 817264 35867 817320
rect 35788 817262 35867 817264
rect 35801 817259 35867 817262
rect 50337 816914 50403 816917
rect 41492 816912 50403 816914
rect 41492 816856 50342 816912
rect 50398 816856 50403 816912
rect 41492 816854 50403 816856
rect 50337 816851 50403 816854
rect 35801 816506 35867 816509
rect 651465 816506 651531 816509
rect 35788 816504 35867 816506
rect 35788 816448 35806 816504
rect 35862 816448 35867 816504
rect 35788 816446 35867 816448
rect 650164 816504 651531 816506
rect 650164 816448 651470 816504
rect 651526 816448 651531 816504
rect 650164 816446 651531 816448
rect 35801 816443 35867 816446
rect 651465 816443 651531 816446
rect 44357 816098 44423 816101
rect 41492 816096 44423 816098
rect 41492 816040 44362 816096
rect 44418 816040 44423 816096
rect 41492 816038 44423 816040
rect 44357 816035 44423 816038
rect 44633 815690 44699 815693
rect 41492 815688 44699 815690
rect 41492 815632 44638 815688
rect 44694 815632 44699 815688
rect 41492 815630 44699 815632
rect 44633 815627 44699 815630
rect 44817 815282 44883 815285
rect 41492 815280 44883 815282
rect 41492 815224 44822 815280
rect 44878 815224 44883 815280
rect 41492 815222 44883 815224
rect 44817 815219 44883 815222
rect 35801 814874 35867 814877
rect 35788 814872 35867 814874
rect 35788 814816 35806 814872
rect 35862 814816 35867 814872
rect 35788 814814 35867 814816
rect 35801 814811 35867 814814
rect 44173 814466 44239 814469
rect 41492 814464 44239 814466
rect 41492 814408 44178 814464
rect 44234 814408 44239 814464
rect 41492 814406 44239 814408
rect 44173 814403 44239 814406
rect 39982 814234 39988 814298
rect 40052 814234 40058 814298
rect 39990 814028 40050 814234
rect 45001 813650 45067 813653
rect 41492 813648 45067 813650
rect 41492 813592 45006 813648
rect 45062 813592 45067 813648
rect 41492 813590 45067 813592
rect 45001 813587 45067 813590
rect 41822 813242 41828 813244
rect 41492 813182 41828 813242
rect 41822 813180 41828 813182
rect 41892 813180 41898 813244
rect 41321 812834 41387 812837
rect 41308 812832 41387 812834
rect 41308 812776 41326 812832
rect 41382 812776 41387 812832
rect 41308 812774 41387 812776
rect 41321 812771 41387 812774
rect 40953 812426 41019 812429
rect 40940 812424 41019 812426
rect 40940 812368 40958 812424
rect 41014 812368 41019 812424
rect 40940 812366 41019 812368
rect 40953 812363 41019 812366
rect 41137 812018 41203 812021
rect 41124 812016 41203 812018
rect 41124 811960 41142 812016
rect 41198 811960 41203 812016
rect 41124 811958 41203 811960
rect 41137 811955 41203 811958
rect 35157 811610 35223 811613
rect 35157 811608 35236 811610
rect 35157 811552 35162 811608
rect 35218 811552 35236 811608
rect 35157 811550 35236 811552
rect 35157 811547 35223 811550
rect 35893 811202 35959 811205
rect 35893 811200 35972 811202
rect 35893 811144 35898 811200
rect 35954 811144 35972 811200
rect 35893 811142 35972 811144
rect 35893 811139 35959 811142
rect 43161 810794 43227 810797
rect 41492 810792 43227 810794
rect 41492 810736 43166 810792
rect 43222 810736 43227 810792
rect 41492 810734 43227 810736
rect 43161 810731 43227 810734
rect 44541 810386 44607 810389
rect 41492 810384 44607 810386
rect 41492 810328 44546 810384
rect 44602 810328 44607 810384
rect 41492 810326 44607 810328
rect 44541 810323 44607 810326
rect 42793 809978 42859 809981
rect 41492 809976 42859 809978
rect 41492 809920 42798 809976
rect 42854 809920 42859 809976
rect 41492 809918 42859 809920
rect 42793 809915 42859 809918
rect 43897 809570 43963 809573
rect 41492 809568 43963 809570
rect 41492 809512 43902 809568
rect 43958 809512 43963 809568
rect 41492 809510 43963 809512
rect 43897 809507 43963 809510
rect 41822 809162 41828 809164
rect 41492 809102 41828 809162
rect 41822 809100 41828 809102
rect 41892 809100 41898 809164
rect 41781 808754 41847 808757
rect 41492 808752 41847 808754
rect 41492 808696 41786 808752
rect 41842 808696 41847 808752
rect 41492 808694 41847 808696
rect 41781 808691 41847 808694
rect 40769 808346 40835 808349
rect 40756 808344 40835 808346
rect 40756 808288 40774 808344
rect 40830 808288 40835 808344
rect 40756 808286 40835 808288
rect 40769 808283 40835 808286
rect 45185 807938 45251 807941
rect 41492 807936 45251 807938
rect 41492 807880 45190 807936
rect 45246 807880 45251 807936
rect 41492 807878 45251 807880
rect 45185 807875 45251 807878
rect 42977 807530 43043 807533
rect 41308 807528 43043 807530
rect 41308 807472 42982 807528
rect 43038 807472 43043 807528
rect 41308 807470 43043 807472
rect 42977 807467 43043 807470
rect 41462 806714 41522 807092
rect 42333 806714 42399 806717
rect 41462 806712 42399 806714
rect 41462 806684 42338 806712
rect 41492 806656 42338 806684
rect 42394 806656 42399 806712
rect 41492 806654 42399 806656
rect 42333 806651 42399 806654
rect 62113 806578 62179 806581
rect 62113 806576 64492 806578
rect 62113 806520 62118 806576
rect 62174 806520 64492 806576
rect 62113 806518 64492 806520
rect 62113 806515 62179 806518
rect 43713 806306 43779 806309
rect 41492 806304 43779 806306
rect 41492 806248 43718 806304
rect 43774 806248 43779 806304
rect 41492 806246 43779 806248
rect 43713 806243 43779 806246
rect 40902 805428 40908 805492
rect 40972 805490 40978 805492
rect 41822 805490 41828 805492
rect 40972 805430 41828 805490
rect 40972 805428 40978 805430
rect 41822 805428 41828 805430
rect 41892 805428 41898 805492
rect 40585 805220 40651 805221
rect 40534 805218 40540 805220
rect 40494 805158 40540 805218
rect 40604 805216 40651 805220
rect 40646 805160 40651 805216
rect 40534 805156 40540 805158
rect 40604 805156 40651 805160
rect 40585 805155 40651 805156
rect 40769 805084 40835 805085
rect 40718 805020 40724 805084
rect 40788 805082 40835 805084
rect 40788 805080 40880 805082
rect 40830 805024 40880 805080
rect 40788 805022 40880 805024
rect 40788 805020 40835 805022
rect 40769 805019 40835 805020
rect 40953 804810 41019 804813
rect 41638 804810 41644 804812
rect 40953 804808 41644 804810
rect 40953 804752 40958 804808
rect 41014 804752 41644 804808
rect 40953 804750 41644 804752
rect 40953 804747 41019 804750
rect 41638 804748 41644 804750
rect 41708 804748 41714 804812
rect 41137 804538 41203 804541
rect 42006 804538 42012 804540
rect 41137 804536 42012 804538
rect 41137 804480 41142 804536
rect 41198 804480 42012 804536
rect 41137 804478 42012 804480
rect 41137 804475 41203 804478
rect 42006 804476 42012 804478
rect 42076 804476 42082 804540
rect 651465 803314 651531 803317
rect 650164 803312 651531 803314
rect 650164 803256 651470 803312
rect 651526 803256 651531 803312
rect 650164 803254 651531 803256
rect 651465 803251 651531 803254
rect 41689 802498 41755 802501
rect 42609 802498 42675 802501
rect 41689 802496 42675 802498
rect 41689 802440 41694 802496
rect 41750 802440 42614 802496
rect 42670 802440 42675 802496
rect 41689 802438 42675 802440
rect 41689 802435 41755 802438
rect 42609 802435 42675 802438
rect 41781 800320 41847 800325
rect 41781 800264 41786 800320
rect 41842 800264 41847 800320
rect 41781 800259 41847 800264
rect 41784 799917 41844 800259
rect 41781 799912 41847 799917
rect 41781 799856 41786 799912
rect 41842 799856 41847 799912
rect 41781 799851 41847 799856
rect 53097 799234 53163 799237
rect 51030 799232 53163 799234
rect 51030 799176 53102 799232
rect 53158 799176 53163 799232
rect 51030 799174 53163 799176
rect 51030 799098 51090 799174
rect 53097 799171 53163 799174
rect 42428 799038 51090 799098
rect 42241 798964 42307 798965
rect 42190 798962 42196 798964
rect 42150 798902 42196 798962
rect 42260 798960 42307 798964
rect 42302 798904 42307 798960
rect 42190 798900 42196 798902
rect 42260 798900 42307 798904
rect 42241 798899 42307 798900
rect 42428 798149 42488 799038
rect 42425 798144 42491 798149
rect 42425 798088 42430 798144
rect 42486 798088 42491 798144
rect 42425 798083 42491 798088
rect 42149 797876 42215 797877
rect 42149 797874 42196 797876
rect 42104 797872 42196 797874
rect 42104 797816 42154 797872
rect 42104 797814 42196 797816
rect 42149 797812 42196 797814
rect 42260 797812 42266 797876
rect 42149 797811 42215 797812
rect 43897 797738 43963 797741
rect 42382 797736 43963 797738
rect 42382 797680 43902 797736
rect 43958 797680 43963 797736
rect 42382 797678 43963 797680
rect 42382 797197 42442 797678
rect 43897 797675 43963 797678
rect 42333 797192 42442 797197
rect 42333 797136 42338 797192
rect 42394 797136 42442 797192
rect 42333 797134 42442 797136
rect 42333 797131 42399 797134
rect 674833 796922 674899 796925
rect 675201 796922 675267 796925
rect 674833 796920 675267 796922
rect 674833 796864 674838 796920
rect 674894 796864 675206 796920
rect 675262 796864 675267 796920
rect 674833 796862 675267 796864
rect 674833 796859 674899 796862
rect 675201 796859 675267 796862
rect 42425 796786 42491 796789
rect 45185 796786 45251 796789
rect 42425 796784 45251 796786
rect 42425 796728 42430 796784
rect 42486 796728 45190 796784
rect 45246 796728 45251 796784
rect 42425 796726 45251 796728
rect 42425 796723 42491 796726
rect 45185 796723 45251 796726
rect 40718 794956 40724 795020
rect 40788 795018 40794 795020
rect 40788 794958 42258 795018
rect 40788 794956 40794 794958
rect 42198 794882 42258 794958
rect 42425 794882 42491 794885
rect 42198 794880 42491 794882
rect 42198 794824 42430 794880
rect 42486 794824 42491 794880
rect 42198 794822 42491 794824
rect 42425 794819 42491 794822
rect 40902 794140 40908 794204
rect 40972 794202 40978 794204
rect 41781 794202 41847 794205
rect 40972 794200 41847 794202
rect 40972 794144 41786 794200
rect 41842 794144 41847 794200
rect 40972 794142 41847 794144
rect 40972 794140 40978 794142
rect 41781 794139 41847 794142
rect 62941 793658 63007 793661
rect 62941 793656 64492 793658
rect 62941 793600 62946 793656
rect 63002 793600 64492 793656
rect 62941 793598 64492 793600
rect 62941 793595 63007 793598
rect 40534 792508 40540 792572
rect 40604 792570 40610 792572
rect 42241 792570 42307 792573
rect 40604 792568 42307 792570
rect 40604 792512 42246 792568
rect 42302 792512 42307 792568
rect 40604 792510 42307 792512
rect 40604 792508 40610 792510
rect 42241 792507 42307 792510
rect 651465 789986 651531 789989
rect 650164 789984 651531 789986
rect 650164 789928 651470 789984
rect 651526 789928 651531 789984
rect 650164 789926 651531 789928
rect 651465 789923 651531 789926
rect 669589 789442 669655 789445
rect 675201 789442 675267 789445
rect 669589 789440 675267 789442
rect 669589 789384 669594 789440
rect 669650 789384 675206 789440
rect 675262 789384 675267 789440
rect 669589 789382 675267 789384
rect 669589 789379 669655 789382
rect 675201 789379 675267 789382
rect 42149 789306 42215 789309
rect 44541 789306 44607 789309
rect 42149 789304 44607 789306
rect 42149 789248 42154 789304
rect 42210 789248 44546 789304
rect 44602 789248 44607 789304
rect 42149 789246 44607 789248
rect 42149 789243 42215 789246
rect 44541 789243 44607 789246
rect 41638 788972 41644 789036
rect 41708 789034 41714 789036
rect 42701 789034 42767 789037
rect 41708 789032 42767 789034
rect 41708 788976 42706 789032
rect 42762 788976 42767 789032
rect 41708 788974 42767 788976
rect 41708 788972 41714 788974
rect 42701 788971 42767 788974
rect 41781 788628 41847 788629
rect 41781 788624 41828 788628
rect 41892 788626 41898 788628
rect 42793 788626 42859 788629
rect 62757 788626 62823 788629
rect 41781 788568 41786 788624
rect 41781 788564 41828 788568
rect 41892 788566 41938 788626
rect 42793 788624 62823 788626
rect 42793 788568 42798 788624
rect 42854 788568 62762 788624
rect 62818 788568 62823 788624
rect 42793 788566 62823 788568
rect 41892 788564 41898 788566
rect 41781 788563 41847 788564
rect 42793 788563 42859 788566
rect 62757 788563 62823 788566
rect 42241 788218 42307 788221
rect 43161 788218 43227 788221
rect 42241 788216 43227 788218
rect 42241 788160 42246 788216
rect 42302 788160 43166 788216
rect 43222 788160 43227 788216
rect 42241 788158 43227 788160
rect 42241 788155 42307 788158
rect 43161 788155 43227 788158
rect 674465 788082 674531 788085
rect 675385 788082 675451 788085
rect 674465 788080 675451 788082
rect 674465 788024 674470 788080
rect 674526 788024 675390 788080
rect 675446 788024 675451 788080
rect 674465 788022 675451 788024
rect 674465 788019 674531 788022
rect 675385 788019 675451 788022
rect 41454 786796 41460 786860
rect 41524 786858 41530 786860
rect 41781 786858 41847 786861
rect 41524 786856 41847 786858
rect 41524 786800 41786 786856
rect 41842 786800 41847 786856
rect 41524 786798 41847 786800
rect 41524 786796 41530 786798
rect 41781 786795 41847 786798
rect 667749 786722 667815 786725
rect 675293 786722 675359 786725
rect 667749 786720 675359 786722
rect 667749 786664 667754 786720
rect 667810 786664 675298 786720
rect 675354 786664 675359 786720
rect 667749 786662 675359 786664
rect 667749 786659 667815 786662
rect 675293 786659 675359 786662
rect 672349 784410 672415 784413
rect 675385 784410 675451 784413
rect 672349 784408 675451 784410
rect 672349 784352 672354 784408
rect 672410 784352 675390 784408
rect 675446 784352 675451 784408
rect 672349 784350 675451 784352
rect 672349 784347 672415 784350
rect 675385 784347 675451 784350
rect 674833 784138 674899 784141
rect 675293 784138 675359 784141
rect 674833 784136 675359 784138
rect 674833 784080 674838 784136
rect 674894 784080 675298 784136
rect 675354 784080 675359 784136
rect 674833 784078 675359 784080
rect 674833 784075 674899 784078
rect 675293 784075 675359 784078
rect 668393 783866 668459 783869
rect 675477 783866 675543 783869
rect 668393 783864 675543 783866
rect 668393 783808 668398 783864
rect 668454 783808 675482 783864
rect 675538 783808 675543 783864
rect 668393 783806 675543 783808
rect 668393 783803 668459 783806
rect 675477 783803 675543 783806
rect 670325 783050 670391 783053
rect 675477 783050 675543 783053
rect 670325 783048 675543 783050
rect 670325 782992 670330 783048
rect 670386 782992 675482 783048
rect 675538 782992 675543 783048
rect 670325 782990 675543 782992
rect 670325 782987 670391 782990
rect 675477 782987 675543 782990
rect 670141 780738 670207 780741
rect 675477 780738 675543 780741
rect 670141 780736 675543 780738
rect 670141 780680 670146 780736
rect 670202 780680 675482 780736
rect 675538 780680 675543 780736
rect 670141 780678 675543 780680
rect 670141 780675 670207 780678
rect 675477 780675 675543 780678
rect 62757 780466 62823 780469
rect 62757 780464 64492 780466
rect 62757 780408 62762 780464
rect 62818 780408 64492 780464
rect 62757 780406 64492 780408
rect 62757 780403 62823 780406
rect 674281 780058 674347 780061
rect 675477 780058 675543 780061
rect 674281 780056 675543 780058
rect 674281 780000 674286 780056
rect 674342 780000 675482 780056
rect 675538 780000 675543 780056
rect 674281 779998 675543 780000
rect 674281 779995 674347 779998
rect 675477 779995 675543 779998
rect 673729 779378 673795 779381
rect 675477 779378 675543 779381
rect 673729 779376 675543 779378
rect 673729 779320 673734 779376
rect 673790 779320 675482 779376
rect 675538 779320 675543 779376
rect 673729 779318 675543 779320
rect 673729 779315 673795 779318
rect 675477 779315 675543 779318
rect 660297 778970 660363 778973
rect 674833 778970 674899 778973
rect 660297 778968 674899 778970
rect 660297 778912 660302 778968
rect 660358 778912 674838 778968
rect 674894 778912 674899 778968
rect 660297 778910 674899 778912
rect 660297 778907 660363 778910
rect 674833 778907 674899 778910
rect 670969 778698 671035 778701
rect 675477 778698 675543 778701
rect 670969 778696 675543 778698
rect 670969 778640 670974 778696
rect 671030 778640 675482 778696
rect 675538 778640 675543 778696
rect 670969 778638 675543 778640
rect 670969 778635 671035 778638
rect 675477 778635 675543 778638
rect 673545 777474 673611 777477
rect 675477 777474 675543 777477
rect 673545 777472 675543 777474
rect 673545 777416 673550 777472
rect 673606 777416 675482 777472
rect 675538 777416 675543 777472
rect 673545 777414 675543 777416
rect 673545 777411 673611 777414
rect 675477 777411 675543 777414
rect 666277 777066 666343 777069
rect 675702 777066 675708 777068
rect 666277 777064 675708 777066
rect 666277 777008 666282 777064
rect 666338 777008 675708 777064
rect 666277 777006 675708 777008
rect 666277 777003 666343 777006
rect 675702 777004 675708 777006
rect 675772 777004 675778 777068
rect 651465 776658 651531 776661
rect 650164 776656 651531 776658
rect 650164 776600 651470 776656
rect 651526 776600 651531 776656
rect 650164 776598 651531 776600
rect 651465 776595 651531 776598
rect 674833 776522 674899 776525
rect 675477 776522 675543 776525
rect 674833 776520 675543 776522
rect 674833 776464 674838 776520
rect 674894 776464 675482 776520
rect 675538 776464 675543 776520
rect 674833 776462 675543 776464
rect 674833 776459 674899 776462
rect 675477 776459 675543 776462
rect 674833 775842 674899 775845
rect 675477 775842 675543 775845
rect 674833 775840 675543 775842
rect 674833 775784 674838 775840
rect 674894 775784 675482 775840
rect 675538 775784 675543 775840
rect 674833 775782 675543 775784
rect 674833 775779 674899 775782
rect 675477 775779 675543 775782
rect 675661 775708 675727 775709
rect 675661 775704 675708 775708
rect 675772 775706 675778 775708
rect 675661 775648 675666 775704
rect 675661 775644 675708 775648
rect 675772 775646 675818 775706
rect 675772 775644 675778 775646
rect 675661 775643 675727 775644
rect 675017 774890 675083 774893
rect 676806 774890 676812 774892
rect 675017 774888 676812 774890
rect 675017 774832 675022 774888
rect 675078 774832 676812 774888
rect 675017 774830 676812 774832
rect 675017 774827 675083 774830
rect 676806 774828 676812 774830
rect 676876 774828 676882 774892
rect 41462 774346 41522 774452
rect 54477 774346 54543 774349
rect 41462 774344 54543 774346
rect 41462 774288 54482 774344
rect 54538 774288 54543 774344
rect 41462 774286 54543 774288
rect 54477 774283 54543 774286
rect 41462 773938 41522 774044
rect 41462 773878 45570 773938
rect 35758 773533 35818 773636
rect 35758 773528 35867 773533
rect 35758 773472 35806 773528
rect 35862 773472 35867 773528
rect 35758 773470 35867 773472
rect 35801 773467 35867 773470
rect 44357 773258 44423 773261
rect 41492 773256 44423 773258
rect 41492 773200 44362 773256
rect 44418 773200 44423 773256
rect 41492 773198 44423 773200
rect 44357 773195 44423 773198
rect 44633 772850 44699 772853
rect 41492 772848 44699 772850
rect 41492 772792 44638 772848
rect 44694 772792 44699 772848
rect 41492 772790 44699 772792
rect 45510 772850 45570 773878
rect 668945 773802 669011 773805
rect 675477 773802 675543 773805
rect 668945 773800 675543 773802
rect 668945 773744 668950 773800
rect 669006 773744 675482 773800
rect 675538 773744 675543 773800
rect 668945 773742 675543 773744
rect 668945 773739 669011 773742
rect 675477 773739 675543 773742
rect 55857 772850 55923 772853
rect 45510 772848 55923 772850
rect 45510 772792 55862 772848
rect 55918 772792 55923 772848
rect 45510 772790 55923 772792
rect 44633 772787 44699 772790
rect 55857 772787 55923 772790
rect 676070 772652 676076 772716
rect 676140 772714 676146 772716
rect 682377 772714 682443 772717
rect 676140 772712 682443 772714
rect 676140 772656 682382 772712
rect 682438 772656 682443 772712
rect 676140 772654 682443 772656
rect 676140 772652 676146 772654
rect 682377 772651 682443 772654
rect 44817 772442 44883 772445
rect 41492 772440 44883 772442
rect 41492 772384 44822 772440
rect 44878 772384 44883 772440
rect 41492 772382 44883 772384
rect 44817 772379 44883 772382
rect 44173 772034 44239 772037
rect 41492 772032 44239 772034
rect 41492 771976 44178 772032
rect 44234 771976 44239 772032
rect 41492 771974 44239 771976
rect 44173 771971 44239 771974
rect 673913 772034 673979 772037
rect 683205 772034 683271 772037
rect 673913 772032 683271 772034
rect 673913 771976 673918 772032
rect 673974 771976 683210 772032
rect 683266 771976 683271 772032
rect 673913 771974 683271 771976
rect 673913 771971 673979 771974
rect 683205 771971 683271 771974
rect 44357 771626 44423 771629
rect 41492 771624 44423 771626
rect 41492 771568 44362 771624
rect 44418 771568 44423 771624
rect 41492 771566 44423 771568
rect 44357 771563 44423 771566
rect 44357 771218 44423 771221
rect 41492 771216 44423 771218
rect 41492 771160 44362 771216
rect 44418 771160 44423 771216
rect 41492 771158 44423 771160
rect 44357 771155 44423 771158
rect 673862 770884 673868 770948
rect 673932 770946 673938 770948
rect 683389 770946 683455 770949
rect 673932 770944 683455 770946
rect 673932 770888 683394 770944
rect 683450 770888 683455 770944
rect 673932 770886 683455 770888
rect 673932 770884 673938 770886
rect 683389 770883 683455 770886
rect 45001 770810 45067 770813
rect 41492 770808 45067 770810
rect 41492 770752 45006 770808
rect 45062 770752 45067 770808
rect 41492 770750 45067 770752
rect 45001 770747 45067 770750
rect 672165 770674 672231 770677
rect 683573 770674 683639 770677
rect 672165 770672 683639 770674
rect 672165 770616 672170 770672
rect 672226 770616 683578 770672
rect 683634 770616 683639 770672
rect 672165 770614 683639 770616
rect 672165 770611 672231 770614
rect 683573 770611 683639 770614
rect 45093 770402 45159 770405
rect 41492 770400 45159 770402
rect 41492 770344 45098 770400
rect 45154 770344 45159 770400
rect 41492 770342 45159 770344
rect 45093 770339 45159 770342
rect 41462 769860 41522 769964
rect 41454 769796 41460 769860
rect 41524 769796 41530 769860
rect 35574 769453 35634 769556
rect 35574 769448 35683 769453
rect 35574 769392 35622 769448
rect 35678 769392 35683 769448
rect 35574 769390 35683 769392
rect 35617 769387 35683 769390
rect 35390 769045 35450 769148
rect 35390 769040 35499 769045
rect 35801 769042 35867 769045
rect 35390 768984 35438 769040
rect 35494 768984 35499 769040
rect 35390 768982 35499 768984
rect 35433 768979 35499 768982
rect 35758 769040 35867 769042
rect 35758 768984 35806 769040
rect 35862 768984 35867 769040
rect 35758 768979 35867 768984
rect 35758 768740 35818 768979
rect 30974 768229 31034 768332
rect 30974 768224 31083 768229
rect 30974 768168 31022 768224
rect 31078 768168 31083 768224
rect 30974 768166 31083 768168
rect 31017 768163 31083 768166
rect 674833 768226 674899 768229
rect 676121 768226 676187 768229
rect 674833 768224 676187 768226
rect 674833 768168 674838 768224
rect 674894 768168 676126 768224
rect 676182 768168 676187 768224
rect 674833 768166 676187 768168
rect 674833 768163 674899 768166
rect 676121 768163 676187 768166
rect 35758 767821 35818 767924
rect 35758 767816 35867 767821
rect 35758 767760 35806 767816
rect 35862 767760 35867 767816
rect 35758 767758 35867 767760
rect 35801 767755 35867 767758
rect 35758 767413 35818 767516
rect 35758 767408 35867 767413
rect 35758 767352 35806 767408
rect 35862 767352 35867 767408
rect 35758 767350 35867 767352
rect 35801 767347 35867 767350
rect 62113 767410 62179 767413
rect 62113 767408 64492 767410
rect 62113 767352 62118 767408
rect 62174 767352 64492 767408
rect 62113 767350 64492 767352
rect 62113 767347 62179 767350
rect 35206 767005 35266 767108
rect 35157 767000 35266 767005
rect 35157 766944 35162 767000
rect 35218 766944 35266 767000
rect 35157 766942 35266 766944
rect 35157 766939 35223 766942
rect 44817 766730 44883 766733
rect 41492 766728 44883 766730
rect 41492 766672 44822 766728
rect 44878 766672 44883 766728
rect 41492 766670 44883 766672
rect 44817 766667 44883 766670
rect 675201 766594 675267 766597
rect 676121 766596 676187 766597
rect 675886 766594 675892 766596
rect 675201 766592 675892 766594
rect 675201 766536 675206 766592
rect 675262 766536 675892 766592
rect 675201 766534 675892 766536
rect 675201 766531 675267 766534
rect 675886 766532 675892 766534
rect 675956 766532 675962 766596
rect 676070 766532 676076 766596
rect 676140 766594 676187 766596
rect 676140 766592 676232 766594
rect 676182 766536 676232 766592
rect 676140 766534 676232 766536
rect 676140 766532 676187 766534
rect 676121 766531 676187 766532
rect 43161 766322 43227 766325
rect 41492 766320 43227 766322
rect 41492 766264 43166 766320
rect 43222 766264 43227 766320
rect 41492 766262 43227 766264
rect 43161 766259 43227 766262
rect 40910 765780 40970 765884
rect 40902 765716 40908 765780
rect 40972 765716 40978 765780
rect 41321 765778 41387 765781
rect 42241 765778 42307 765781
rect 41321 765776 42307 765778
rect 41321 765720 41326 765776
rect 41382 765720 42246 765776
rect 42302 765720 42307 765776
rect 41321 765718 42307 765720
rect 41321 765715 41387 765718
rect 42241 765715 42307 765718
rect 40542 765372 40602 765476
rect 40534 765308 40540 765372
rect 40604 765308 40610 765372
rect 40726 764964 40786 765068
rect 40718 764900 40724 764964
rect 40788 764900 40794 764964
rect 45277 764826 45343 764829
rect 41462 764824 45343 764826
rect 41462 764768 45282 764824
rect 45338 764768 45343 764824
rect 41462 764766 45343 764768
rect 41462 764660 41522 764766
rect 45277 764763 45343 764766
rect 40033 764554 40099 764557
rect 41638 764554 41644 764556
rect 40033 764552 41644 764554
rect 40033 764496 40038 764552
rect 40094 764496 41644 764552
rect 40033 764494 41644 764496
rect 40033 764491 40099 764494
rect 41638 764492 41644 764494
rect 41708 764492 41714 764556
rect 45553 764282 45619 764285
rect 41492 764280 45619 764282
rect 41492 764224 45558 764280
rect 45614 764224 45619 764280
rect 41492 764222 45619 764224
rect 45553 764219 45619 764222
rect 37046 763333 37106 763844
rect 37046 763328 37155 763333
rect 651465 763330 651531 763333
rect 37046 763272 37094 763328
rect 37150 763272 37155 763328
rect 37046 763270 37155 763272
rect 650164 763328 651531 763330
rect 650164 763272 651470 763328
rect 651526 763272 651531 763328
rect 650164 763270 651531 763272
rect 37089 763267 37155 763270
rect 651465 763267 651531 763270
rect 46381 763058 46447 763061
rect 41492 763056 46447 763058
rect 41492 763000 46386 763056
rect 46442 763000 46447 763056
rect 41492 762998 46447 763000
rect 46381 762995 46447 762998
rect 671337 763058 671403 763061
rect 676029 763058 676095 763061
rect 671337 763056 676095 763058
rect 671337 763000 671342 763056
rect 671398 763000 676034 763056
rect 676090 763000 676095 763056
rect 671337 762998 676095 763000
rect 671337 762995 671403 762998
rect 676029 762995 676095 762998
rect 677041 761972 677107 761973
rect 676990 761908 676996 761972
rect 677060 761970 677107 761972
rect 677060 761968 677152 761970
rect 677102 761912 677152 761968
rect 677060 761910 677152 761912
rect 677060 761908 677107 761910
rect 677041 761907 677107 761908
rect 676765 761836 676831 761837
rect 676765 761832 676812 761836
rect 676876 761834 676882 761836
rect 676765 761776 676770 761832
rect 676765 761772 676812 761776
rect 676876 761774 676922 761834
rect 676876 761772 676882 761774
rect 676765 761771 676831 761772
rect 663750 761502 676292 761562
rect 663057 760882 663123 760885
rect 663750 760882 663810 761502
rect 663057 760880 663810 760882
rect 663057 760824 663062 760880
rect 663118 760824 663810 760880
rect 663057 760822 663810 760824
rect 669270 761094 676292 761154
rect 663057 760819 663123 760822
rect 661677 760474 661743 760477
rect 669270 760474 669330 761094
rect 676029 760746 676095 760749
rect 676029 760744 676292 760746
rect 676029 760688 676034 760744
rect 676090 760688 676292 760744
rect 676029 760686 676292 760688
rect 676029 760683 676095 760686
rect 661677 760472 669330 760474
rect 661677 760416 661682 760472
rect 661738 760416 669330 760472
rect 661677 760414 669330 760416
rect 661677 760411 661743 760414
rect 672717 760338 672783 760341
rect 672717 760336 676292 760338
rect 672717 760280 672722 760336
rect 672778 760280 676292 760336
rect 672717 760278 676292 760280
rect 672717 760275 672783 760278
rect 672717 759930 672783 759933
rect 672717 759928 676292 759930
rect 672717 759872 672722 759928
rect 672778 759872 676292 759928
rect 672717 759870 676292 759872
rect 672717 759867 672783 759870
rect 683573 759522 683639 759525
rect 683573 759520 683652 759522
rect 683573 759464 683578 759520
rect 683634 759464 683652 759520
rect 683573 759462 683652 759464
rect 683573 759459 683639 759462
rect 39297 759114 39363 759117
rect 42333 759114 42399 759117
rect 39297 759112 42399 759114
rect 39297 759056 39302 759112
rect 39358 759056 42338 759112
rect 42394 759056 42399 759112
rect 39297 759054 42399 759056
rect 39297 759051 39363 759054
rect 42333 759051 42399 759054
rect 673177 759114 673243 759117
rect 673177 759112 676292 759114
rect 673177 759056 673182 759112
rect 673238 759056 676292 759112
rect 673177 759054 676292 759056
rect 673177 759051 673243 759054
rect 42057 758706 42123 758709
rect 42374 758706 42380 758708
rect 42057 758704 42380 758706
rect 42057 758648 42062 758704
rect 42118 758648 42380 758704
rect 42057 758646 42380 758648
rect 42057 758643 42123 758646
rect 42374 758644 42380 758646
rect 42444 758644 42450 758708
rect 671797 758706 671863 758709
rect 671797 758704 676292 758706
rect 671797 758648 671802 758704
rect 671858 758648 676292 758704
rect 671797 758646 676292 758648
rect 671797 758643 671863 758646
rect 40585 758298 40651 758301
rect 42517 758298 42583 758301
rect 40585 758296 42583 758298
rect 40585 758240 40590 758296
rect 40646 758240 42522 758296
rect 42578 758240 42583 758296
rect 40585 758238 42583 758240
rect 40585 758235 40651 758238
rect 42517 758235 42583 758238
rect 671521 758298 671587 758301
rect 671521 758296 676292 758298
rect 671521 758240 671526 758296
rect 671582 758240 676292 758296
rect 671521 758238 676292 758240
rect 671521 758235 671587 758238
rect 671705 757890 671771 757893
rect 671705 757888 676292 757890
rect 671705 757832 671710 757888
rect 671766 757832 676292 757888
rect 671705 757830 676292 757832
rect 671705 757827 671771 757830
rect 36537 757754 36603 757757
rect 41822 757754 41828 757756
rect 36537 757752 41828 757754
rect 36537 757696 36542 757752
rect 36598 757696 41828 757752
rect 36537 757694 41828 757696
rect 36537 757691 36603 757694
rect 41822 757692 41828 757694
rect 41892 757692 41898 757756
rect 671705 757482 671771 757485
rect 671705 757480 676292 757482
rect 671705 757424 671710 757480
rect 671766 757424 676292 757480
rect 671705 757422 676292 757424
rect 671705 757419 671771 757422
rect 40309 757348 40375 757349
rect 40309 757346 40356 757348
rect 40264 757344 40356 757346
rect 40264 757288 40314 757344
rect 40264 757286 40356 757288
rect 40309 757284 40356 757286
rect 40420 757284 40426 757348
rect 40861 757346 40927 757349
rect 40861 757344 40970 757346
rect 40861 757288 40866 757344
rect 40922 757288 40970 757344
rect 40309 757283 40375 757284
rect 40861 757283 40970 757288
rect 40910 756666 40970 757283
rect 674649 757210 674715 757213
rect 676029 757210 676095 757213
rect 674649 757208 676095 757210
rect 674649 757152 674654 757208
rect 674710 757152 676034 757208
rect 676090 757152 676095 757208
rect 674649 757150 676095 757152
rect 674649 757147 674715 757150
rect 676029 757147 676095 757150
rect 682377 757074 682443 757077
rect 682364 757072 682443 757074
rect 682364 757016 682382 757072
rect 682438 757016 682443 757072
rect 682364 757014 682443 757016
rect 682377 757011 682443 757014
rect 41781 756666 41847 756669
rect 683297 756666 683363 756669
rect 40910 756664 41847 756666
rect 40910 756608 41786 756664
rect 41842 756608 41847 756664
rect 40910 756606 41847 756608
rect 683284 756664 683363 756666
rect 683284 756608 683302 756664
rect 683358 756608 683363 756664
rect 683284 756606 683363 756608
rect 41781 756603 41847 756606
rect 683297 756603 683363 756606
rect 669270 756198 676292 756258
rect 669270 755173 669330 756198
rect 675845 755850 675911 755853
rect 675845 755848 676292 755850
rect 675845 755792 675850 755848
rect 675906 755792 676292 755848
rect 675845 755790 676292 755792
rect 675845 755787 675911 755790
rect 672993 755442 673059 755445
rect 672993 755440 676292 755442
rect 672993 755384 672998 755440
rect 673054 755384 676292 755440
rect 672993 755382 676292 755384
rect 672993 755379 673059 755382
rect 669221 755168 669330 755173
rect 669221 755112 669226 755168
rect 669282 755112 669330 755168
rect 669221 755110 669330 755112
rect 669221 755107 669287 755110
rect 676765 755034 676831 755037
rect 676765 755032 676844 755034
rect 676765 754976 676770 755032
rect 676826 754976 676844 755032
rect 676765 754974 676844 754976
rect 676765 754971 676831 754974
rect 42333 754900 42399 754901
rect 40902 754836 40908 754900
rect 40972 754898 40978 754900
rect 42006 754898 42012 754900
rect 40972 754838 42012 754898
rect 40972 754836 40978 754838
rect 42006 754836 42012 754838
rect 42076 754836 42082 754900
rect 42333 754896 42380 754900
rect 42444 754898 42450 754900
rect 42333 754840 42338 754896
rect 42333 754836 42380 754840
rect 42444 754838 42490 754898
rect 42444 754836 42450 754838
rect 42333 754835 42399 754836
rect 40350 754564 40356 754628
rect 40420 754626 40426 754628
rect 42793 754626 42859 754629
rect 677041 754626 677107 754629
rect 40420 754624 42859 754626
rect 40420 754568 42798 754624
rect 42854 754568 42859 754624
rect 40420 754566 42859 754568
rect 677028 754624 677107 754626
rect 677028 754568 677046 754624
rect 677102 754568 677107 754624
rect 677028 754566 677107 754568
rect 40420 754564 40426 754566
rect 42793 754563 42859 754566
rect 677041 754563 677107 754566
rect 62113 754354 62179 754357
rect 62113 754352 64492 754354
rect 62113 754296 62118 754352
rect 62174 754296 64492 754352
rect 62113 754294 64492 754296
rect 62113 754291 62179 754294
rect 672533 754218 672599 754221
rect 672533 754216 676292 754218
rect 672533 754160 672538 754216
rect 672594 754160 676292 754216
rect 672533 754158 676292 754160
rect 672533 754155 672599 754158
rect 42057 754082 42123 754085
rect 46197 754082 46263 754085
rect 42057 754080 46263 754082
rect 42057 754024 42062 754080
rect 42118 754024 46202 754080
rect 46258 754024 46263 754080
rect 42057 754022 46263 754024
rect 42057 754019 42123 754022
rect 46197 754019 46263 754022
rect 683481 753810 683547 753813
rect 683468 753808 683547 753810
rect 683468 753752 683486 753808
rect 683542 753752 683547 753808
rect 683468 753750 683547 753752
rect 683481 753747 683547 753750
rect 42333 753674 42399 753677
rect 45277 753674 45343 753677
rect 42333 753672 45343 753674
rect 42333 753616 42338 753672
rect 42394 753616 45282 753672
rect 45338 753616 45343 753672
rect 42333 753614 45343 753616
rect 42333 753611 42399 753614
rect 45277 753611 45343 753614
rect 669270 753342 676292 753402
rect 42057 752994 42123 752997
rect 43161 752994 43227 752997
rect 42057 752992 43227 752994
rect 42057 752936 42062 752992
rect 42118 752936 43166 752992
rect 43222 752936 43227 752992
rect 42057 752934 43227 752936
rect 42057 752931 42123 752934
rect 43161 752931 43227 752934
rect 668209 752314 668275 752317
rect 669270 752314 669330 753342
rect 683113 752994 683179 752997
rect 683100 752992 683179 752994
rect 683100 752936 683118 752992
rect 683174 752936 683179 752992
rect 683100 752934 683179 752936
rect 683113 752931 683179 752934
rect 671153 752586 671219 752589
rect 671153 752584 676292 752586
rect 671153 752528 671158 752584
rect 671214 752528 676292 752584
rect 671153 752526 676292 752528
rect 671153 752523 671219 752526
rect 668209 752312 669330 752314
rect 668209 752256 668214 752312
rect 668270 752256 669330 752312
rect 668209 752254 669330 752256
rect 668209 752251 668275 752254
rect 673913 752178 673979 752181
rect 673913 752176 676292 752178
rect 673913 752120 673918 752176
rect 673974 752120 676292 752176
rect 673913 752118 676292 752120
rect 673913 752115 673979 752118
rect 670601 751770 670667 751773
rect 670601 751768 676292 751770
rect 670601 751712 670606 751768
rect 670662 751712 676292 751768
rect 670601 751710 676292 751712
rect 670601 751707 670667 751710
rect 672901 751362 672967 751365
rect 672901 751360 676292 751362
rect 672901 751304 672906 751360
rect 672962 751304 676292 751360
rect 672901 751302 676292 751304
rect 672901 751299 672967 751302
rect 41965 751092 42031 751093
rect 41965 751088 42012 751092
rect 42076 751090 42082 751092
rect 41965 751032 41970 751088
rect 41965 751028 42012 751032
rect 42076 751030 42122 751090
rect 42076 751028 42082 751030
rect 41965 751027 42031 751028
rect 669773 750954 669839 750957
rect 669773 750952 676292 750954
rect 669773 750896 669778 750952
rect 669834 750924 676292 750952
rect 669834 750896 676322 750924
rect 669773 750894 676322 750896
rect 669773 750891 669839 750894
rect 676262 750516 676322 750894
rect 40718 750348 40724 750412
rect 40788 750410 40794 750412
rect 41781 750410 41847 750413
rect 40788 750408 41847 750410
rect 40788 750352 41786 750408
rect 41842 750352 41847 750408
rect 40788 750350 41847 750352
rect 40788 750348 40794 750350
rect 41781 750347 41847 750350
rect 651465 750138 651531 750141
rect 650164 750136 651531 750138
rect 650164 750080 651470 750136
rect 651526 750080 651531 750136
rect 650164 750078 651531 750080
rect 651465 750075 651531 750078
rect 670785 750138 670851 750141
rect 670785 750136 676292 750138
rect 670785 750080 670790 750136
rect 670846 750080 676292 750136
rect 670785 750078 676292 750080
rect 670785 750075 670851 750078
rect 40534 747356 40540 747420
rect 40604 747418 40610 747420
rect 41781 747418 41847 747421
rect 40604 747416 41847 747418
rect 40604 747360 41786 747416
rect 41842 747360 41847 747416
rect 40604 747358 41847 747360
rect 40604 747356 40610 747358
rect 41781 747355 41847 747358
rect 42149 746738 42215 746741
rect 44817 746738 44883 746741
rect 42149 746736 44883 746738
rect 42149 746680 42154 746736
rect 42210 746680 44822 746736
rect 44878 746680 44883 746736
rect 42149 746678 44883 746680
rect 42149 746675 42215 746678
rect 44817 746675 44883 746678
rect 42149 746058 42215 746061
rect 42701 746058 42767 746061
rect 42149 746056 42767 746058
rect 42149 746000 42154 746056
rect 42210 746000 42706 746056
rect 42762 746000 42767 746056
rect 42149 745998 42767 746000
rect 42149 745995 42215 745998
rect 42701 745995 42767 745998
rect 41822 745316 41828 745380
rect 41892 745378 41898 745380
rect 42241 745378 42307 745381
rect 41892 745376 42307 745378
rect 41892 745320 42246 745376
rect 42302 745320 42307 745376
rect 41892 745318 42307 745320
rect 41892 745316 41898 745318
rect 42241 745315 42307 745318
rect 41638 744364 41644 744428
rect 41708 744426 41714 744428
rect 42609 744426 42675 744429
rect 41708 744424 42675 744426
rect 41708 744368 42614 744424
rect 42670 744368 42675 744424
rect 41708 744366 42675 744368
rect 41708 744364 41714 744366
rect 42609 744363 42675 744366
rect 41454 743684 41460 743748
rect 41524 743746 41530 743748
rect 41781 743746 41847 743749
rect 41524 743744 41847 743746
rect 41524 743688 41786 743744
rect 41842 743688 41847 743744
rect 41524 743686 41847 743688
rect 41524 743684 41530 743686
rect 41781 743683 41847 743686
rect 667565 743202 667631 743205
rect 675109 743202 675175 743205
rect 667565 743200 675175 743202
rect 667565 743144 667570 743200
rect 667626 743144 675114 743200
rect 675170 743144 675175 743200
rect 667565 743142 675175 743144
rect 667565 743139 667631 743142
rect 675109 743139 675175 743142
rect 42609 743066 42675 743069
rect 62757 743066 62823 743069
rect 42609 743064 62823 743066
rect 42609 743008 42614 743064
rect 42670 743008 62762 743064
rect 62818 743008 62823 743064
rect 42609 743006 62823 743008
rect 42609 743003 42675 743006
rect 62757 743003 62823 743006
rect 666461 742794 666527 742797
rect 674925 742794 674991 742797
rect 666461 742792 674991 742794
rect 666461 742736 666466 742792
rect 666522 742736 674930 742792
rect 674986 742736 674991 742792
rect 666461 742734 674991 742736
rect 666461 742731 666527 742734
rect 674925 742731 674991 742734
rect 674414 742460 674420 742524
rect 674484 742522 674490 742524
rect 675385 742522 675451 742525
rect 674484 742520 675451 742522
rect 674484 742464 675390 742520
rect 675446 742464 675451 742520
rect 674484 742462 675451 742464
rect 674484 742460 674490 742462
rect 675385 742459 675451 742462
rect 42425 741706 42491 741709
rect 62941 741706 63007 741709
rect 42425 741704 63007 741706
rect 42425 741648 42430 741704
rect 42486 741648 62946 741704
rect 63002 741648 63007 741704
rect 42425 741646 63007 741648
rect 42425 741643 42491 741646
rect 62941 741643 63007 741646
rect 674230 741508 674236 741572
rect 674300 741570 674306 741572
rect 675109 741570 675175 741573
rect 674300 741568 675175 741570
rect 674300 741512 675114 741568
rect 675170 741512 675175 741568
rect 674300 741510 675175 741512
rect 674300 741508 674306 741510
rect 675109 741507 675175 741510
rect 62113 741298 62179 741301
rect 62113 741296 64492 741298
rect 62113 741240 62118 741296
rect 62174 741240 64492 741296
rect 62113 741238 64492 741240
rect 62113 741235 62179 741238
rect 669405 741162 669471 741165
rect 674925 741162 674991 741165
rect 669405 741160 674991 741162
rect 669405 741104 669410 741160
rect 669466 741104 674930 741160
rect 674986 741104 674991 741160
rect 669405 741102 674991 741104
rect 669405 741099 669471 741102
rect 674925 741099 674991 741102
rect 674598 739604 674604 739668
rect 674668 739666 674674 739668
rect 675109 739666 675175 739669
rect 674668 739664 675175 739666
rect 674668 739608 675114 739664
rect 675170 739608 675175 739664
rect 674668 739606 675175 739608
rect 674668 739604 674674 739606
rect 675109 739603 675175 739606
rect 669773 738578 669839 738581
rect 675017 738578 675083 738581
rect 669773 738576 675083 738578
rect 669773 738520 669778 738576
rect 669834 738520 675022 738576
rect 675078 738520 675083 738576
rect 669773 738518 675083 738520
rect 669773 738515 669839 738518
rect 675017 738515 675083 738518
rect 675201 738374 675267 738377
rect 675158 738372 675267 738374
rect 675158 738316 675206 738372
rect 675262 738316 675267 738372
rect 675158 738311 675267 738316
rect 672533 738306 672599 738309
rect 675158 738306 675218 738311
rect 672533 738304 675218 738306
rect 672533 738248 672538 738304
rect 672594 738248 675218 738304
rect 672533 738246 675218 738248
rect 672533 738243 672599 738246
rect 671153 737082 671219 737085
rect 675109 737082 675175 737085
rect 671153 737080 675175 737082
rect 671153 737024 671158 737080
rect 671214 737024 675114 737080
rect 675170 737024 675175 737080
rect 671153 737022 675175 737024
rect 671153 737019 671219 737022
rect 675109 737019 675175 737022
rect 652569 736810 652635 736813
rect 650164 736808 652635 736810
rect 650164 736752 652574 736808
rect 652630 736752 652635 736808
rect 650164 736750 652635 736752
rect 652569 736747 652635 736750
rect 668761 734362 668827 734365
rect 674925 734362 674991 734365
rect 668761 734360 674991 734362
rect 668761 734304 668766 734360
rect 668822 734304 674930 734360
rect 674986 734304 674991 734360
rect 668761 734302 674991 734304
rect 668761 734299 668827 734302
rect 674925 734299 674991 734302
rect 672165 733682 672231 733685
rect 675109 733682 675175 733685
rect 672165 733680 675175 733682
rect 672165 733624 672170 733680
rect 672226 733624 675114 733680
rect 675170 733624 675175 733680
rect 672165 733622 675175 733624
rect 672165 733619 672231 733622
rect 675109 733619 675175 733622
rect 668209 733410 668275 733413
rect 675109 733410 675175 733413
rect 668209 733408 675175 733410
rect 668209 733352 668214 733408
rect 668270 733352 675114 733408
rect 675170 733352 675175 733408
rect 668209 733350 675175 733352
rect 668209 733347 668275 733350
rect 675109 733347 675175 733350
rect 671981 732868 672047 732869
rect 673361 732868 673427 732869
rect 671981 732864 672028 732868
rect 672092 732866 672098 732868
rect 673310 732866 673316 732868
rect 671981 732808 671986 732864
rect 671981 732804 672028 732808
rect 672092 732806 672138 732866
rect 673270 732806 673316 732866
rect 673380 732864 673427 732868
rect 673422 732808 673427 732864
rect 672092 732804 672098 732806
rect 673310 732804 673316 732806
rect 673380 732804 673427 732808
rect 671981 732803 672047 732804
rect 673361 732803 673427 732804
rect 668761 731506 668827 731509
rect 675109 731506 675175 731509
rect 668761 731504 675175 731506
rect 668761 731448 668766 731504
rect 668822 731448 675114 731504
rect 675170 731448 675175 731504
rect 668761 731446 675175 731448
rect 668761 731443 668827 731446
rect 675109 731443 675175 731446
rect 35617 731370 35683 731373
rect 35604 731368 35683 731370
rect 35604 731312 35622 731368
rect 35678 731312 35683 731368
rect 35604 731310 35683 731312
rect 35617 731307 35683 731310
rect 35801 730962 35867 730965
rect 35788 730960 35867 730962
rect 35788 730904 35806 730960
rect 35862 730904 35867 730960
rect 35788 730902 35867 730904
rect 35801 730899 35867 730902
rect 50337 730554 50403 730557
rect 41492 730552 50403 730554
rect 41492 730496 50342 730552
rect 50398 730496 50403 730552
rect 41492 730494 50403 730496
rect 50337 730491 50403 730494
rect 671061 730554 671127 730557
rect 675477 730554 675543 730557
rect 671061 730552 675543 730554
rect 671061 730496 671066 730552
rect 671122 730496 675482 730552
rect 675538 730496 675543 730552
rect 671061 730494 675543 730496
rect 671061 730491 671127 730494
rect 675477 730491 675543 730494
rect 44633 730146 44699 730149
rect 41492 730144 44699 730146
rect 41492 730088 44638 730144
rect 44694 730088 44699 730144
rect 41492 730086 44699 730088
rect 44633 730083 44699 730086
rect 673361 730146 673427 730149
rect 675293 730146 675359 730149
rect 673361 730144 675359 730146
rect 673361 730088 673366 730144
rect 673422 730088 675298 730144
rect 675354 730088 675359 730144
rect 673361 730086 675359 730088
rect 673361 730083 673427 730086
rect 675293 730083 675359 730086
rect 675886 729948 675892 730012
rect 675956 730010 675962 730012
rect 676806 730010 676812 730012
rect 675956 729950 676812 730010
rect 675956 729948 675962 729950
rect 676806 729948 676812 729950
rect 676876 729948 676882 730012
rect 44541 729738 44607 729741
rect 41492 729736 44607 729738
rect 41492 729680 44546 729736
rect 44602 729680 44607 729736
rect 41492 729678 44607 729680
rect 44541 729675 44607 729678
rect 44173 729330 44239 729333
rect 41492 729328 44239 729330
rect 41492 729272 44178 729328
rect 44234 729272 44239 729328
rect 41492 729270 44239 729272
rect 44173 729267 44239 729270
rect 44909 728922 44975 728925
rect 41492 728920 44975 728922
rect 41492 728864 44914 728920
rect 44970 728864 44975 728920
rect 41492 728862 44975 728864
rect 44909 728859 44975 728862
rect 44357 728514 44423 728517
rect 673361 728516 673427 728517
rect 41492 728512 44423 728514
rect 41492 728456 44362 728512
rect 44418 728456 44423 728512
rect 41492 728454 44423 728456
rect 44357 728451 44423 728454
rect 673310 728452 673316 728516
rect 673380 728514 673427 728516
rect 673380 728512 673472 728514
rect 673422 728456 673472 728512
rect 673380 728454 673472 728456
rect 673380 728452 673427 728454
rect 673361 728451 673427 728452
rect 62757 728242 62823 728245
rect 62757 728240 64492 728242
rect 62757 728184 62762 728240
rect 62818 728184 64492 728240
rect 62757 728182 64492 728184
rect 62757 728179 62823 728182
rect 672022 728180 672028 728244
rect 672092 728242 672098 728244
rect 673821 728242 673887 728245
rect 672092 728240 673887 728242
rect 672092 728184 673826 728240
rect 673882 728184 673887 728240
rect 672092 728182 673887 728184
rect 672092 728180 672098 728182
rect 673821 728179 673887 728182
rect 45277 728106 45343 728109
rect 41492 728104 45343 728106
rect 41492 728048 45282 728104
rect 45338 728048 45343 728104
rect 41492 728046 45343 728048
rect 45277 728043 45343 728046
rect 670785 727970 670851 727973
rect 674143 727970 674209 727973
rect 670785 727968 674209 727970
rect 670785 727912 670790 727968
rect 670846 727912 674148 727968
rect 674204 727912 674209 727968
rect 670785 727910 674209 727912
rect 670785 727907 670851 727910
rect 674143 727907 674209 727910
rect 45093 727698 45159 727701
rect 41492 727696 45159 727698
rect 41492 727640 45098 727696
rect 45154 727640 45159 727696
rect 41492 727638 45159 727640
rect 45093 727635 45159 727638
rect 673821 727698 673887 727701
rect 674741 727698 674807 727701
rect 673821 727696 674807 727698
rect 673821 727640 673826 727696
rect 673882 727640 674746 727696
rect 674802 727640 674807 727696
rect 673821 727638 674807 727640
rect 673821 727635 673887 727638
rect 674741 727635 674807 727638
rect 44265 727290 44331 727293
rect 41492 727288 44331 727290
rect 41492 727232 44270 727288
rect 44326 727232 44331 727288
rect 41492 727230 44331 727232
rect 44265 727227 44331 727230
rect 41822 726882 41828 726884
rect 41492 726822 41828 726882
rect 41822 726820 41828 726822
rect 41892 726820 41898 726884
rect 674281 726882 674347 726885
rect 683481 726882 683547 726885
rect 674281 726880 683547 726882
rect 674281 726824 674286 726880
rect 674342 726824 683486 726880
rect 683542 726824 683547 726880
rect 674281 726822 683547 726824
rect 674281 726819 674347 726822
rect 683481 726819 683547 726822
rect 674005 726610 674071 726613
rect 674557 726610 674623 726613
rect 674005 726608 674114 726610
rect 674005 726552 674010 726608
rect 674066 726552 674114 726608
rect 674005 726547 674114 726552
rect 674557 726608 678990 726610
rect 674557 726552 674562 726608
rect 674618 726552 678990 726608
rect 674557 726550 678990 726552
rect 674557 726547 674623 726550
rect 41321 726474 41387 726477
rect 41308 726472 41387 726474
rect 41308 726416 41326 726472
rect 41382 726416 41387 726472
rect 41308 726414 41387 726416
rect 41321 726411 41387 726414
rect 41137 726066 41203 726069
rect 41124 726064 41203 726066
rect 41124 726008 41142 726064
rect 41198 726008 41203 726064
rect 41124 726006 41203 726008
rect 41137 726003 41203 726006
rect 41321 725658 41387 725661
rect 41308 725656 41387 725658
rect 41308 725600 41326 725656
rect 41382 725600 41387 725656
rect 41308 725598 41387 725600
rect 41321 725595 41387 725598
rect 674054 725522 674114 726547
rect 678930 726474 678990 726550
rect 683665 726474 683731 726477
rect 678930 726472 683731 726474
rect 678930 726416 683670 726472
rect 683726 726416 683731 726472
rect 678930 726414 683731 726416
rect 683665 726411 683731 726414
rect 676070 725732 676076 725796
rect 676140 725794 676146 725796
rect 682377 725794 682443 725797
rect 676140 725792 682443 725794
rect 676140 725736 682382 725792
rect 682438 725736 682443 725792
rect 676140 725734 682443 725736
rect 676140 725732 676146 725734
rect 682377 725731 682443 725734
rect 683113 725522 683179 725525
rect 674054 725520 683179 725522
rect 674054 725464 683118 725520
rect 683174 725464 683179 725520
rect 674054 725462 683179 725464
rect 683113 725459 683179 725462
rect 31017 725250 31083 725253
rect 31004 725248 31083 725250
rect 31004 725192 31022 725248
rect 31078 725192 31083 725248
rect 31004 725190 31083 725192
rect 31017 725187 31083 725190
rect 36537 724842 36603 724845
rect 36524 724840 36603 724842
rect 36524 724784 36542 724840
rect 36598 724784 36603 724840
rect 36524 724782 36603 724784
rect 36537 724779 36603 724782
rect 40677 724434 40743 724437
rect 40677 724432 40756 724434
rect 40677 724376 40682 724432
rect 40738 724376 40756 724432
rect 40677 724374 40756 724376
rect 40677 724371 40743 724374
rect 677317 724298 677383 724301
rect 676170 724296 677383 724298
rect 676170 724240 677322 724296
rect 677378 724240 677383 724296
rect 676170 724238 677383 724240
rect 673545 724162 673611 724165
rect 676170 724162 676230 724238
rect 677317 724235 677383 724238
rect 673545 724160 676230 724162
rect 673545 724104 673550 724160
rect 673606 724104 676230 724160
rect 673545 724102 676230 724104
rect 673545 724099 673611 724102
rect 33041 724026 33107 724029
rect 33028 724024 33107 724026
rect 33028 723968 33046 724024
rect 33102 723968 33107 724024
rect 33028 723966 33107 723968
rect 33041 723963 33107 723966
rect 43161 723618 43227 723621
rect 41492 723616 43227 723618
rect 41492 723560 43166 723616
rect 43222 723560 43227 723616
rect 41492 723558 43227 723560
rect 43161 723555 43227 723558
rect 651465 723482 651531 723485
rect 650164 723480 651531 723482
rect 650164 723424 651470 723480
rect 651526 723424 651531 723480
rect 650164 723422 651531 723424
rect 651465 723419 651531 723422
rect 33777 723210 33843 723213
rect 33764 723208 33843 723210
rect 33764 723152 33782 723208
rect 33838 723152 33843 723208
rect 33764 723150 33843 723152
rect 33777 723147 33843 723150
rect 45093 722802 45159 722805
rect 41492 722800 45159 722802
rect 41492 722744 45098 722800
rect 45154 722744 45159 722800
rect 41492 722742 45159 722744
rect 45093 722739 45159 722742
rect 41873 722394 41939 722397
rect 41492 722392 41939 722394
rect 41492 722336 41878 722392
rect 41934 722336 41939 722392
rect 41492 722334 41939 722336
rect 41873 722331 41939 722334
rect 40726 721772 40786 721956
rect 40718 721708 40724 721772
rect 40788 721708 40794 721772
rect 41137 721770 41203 721773
rect 41638 721770 41644 721772
rect 41137 721768 41644 721770
rect 41137 721712 41142 721768
rect 41198 721712 41644 721768
rect 41137 721710 41644 721712
rect 41137 721707 41203 721710
rect 41638 721708 41644 721710
rect 41708 721708 41714 721772
rect 43897 721578 43963 721581
rect 41492 721576 43963 721578
rect 41492 721520 43902 721576
rect 43958 721520 43963 721576
rect 41492 721518 43963 721520
rect 43897 721515 43963 721518
rect 44725 721170 44791 721173
rect 41492 721168 44791 721170
rect 41492 721112 44730 721168
rect 44786 721112 44791 721168
rect 41492 721110 44791 721112
rect 44725 721107 44791 721110
rect 40033 720354 40099 720357
rect 40020 720352 40099 720354
rect 40020 720296 40038 720352
rect 40094 720296 40099 720352
rect 40020 720294 40099 720296
rect 40033 720291 40099 720294
rect 46933 719946 46999 719949
rect 41492 719944 46999 719946
rect 41492 719888 46938 719944
rect 46994 719888 46999 719944
rect 41492 719886 46999 719888
rect 46933 719883 46999 719886
rect 41689 719266 41755 719269
rect 42517 719266 42583 719269
rect 41689 719264 42583 719266
rect 41689 719208 41694 719264
rect 41750 719208 42522 719264
rect 42578 719208 42583 719264
rect 41689 719206 42583 719208
rect 41689 719203 41755 719206
rect 42517 719203 42583 719206
rect 40534 718524 40540 718588
rect 40604 718586 40610 718588
rect 41873 718586 41939 718589
rect 40604 718584 41939 718586
rect 40604 718528 41878 718584
rect 41934 718528 41939 718584
rect 40604 718526 41939 718528
rect 40604 718524 40610 718526
rect 41873 718523 41939 718526
rect 42149 718314 42215 718317
rect 42558 718314 42564 718316
rect 42149 718312 42564 718314
rect 42149 718256 42154 718312
rect 42210 718256 42564 718312
rect 42149 718254 42564 718256
rect 42149 718251 42215 718254
rect 42558 718252 42564 718254
rect 42628 718252 42634 718316
rect 652017 718314 652083 718317
rect 676029 718314 676095 718317
rect 652017 718312 676095 718314
rect 652017 718256 652022 718312
rect 652078 718256 676034 718312
rect 676090 718256 676095 718312
rect 652017 718254 676095 718256
rect 652017 718251 652083 718254
rect 676029 718251 676095 718254
rect 664437 716546 664503 716549
rect 664437 716544 676292 716546
rect 664437 716488 664442 716544
rect 664498 716488 676292 716544
rect 664437 716486 676292 716488
rect 664437 716483 664503 716486
rect 663750 716078 676292 716138
rect 658917 716002 658983 716005
rect 663750 716002 663810 716078
rect 658917 716000 663810 716002
rect 658917 715944 658922 716000
rect 658978 715944 663810 716000
rect 658917 715942 663810 715944
rect 658917 715939 658983 715942
rect 676029 715730 676095 715733
rect 676029 715728 676292 715730
rect 676029 715672 676034 715728
rect 676090 715672 676292 715728
rect 676029 715670 676292 715672
rect 676029 715667 676095 715670
rect 40217 715594 40283 715597
rect 42701 715594 42767 715597
rect 40217 715592 42767 715594
rect 40217 715536 40222 715592
rect 40278 715536 42706 715592
rect 42762 715536 42767 715592
rect 40217 715534 42767 715536
rect 40217 715531 40283 715534
rect 42701 715531 42767 715534
rect 62113 715322 62179 715325
rect 672809 715322 672875 715325
rect 62113 715320 64492 715322
rect 62113 715264 62118 715320
rect 62174 715264 64492 715320
rect 62113 715262 64492 715264
rect 672809 715320 676292 715322
rect 672809 715264 672814 715320
rect 672870 715264 676292 715320
rect 672809 715262 676292 715264
rect 62113 715259 62179 715262
rect 672809 715259 672875 715262
rect 39849 715186 39915 715189
rect 42333 715186 42399 715189
rect 39849 715184 42399 715186
rect 39849 715128 39854 715184
rect 39910 715128 42338 715184
rect 42394 715128 42399 715184
rect 39849 715126 42399 715128
rect 39849 715123 39915 715126
rect 42333 715123 42399 715126
rect 672809 714914 672875 714917
rect 672809 714912 676292 714914
rect 672809 714856 672814 714912
rect 672870 714856 676292 714912
rect 672809 714854 676292 714856
rect 672809 714851 672875 714854
rect 40677 714778 40743 714781
rect 42057 714780 42123 714781
rect 41822 714778 41828 714780
rect 40677 714776 41828 714778
rect 40677 714720 40682 714776
rect 40738 714720 41828 714776
rect 40677 714718 41828 714720
rect 40677 714715 40743 714718
rect 41822 714716 41828 714718
rect 41892 714716 41898 714780
rect 42006 714716 42012 714780
rect 42076 714778 42123 714780
rect 42076 714776 42168 714778
rect 42118 714720 42168 714776
rect 42076 714718 42168 714720
rect 42076 714716 42123 714718
rect 42057 714715 42123 714716
rect 40033 714506 40099 714509
rect 42057 714506 42123 714509
rect 40033 714504 42123 714506
rect 40033 714448 40038 714504
rect 40094 714448 42062 714504
rect 42118 714448 42123 714504
rect 40033 714446 42123 714448
rect 40033 714443 40099 714446
rect 42057 714443 42123 714446
rect 673177 714506 673243 714509
rect 673177 714504 676292 714506
rect 673177 714448 673182 714504
rect 673238 714448 676292 714504
rect 673177 714446 676292 714448
rect 673177 714443 673243 714446
rect 41505 714234 41571 714237
rect 42374 714234 42380 714236
rect 41505 714232 42380 714234
rect 41505 714176 41510 714232
rect 41566 714176 42380 714232
rect 41505 714174 42380 714176
rect 41505 714171 41571 714174
rect 42374 714172 42380 714174
rect 42444 714172 42450 714236
rect 672993 714098 673059 714101
rect 672993 714096 676292 714098
rect 672993 714040 672998 714096
rect 673054 714040 676292 714096
rect 672993 714038 676292 714040
rect 672993 714035 673059 714038
rect 671521 713690 671587 713693
rect 671521 713688 676292 713690
rect 671521 713632 671526 713688
rect 671582 713632 676292 713688
rect 671521 713630 676292 713632
rect 671521 713627 671587 713630
rect 41965 713420 42031 713421
rect 41965 713416 42012 713420
rect 42076 713418 42082 713420
rect 41965 713360 41970 713416
rect 41965 713356 42012 713360
rect 42076 713358 42122 713418
rect 42076 713356 42082 713358
rect 41965 713355 42031 713356
rect 671521 713282 671587 713285
rect 671521 713280 676292 713282
rect 671521 713224 671526 713280
rect 671582 713224 676292 713280
rect 671521 713222 676292 713224
rect 671521 713219 671587 713222
rect 671705 712874 671771 712877
rect 671705 712872 676292 712874
rect 671705 712816 671710 712872
rect 671766 712816 676292 712872
rect 671705 712814 676292 712816
rect 671705 712811 671771 712814
rect 670785 712466 670851 712469
rect 670785 712464 676292 712466
rect 670785 712408 670790 712464
rect 670846 712408 676292 712464
rect 670785 712406 676292 712408
rect 670785 712403 670851 712406
rect 675886 711996 675892 712060
rect 675956 712058 675962 712060
rect 675956 711998 676292 712058
rect 675956 711996 675962 711998
rect 42149 711650 42215 711653
rect 42558 711650 42564 711652
rect 42149 711648 42564 711650
rect 42149 711592 42154 711648
rect 42210 711592 42564 711648
rect 42149 711590 42564 711592
rect 42149 711587 42215 711590
rect 42558 711588 42564 711590
rect 42628 711588 42634 711652
rect 682377 711650 682443 711653
rect 682364 711648 682443 711650
rect 682364 711592 682382 711648
rect 682438 711592 682443 711648
rect 682364 711590 682443 711592
rect 682377 711587 682443 711590
rect 683665 711242 683731 711245
rect 683652 711240 683731 711242
rect 683652 711184 683670 711240
rect 683726 711184 683731 711240
rect 683652 711182 683731 711184
rect 683665 711179 683731 711182
rect 42149 710834 42215 710837
rect 47577 710834 47643 710837
rect 42149 710832 47643 710834
rect 42149 710776 42154 710832
rect 42210 710776 47582 710832
rect 47638 710776 47643 710832
rect 42149 710774 47643 710776
rect 42149 710771 42215 710774
rect 47577 710771 47643 710774
rect 667749 710834 667815 710837
rect 667749 710832 676292 710834
rect 667749 710776 667754 710832
rect 667810 710776 676292 710832
rect 667749 710774 676292 710776
rect 667749 710771 667815 710774
rect 670141 710426 670207 710429
rect 670141 710424 676292 710426
rect 670141 710368 670146 710424
rect 670202 710368 676292 710424
rect 670141 710366 676292 710368
rect 670141 710363 670207 710366
rect 652569 710290 652635 710293
rect 650164 710288 652635 710290
rect 650164 710232 652574 710288
rect 652630 710232 652635 710288
rect 650164 710230 652635 710232
rect 652569 710227 652635 710230
rect 668945 710018 669011 710021
rect 668945 710016 676292 710018
rect 668945 709960 668950 710016
rect 669006 709960 676292 710016
rect 668945 709958 676292 709960
rect 668945 709955 669011 709958
rect 669589 709610 669655 709613
rect 669589 709608 676292 709610
rect 669589 709552 669594 709608
rect 669650 709552 676292 709608
rect 669589 709550 676292 709552
rect 669589 709547 669655 709550
rect 40534 709140 40540 709204
rect 40604 709202 40610 709204
rect 42241 709202 42307 709205
rect 40604 709200 42307 709202
rect 40604 709144 42246 709200
rect 42302 709144 42307 709200
rect 40604 709142 42307 709144
rect 40604 709140 40610 709142
rect 42241 709139 42307 709142
rect 672349 709202 672415 709205
rect 672349 709200 676292 709202
rect 672349 709144 672354 709200
rect 672410 709144 676292 709200
rect 672349 709142 676292 709144
rect 672349 709139 672415 709142
rect 668393 708794 668459 708797
rect 668393 708792 676292 708794
rect 668393 708736 668398 708792
rect 668454 708736 676292 708792
rect 668393 708734 676292 708736
rect 668393 708731 668459 708734
rect 42149 708522 42215 708525
rect 43897 708522 43963 708525
rect 42149 708520 43963 708522
rect 42149 708464 42154 708520
rect 42210 708464 43902 708520
rect 43958 708464 43963 708520
rect 42149 708462 43963 708464
rect 42149 708459 42215 708462
rect 43897 708459 43963 708462
rect 683113 708386 683179 708389
rect 683100 708384 683179 708386
rect 683100 708328 683118 708384
rect 683174 708328 683179 708384
rect 683100 708326 683179 708328
rect 683113 708323 683179 708326
rect 683297 707978 683363 707981
rect 683284 707976 683363 707978
rect 683284 707920 683302 707976
rect 683358 707920 683363 707976
rect 683284 707918 683363 707920
rect 683297 707915 683363 707918
rect 42057 707706 42123 707709
rect 45093 707706 45159 707709
rect 42057 707704 45159 707706
rect 42057 707648 42062 707704
rect 42118 707648 45098 707704
rect 45154 707648 45159 707704
rect 42057 707646 45159 707648
rect 42057 707643 42123 707646
rect 45093 707643 45159 707646
rect 670325 707570 670391 707573
rect 670325 707568 676292 707570
rect 670325 707512 670330 707568
rect 670386 707512 676292 707568
rect 670325 707510 676292 707512
rect 670325 707507 670391 707510
rect 40718 707372 40724 707436
rect 40788 707434 40794 707436
rect 41781 707434 41847 707437
rect 40788 707432 41847 707434
rect 40788 707376 41786 707432
rect 41842 707376 41847 707432
rect 40788 707374 41847 707376
rect 40788 707372 40794 707374
rect 41781 707371 41847 707374
rect 683481 707162 683547 707165
rect 683468 707160 683547 707162
rect 683468 707104 683486 707160
rect 683542 707104 683547 707160
rect 683468 707102 683547 707104
rect 683481 707099 683547 707102
rect 670969 706754 671035 706757
rect 670969 706752 676292 706754
rect 670969 706696 670974 706752
rect 671030 706696 676292 706752
rect 670969 706694 676292 706696
rect 670969 706691 671035 706694
rect 42057 706618 42123 706621
rect 42374 706618 42380 706620
rect 42057 706616 42380 706618
rect 42057 706560 42062 706616
rect 42118 706560 42380 706616
rect 42057 706558 42380 706560
rect 42057 706555 42123 706558
rect 42374 706556 42380 706558
rect 42444 706556 42450 706620
rect 674373 706346 674439 706349
rect 674373 706344 676292 706346
rect 674373 706288 674378 706344
rect 674434 706288 676292 706344
rect 674373 706286 676292 706288
rect 674373 706283 674439 706286
rect 666277 705530 666343 705533
rect 676262 705530 676322 705908
rect 666277 705528 676322 705530
rect 666277 705472 666282 705528
rect 666338 705500 676322 705528
rect 666338 705472 676292 705500
rect 666277 705470 676292 705472
rect 666277 705467 666343 705470
rect 42241 705258 42307 705261
rect 43161 705258 43227 705261
rect 42241 705256 43227 705258
rect 42241 705200 42246 705256
rect 42302 705200 43166 705256
rect 43222 705200 43227 705256
rect 42241 705198 43227 705200
rect 42241 705195 42307 705198
rect 43161 705195 43227 705198
rect 669221 705122 669287 705125
rect 669221 705120 676292 705122
rect 669221 705064 669226 705120
rect 669282 705064 676292 705120
rect 669221 705062 676292 705064
rect 669221 705059 669287 705062
rect 42241 704032 42307 704037
rect 42241 703976 42246 704032
rect 42302 703976 42307 704032
rect 42241 703971 42307 703976
rect 42244 703629 42304 703971
rect 42241 703624 42307 703629
rect 42241 703568 42246 703624
rect 42302 703568 42307 703624
rect 42241 703563 42307 703568
rect 42057 703082 42123 703085
rect 42793 703082 42859 703085
rect 42057 703080 42859 703082
rect 42057 703024 42062 703080
rect 42118 703024 42798 703080
rect 42854 703024 42859 703080
rect 42057 703022 42859 703024
rect 42057 703019 42123 703022
rect 42793 703019 42859 703022
rect 62113 702266 62179 702269
rect 62113 702264 64492 702266
rect 62113 702208 62118 702264
rect 62174 702208 64492 702264
rect 62113 702206 64492 702208
rect 62113 702203 62179 702206
rect 41638 702068 41644 702132
rect 41708 702130 41714 702132
rect 42609 702130 42675 702133
rect 41708 702128 42675 702130
rect 41708 702072 42614 702128
rect 42670 702072 42675 702128
rect 41708 702070 42675 702072
rect 41708 702068 41714 702070
rect 42609 702067 42675 702070
rect 41454 701796 41460 701860
rect 41524 701858 41530 701860
rect 42241 701858 42307 701861
rect 41524 701856 42307 701858
rect 41524 701800 42246 701856
rect 42302 701800 42307 701856
rect 41524 701798 42307 701800
rect 41524 701796 41530 701798
rect 42241 701795 42307 701798
rect 41822 701524 41828 701588
rect 41892 701586 41898 701588
rect 42425 701586 42491 701589
rect 41892 701584 42491 701586
rect 41892 701528 42430 701584
rect 42486 701528 42491 701584
rect 41892 701526 42491 701528
rect 41892 701524 41898 701526
rect 42425 701523 42491 701526
rect 670601 699818 670667 699821
rect 674925 699818 674991 699821
rect 670601 699816 674991 699818
rect 670601 699760 670606 699816
rect 670662 699760 674930 699816
rect 674986 699760 674991 699816
rect 670601 699758 674991 699760
rect 670601 699755 670667 699758
rect 674925 699755 674991 699758
rect 673177 698322 673243 698325
rect 675109 698322 675175 698325
rect 673177 698320 675175 698322
rect 673177 698264 673182 698320
rect 673238 698264 675114 698320
rect 675170 698264 675175 698320
rect 673177 698262 675175 698264
rect 673177 698259 673243 698262
rect 675109 698259 675175 698262
rect 41689 697914 41755 697917
rect 62757 697914 62823 697917
rect 41689 697912 62823 697914
rect 41689 697856 41694 697912
rect 41750 697856 62762 697912
rect 62818 697856 62823 697912
rect 41689 697854 62823 697856
rect 41689 697851 41755 697854
rect 62757 697851 62823 697854
rect 652385 696962 652451 696965
rect 650164 696960 652451 696962
rect 650164 696904 652390 696960
rect 652446 696904 652451 696960
rect 650164 696902 652451 696904
rect 652385 696899 652451 696902
rect 675385 696828 675451 696829
rect 675334 696826 675340 696828
rect 675294 696766 675340 696826
rect 675404 696824 675451 696828
rect 675446 696768 675451 696824
rect 675334 696764 675340 696766
rect 675404 696764 675451 696768
rect 675385 696763 675451 696764
rect 669589 695194 669655 695197
rect 675109 695194 675175 695197
rect 669589 695192 675175 695194
rect 669589 695136 669594 695192
rect 669650 695136 675114 695192
rect 675170 695136 675175 695192
rect 669589 695134 675175 695136
rect 669589 695131 669655 695134
rect 675109 695131 675175 695134
rect 675661 694378 675727 694381
rect 675661 694376 675954 694378
rect 675661 694320 675666 694376
rect 675722 694320 675954 694376
rect 675661 694318 675954 694320
rect 675661 694315 675727 694318
rect 675894 694106 675954 694318
rect 676990 694106 676996 694108
rect 675894 694046 676996 694106
rect 676990 694044 676996 694046
rect 677060 694044 677066 694108
rect 668393 693290 668459 693293
rect 674925 693290 674991 693293
rect 668393 693288 674991 693290
rect 668393 693232 668398 693288
rect 668454 693232 674930 693288
rect 674986 693232 674991 693288
rect 668393 693230 674991 693232
rect 668393 693227 668459 693230
rect 674925 693227 674991 693230
rect 674005 693018 674071 693021
rect 675109 693018 675175 693021
rect 674005 693016 675175 693018
rect 674005 692960 674010 693016
rect 674066 692960 675114 693016
rect 675170 692960 675175 693016
rect 674005 692958 675175 692960
rect 674005 692955 674071 692958
rect 675109 692955 675175 692958
rect 35617 691386 35683 691389
rect 51717 691386 51783 691389
rect 35617 691384 51783 691386
rect 35617 691328 35622 691384
rect 35678 691328 51722 691384
rect 51778 691328 51783 691384
rect 35617 691326 51783 691328
rect 35617 691323 35683 691326
rect 51717 691323 51783 691326
rect 674189 690162 674255 690165
rect 675385 690162 675451 690165
rect 674189 690160 675451 690162
rect 674189 690104 674194 690160
rect 674250 690104 675390 690160
rect 675446 690104 675451 690160
rect 674189 690102 675451 690104
rect 674189 690099 674255 690102
rect 675385 690099 675451 690102
rect 673545 689618 673611 689621
rect 675293 689618 675359 689621
rect 673545 689616 675359 689618
rect 673545 689560 673550 689616
rect 673606 689560 675298 689616
rect 675354 689560 675359 689616
rect 673545 689558 675359 689560
rect 673545 689555 673611 689558
rect 675293 689555 675359 689558
rect 663057 689346 663123 689349
rect 663057 689344 675172 689346
rect 663057 689288 663062 689344
rect 663118 689288 675172 689344
rect 663057 689286 675172 689288
rect 663057 689283 663123 689286
rect 62113 689210 62179 689213
rect 62113 689208 64492 689210
rect 62113 689152 62118 689208
rect 62174 689152 64492 689208
rect 62113 689150 64492 689152
rect 62113 689147 62179 689150
rect 667749 688938 667815 688941
rect 674925 688938 674991 688941
rect 667749 688936 674991 688938
rect 667749 688880 667754 688936
rect 667810 688880 674930 688936
rect 674986 688880 674991 688936
rect 667749 688878 674991 688880
rect 675112 688938 675172 689286
rect 675293 688938 675359 688941
rect 675112 688936 675359 688938
rect 675112 688880 675298 688936
rect 675354 688880 675359 688936
rect 675112 688878 675359 688880
rect 667749 688875 667815 688878
rect 674925 688875 674991 688878
rect 675293 688875 675359 688878
rect 671981 688666 672047 688669
rect 675109 688666 675175 688669
rect 671981 688664 675175 688666
rect 671981 688608 671986 688664
rect 672042 688608 675114 688664
rect 675170 688608 675175 688664
rect 671981 688606 675175 688608
rect 671981 688603 672047 688606
rect 675109 688603 675175 688606
rect 54477 688122 54543 688125
rect 41492 688120 54543 688122
rect 41492 688064 54482 688120
rect 54538 688064 54543 688120
rect 41492 688062 54543 688064
rect 54477 688059 54543 688062
rect 35801 687714 35867 687717
rect 35788 687712 35867 687714
rect 35788 687656 35806 687712
rect 35862 687656 35867 687712
rect 35788 687654 35867 687656
rect 35801 687651 35867 687654
rect 670325 687442 670391 687445
rect 675477 687442 675543 687445
rect 670325 687440 675543 687442
rect 670325 687384 670330 687440
rect 670386 687384 675482 687440
rect 675538 687384 675543 687440
rect 670325 687382 675543 687384
rect 670325 687379 670391 687382
rect 675477 687379 675543 687382
rect 35617 687306 35683 687309
rect 35604 687304 35683 687306
rect 35604 687248 35622 687304
rect 35678 687248 35683 687304
rect 35604 687246 35683 687248
rect 35617 687243 35683 687246
rect 44541 686898 44607 686901
rect 41492 686896 44607 686898
rect 41492 686840 44546 686896
rect 44602 686840 44607 686896
rect 41492 686838 44607 686840
rect 44541 686835 44607 686838
rect 44541 686490 44607 686493
rect 41492 686488 44607 686490
rect 41492 686432 44546 686488
rect 44602 686432 44607 686488
rect 41492 686430 44607 686432
rect 44541 686427 44607 686430
rect 674833 686490 674899 686493
rect 675334 686490 675340 686492
rect 674833 686488 675340 686490
rect 674833 686432 674838 686488
rect 674894 686432 675340 686488
rect 674833 686430 675340 686432
rect 674833 686427 674899 686430
rect 675334 686428 675340 686430
rect 675404 686428 675410 686492
rect 44909 686082 44975 686085
rect 41492 686080 44975 686082
rect 41492 686024 44914 686080
rect 44970 686024 44975 686080
rect 41492 686022 44975 686024
rect 44909 686019 44975 686022
rect 672993 685810 673059 685813
rect 675477 685810 675543 685813
rect 672993 685808 675543 685810
rect 672993 685752 672998 685808
rect 673054 685752 675482 685808
rect 675538 685752 675543 685808
rect 672993 685750 675543 685752
rect 672993 685747 673059 685750
rect 675477 685747 675543 685750
rect 45093 685674 45159 685677
rect 41492 685672 45159 685674
rect 41492 685616 45098 685672
rect 45154 685616 45159 685672
rect 41492 685614 45159 685616
rect 45093 685611 45159 685614
rect 670969 685538 671035 685541
rect 675201 685538 675267 685541
rect 670969 685536 675267 685538
rect 670969 685480 670974 685536
rect 671030 685480 675206 685536
rect 675262 685480 675267 685536
rect 670969 685478 675267 685480
rect 670969 685475 671035 685478
rect 675201 685475 675267 685478
rect 45277 685266 45343 685269
rect 41492 685264 45343 685266
rect 41492 685208 45282 685264
rect 45338 685208 45343 685264
rect 41492 685206 45343 685208
rect 45277 685203 45343 685206
rect 44909 684858 44975 684861
rect 41492 684856 44975 684858
rect 41492 684800 44914 684856
rect 44970 684800 44975 684856
rect 41492 684798 44975 684800
rect 44909 684795 44975 684798
rect 44265 684450 44331 684453
rect 41492 684448 44331 684450
rect 41492 684392 44270 684448
rect 44326 684392 44331 684448
rect 41492 684390 44331 684392
rect 44265 684387 44331 684390
rect 44357 684042 44423 684045
rect 41492 684040 44423 684042
rect 41492 683984 44362 684040
rect 44418 683984 44423 684040
rect 41492 683982 44423 683984
rect 44357 683979 44423 683982
rect 41822 683634 41828 683636
rect 41492 683574 41828 683634
rect 41822 683572 41828 683574
rect 41892 683572 41898 683636
rect 652017 683634 652083 683637
rect 650164 683632 652083 683634
rect 650164 683576 652022 683632
rect 652078 683576 652083 683632
rect 650164 683574 652083 683576
rect 652017 683571 652083 683574
rect 35801 683226 35867 683229
rect 35788 683224 35867 683226
rect 35788 683168 35806 683224
rect 35862 683168 35867 683224
rect 35788 683166 35867 683168
rect 35801 683163 35867 683166
rect 35433 682818 35499 682821
rect 35420 682816 35499 682818
rect 35420 682760 35438 682816
rect 35494 682760 35499 682816
rect 35420 682758 35499 682760
rect 35433 682755 35499 682758
rect 674414 682620 674420 682684
rect 674484 682682 674490 682684
rect 683205 682682 683271 682685
rect 674484 682680 683271 682682
rect 674484 682624 683210 682680
rect 683266 682624 683271 682680
rect 674484 682622 683271 682624
rect 674484 682620 674490 682622
rect 683205 682619 683271 682622
rect 35617 682410 35683 682413
rect 35604 682408 35683 682410
rect 35604 682352 35622 682408
rect 35678 682352 35683 682408
rect 35604 682350 35683 682352
rect 35617 682347 35683 682350
rect 674230 682348 674236 682412
rect 674300 682410 674306 682412
rect 683665 682410 683731 682413
rect 674300 682408 683731 682410
rect 674300 682352 683670 682408
rect 683726 682352 683731 682408
rect 674300 682350 683731 682352
rect 674300 682348 674306 682350
rect 683665 682347 683731 682350
rect 35801 682002 35867 682005
rect 35788 682000 35867 682002
rect 35788 681944 35806 682000
rect 35862 681944 35867 682000
rect 35788 681942 35867 681944
rect 35801 681939 35867 681942
rect 35617 681594 35683 681597
rect 35604 681592 35683 681594
rect 35604 681536 35622 681592
rect 35678 681536 35683 681592
rect 35604 681534 35683 681536
rect 35617 681531 35683 681534
rect 35801 681186 35867 681189
rect 35788 681184 35867 681186
rect 35788 681128 35806 681184
rect 35862 681128 35867 681184
rect 35788 681126 35867 681128
rect 35801 681123 35867 681126
rect 41781 681052 41847 681053
rect 41781 681050 41828 681052
rect 41736 681048 41828 681050
rect 41736 680992 41786 681048
rect 41736 680990 41828 680992
rect 41781 680988 41828 680990
rect 41892 680988 41898 681052
rect 673729 681050 673795 681053
rect 683481 681050 683547 681053
rect 673729 681048 683547 681050
rect 673729 680992 673734 681048
rect 673790 680992 683486 681048
rect 683542 680992 683547 681048
rect 673729 680990 683547 680992
rect 41781 680987 41847 680988
rect 673729 680987 673795 680990
rect 683481 680987 683547 680990
rect 35157 680778 35223 680781
rect 35157 680776 35236 680778
rect 35157 680720 35162 680776
rect 35218 680720 35236 680776
rect 35157 680718 35236 680720
rect 35157 680715 35223 680718
rect 44173 680370 44239 680373
rect 41492 680368 44239 680370
rect 41492 680312 44178 680368
rect 44234 680312 44239 680368
rect 41492 680310 44239 680312
rect 44173 680307 44239 680310
rect 42793 679962 42859 679965
rect 41492 679960 42859 679962
rect 41492 679904 42798 679960
rect 42854 679904 42859 679960
rect 41492 679902 42859 679904
rect 42793 679899 42859 679902
rect 45185 679554 45251 679557
rect 41492 679552 45251 679554
rect 41492 679496 45190 679552
rect 45246 679496 45251 679552
rect 41492 679494 45251 679496
rect 45185 679491 45251 679494
rect 43161 679146 43227 679149
rect 41492 679144 43227 679146
rect 41492 679088 43166 679144
rect 43222 679088 43227 679144
rect 41492 679086 43227 679088
rect 43161 679083 43227 679086
rect 40534 678928 40540 678992
rect 40604 678928 40610 678992
rect 40718 678928 40724 678992
rect 40788 678990 40794 678992
rect 40788 678930 41844 678990
rect 40788 678928 40794 678930
rect 40542 678708 40602 678928
rect 41784 678330 41844 678930
rect 41492 678270 41844 678330
rect 47209 677922 47275 677925
rect 41492 677920 47275 677922
rect 41492 677864 47214 677920
rect 47270 677864 47275 677920
rect 41492 677862 47275 677864
rect 47209 677859 47275 677862
rect 39990 677109 40050 677484
rect 39941 677104 40050 677109
rect 39941 677048 39946 677104
rect 40002 677076 40050 677104
rect 40002 677048 40020 677076
rect 39941 677046 40020 677048
rect 39941 677043 40007 677046
rect 45737 676698 45803 676701
rect 41492 676696 45803 676698
rect 41492 676640 45742 676696
rect 45798 676640 45803 676696
rect 41492 676638 45803 676640
rect 45737 676635 45803 676638
rect 62113 676154 62179 676157
rect 62113 676152 64492 676154
rect 62113 676096 62118 676152
rect 62174 676096 64492 676152
rect 62113 676094 64492 676096
rect 62113 676091 62179 676094
rect 42374 674188 42380 674252
rect 42444 674250 42450 674252
rect 42609 674250 42675 674253
rect 42444 674248 42675 674250
rect 42444 674192 42614 674248
rect 42670 674192 42675 674248
rect 42444 674190 42675 674192
rect 42444 674188 42450 674190
rect 42609 674187 42675 674190
rect 669957 673162 670023 673165
rect 676489 673162 676555 673165
rect 669957 673160 676555 673162
rect 669957 673104 669962 673160
rect 670018 673104 676494 673160
rect 676550 673104 676555 673160
rect 669957 673102 676555 673104
rect 669957 673099 670023 673102
rect 676489 673099 676555 673102
rect 39941 672482 40007 672485
rect 42241 672482 42307 672485
rect 39941 672480 42307 672482
rect 39941 672424 39946 672480
rect 40002 672424 42246 672480
rect 42302 672424 42307 672480
rect 39941 672422 42307 672424
rect 39941 672419 40007 672422
rect 42241 672419 42307 672422
rect 42425 672482 42491 672485
rect 42425 672480 42856 672482
rect 42425 672424 42430 672480
rect 42486 672424 42856 672480
rect 42425 672422 42856 672424
rect 42425 672419 42491 672422
rect 42796 672213 42856 672422
rect 38929 672210 38995 672213
rect 42517 672210 42583 672213
rect 38929 672208 42583 672210
rect 38929 672152 38934 672208
rect 38990 672152 42522 672208
rect 42578 672152 42583 672208
rect 38929 672150 42583 672152
rect 38929 672147 38995 672150
rect 42517 672147 42583 672150
rect 42793 672208 42859 672213
rect 42793 672152 42798 672208
rect 42854 672152 42859 672208
rect 42793 672147 42859 672152
rect 39573 671258 39639 671261
rect 40350 671258 40356 671260
rect 39573 671256 40356 671258
rect 39573 671200 39578 671256
rect 39634 671200 40356 671256
rect 39573 671198 40356 671200
rect 39573 671195 39639 671198
rect 40350 671196 40356 671198
rect 40420 671196 40426 671260
rect 41505 671258 41571 671261
rect 42006 671258 42012 671260
rect 41505 671256 42012 671258
rect 41505 671200 41510 671256
rect 41566 671200 42012 671256
rect 41505 671198 42012 671200
rect 41505 671195 41571 671198
rect 42006 671196 42012 671198
rect 42076 671196 42082 671260
rect 667197 671122 667263 671125
rect 676262 671122 676322 671364
rect 676489 671122 676555 671125
rect 667197 671120 676322 671122
rect 667197 671064 667202 671120
rect 667258 671064 676322 671120
rect 667197 671062 676322 671064
rect 676446 671120 676555 671122
rect 676446 671064 676494 671120
rect 676550 671064 676555 671120
rect 667197 671059 667263 671062
rect 676446 671059 676555 671064
rect 37917 670986 37983 670989
rect 41822 670986 41828 670988
rect 37917 670984 41828 670986
rect 37917 670928 37922 670984
rect 37978 670928 41828 670984
rect 37917 670926 41828 670928
rect 37917 670923 37983 670926
rect 41822 670924 41828 670926
rect 41892 670924 41898 670988
rect 676446 670956 676506 671059
rect 668577 670578 668643 670581
rect 668577 670576 676292 670578
rect 668577 670520 668582 670576
rect 668638 670520 676292 670576
rect 668577 670518 676292 670520
rect 668577 670515 668643 670518
rect 651465 670442 651531 670445
rect 650164 670440 651531 670442
rect 650164 670384 651470 670440
rect 651526 670384 651531 670440
rect 650164 670382 651531 670384
rect 651465 670379 651531 670382
rect 40350 670244 40356 670308
rect 40420 670306 40426 670308
rect 41781 670306 41847 670309
rect 40420 670304 41847 670306
rect 40420 670248 41786 670304
rect 41842 670248 41847 670304
rect 40420 670246 41847 670248
rect 40420 670244 40426 670246
rect 41781 670243 41847 670246
rect 672441 670306 672507 670309
rect 676489 670306 676555 670309
rect 672441 670304 676555 670306
rect 672441 670248 672446 670304
rect 672502 670248 676494 670304
rect 676550 670248 676555 670304
rect 672441 670246 676555 670248
rect 672441 670243 672507 670246
rect 676489 670243 676555 670246
rect 672809 669898 672875 669901
rect 676262 669898 676322 670140
rect 672809 669896 676322 669898
rect 672809 669840 672814 669896
rect 672870 669840 676322 669896
rect 672809 669838 676322 669840
rect 672809 669835 672875 669838
rect 672809 669490 672875 669493
rect 676262 669490 676322 669732
rect 676489 669490 676555 669493
rect 672809 669488 676322 669490
rect 672809 669432 672814 669488
rect 672870 669432 676322 669488
rect 672809 669430 676322 669432
rect 676446 669488 676555 669490
rect 676446 669432 676494 669488
rect 676550 669432 676555 669488
rect 672809 669427 672875 669430
rect 676446 669427 676555 669432
rect 42190 669292 42196 669356
rect 42260 669354 42266 669356
rect 48957 669354 49023 669357
rect 42260 669352 49023 669354
rect 42260 669296 48962 669352
rect 49018 669296 49023 669352
rect 676446 669324 676506 669427
rect 42260 669294 49023 669296
rect 42260 669292 42266 669294
rect 48957 669291 49023 669294
rect 672441 668946 672507 668949
rect 672441 668944 676292 668946
rect 672441 668888 672446 668944
rect 672502 668888 676292 668944
rect 672441 668886 676292 668888
rect 672441 668883 672507 668886
rect 41965 668538 42031 668541
rect 42374 668538 42380 668540
rect 41965 668536 42380 668538
rect 41965 668480 41970 668536
rect 42026 668480 42380 668536
rect 41965 668478 42380 668480
rect 41965 668475 42031 668478
rect 42374 668476 42380 668478
rect 42444 668476 42450 668540
rect 671613 668538 671679 668541
rect 671613 668536 676292 668538
rect 671613 668480 671618 668536
rect 671674 668480 676292 668536
rect 671613 668478 676292 668480
rect 671613 668475 671679 668478
rect 671797 668130 671863 668133
rect 671797 668128 676292 668130
rect 671797 668072 671802 668128
rect 671858 668072 676292 668128
rect 671797 668070 676292 668072
rect 671797 668067 671863 668070
rect 42190 667994 42196 667996
rect 41830 667934 42196 667994
rect 41830 667725 41890 667934
rect 42190 667932 42196 667934
rect 42260 667932 42266 667996
rect 41830 667720 41939 667725
rect 41830 667664 41878 667720
rect 41934 667664 41939 667720
rect 41830 667662 41939 667664
rect 41873 667659 41939 667662
rect 670785 667722 670851 667725
rect 670785 667720 676292 667722
rect 670785 667664 670790 667720
rect 670846 667664 676292 667720
rect 670785 667662 676292 667664
rect 670785 667659 670851 667662
rect 42006 667252 42012 667316
rect 42076 667314 42082 667316
rect 42793 667314 42859 667317
rect 42076 667312 42859 667314
rect 42076 667256 42798 667312
rect 42854 667256 42859 667312
rect 42076 667254 42859 667256
rect 42076 667252 42082 667254
rect 42793 667251 42859 667254
rect 671521 667314 671587 667317
rect 671521 667312 676292 667314
rect 671521 667256 671526 667312
rect 671582 667256 676292 667312
rect 671521 667254 676292 667256
rect 671521 667251 671587 667254
rect 683665 667042 683731 667045
rect 683622 667040 683731 667042
rect 683622 666984 683670 667040
rect 683726 666984 683731 667040
rect 683622 666979 683731 666984
rect 683622 666876 683682 666979
rect 673361 666498 673427 666501
rect 673361 666496 676292 666498
rect 673361 666440 673366 666496
rect 673422 666440 676292 666496
rect 673361 666438 676292 666440
rect 673361 666435 673427 666438
rect 669773 666226 669839 666229
rect 676489 666226 676555 666229
rect 669773 666224 676555 666226
rect 669773 666168 669778 666224
rect 669834 666168 676494 666224
rect 676550 666168 676555 666224
rect 669773 666166 676555 666168
rect 669773 666163 669839 666166
rect 676489 666163 676555 666166
rect 667565 665954 667631 665957
rect 676262 665954 676322 666060
rect 667565 665952 676322 665954
rect 667565 665896 667570 665952
rect 667626 665896 676322 665952
rect 667565 665894 676322 665896
rect 667565 665891 667631 665894
rect 40718 665348 40724 665412
rect 40788 665410 40794 665412
rect 42149 665410 42215 665413
rect 40788 665408 42215 665410
rect 40788 665352 42154 665408
rect 42210 665352 42215 665408
rect 40788 665350 42215 665352
rect 40788 665348 40794 665350
rect 42149 665347 42215 665350
rect 666461 665410 666527 665413
rect 676262 665410 676322 665652
rect 676489 665410 676555 665413
rect 666461 665408 676322 665410
rect 666461 665352 666466 665408
rect 666522 665352 676322 665408
rect 666461 665350 676322 665352
rect 676446 665408 676555 665410
rect 676446 665352 676494 665408
rect 676550 665352 676555 665408
rect 666461 665347 666527 665350
rect 676446 665347 676555 665352
rect 676446 665244 676506 665347
rect 42149 664866 42215 664869
rect 45185 664866 45251 664869
rect 42149 664864 45251 664866
rect 42149 664808 42154 664864
rect 42210 664808 45190 664864
rect 45246 664808 45251 664864
rect 42149 664806 45251 664808
rect 42149 664803 42215 664806
rect 45185 664803 45251 664806
rect 668761 664594 668827 664597
rect 676262 664594 676322 664836
rect 668761 664592 676322 664594
rect 668761 664536 668766 664592
rect 668822 664536 676322 664592
rect 668761 664534 676322 664536
rect 683205 664594 683271 664597
rect 683205 664592 683314 664594
rect 683205 664536 683210 664592
rect 683266 664536 683314 664592
rect 668761 664531 668827 664534
rect 683205 664531 683314 664536
rect 683254 664428 683314 664531
rect 40534 664124 40540 664188
rect 40604 664186 40610 664188
rect 41781 664186 41847 664189
rect 40604 664184 41847 664186
rect 40604 664128 41786 664184
rect 41842 664128 41847 664184
rect 40604 664126 41847 664128
rect 40604 664124 40610 664126
rect 41781 664123 41847 664126
rect 42241 664050 42307 664053
rect 42793 664050 42859 664053
rect 42241 664048 42859 664050
rect 42241 663992 42246 664048
rect 42302 663992 42798 664048
rect 42854 663992 42859 664048
rect 42241 663990 42859 663992
rect 42241 663987 42307 663990
rect 42793 663987 42859 663990
rect 674782 663988 674788 664052
rect 674852 664050 674858 664052
rect 674852 663990 676292 664050
rect 674852 663988 674858 663990
rect 42701 663778 42767 663781
rect 43161 663778 43227 663781
rect 42701 663776 43227 663778
rect 42701 663720 42706 663776
rect 42762 663720 43166 663776
rect 43222 663720 43227 663776
rect 42701 663718 43227 663720
rect 42701 663715 42767 663718
rect 43161 663715 43227 663718
rect 669405 663642 669471 663645
rect 669405 663640 676292 663642
rect 669405 663584 669410 663640
rect 669466 663584 676292 663640
rect 669405 663582 676292 663584
rect 669405 663579 669471 663582
rect 62113 663098 62179 663101
rect 62113 663096 64492 663098
rect 62113 663040 62118 663096
rect 62174 663040 64492 663096
rect 62113 663038 64492 663040
rect 62113 663035 62179 663038
rect 676262 662962 676322 663204
rect 683481 662962 683547 662965
rect 669270 662902 676322 662962
rect 683438 662960 683547 662962
rect 683438 662904 683486 662960
rect 683542 662904 683547 662960
rect 42057 662826 42123 662829
rect 44173 662826 44239 662829
rect 42057 662824 44239 662826
rect 42057 662768 42062 662824
rect 42118 662768 44178 662824
rect 44234 662768 44239 662824
rect 42057 662766 44239 662768
rect 42057 662763 42123 662766
rect 44173 662763 44239 662766
rect 668209 662554 668275 662557
rect 669270 662554 669330 662902
rect 683438 662899 683547 662904
rect 683438 662796 683498 662899
rect 668209 662552 669330 662554
rect 668209 662496 668214 662552
rect 668270 662496 669330 662552
rect 668209 662494 669330 662496
rect 668209 662491 668275 662494
rect 671153 662416 671219 662421
rect 671153 662360 671158 662416
rect 671214 662360 671219 662416
rect 671153 662355 671219 662360
rect 672625 662418 672691 662421
rect 672625 662416 676292 662418
rect 672625 662360 672630 662416
rect 672686 662360 676292 662416
rect 672625 662358 676292 662360
rect 672625 662355 672691 662358
rect 671156 662146 671216 662355
rect 671156 662086 676322 662146
rect 676262 661980 676322 662086
rect 672165 661602 672231 661605
rect 672165 661600 676292 661602
rect 672165 661544 672170 661600
rect 672226 661544 676292 661600
rect 672165 661542 676292 661544
rect 672165 661539 672231 661542
rect 672625 661194 672691 661197
rect 672625 661192 676292 661194
rect 672625 661136 672630 661192
rect 672686 661136 676292 661192
rect 672625 661134 676292 661136
rect 672625 661131 672691 661134
rect 42057 661058 42123 661061
rect 42701 661058 42767 661061
rect 42057 661056 42767 661058
rect 42057 661000 42062 661056
rect 42118 661000 42706 661056
rect 42762 661000 42767 661056
rect 42057 660998 42767 661000
rect 42057 660995 42123 660998
rect 42701 660995 42767 660998
rect 41454 660724 41460 660788
rect 41524 660786 41530 660788
rect 42701 660786 42767 660789
rect 41524 660784 42767 660786
rect 41524 660728 42706 660784
rect 42762 660728 42767 660784
rect 41524 660726 42767 660728
rect 41524 660724 41530 660726
rect 42701 660723 42767 660726
rect 673361 660786 673427 660789
rect 673361 660784 676292 660786
rect 673361 660728 673366 660784
rect 673422 660756 676292 660784
rect 673422 660728 676322 660756
rect 673361 660726 676322 660728
rect 673361 660723 673427 660726
rect 676262 660348 676322 660726
rect 673361 659970 673427 659973
rect 673361 659968 676292 659970
rect 673361 659912 673366 659968
rect 673422 659912 676292 659968
rect 673361 659910 676292 659912
rect 673361 659907 673427 659910
rect 41638 658548 41644 658612
rect 41708 658610 41714 658612
rect 42425 658610 42491 658613
rect 41708 658608 42491 658610
rect 41708 658552 42430 658608
rect 42486 658552 42491 658608
rect 41708 658550 42491 658552
rect 41708 658548 41714 658550
rect 42425 658547 42491 658550
rect 41822 658276 41828 658340
rect 41892 658338 41898 658340
rect 42241 658338 42307 658341
rect 41892 658336 42307 658338
rect 41892 658280 42246 658336
rect 42302 658280 42307 658336
rect 41892 658278 42307 658280
rect 41892 658276 41898 658278
rect 42241 658275 42307 658278
rect 42057 657386 42123 657389
rect 42609 657386 42675 657389
rect 42057 657384 42675 657386
rect 42057 657328 42062 657384
rect 42118 657328 42614 657384
rect 42670 657328 42675 657384
rect 42057 657326 42675 657328
rect 42057 657323 42123 657326
rect 42609 657323 42675 657326
rect 651465 657114 651531 657117
rect 650164 657112 651531 657114
rect 650164 657056 651470 657112
rect 651526 657056 651531 657112
rect 650164 657054 651531 657056
rect 651465 657051 651531 657054
rect 668209 654258 668275 654261
rect 675385 654258 675451 654261
rect 668209 654256 675451 654258
rect 668209 654200 668214 654256
rect 668270 654200 675390 654256
rect 675446 654200 675451 654256
rect 668209 654198 675451 654200
rect 668209 654195 668275 654198
rect 675385 654195 675451 654198
rect 44214 653108 44220 653172
rect 44284 653170 44290 653172
rect 44725 653170 44791 653173
rect 44284 653168 44791 653170
rect 44284 653112 44730 653168
rect 44786 653112 44791 653168
rect 44284 653110 44791 653112
rect 44284 653108 44290 653110
rect 44725 653107 44791 653110
rect 675334 652836 675340 652900
rect 675404 652898 675410 652900
rect 675569 652898 675635 652901
rect 675404 652896 675635 652898
rect 675404 652840 675574 652896
rect 675630 652840 675635 652896
rect 675404 652838 675635 652840
rect 675404 652836 675410 652838
rect 675569 652835 675635 652838
rect 675017 651538 675083 651541
rect 675385 651538 675451 651541
rect 675017 651536 675451 651538
rect 675017 651480 675022 651536
rect 675078 651480 675390 651536
rect 675446 651480 675451 651536
rect 675017 651478 675451 651480
rect 675017 651475 675083 651478
rect 675385 651475 675451 651478
rect 674782 650116 674788 650180
rect 674852 650178 674858 650180
rect 675201 650178 675267 650181
rect 674852 650176 675267 650178
rect 674852 650120 675206 650176
rect 675262 650120 675267 650176
rect 674852 650118 675267 650120
rect 674852 650116 674858 650118
rect 675201 650115 675267 650118
rect 62113 650042 62179 650045
rect 62113 650040 64492 650042
rect 62113 649984 62118 650040
rect 62174 649984 64492 650040
rect 62113 649982 64492 649984
rect 62113 649979 62179 649982
rect 674557 648954 674623 648957
rect 675385 648954 675451 648957
rect 674557 648952 675451 648954
rect 674557 648896 674562 648952
rect 674618 648896 675390 648952
rect 675446 648896 675451 648952
rect 674557 648894 675451 648896
rect 674557 648891 674623 648894
rect 675385 648891 675451 648894
rect 669037 648682 669103 648685
rect 675477 648682 675543 648685
rect 669037 648680 675543 648682
rect 669037 648624 669042 648680
rect 669098 648624 675482 648680
rect 675538 648624 675543 648680
rect 669037 648622 675543 648624
rect 669037 648619 669103 648622
rect 675477 648619 675543 648622
rect 669957 648138 670023 648141
rect 675518 648138 675524 648140
rect 669957 648136 675524 648138
rect 669957 648080 669962 648136
rect 670018 648080 675524 648136
rect 669957 648078 675524 648080
rect 669957 648075 670023 648078
rect 675518 648076 675524 648078
rect 675588 648076 675594 648140
rect 673729 647866 673795 647869
rect 675477 647866 675543 647869
rect 673729 647864 675543 647866
rect 673729 647808 673734 647864
rect 673790 647808 675482 647864
rect 675538 647808 675543 647864
rect 673729 647806 675543 647808
rect 673729 647803 673795 647806
rect 675477 647803 675543 647806
rect 674833 647596 674899 647597
rect 674782 647532 674788 647596
rect 674852 647594 674899 647596
rect 674852 647592 674944 647594
rect 674894 647536 674944 647592
rect 674852 647534 674944 647536
rect 674852 647532 674899 647534
rect 674833 647531 674899 647532
rect 675518 647458 675524 647460
rect 675296 647398 675524 647458
rect 675296 647253 675356 647398
rect 675518 647396 675524 647398
rect 675588 647396 675594 647460
rect 675293 647248 675359 647253
rect 675293 647192 675298 647248
rect 675354 647192 675359 647248
rect 675293 647187 675359 647192
rect 35801 646778 35867 646781
rect 35801 646776 35910 646778
rect 35801 646720 35806 646776
rect 35862 646720 35910 646776
rect 35801 646715 35910 646720
rect 35850 646642 35910 646715
rect 51717 646642 51783 646645
rect 35850 646640 51783 646642
rect 35850 646584 51722 646640
rect 51778 646584 51783 646640
rect 35850 646582 51783 646584
rect 51717 646579 51783 646582
rect 675293 646098 675359 646101
rect 675293 646096 675816 646098
rect 675293 646040 675298 646096
rect 675354 646040 675816 646096
rect 675293 646038 675816 646040
rect 675293 646035 675359 646038
rect 675150 645764 675156 645828
rect 675220 645826 675226 645828
rect 675477 645826 675543 645829
rect 675220 645824 675543 645826
rect 675220 645768 675482 645824
rect 675538 645768 675543 645824
rect 675220 645766 675543 645768
rect 675220 645764 675226 645766
rect 675477 645763 675543 645766
rect 675756 645557 675816 646038
rect 675753 645552 675819 645557
rect 675753 645496 675758 645552
rect 675814 645496 675819 645552
rect 675753 645491 675819 645496
rect 669773 645418 669839 645421
rect 675477 645418 675543 645421
rect 669773 645416 675543 645418
rect 669773 645360 669778 645416
rect 669834 645360 675482 645416
rect 675538 645360 675543 645416
rect 669773 645358 675543 645360
rect 669773 645355 669839 645358
rect 675477 645355 675543 645358
rect 674046 645084 674052 645148
rect 674116 645146 674122 645148
rect 674465 645146 674531 645149
rect 674116 645144 674531 645146
rect 674116 645088 674470 645144
rect 674526 645088 674531 645144
rect 674116 645086 674531 645088
rect 674116 645084 674122 645086
rect 674465 645083 674531 645086
rect 35801 644738 35867 644741
rect 35758 644736 35867 644738
rect 35758 644680 35806 644736
rect 35862 644680 35867 644736
rect 35758 644675 35867 644680
rect 41462 644738 41522 644912
rect 53097 644738 53163 644741
rect 41462 644736 53163 644738
rect 41462 644680 53102 644736
rect 53158 644680 53163 644736
rect 41462 644678 53163 644680
rect 53097 644675 53163 644678
rect 35758 644504 35818 644675
rect 674966 644268 674972 644332
rect 675036 644330 675042 644332
rect 675293 644330 675359 644333
rect 675036 644328 675359 644330
rect 675036 644272 675298 644328
rect 675354 644272 675359 644328
rect 675036 644270 675359 644272
rect 675036 644268 675042 644270
rect 675293 644267 675359 644270
rect 675753 644330 675819 644333
rect 676806 644330 676812 644332
rect 675753 644328 676812 644330
rect 675753 644272 675758 644328
rect 675814 644272 676812 644328
rect 675753 644270 676812 644272
rect 675753 644267 675819 644270
rect 676806 644268 676812 644270
rect 676876 644268 676882 644332
rect 41462 643922 41522 644096
rect 674925 644058 674991 644061
rect 675518 644058 675524 644060
rect 674925 644056 675524 644058
rect 674925 644000 674930 644056
rect 674986 644000 675524 644056
rect 674925 643998 675524 644000
rect 674925 643995 674991 643998
rect 675518 643996 675524 643998
rect 675588 643996 675594 644060
rect 41462 643862 55230 643922
rect 41462 643650 41522 643688
rect 45369 643650 45435 643653
rect 41462 643648 45435 643650
rect 41462 643592 45374 643648
rect 45430 643592 45435 643648
rect 41462 643590 45435 643592
rect 45369 643587 45435 643590
rect 44541 643378 44607 643381
rect 41462 643376 44607 643378
rect 41462 643320 44546 643376
rect 44602 643320 44607 643376
rect 41462 643318 44607 643320
rect 41462 643280 41522 643318
rect 44541 643315 44607 643318
rect 55170 643242 55230 643862
rect 651465 643786 651531 643789
rect 650164 643784 651531 643786
rect 650164 643728 651470 643784
rect 651526 643728 651531 643784
rect 650164 643726 651531 643728
rect 651465 643723 651531 643726
rect 661861 643786 661927 643789
rect 675109 643786 675175 643789
rect 661861 643784 675175 643786
rect 661861 643728 661866 643784
rect 661922 643728 675114 643784
rect 675170 643728 675175 643784
rect 661861 643726 675175 643728
rect 661861 643723 661927 643726
rect 675109 643723 675175 643726
rect 671470 643452 671476 643516
rect 671540 643514 671546 643516
rect 675477 643514 675543 643517
rect 671540 643512 675543 643514
rect 671540 643456 675482 643512
rect 675538 643456 675543 643512
rect 671540 643454 675543 643456
rect 671540 643452 671546 643454
rect 675477 643451 675543 643454
rect 55857 643242 55923 643245
rect 55170 643240 55923 643242
rect 55170 643184 55862 643240
rect 55918 643184 55923 643240
rect 55170 643182 55923 643184
rect 55857 643179 55923 643182
rect 45093 643106 45159 643109
rect 41462 643104 45159 643106
rect 41462 643048 45098 643104
rect 45154 643048 45159 643104
rect 41462 643046 45159 643048
rect 41462 642872 41522 643046
rect 45093 643043 45159 643046
rect 44725 642562 44791 642565
rect 41462 642560 44791 642562
rect 41462 642504 44730 642560
rect 44786 642504 44791 642560
rect 41462 642502 44791 642504
rect 41462 642464 41522 642502
rect 44725 642499 44791 642502
rect 44909 642290 44975 642293
rect 41462 642288 44975 642290
rect 41462 642232 44914 642288
rect 44970 642232 44975 642288
rect 41462 642230 44975 642232
rect 41462 642056 41522 642230
rect 44909 642227 44975 642230
rect 674189 641746 674255 641749
rect 675293 641746 675359 641749
rect 674189 641744 675359 641746
rect 674189 641688 674194 641744
rect 674250 641688 675298 641744
rect 675354 641688 675359 641744
rect 674189 641686 675359 641688
rect 674189 641683 674255 641686
rect 675293 641683 675359 641686
rect 41781 641678 41847 641681
rect 41492 641676 41847 641678
rect 41492 641620 41786 641676
rect 41842 641620 41847 641676
rect 41492 641618 41847 641620
rect 41781 641615 41847 641618
rect 44357 641474 44423 641477
rect 41462 641472 44423 641474
rect 41462 641416 44362 641472
rect 44418 641416 44423 641472
rect 41462 641414 44423 641416
rect 41462 641240 41522 641414
rect 44357 641411 44423 641414
rect 41781 641202 41847 641205
rect 45277 641202 45343 641205
rect 41781 641200 45343 641202
rect 41781 641144 41786 641200
rect 41842 641144 45282 641200
rect 45338 641144 45343 641200
rect 41781 641142 45343 641144
rect 41781 641139 41847 641142
rect 45277 641139 45343 641142
rect 44909 640930 44975 640933
rect 41462 640928 44975 640930
rect 41462 640872 44914 640928
rect 44970 640872 44975 640928
rect 41462 640870 44975 640872
rect 41462 640832 41522 640870
rect 44909 640867 44975 640870
rect 674925 640796 674991 640797
rect 674925 640794 674972 640796
rect 674880 640792 674972 640794
rect 674880 640736 674930 640792
rect 674880 640734 674972 640736
rect 674925 640732 674972 640734
rect 675036 640732 675042 640796
rect 674925 640731 674991 640732
rect 41638 640658 41644 640660
rect 41462 640598 41644 640658
rect 41462 640424 41522 640598
rect 41638 640596 41644 640598
rect 41708 640596 41714 640660
rect 671153 640522 671219 640525
rect 675385 640522 675451 640525
rect 671153 640520 675451 640522
rect 671153 640464 671158 640520
rect 671214 640464 675390 640520
rect 675446 640464 675451 640520
rect 671153 640462 675451 640464
rect 671153 640459 671219 640462
rect 675385 640459 675451 640462
rect 675518 640188 675524 640252
rect 675588 640250 675594 640252
rect 676622 640250 676628 640252
rect 675588 640190 676628 640250
rect 675588 640188 675594 640190
rect 676622 640188 676628 640190
rect 676692 640188 676698 640252
rect 35758 639845 35818 640016
rect 35758 639840 35867 639845
rect 35758 639784 35806 639840
rect 35862 639784 35867 639840
rect 35758 639782 35867 639784
rect 35801 639779 35867 639782
rect 41462 639436 41522 639608
rect 41454 639372 41460 639436
rect 41524 639372 41530 639436
rect 35758 639029 35818 639200
rect 35758 639024 35867 639029
rect 35758 638968 35806 639024
rect 35862 638968 35867 639024
rect 35758 638966 35867 638968
rect 35801 638963 35867 638966
rect 35758 638621 35818 638792
rect 672349 638754 672415 638757
rect 675477 638754 675543 638757
rect 672349 638752 675543 638754
rect 672349 638696 672354 638752
rect 672410 638696 675482 638752
rect 675538 638696 675543 638752
rect 672349 638694 675543 638696
rect 672349 638691 672415 638694
rect 675477 638691 675543 638694
rect 35758 638616 35867 638621
rect 35758 638560 35806 638616
rect 35862 638560 35867 638616
rect 35758 638558 35867 638560
rect 35801 638555 35867 638558
rect 32446 638213 32506 638384
rect 32397 638208 32506 638213
rect 32397 638152 32402 638208
rect 32458 638152 32506 638208
rect 32397 638150 32506 638152
rect 32397 638147 32463 638150
rect 41965 638074 42031 638077
rect 47393 638074 47459 638077
rect 41965 638072 47459 638074
rect 41965 638016 41970 638072
rect 42026 638016 47398 638072
rect 47454 638016 47459 638072
rect 41965 638014 47459 638016
rect 41965 638011 42031 638014
rect 47393 638011 47459 638014
rect 675150 638012 675156 638076
rect 675220 638074 675226 638076
rect 675385 638074 675451 638077
rect 675220 638072 675451 638074
rect 675220 638016 675390 638072
rect 675446 638016 675451 638072
rect 675220 638014 675451 638016
rect 675220 638012 675226 638014
rect 675385 638011 675451 638014
rect 41462 637802 41522 637976
rect 676622 637876 676628 637940
rect 676692 637938 676698 637940
rect 677501 637938 677567 637941
rect 676692 637936 677567 637938
rect 676692 637880 677506 637936
rect 677562 637880 677567 637936
rect 676692 637878 677567 637880
rect 676692 637876 676698 637878
rect 677501 637875 677567 637878
rect 46013 637802 46079 637805
rect 41462 637800 46079 637802
rect 41462 637744 46018 637800
rect 46074 637744 46079 637800
rect 41462 637742 46079 637744
rect 46013 637739 46079 637742
rect 675334 637604 675340 637668
rect 675404 637666 675410 637668
rect 675753 637666 675819 637669
rect 675404 637664 675819 637666
rect 675404 637608 675758 637664
rect 675814 637608 675819 637664
rect 675404 637606 675819 637608
rect 675404 637604 675410 637606
rect 675753 637603 675819 637606
rect 41965 637598 42031 637601
rect 41492 637596 42031 637598
rect 41492 637540 41970 637596
rect 42026 637540 42031 637596
rect 41492 637538 42031 637540
rect 41965 637535 42031 637538
rect 40033 637394 40099 637397
rect 41822 637394 41828 637396
rect 40033 637392 41828 637394
rect 40033 637336 40038 637392
rect 40094 637336 41828 637392
rect 40033 637334 41828 637336
rect 40033 637331 40099 637334
rect 41822 637332 41828 637334
rect 41892 637332 41898 637396
rect 41462 636986 41522 637160
rect 62113 637122 62179 637125
rect 62113 637120 64492 637122
rect 62113 637064 62118 637120
rect 62174 637064 64492 637120
rect 62113 637062 64492 637064
rect 62113 637059 62179 637062
rect 46197 636986 46263 636989
rect 41462 636984 46263 636986
rect 41462 636928 46202 636984
rect 46258 636928 46263 636984
rect 41462 636926 46263 636928
rect 46197 636923 46263 636926
rect 673545 636850 673611 636853
rect 683389 636850 683455 636853
rect 673545 636848 683455 636850
rect 673545 636792 673550 636848
rect 673606 636792 683394 636848
rect 683450 636792 683455 636848
rect 673545 636790 683455 636792
rect 673545 636787 673611 636790
rect 683389 636787 683455 636790
rect 41462 636578 41522 636752
rect 44173 636578 44239 636581
rect 41462 636576 44239 636578
rect 41462 636520 44178 636576
rect 44234 636520 44239 636576
rect 41462 636518 44239 636520
rect 44173 636515 44239 636518
rect 41462 636306 41522 636344
rect 43161 636306 43227 636309
rect 41462 636304 43227 636306
rect 41462 636248 43166 636304
rect 43222 636248 43227 636304
rect 41462 636246 43227 636248
rect 43161 636243 43227 636246
rect 41462 635762 41522 635936
rect 44909 635762 44975 635765
rect 41462 635760 44975 635762
rect 41462 635704 44914 635760
rect 44970 635704 44975 635760
rect 41462 635702 44975 635704
rect 44909 635699 44975 635702
rect 41462 635354 41522 635528
rect 672165 635490 672231 635493
rect 683205 635490 683271 635493
rect 672165 635488 683271 635490
rect 672165 635432 672170 635488
rect 672226 635432 683210 635488
rect 683266 635432 683271 635488
rect 672165 635430 683271 635432
rect 672165 635427 672231 635430
rect 683205 635427 683271 635430
rect 43897 635354 43963 635357
rect 41462 635352 43963 635354
rect 41462 635296 43902 635352
rect 43958 635296 43963 635352
rect 41462 635294 43963 635296
rect 43897 635291 43963 635294
rect 40726 634948 40786 635120
rect 40718 634884 40724 634948
rect 40788 634884 40794 634948
rect 40542 634540 40602 634712
rect 40534 634476 40540 634540
rect 40604 634476 40610 634540
rect 41462 633858 41522 634304
rect 42333 633858 42399 633861
rect 41462 633856 42399 633858
rect 41462 633800 42338 633856
rect 42394 633800 42399 633856
rect 41462 633798 42399 633800
rect 42333 633795 42399 633798
rect 41462 633450 41522 633488
rect 45369 633450 45435 633453
rect 41462 633448 45435 633450
rect 41462 633392 45374 633448
rect 45430 633392 45435 633448
rect 41462 633390 45435 633392
rect 45369 633387 45435 633390
rect 674925 631410 674991 631413
rect 675334 631410 675340 631412
rect 674925 631408 675340 631410
rect 674925 631352 674930 631408
rect 674986 631352 675340 631408
rect 674925 631350 675340 631352
rect 674925 631347 674991 631350
rect 675334 631348 675340 631350
rect 675404 631348 675410 631412
rect 675753 631410 675819 631413
rect 676070 631410 676076 631412
rect 675753 631408 676076 631410
rect 675753 631352 675758 631408
rect 675814 631352 676076 631408
rect 675753 631350 676076 631352
rect 675753 631347 675819 631350
rect 676070 631348 676076 631350
rect 676140 631348 676146 631412
rect 651465 630594 651531 630597
rect 650164 630592 651531 630594
rect 650164 630536 651470 630592
rect 651526 630536 651531 630592
rect 650164 630534 651531 630536
rect 651465 630531 651531 630534
rect 671521 627874 671587 627877
rect 675845 627874 675911 627877
rect 671521 627872 675911 627874
rect 671521 627816 671526 627872
rect 671582 627816 675850 627872
rect 675906 627816 675911 627872
rect 671521 627814 675911 627816
rect 671521 627811 671587 627814
rect 675845 627811 675911 627814
rect 41413 627738 41479 627741
rect 41822 627738 41828 627740
rect 41413 627736 41828 627738
rect 41413 627680 41418 627736
rect 41474 627680 41828 627736
rect 41413 627678 41828 627680
rect 41413 627675 41479 627678
rect 41822 627676 41828 627678
rect 41892 627676 41898 627740
rect 42701 627330 42767 627333
rect 50337 627330 50403 627333
rect 42701 627328 50403 627330
rect 42701 627272 42706 627328
rect 42762 627272 50342 627328
rect 50398 627272 50403 627328
rect 42701 627270 50403 627272
rect 42701 627267 42767 627270
rect 50337 627267 50403 627270
rect 665817 626106 665883 626109
rect 676262 626106 676322 626348
rect 665817 626104 676322 626106
rect 665817 626048 665822 626104
rect 665878 626048 676322 626104
rect 665817 626046 676322 626048
rect 665817 626043 665883 626046
rect 676262 625698 676322 625940
rect 676489 625698 676555 625701
rect 669270 625638 676322 625698
rect 676446 625696 676555 625698
rect 676446 625640 676494 625696
rect 676550 625640 676555 625696
rect 660297 625290 660363 625293
rect 669270 625290 669330 625638
rect 676446 625635 676555 625640
rect 676446 625532 676506 625635
rect 660297 625288 669330 625290
rect 660297 625232 660302 625288
rect 660358 625232 669330 625288
rect 660297 625230 669330 625232
rect 660297 625227 660363 625230
rect 673545 625154 673611 625157
rect 673545 625152 676292 625154
rect 673545 625096 673550 625152
rect 673606 625096 676292 625152
rect 673545 625094 676292 625096
rect 673545 625091 673611 625094
rect 674373 624882 674439 624885
rect 683389 624882 683455 624885
rect 674373 624880 683455 624882
rect 674373 624824 674378 624880
rect 674434 624824 683394 624880
rect 683450 624824 683455 624880
rect 674373 624822 683455 624824
rect 674373 624819 674439 624822
rect 683389 624819 683455 624822
rect 42425 624610 42491 624613
rect 43161 624610 43227 624613
rect 42425 624608 43227 624610
rect 42425 624552 42430 624608
rect 42486 624552 43166 624608
rect 43222 624552 43227 624608
rect 42425 624550 43227 624552
rect 42425 624547 42491 624550
rect 43161 624547 43227 624550
rect 671797 624474 671863 624477
rect 676446 624474 676506 624716
rect 671797 624472 676506 624474
rect 671797 624416 671802 624472
rect 671858 624416 676506 624472
rect 671797 624414 676506 624416
rect 683205 624474 683271 624477
rect 683205 624472 683314 624474
rect 683205 624416 683210 624472
rect 683266 624416 683314 624472
rect 671797 624411 671863 624414
rect 683205 624411 683314 624416
rect 683254 624308 683314 624411
rect 62113 624066 62179 624069
rect 62113 624064 64492 624066
rect 62113 624008 62118 624064
rect 62174 624008 64492 624064
rect 62113 624006 64492 624008
rect 62113 624003 62179 624006
rect 670785 623930 670851 623933
rect 670785 623928 676292 623930
rect 670785 623872 670790 623928
rect 670846 623872 676292 623928
rect 670785 623870 676292 623872
rect 670785 623867 670851 623870
rect 40718 623732 40724 623796
rect 40788 623794 40794 623796
rect 42241 623794 42307 623797
rect 40788 623792 42307 623794
rect 40788 623736 42246 623792
rect 42302 623736 42307 623792
rect 40788 623734 42307 623736
rect 40788 623732 40794 623734
rect 42241 623731 42307 623734
rect 671613 623522 671679 623525
rect 671613 623520 676292 623522
rect 671613 623464 671618 623520
rect 671674 623464 676292 623520
rect 671613 623462 676292 623464
rect 671613 623459 671679 623462
rect 42057 623386 42123 623389
rect 44265 623386 44331 623389
rect 42057 623384 44331 623386
rect 42057 623328 42062 623384
rect 42118 623328 44270 623384
rect 44326 623328 44331 623384
rect 42057 623326 44331 623328
rect 42057 623323 42123 623326
rect 44265 623323 44331 623326
rect 671705 623114 671771 623117
rect 671705 623112 676292 623114
rect 671705 623056 671710 623112
rect 671766 623056 676292 623112
rect 671705 623054 676292 623056
rect 671705 623051 671771 623054
rect 671521 622706 671587 622709
rect 671521 622704 676292 622706
rect 671521 622648 671526 622704
rect 671582 622648 676292 622704
rect 671521 622646 676292 622648
rect 671521 622643 671587 622646
rect 673177 622298 673243 622301
rect 673177 622296 676292 622298
rect 673177 622240 673182 622296
rect 673238 622240 676292 622296
rect 673177 622238 676292 622240
rect 673177 622235 673243 622238
rect 677501 622026 677567 622029
rect 677501 622024 677610 622026
rect 677501 621968 677506 622024
rect 677562 621968 677610 622024
rect 677501 621963 677610 621968
rect 677550 621860 677610 621963
rect 672993 621618 673059 621621
rect 676489 621618 676555 621621
rect 672993 621616 676555 621618
rect 672993 621560 672998 621616
rect 673054 621560 676494 621616
rect 676550 621560 676555 621616
rect 672993 621558 676555 621560
rect 672993 621555 673059 621558
rect 676489 621555 676555 621558
rect 667749 621210 667815 621213
rect 676262 621210 676322 621452
rect 676489 621210 676555 621213
rect 667749 621208 676322 621210
rect 667749 621152 667754 621208
rect 667810 621152 676322 621208
rect 667749 621150 676322 621152
rect 676446 621208 676555 621210
rect 676446 621152 676494 621208
rect 676550 621152 676555 621208
rect 667749 621147 667815 621150
rect 676446 621147 676555 621152
rect 676446 621044 676506 621147
rect 42057 620938 42123 620941
rect 43897 620938 43963 620941
rect 42057 620936 43963 620938
rect 42057 620880 42062 620936
rect 42118 620880 43902 620936
rect 43958 620880 43963 620936
rect 42057 620878 43963 620880
rect 42057 620875 42123 620878
rect 43897 620875 43963 620878
rect 42241 620666 42307 620669
rect 44081 620666 44147 620669
rect 42241 620664 44147 620666
rect 42241 620608 42246 620664
rect 42302 620608 44086 620664
rect 44142 620608 44147 620664
rect 42241 620606 44147 620608
rect 42241 620603 42307 620606
rect 44081 620603 44147 620606
rect 669589 620666 669655 620669
rect 669589 620664 676292 620666
rect 669589 620608 669594 620664
rect 669650 620608 676292 620664
rect 669589 620606 676292 620608
rect 669589 620603 669655 620606
rect 42425 620394 42491 620397
rect 47393 620394 47459 620397
rect 42425 620392 47459 620394
rect 42425 620336 42430 620392
rect 42486 620336 47398 620392
rect 47454 620336 47459 620392
rect 42425 620334 47459 620336
rect 42425 620331 42491 620334
rect 47393 620331 47459 620334
rect 41781 620260 41847 620261
rect 41781 620256 41828 620260
rect 41892 620258 41898 620260
rect 668393 620258 668459 620261
rect 41781 620200 41786 620256
rect 41781 620196 41828 620200
rect 41892 620198 41938 620258
rect 668393 620256 676292 620258
rect 668393 620200 668398 620256
rect 668454 620200 676292 620256
rect 668393 620198 676292 620200
rect 41892 620196 41898 620198
rect 41781 620195 41847 620196
rect 668393 620195 668459 620198
rect 40534 619924 40540 619988
rect 40604 619986 40610 619988
rect 42701 619986 42767 619989
rect 40604 619984 42767 619986
rect 40604 619928 42706 619984
rect 42762 619928 42767 619984
rect 40604 619926 42767 619928
rect 40604 619924 40610 619926
rect 42701 619923 42767 619926
rect 672165 619850 672231 619853
rect 672165 619848 676292 619850
rect 672165 619792 672170 619848
rect 672226 619792 676292 619848
rect 672165 619790 676292 619792
rect 672165 619787 672231 619790
rect 670601 619442 670667 619445
rect 670601 619440 676292 619442
rect 670601 619384 670606 619440
rect 670662 619384 676292 619440
rect 670601 619382 676292 619384
rect 670601 619379 670667 619382
rect 676990 619108 676996 619172
rect 677060 619108 677066 619172
rect 42425 619034 42491 619037
rect 46197 619034 46263 619037
rect 42425 619032 46263 619034
rect 42425 618976 42430 619032
rect 42486 618976 46202 619032
rect 46258 618976 46263 619032
rect 676998 619004 677058 619108
rect 42425 618974 46263 618976
rect 42425 618971 42491 618974
rect 46197 618971 46263 618974
rect 674741 618626 674807 618629
rect 674741 618624 676292 618626
rect 674741 618568 674746 618624
rect 674802 618568 676292 618624
rect 674741 618566 676292 618568
rect 674741 618563 674807 618566
rect 670325 618218 670391 618221
rect 670325 618216 676292 618218
rect 670325 618160 670330 618216
rect 670386 618160 676292 618216
rect 670325 618158 676292 618160
rect 670325 618155 670391 618158
rect 683573 617946 683639 617949
rect 683573 617944 683682 617946
rect 683573 617888 683578 617944
rect 683634 617888 683682 617944
rect 683573 617883 683682 617888
rect 683622 617780 683682 617883
rect 673913 617402 673979 617405
rect 673913 617400 676292 617402
rect 673913 617344 673918 617400
rect 673974 617344 676292 617400
rect 673913 617342 676292 617344
rect 673913 617339 673979 617342
rect 651465 617266 651531 617269
rect 650164 617264 651531 617266
rect 650164 617208 651470 617264
rect 651526 617208 651531 617264
rect 650164 617206 651531 617208
rect 651465 617203 651531 617206
rect 683389 617130 683455 617133
rect 683389 617128 683498 617130
rect 683389 617072 683394 617128
rect 683450 617072 683498 617128
rect 683389 617067 683498 617072
rect 683438 616964 683498 617067
rect 672165 616722 672231 616725
rect 672165 616720 676322 616722
rect 672165 616664 672170 616720
rect 672226 616664 676322 616720
rect 672165 616662 676322 616664
rect 672165 616659 672231 616662
rect 676262 616556 676322 616662
rect 673862 616116 673868 616180
rect 673932 616178 673938 616180
rect 673932 616118 676292 616178
rect 673932 616116 673938 616118
rect 42057 615908 42123 615909
rect 42006 615906 42012 615908
rect 41966 615846 42012 615906
rect 42076 615904 42123 615908
rect 42118 615848 42123 615904
rect 42006 615844 42012 615846
rect 42076 615844 42123 615848
rect 42057 615843 42123 615844
rect 672901 615770 672967 615773
rect 672901 615768 676292 615770
rect 672901 615712 672906 615768
rect 672962 615740 676292 615768
rect 672962 615712 676322 615740
rect 672901 615710 676322 615712
rect 672901 615707 672967 615710
rect 46013 615634 46079 615637
rect 42704 615632 46079 615634
rect 42704 615576 46018 615632
rect 46074 615576 46079 615632
rect 42704 615574 46079 615576
rect 41454 615436 41460 615500
rect 41524 615498 41530 615500
rect 42425 615498 42491 615501
rect 41524 615496 42491 615498
rect 41524 615440 42430 615496
rect 42486 615440 42491 615496
rect 41524 615438 42491 615440
rect 41524 615436 41530 615438
rect 42425 615435 42491 615438
rect 42057 615226 42123 615229
rect 42704 615226 42764 615574
rect 46013 615571 46079 615574
rect 676262 615332 676322 615710
rect 42057 615224 42764 615226
rect 42057 615168 42062 615224
rect 42118 615168 42764 615224
rect 42057 615166 42764 615168
rect 42057 615163 42123 615166
rect 671981 614954 672047 614957
rect 671981 614952 676292 614954
rect 671981 614896 671986 614952
rect 672042 614896 676292 614952
rect 671981 614894 676292 614896
rect 671981 614891 672047 614894
rect 41873 614140 41939 614141
rect 41822 614138 41828 614140
rect 41782 614078 41828 614138
rect 41892 614136 41939 614140
rect 44173 614140 44239 614141
rect 44173 614138 44220 614140
rect 41934 614080 41939 614136
rect 41822 614076 41828 614078
rect 41892 614076 41939 614080
rect 44128 614136 44220 614138
rect 44128 614080 44178 614136
rect 44128 614078 44220 614080
rect 41873 614075 41939 614076
rect 44173 614076 44220 614078
rect 44284 614076 44290 614140
rect 44173 614075 44239 614076
rect 42977 612370 43043 612373
rect 43575 612370 43641 612373
rect 42977 612368 43641 612370
rect 42977 612312 42982 612368
rect 43038 612312 43580 612368
rect 43636 612312 43641 612368
rect 42977 612310 43641 612312
rect 42977 612307 43043 612310
rect 43575 612307 43641 612310
rect 42701 611010 42767 611013
rect 44265 611010 44331 611013
rect 42701 611008 44331 611010
rect 42701 610952 42706 611008
rect 42762 610952 44270 611008
rect 44326 610952 44331 611008
rect 42701 610950 44331 610952
rect 42701 610947 42767 610950
rect 44265 610947 44331 610950
rect 62113 611010 62179 611013
rect 62113 611008 64492 611010
rect 62113 610952 62118 611008
rect 62174 610952 64492 611008
rect 62113 610950 64492 610952
rect 62113 610947 62179 610950
rect 675477 608292 675543 608293
rect 675477 608288 675524 608292
rect 675588 608290 675594 608292
rect 675477 608232 675482 608288
rect 675477 608228 675524 608232
rect 675588 608230 675634 608290
rect 675588 608228 675594 608230
rect 675477 608227 675543 608228
rect 670601 608018 670667 608021
rect 675477 608018 675543 608021
rect 670601 608016 675543 608018
rect 670601 607960 670606 608016
rect 670662 607960 675482 608016
rect 675538 607960 675543 608016
rect 670601 607958 675543 607960
rect 670601 607955 670667 607958
rect 675477 607955 675543 607958
rect 674373 606522 674439 606525
rect 675477 606522 675543 606525
rect 674373 606520 675543 606522
rect 674373 606464 674378 606520
rect 674434 606464 675482 606520
rect 675538 606464 675543 606520
rect 674373 606462 675543 606464
rect 674373 606459 674439 606462
rect 675477 606459 675543 606462
rect 672165 604754 672231 604757
rect 675477 604754 675543 604757
rect 672165 604752 675543 604754
rect 672165 604696 672170 604752
rect 672226 604696 675482 604752
rect 675538 604696 675543 604752
rect 672165 604694 675543 604696
rect 672165 604691 672231 604694
rect 675477 604691 675543 604694
rect 672533 604346 672599 604349
rect 675477 604346 675543 604349
rect 672533 604344 675543 604346
rect 672533 604288 672538 604344
rect 672594 604288 675482 604344
rect 675538 604288 675543 604344
rect 672533 604286 675543 604288
rect 672533 604283 672599 604286
rect 675477 604283 675543 604286
rect 651465 603938 651531 603941
rect 650164 603936 651531 603938
rect 650164 603880 651470 603936
rect 651526 603880 651531 603936
rect 650164 603878 651531 603880
rect 651465 603875 651531 603878
rect 673545 603530 673611 603533
rect 675477 603530 675543 603533
rect 673545 603528 675543 603530
rect 673545 603472 673550 603528
rect 673606 603472 675482 603528
rect 675538 603472 675543 603528
rect 673545 603470 675543 603472
rect 673545 603467 673611 603470
rect 675477 603467 675543 603470
rect 666461 603122 666527 603125
rect 674833 603122 674899 603125
rect 666461 603120 674899 603122
rect 666461 603064 666466 603120
rect 666522 603064 674838 603120
rect 674894 603064 674899 603120
rect 666461 603062 674899 603064
rect 666461 603059 666527 603062
rect 674833 603059 674899 603062
rect 674414 602788 674420 602852
rect 674484 602850 674490 602852
rect 675477 602850 675543 602853
rect 674484 602848 675543 602850
rect 674484 602792 675482 602848
rect 675538 602792 675543 602848
rect 674484 602790 675543 602792
rect 674484 602788 674490 602790
rect 675477 602787 675543 602790
rect 51717 601762 51783 601765
rect 41492 601760 51783 601762
rect 41492 601704 51722 601760
rect 51778 601704 51783 601760
rect 41492 601702 51783 601704
rect 51717 601699 51783 601702
rect 668393 601762 668459 601765
rect 675017 601762 675083 601765
rect 668393 601760 675083 601762
rect 668393 601704 668398 601760
rect 668454 601704 675022 601760
rect 675078 601704 675083 601760
rect 668393 601702 675083 601704
rect 668393 601699 668459 601702
rect 675017 601699 675083 601702
rect 48957 601354 49023 601357
rect 41492 601352 49023 601354
rect 41492 601296 48962 601352
rect 49018 601296 49023 601352
rect 41492 601294 49023 601296
rect 48957 601291 49023 601294
rect 674833 601082 674899 601085
rect 675477 601082 675543 601085
rect 674833 601080 675543 601082
rect 674833 601024 674838 601080
rect 674894 601024 675482 601080
rect 675538 601024 675543 601080
rect 674833 601022 675543 601024
rect 674833 601019 674899 601022
rect 675477 601019 675543 601022
rect 54477 600946 54543 600949
rect 41492 600944 54543 600946
rect 41492 600888 54482 600944
rect 54538 600888 54543 600944
rect 41492 600886 54543 600888
rect 54477 600883 54543 600886
rect 44541 600538 44607 600541
rect 41492 600536 44607 600538
rect 41492 600480 44546 600536
rect 44602 600480 44607 600536
rect 41492 600478 44607 600480
rect 44541 600475 44607 600478
rect 675017 600538 675083 600541
rect 675477 600538 675543 600541
rect 675017 600536 675543 600538
rect 675017 600480 675022 600536
rect 675078 600480 675482 600536
rect 675538 600480 675543 600536
rect 675017 600478 675543 600480
rect 675017 600475 675083 600478
rect 675477 600475 675543 600478
rect 44633 600130 44699 600133
rect 41492 600128 44699 600130
rect 41492 600072 44638 600128
rect 44694 600072 44699 600128
rect 41492 600070 44699 600072
rect 44633 600067 44699 600070
rect 44817 599722 44883 599725
rect 41492 599720 44883 599722
rect 41492 599664 44822 599720
rect 44878 599664 44883 599720
rect 41492 599662 44883 599664
rect 44817 599659 44883 599662
rect 660297 599586 660363 599589
rect 674005 599586 674071 599589
rect 660297 599584 663810 599586
rect 660297 599528 660302 599584
rect 660358 599528 663810 599584
rect 660297 599526 663810 599528
rect 660297 599523 660363 599526
rect 44817 599314 44883 599317
rect 41492 599312 44883 599314
rect 41492 599256 44822 599312
rect 44878 599256 44883 599312
rect 41492 599254 44883 599256
rect 44817 599251 44883 599254
rect 663750 599042 663810 599526
rect 674005 599584 675770 599586
rect 674005 599528 674010 599584
rect 674066 599528 675770 599584
rect 674005 599526 675770 599528
rect 674005 599523 674071 599526
rect 674005 599314 674071 599317
rect 675477 599314 675543 599317
rect 674005 599312 675543 599314
rect 674005 599256 674010 599312
rect 674066 599256 675482 599312
rect 675538 599256 675543 599312
rect 674005 599254 675543 599256
rect 674005 599251 674071 599254
rect 675477 599251 675543 599254
rect 675710 599181 675770 599526
rect 675661 599176 675770 599181
rect 675661 599120 675666 599176
rect 675722 599120 675770 599176
rect 675661 599118 675770 599120
rect 675661 599115 675727 599118
rect 675017 599042 675083 599045
rect 663750 599040 675083 599042
rect 663750 598984 675022 599040
rect 675078 598984 675083 599040
rect 663750 598982 675083 598984
rect 675017 598979 675083 598982
rect 45185 598906 45251 598909
rect 41492 598904 45251 598906
rect 41492 598848 45190 598904
rect 45246 598848 45251 598904
rect 41492 598846 45251 598848
rect 45185 598843 45251 598846
rect 45185 598498 45251 598501
rect 41492 598496 45251 598498
rect 41492 598440 45190 598496
rect 45246 598440 45251 598496
rect 41492 598438 45251 598440
rect 45185 598435 45251 598438
rect 45001 598090 45067 598093
rect 41492 598088 45067 598090
rect 41492 598032 45006 598088
rect 45062 598032 45067 598088
rect 41492 598030 45067 598032
rect 45001 598027 45067 598030
rect 670325 598090 670391 598093
rect 675477 598090 675543 598093
rect 670325 598088 675543 598090
rect 670325 598032 670330 598088
rect 670386 598032 675482 598088
rect 675538 598032 675543 598088
rect 670325 598030 675543 598032
rect 670325 598027 670391 598030
rect 675477 598027 675543 598030
rect 62113 597954 62179 597957
rect 62113 597952 64492 597954
rect 62113 597896 62118 597952
rect 62174 597896 64492 597952
rect 62113 597894 64492 597896
rect 62113 597891 62179 597894
rect 41492 597622 42994 597682
rect 40309 597274 40375 597277
rect 40309 597272 40388 597274
rect 40309 597216 40314 597272
rect 40370 597216 40388 597272
rect 40309 597214 40388 597216
rect 40309 597211 40375 597214
rect 42934 597005 42994 597622
rect 42934 597000 43043 597005
rect 42934 596944 42982 597000
rect 43038 596944 43043 597000
rect 42934 596942 43043 596944
rect 42977 596939 43043 596942
rect 42609 596866 42675 596869
rect 41492 596864 42675 596866
rect 41492 596808 42614 596864
rect 42670 596808 42675 596864
rect 41492 596806 42675 596808
rect 42609 596803 42675 596806
rect 675017 596866 675083 596869
rect 675477 596866 675543 596869
rect 675017 596864 675543 596866
rect 675017 596808 675022 596864
rect 675078 596808 675482 596864
rect 675538 596808 675543 596864
rect 675017 596806 675543 596808
rect 675017 596803 675083 596806
rect 675477 596803 675543 596806
rect 40910 596223 40970 596428
rect 40861 596218 40970 596223
rect 41137 596220 41203 596223
rect 40861 596162 40866 596218
rect 40922 596162 40970 596218
rect 40861 596160 40970 596162
rect 41094 596218 41203 596220
rect 41094 596162 41142 596218
rect 41198 596162 41203 596218
rect 40861 596157 40927 596160
rect 41094 596157 41203 596162
rect 41094 596020 41154 596157
rect 41781 596052 41847 596053
rect 41781 596048 41828 596052
rect 41892 596050 41898 596052
rect 41781 595992 41786 596048
rect 41781 595988 41828 595992
rect 41892 595990 41938 596050
rect 41892 595988 41898 595990
rect 41781 595987 41847 595988
rect 32397 595642 32463 595645
rect 673637 595642 673703 595645
rect 674782 595642 674788 595644
rect 32397 595640 32476 595642
rect 32397 595584 32402 595640
rect 32458 595584 32476 595640
rect 32397 595582 32476 595584
rect 673637 595640 674788 595642
rect 673637 595584 673642 595640
rect 673698 595584 674788 595640
rect 673637 595582 674788 595584
rect 32397 595579 32463 595582
rect 673637 595579 673703 595582
rect 674782 595580 674788 595582
rect 674852 595580 674858 595644
rect 674925 595506 674991 595509
rect 675385 595506 675451 595509
rect 674925 595504 675451 595506
rect 674925 595448 674930 595504
rect 674986 595448 675390 595504
rect 675446 595448 675451 595504
rect 674925 595446 675451 595448
rect 674925 595443 674991 595446
rect 675385 595443 675451 595446
rect 673678 595308 673684 595372
rect 673748 595370 673754 595372
rect 674005 595370 674071 595373
rect 673748 595368 674071 595370
rect 673748 595312 674010 595368
rect 674066 595312 674071 595368
rect 673748 595310 674071 595312
rect 673748 595308 673754 595310
rect 674005 595307 674071 595310
rect 36537 595234 36603 595237
rect 36524 595232 36603 595234
rect 36524 595176 36542 595232
rect 36598 595176 36603 595232
rect 36524 595174 36603 595176
rect 36537 595171 36603 595174
rect 41689 594962 41755 594965
rect 42006 594962 42012 594964
rect 41689 594960 42012 594962
rect 41689 594904 41694 594960
rect 41750 594904 42012 594960
rect 41689 594902 42012 594904
rect 41689 594899 41755 594902
rect 42006 594900 42012 594902
rect 42076 594900 42082 594964
rect 37917 594826 37983 594829
rect 671245 594826 671311 594829
rect 675477 594826 675543 594829
rect 37917 594824 37996 594826
rect 37917 594768 37922 594824
rect 37978 594768 37996 594824
rect 37917 594766 37996 594768
rect 671245 594824 675543 594826
rect 671245 594768 671250 594824
rect 671306 594768 675482 594824
rect 675538 594768 675543 594824
rect 671245 594766 675543 594768
rect 37917 594763 37983 594766
rect 671245 594763 671311 594766
rect 675477 594763 675543 594766
rect 35157 594418 35223 594421
rect 35157 594416 35236 594418
rect 35157 594360 35162 594416
rect 35218 594360 35236 594416
rect 35157 594358 35236 594360
rect 35157 594355 35223 594358
rect 42793 594010 42859 594013
rect 41492 594008 42859 594010
rect 41492 593952 42798 594008
rect 42854 593952 42859 594008
rect 41492 593950 42859 593952
rect 42793 593947 42859 593950
rect 668853 593738 668919 593741
rect 675385 593738 675451 593741
rect 668853 593736 675451 593738
rect 668853 593680 668858 593736
rect 668914 593680 675390 593736
rect 675446 593680 675451 593736
rect 668853 593678 675451 593680
rect 668853 593675 668919 593678
rect 675385 593675 675451 593678
rect 41781 593602 41847 593605
rect 41492 593600 41847 593602
rect 41492 593544 41786 593600
rect 41842 593544 41847 593600
rect 41492 593542 41847 593544
rect 41781 593539 41847 593542
rect 676070 593404 676076 593468
rect 676140 593466 676146 593468
rect 676990 593466 676996 593468
rect 676140 593406 676996 593466
rect 676140 593404 676146 593406
rect 676990 593404 676996 593406
rect 677060 593404 677066 593468
rect 41781 593194 41847 593197
rect 41492 593192 41847 593194
rect 41492 593136 41786 593192
rect 41842 593136 41847 593192
rect 41492 593134 41847 593136
rect 41781 593131 41847 593134
rect 674281 592922 674347 592925
rect 683297 592922 683363 592925
rect 674281 592920 683363 592922
rect 674281 592864 674286 592920
rect 674342 592864 683302 592920
rect 683358 592864 683363 592920
rect 674281 592862 683363 592864
rect 674281 592859 674347 592862
rect 683297 592859 683363 592862
rect 41781 592786 41847 592789
rect 41492 592784 41847 592786
rect 41492 592728 41786 592784
rect 41842 592728 41847 592784
rect 41492 592726 41847 592728
rect 41781 592723 41847 592726
rect 674649 592650 674715 592653
rect 683481 592650 683547 592653
rect 674649 592648 683547 592650
rect 674649 592592 674654 592648
rect 674710 592592 683486 592648
rect 683542 592592 683547 592648
rect 674649 592590 683547 592592
rect 674649 592587 674715 592590
rect 683481 592587 683547 592590
rect 40718 592350 40724 592414
rect 40788 592350 40794 592414
rect 40726 592348 40786 592350
rect 675334 592316 675340 592380
rect 675404 592378 675410 592380
rect 675753 592378 675819 592381
rect 675404 592376 675819 592378
rect 675404 592320 675758 592376
rect 675814 592320 675819 592376
rect 675404 592318 675819 592320
rect 675404 592316 675410 592318
rect 675753 592315 675819 592318
rect 675569 592108 675635 592109
rect 675518 592106 675524 592108
rect 675478 592046 675524 592106
rect 675588 592104 675635 592108
rect 675630 592048 675635 592104
rect 675518 592044 675524 592046
rect 675588 592044 675635 592048
rect 675569 592043 675635 592044
rect 44449 591970 44515 591973
rect 41492 591968 44515 591970
rect 41492 591912 44454 591968
rect 44510 591912 44515 591968
rect 41492 591910 44515 591912
rect 44449 591907 44515 591910
rect 673678 591636 673684 591700
rect 673748 591698 673754 591700
rect 673913 591698 673979 591701
rect 673748 591696 673979 591698
rect 673748 591640 673918 591696
rect 673974 591640 673979 591696
rect 673748 591638 673979 591640
rect 673748 591636 673754 591638
rect 673913 591635 673979 591638
rect 43846 591562 43852 591564
rect 41492 591502 43852 591562
rect 43846 591500 43852 591502
rect 43916 591500 43922 591564
rect 674782 591364 674788 591428
rect 674852 591426 674858 591428
rect 683757 591426 683823 591429
rect 674852 591424 683823 591426
rect 674852 591368 683762 591424
rect 683818 591368 683823 591424
rect 674852 591366 683823 591368
rect 674852 591364 674858 591366
rect 683757 591363 683823 591366
rect 39990 590749 40050 591124
rect 39941 590744 40050 590749
rect 651465 590746 651531 590749
rect 39941 590688 39946 590744
rect 40002 590716 40050 590744
rect 650164 590744 651531 590746
rect 40002 590688 40020 590716
rect 39941 590686 40020 590688
rect 650164 590688 651470 590744
rect 651526 590688 651531 590744
rect 650164 590686 651531 590688
rect 39941 590683 40007 590686
rect 651465 590683 651531 590686
rect 43437 590338 43503 590341
rect 41492 590336 43503 590338
rect 41492 590280 43442 590336
rect 43498 590280 43503 590336
rect 41492 590278 43503 590280
rect 43437 590275 43503 590278
rect 40953 589660 41019 589661
rect 40902 589658 40908 589660
rect 40862 589598 40908 589658
rect 40972 589656 41019 589660
rect 41014 589600 41019 589656
rect 40902 589596 40908 589598
rect 40972 589596 41019 589600
rect 40953 589595 41019 589596
rect 40534 589324 40540 589388
rect 40604 589386 40610 589388
rect 41781 589386 41847 589389
rect 40604 589384 41847 589386
rect 40604 589328 41786 589384
rect 41842 589328 41847 589384
rect 40604 589326 41847 589328
rect 40604 589324 40610 589326
rect 41781 589323 41847 589326
rect 41454 587148 41460 587212
rect 41524 587210 41530 587212
rect 42006 587210 42012 587212
rect 41524 587150 42012 587210
rect 41524 587148 41530 587150
rect 42006 587148 42012 587150
rect 42076 587148 42082 587212
rect 675569 586258 675635 586261
rect 676070 586258 676076 586260
rect 675569 586256 676076 586258
rect 675569 586200 675574 586256
rect 675630 586200 676076 586256
rect 675569 586198 676076 586200
rect 675569 586195 675635 586198
rect 676070 586196 676076 586198
rect 676140 586196 676146 586260
rect 42374 586060 42380 586124
rect 42444 586122 42450 586124
rect 42701 586122 42767 586125
rect 42444 586120 42767 586122
rect 42444 586064 42706 586120
rect 42762 586064 42767 586120
rect 42444 586062 42767 586064
rect 42444 586060 42450 586062
rect 42701 586059 42767 586062
rect 39941 585986 40007 585989
rect 42241 585986 42307 585989
rect 39941 585984 42307 585986
rect 39941 585928 39946 585984
rect 40002 585928 42246 585984
rect 42302 585928 42307 585984
rect 39941 585926 42307 585928
rect 39941 585923 40007 585926
rect 42241 585923 42307 585926
rect 40493 585714 40559 585717
rect 42609 585714 42675 585717
rect 40493 585712 42675 585714
rect 40493 585656 40498 585712
rect 40554 585656 42614 585712
rect 42670 585656 42675 585712
rect 40493 585654 42675 585656
rect 40493 585651 40559 585654
rect 42609 585651 42675 585654
rect 41413 585442 41479 585445
rect 42425 585442 42491 585445
rect 41413 585440 42491 585442
rect 41413 585384 41418 585440
rect 41474 585384 42430 585440
rect 42486 585384 42491 585440
rect 41413 585382 42491 585384
rect 41413 585379 41479 585382
rect 42425 585379 42491 585382
rect 37917 585170 37983 585173
rect 41822 585170 41828 585172
rect 37917 585168 41828 585170
rect 37917 585112 37922 585168
rect 37978 585112 41828 585168
rect 37917 585110 41828 585112
rect 37917 585107 37983 585110
rect 41822 585108 41828 585110
rect 41892 585108 41898 585172
rect 39481 584898 39547 584901
rect 42190 584898 42196 584900
rect 39481 584896 42196 584898
rect 39481 584840 39486 584896
rect 39542 584840 42196 584896
rect 39481 584838 42196 584840
rect 39481 584835 39547 584838
rect 42190 584836 42196 584838
rect 42260 584836 42266 584900
rect 62113 584898 62179 584901
rect 62113 584896 64492 584898
rect 62113 584840 62118 584896
rect 62174 584840 64492 584896
rect 62113 584838 64492 584840
rect 62113 584835 62179 584838
rect 40677 584626 40743 584629
rect 41086 584626 41092 584628
rect 40677 584624 41092 584626
rect 40677 584568 40682 584624
rect 40738 584568 41092 584624
rect 40677 584566 41092 584568
rect 40677 584563 40743 584566
rect 41086 584564 41092 584566
rect 41156 584564 41162 584628
rect 652017 582994 652083 582997
rect 676029 582994 676095 582997
rect 652017 582992 676095 582994
rect 652017 582936 652022 582992
rect 652078 582936 676034 582992
rect 676090 582936 676095 582992
rect 652017 582934 676095 582936
rect 652017 582931 652083 582934
rect 676029 582931 676095 582934
rect 47577 582450 47643 582453
rect 42014 582448 47643 582450
rect 42014 582392 47582 582448
rect 47638 582392 47643 582448
rect 42014 582390 47643 582392
rect 42014 581229 42074 582390
rect 47577 582387 47643 582390
rect 42333 581908 42399 581909
rect 42333 581906 42380 581908
rect 42288 581904 42380 581906
rect 42288 581848 42338 581904
rect 42288 581846 42380 581848
rect 42333 581844 42380 581846
rect 42444 581844 42450 581908
rect 42333 581843 42399 581844
rect 42241 581500 42307 581501
rect 42190 581436 42196 581500
rect 42260 581498 42307 581500
rect 42260 581496 42352 581498
rect 42302 581440 42352 581496
rect 42260 581438 42352 581440
rect 42260 581436 42307 581438
rect 42241 581435 42307 581436
rect 42014 581224 42123 581229
rect 42014 581168 42062 581224
rect 42118 581168 42123 581224
rect 42014 581166 42123 581168
rect 42057 581163 42123 581166
rect 44449 581090 44515 581093
rect 42198 581088 44515 581090
rect 42198 581032 44454 581088
rect 44510 581032 44515 581088
rect 42198 581030 44515 581032
rect 42198 580821 42258 581030
rect 44449 581027 44515 581030
rect 661677 581090 661743 581093
rect 661677 581088 676292 581090
rect 661677 581032 661682 581088
rect 661738 581032 676292 581088
rect 661677 581030 676292 581032
rect 661677 581027 661743 581030
rect 42198 580816 42307 580821
rect 42198 580760 42246 580816
rect 42302 580760 42307 580816
rect 42198 580758 42307 580760
rect 42241 580755 42307 580758
rect 676262 580546 676322 580652
rect 669270 580486 676322 580546
rect 41086 580212 41092 580276
rect 41156 580274 41162 580276
rect 41781 580274 41847 580277
rect 41156 580272 41847 580274
rect 41156 580216 41786 580272
rect 41842 580216 41847 580272
rect 41156 580214 41847 580216
rect 41156 580212 41162 580214
rect 41781 580211 41847 580214
rect 664437 579730 664503 579733
rect 669270 579730 669330 580486
rect 676029 580274 676095 580277
rect 676029 580272 676292 580274
rect 676029 580216 676034 580272
rect 676090 580216 676292 580272
rect 676029 580214 676292 580216
rect 676029 580211 676095 580214
rect 671429 579866 671495 579869
rect 671429 579864 676292 579866
rect 671429 579808 671434 579864
rect 671490 579808 676292 579864
rect 671429 579806 676292 579808
rect 671429 579803 671495 579806
rect 664437 579728 669330 579730
rect 664437 579672 664442 579728
rect 664498 579672 669330 579728
rect 664437 579670 669330 579672
rect 664437 579667 664503 579670
rect 671429 579458 671495 579461
rect 671429 579456 676292 579458
rect 671429 579400 671434 579456
rect 671490 579400 676292 579456
rect 671429 579398 676292 579400
rect 671429 579395 671495 579398
rect 670785 579050 670851 579053
rect 670785 579048 676292 579050
rect 670785 578992 670790 579048
rect 670846 578992 676292 579048
rect 670785 578990 676292 578992
rect 670785 578987 670851 578990
rect 670785 578642 670851 578645
rect 670785 578640 676292 578642
rect 670785 578584 670790 578640
rect 670846 578584 676292 578640
rect 670785 578582 676292 578584
rect 670785 578579 670851 578582
rect 40902 578172 40908 578236
rect 40972 578234 40978 578236
rect 41781 578234 41847 578237
rect 40972 578232 41847 578234
rect 40972 578176 41786 578232
rect 41842 578176 41847 578232
rect 40972 578174 41847 578176
rect 40972 578172 40978 578174
rect 41781 578171 41847 578174
rect 671705 578234 671771 578237
rect 671705 578232 676292 578234
rect 671705 578176 671710 578232
rect 671766 578176 676292 578232
rect 671705 578174 676292 578176
rect 671705 578171 671771 578174
rect 670877 577826 670943 577829
rect 670877 577824 676292 577826
rect 670877 577768 670882 577824
rect 670938 577768 676292 577824
rect 670877 577766 676292 577768
rect 670877 577763 670943 577766
rect 40718 577492 40724 577556
rect 40788 577554 40794 577556
rect 41781 577554 41847 577557
rect 40788 577552 41847 577554
rect 40788 577496 41786 577552
rect 41842 577496 41847 577552
rect 40788 577494 41847 577496
rect 40788 577492 40794 577494
rect 41781 577491 41847 577494
rect 651465 577418 651531 577421
rect 650164 577416 651531 577418
rect 650164 577360 651470 577416
rect 651526 577360 651531 577416
rect 650164 577358 651531 577360
rect 651465 577355 651531 577358
rect 673177 577418 673243 577421
rect 673177 577416 676292 577418
rect 673177 577360 673182 577416
rect 673238 577360 676292 577416
rect 673177 577358 676292 577360
rect 673177 577355 673243 577358
rect 672441 577010 672507 577013
rect 672441 577008 676292 577010
rect 672441 576952 672446 577008
rect 672502 576952 676292 577008
rect 672441 576950 676292 576952
rect 672441 576947 672507 576950
rect 40534 576812 40540 576876
rect 40604 576874 40610 576876
rect 42241 576874 42307 576877
rect 40604 576872 42307 576874
rect 40604 576816 42246 576872
rect 42302 576816 42307 576872
rect 40604 576814 42307 576816
rect 40604 576812 40610 576814
rect 42241 576811 42307 576814
rect 675753 576602 675819 576605
rect 675753 576600 676292 576602
rect 675753 576544 675758 576600
rect 675814 576544 676292 576600
rect 675753 576542 676292 576544
rect 675753 576539 675819 576542
rect 42190 576132 42196 576196
rect 42260 576194 42266 576196
rect 42517 576194 42583 576197
rect 42260 576192 42583 576194
rect 42260 576136 42522 576192
rect 42578 576136 42583 576192
rect 42260 576134 42583 576136
rect 42260 576132 42266 576134
rect 42517 576131 42583 576134
rect 671061 576194 671127 576197
rect 671061 576192 676292 576194
rect 671061 576136 671066 576192
rect 671122 576136 676292 576192
rect 671061 576134 676292 576136
rect 671061 576131 671127 576134
rect 676990 575996 676996 576060
rect 677060 575996 677066 576060
rect 676998 575756 677058 575996
rect 682377 575650 682443 575653
rect 682334 575648 682443 575650
rect 682334 575592 682382 575648
rect 682438 575592 682443 575648
rect 682334 575587 682443 575592
rect 682334 575348 682394 575587
rect 669773 574970 669839 574973
rect 669773 574968 676292 574970
rect 669773 574912 669778 574968
rect 669834 574912 676292 574968
rect 669773 574910 676292 574912
rect 669773 574907 669839 574910
rect 672993 574562 673059 574565
rect 672993 574560 676292 574562
rect 672993 574504 672998 574560
rect 673054 574504 676292 574560
rect 672993 574502 676292 574504
rect 672993 574499 673059 574502
rect 668209 574154 668275 574157
rect 668209 574152 676292 574154
rect 668209 574096 668214 574152
rect 668270 574096 676292 574152
rect 668209 574094 676292 574096
rect 668209 574091 668275 574094
rect 683481 574018 683547 574021
rect 683438 574016 683547 574018
rect 683438 573960 683486 574016
rect 683542 573960 683547 574016
rect 683438 573955 683547 573960
rect 683438 573716 683498 573955
rect 42057 573338 42123 573341
rect 42701 573338 42767 573341
rect 42057 573336 42767 573338
rect 42057 573280 42062 573336
rect 42118 573280 42706 573336
rect 42762 573280 42767 573336
rect 42057 573278 42767 573280
rect 42057 573275 42123 573278
rect 42701 573275 42767 573278
rect 669037 573202 669103 573205
rect 676262 573202 676322 573308
rect 683297 573202 683363 573205
rect 669037 573200 676322 573202
rect 669037 573144 669042 573200
rect 669098 573144 676322 573200
rect 669037 573142 676322 573144
rect 683254 573200 683363 573202
rect 683254 573144 683302 573200
rect 683358 573144 683363 573200
rect 669037 573139 669103 573142
rect 683254 573139 683363 573144
rect 683254 572900 683314 573139
rect 676806 572732 676812 572796
rect 676876 572732 676882 572796
rect 41965 572658 42031 572661
rect 42190 572658 42196 572660
rect 41965 572656 42196 572658
rect 41965 572600 41970 572656
rect 42026 572600 42196 572656
rect 41965 572598 42196 572600
rect 41965 572595 42031 572598
rect 42190 572596 42196 572598
rect 42260 572596 42266 572660
rect 676814 572492 676874 572732
rect 683757 572386 683823 572389
rect 683757 572384 683866 572386
rect 683757 572328 683762 572384
rect 683818 572328 683866 572384
rect 683757 572323 683866 572328
rect 41822 572188 41828 572252
rect 41892 572250 41898 572252
rect 42241 572250 42307 572253
rect 41892 572248 42307 572250
rect 41892 572192 42246 572248
rect 42302 572192 42307 572248
rect 41892 572190 42307 572192
rect 41892 572188 41898 572190
rect 42241 572187 42307 572190
rect 683806 572084 683866 572323
rect 41454 571916 41460 571980
rect 41524 571978 41530 571980
rect 42609 571978 42675 571981
rect 41524 571976 42675 571978
rect 41524 571920 42614 571976
rect 42670 571920 42675 571976
rect 41524 571918 42675 571920
rect 41524 571916 41530 571918
rect 42609 571915 42675 571918
rect 62113 571842 62179 571845
rect 62113 571840 64492 571842
rect 62113 571784 62118 571840
rect 62174 571784 64492 571840
rect 62113 571782 64492 571784
rect 62113 571779 62179 571782
rect 669957 571706 670023 571709
rect 669957 571704 676292 571706
rect 669957 571648 669962 571704
rect 670018 571648 676292 571704
rect 669957 571646 676292 571648
rect 669957 571643 670023 571646
rect 671470 571236 671476 571300
rect 671540 571298 671546 571300
rect 671540 571238 676292 571298
rect 671540 571236 671546 571238
rect 41638 570964 41644 571028
rect 41708 571026 41714 571028
rect 42057 571026 42123 571029
rect 41708 571024 42123 571026
rect 41708 570968 42062 571024
rect 42118 570968 42123 571024
rect 41708 570966 42123 570968
rect 41708 570964 41714 570966
rect 42057 570963 42123 570966
rect 669405 570890 669471 570893
rect 669405 570888 676292 570890
rect 669405 570832 669410 570888
rect 669466 570832 676292 570888
rect 669405 570830 676292 570832
rect 669405 570827 669471 570830
rect 683113 570754 683179 570757
rect 683070 570752 683179 570754
rect 683070 570696 683118 570752
rect 683174 570696 683179 570752
rect 683070 570691 683179 570696
rect 683070 570044 683130 570691
rect 671153 569666 671219 569669
rect 671153 569664 676292 569666
rect 671153 569608 671158 569664
rect 671214 569608 676292 569664
rect 671153 569606 676292 569608
rect 671153 569603 671219 569606
rect 42333 569258 42399 569261
rect 62113 569258 62179 569261
rect 42333 569256 62179 569258
rect 42333 569200 42338 569256
rect 42394 569200 62118 569256
rect 62174 569200 62179 569256
rect 42333 569198 62179 569200
rect 42333 569195 42399 569198
rect 62113 569195 62179 569198
rect 668209 564498 668275 564501
rect 675201 564498 675267 564501
rect 668209 564496 675267 564498
rect 668209 564440 668214 564496
rect 668270 564440 675206 564496
rect 675262 564440 675267 564496
rect 668209 564438 675267 564440
rect 668209 564435 668275 564438
rect 675201 564435 675267 564438
rect 651649 564090 651715 564093
rect 650164 564088 651715 564090
rect 650164 564032 651654 564088
rect 651710 564032 651715 564088
rect 650164 564030 651715 564032
rect 651649 564027 651715 564030
rect 675385 563140 675451 563141
rect 675334 563138 675340 563140
rect 675294 563078 675340 563138
rect 675404 563136 675451 563140
rect 675446 563080 675451 563136
rect 675334 563076 675340 563078
rect 675404 563076 675451 563080
rect 675385 563075 675451 563076
rect 675477 561236 675543 561237
rect 675477 561232 675524 561236
rect 675588 561234 675594 561236
rect 675477 561176 675482 561232
rect 675477 561172 675524 561176
rect 675588 561174 675634 561234
rect 675588 561172 675594 561174
rect 675477 561171 675543 561172
rect 669037 559194 669103 559197
rect 669037 559192 669330 559194
rect 669037 559136 669042 559192
rect 669098 559136 669330 559192
rect 669037 559134 669330 559136
rect 669037 559131 669103 559134
rect 62113 558786 62179 558789
rect 669270 558786 669330 559134
rect 672901 559058 672967 559061
rect 675293 559058 675359 559061
rect 672901 559056 675359 559058
rect 672901 559000 672906 559056
rect 672962 559000 675298 559056
rect 675354 559000 675359 559056
rect 672901 558998 675359 559000
rect 672901 558995 672967 558998
rect 675293 558995 675359 558998
rect 675201 558786 675267 558789
rect 62113 558784 64492 558786
rect 62113 558728 62118 558784
rect 62174 558728 64492 558784
rect 62113 558726 64492 558728
rect 669270 558784 675267 558786
rect 669270 558728 675206 558784
rect 675262 558728 675267 558784
rect 669270 558726 675267 558728
rect 62113 558723 62179 558726
rect 675201 558723 675267 558726
rect 42057 558514 42123 558517
rect 41492 558512 42123 558514
rect 41492 558456 42062 558512
rect 42118 558456 42123 558512
rect 41492 558454 42123 558456
rect 42057 558451 42123 558454
rect 674649 558378 674715 558381
rect 675385 558378 675451 558381
rect 674649 558376 675451 558378
rect 674649 558320 674654 558376
rect 674710 558320 675390 558376
rect 675446 558320 675451 558376
rect 674649 558318 675451 558320
rect 674649 558315 674715 558318
rect 675385 558315 675451 558318
rect 35801 558106 35867 558109
rect 35788 558104 35867 558106
rect 35788 558048 35806 558104
rect 35862 558048 35867 558104
rect 35788 558046 35867 558048
rect 35801 558043 35867 558046
rect 48957 557834 49023 557837
rect 41830 557832 49023 557834
rect 41830 557776 48962 557832
rect 49018 557776 49023 557832
rect 41830 557774 49023 557776
rect 41830 557698 41890 557774
rect 48957 557771 49023 557774
rect 41492 557638 41890 557698
rect 42057 557562 42123 557565
rect 51717 557562 51783 557565
rect 42057 557560 51783 557562
rect 42057 557504 42062 557560
rect 42118 557504 51722 557560
rect 51778 557504 51783 557560
rect 42057 557502 51783 557504
rect 42057 557499 42123 557502
rect 51717 557499 51783 557502
rect 44633 557290 44699 557293
rect 41492 557288 44699 557290
rect 41492 557232 44638 557288
rect 44694 557232 44699 557288
rect 41492 557230 44699 557232
rect 44633 557227 44699 557230
rect 45553 556882 45619 556885
rect 41492 556880 45619 556882
rect 41492 556824 45558 556880
rect 45614 556824 45619 556880
rect 41492 556822 45619 556824
rect 45553 556819 45619 556822
rect 44817 556474 44883 556477
rect 41492 556472 44883 556474
rect 41492 556416 44822 556472
rect 44878 556416 44883 556472
rect 41492 556414 44883 556416
rect 44817 556411 44883 556414
rect 669589 556202 669655 556205
rect 675201 556202 675267 556205
rect 669589 556200 675267 556202
rect 669589 556144 669594 556200
rect 669650 556144 675206 556200
rect 675262 556144 675267 556200
rect 669589 556142 675267 556144
rect 669589 556139 669655 556142
rect 675201 556139 675267 556142
rect 44357 556066 44423 556069
rect 41492 556064 44423 556066
rect 41492 556008 44362 556064
rect 44418 556008 44423 556064
rect 41492 556006 44423 556008
rect 44357 556003 44423 556006
rect 45001 555658 45067 555661
rect 41492 555656 45067 555658
rect 41492 555600 45006 555656
rect 45062 555600 45067 555656
rect 41492 555598 45067 555600
rect 45001 555595 45067 555598
rect 44817 555250 44883 555253
rect 41492 555248 44883 555250
rect 41492 555192 44822 555248
rect 44878 555192 44883 555248
rect 41492 555190 44883 555192
rect 44817 555187 44883 555190
rect 671705 555250 671771 555253
rect 675385 555250 675451 555253
rect 671705 555248 675451 555250
rect 671705 555192 671710 555248
rect 671766 555192 675390 555248
rect 675446 555192 675451 555248
rect 671705 555190 675451 555192
rect 671705 555187 671771 555190
rect 675385 555187 675451 555190
rect 35801 554842 35867 554845
rect 35788 554840 35867 554842
rect 35788 554784 35806 554840
rect 35862 554784 35867 554840
rect 35788 554782 35867 554784
rect 35801 554779 35867 554782
rect 675753 554706 675819 554709
rect 676806 554706 676812 554708
rect 675753 554704 676812 554706
rect 675753 554648 675758 554704
rect 675814 554648 676812 554704
rect 675753 554646 676812 554648
rect 675753 554643 675819 554646
rect 676806 554644 676812 554646
rect 676876 554644 676882 554708
rect 44633 554434 44699 554437
rect 41492 554432 44699 554434
rect 41492 554376 44638 554432
rect 44694 554376 44699 554432
rect 41492 554374 44699 554376
rect 44633 554371 44699 554374
rect 35617 554026 35683 554029
rect 35604 554024 35683 554026
rect 35604 553968 35622 554024
rect 35678 553968 35683 554024
rect 35604 553966 35683 553968
rect 35617 553963 35683 553966
rect 658917 554026 658983 554029
rect 658917 554024 669330 554026
rect 658917 553968 658922 554024
rect 658978 553968 669330 554024
rect 658917 553966 669330 553968
rect 658917 553963 658983 553966
rect 35801 553618 35867 553621
rect 35788 553616 35867 553618
rect 35788 553560 35806 553616
rect 35862 553560 35867 553616
rect 35788 553558 35867 553560
rect 35801 553555 35867 553558
rect 669270 553482 669330 553966
rect 669773 553890 669839 553893
rect 675385 553890 675451 553893
rect 669773 553888 675451 553890
rect 669773 553832 669778 553888
rect 669834 553832 675390 553888
rect 675446 553832 675451 553888
rect 669773 553830 675451 553832
rect 669773 553827 669839 553830
rect 675385 553827 675451 553830
rect 675201 553482 675267 553485
rect 669270 553480 675267 553482
rect 669270 553424 675206 553480
rect 675262 553424 675267 553480
rect 669270 553422 675267 553424
rect 675201 553419 675267 553422
rect 40861 553210 40927 553213
rect 41781 553212 41847 553213
rect 40861 553208 40940 553210
rect 40861 553152 40866 553208
rect 40922 553152 40940 553208
rect 40861 553150 40940 553152
rect 41781 553208 41828 553212
rect 41892 553210 41898 553212
rect 41781 553152 41786 553208
rect 40861 553147 40927 553150
rect 41781 553148 41828 553152
rect 41892 553150 41938 553210
rect 41892 553148 41898 553150
rect 41781 553147 41847 553148
rect 41045 552802 41111 552805
rect 41045 552800 41124 552802
rect 41045 552744 41050 552800
rect 41106 552744 41124 552800
rect 41045 552742 41124 552744
rect 41045 552739 41111 552742
rect 42977 552394 43043 552397
rect 41492 552392 43043 552394
rect 41492 552336 42982 552392
rect 43038 552336 43043 552392
rect 41492 552334 43043 552336
rect 42977 552331 43043 552334
rect 674189 552122 674255 552125
rect 675385 552122 675451 552125
rect 674189 552120 675451 552122
rect 674189 552064 674194 552120
rect 674250 552064 675390 552120
rect 675446 552064 675451 552120
rect 674189 552062 675451 552064
rect 674189 552059 674255 552062
rect 675385 552059 675451 552062
rect 33777 551986 33843 551989
rect 41873 551988 41939 551989
rect 33764 551984 33843 551986
rect 33764 551928 33782 551984
rect 33838 551928 33843 551984
rect 33764 551926 33843 551928
rect 33777 551923 33843 551926
rect 41822 551924 41828 551988
rect 41892 551986 41939 551988
rect 41892 551984 41984 551986
rect 41934 551928 41984 551984
rect 41892 551926 41984 551928
rect 41892 551924 41939 551926
rect 41873 551923 41939 551924
rect 45001 551578 45067 551581
rect 41492 551576 45067 551578
rect 41492 551520 45006 551576
rect 45062 551520 45067 551576
rect 41492 551518 45067 551520
rect 45001 551515 45067 551518
rect 41229 551170 41295 551173
rect 41229 551168 41308 551170
rect 41229 551112 41234 551168
rect 41290 551112 41308 551168
rect 41229 551110 41308 551112
rect 41229 551107 41295 551110
rect 651465 550898 651531 550901
rect 650164 550896 651531 550898
rect 650164 550840 651470 550896
rect 651526 550840 651531 550896
rect 650164 550838 651531 550840
rect 651465 550835 651531 550838
rect 45185 550762 45251 550765
rect 41492 550760 45251 550762
rect 41492 550704 45190 550760
rect 45246 550704 45251 550760
rect 41492 550702 45251 550704
rect 45185 550699 45251 550702
rect 675753 550762 675819 550765
rect 677174 550762 677180 550764
rect 675753 550760 677180 550762
rect 675753 550704 675758 550760
rect 675814 550704 677180 550760
rect 675753 550702 677180 550704
rect 675753 550699 675819 550702
rect 677174 550700 677180 550702
rect 677244 550700 677250 550764
rect 42057 550354 42123 550357
rect 41492 550352 42123 550354
rect 41492 550296 42062 550352
rect 42118 550296 42123 550352
rect 41492 550294 42123 550296
rect 42057 550291 42123 550294
rect 42006 549946 42012 549948
rect 41492 549886 42012 549946
rect 42006 549884 42012 549886
rect 42076 549884 42082 549948
rect 675150 549612 675156 549676
rect 675220 549674 675226 549676
rect 675385 549674 675451 549677
rect 675220 549672 675451 549674
rect 675220 549616 675390 549672
rect 675446 549616 675451 549672
rect 675220 549614 675451 549616
rect 675220 549612 675226 549614
rect 675385 549611 675451 549614
rect 43161 549538 43227 549541
rect 41492 549536 43227 549538
rect 41492 549480 43166 549536
rect 43222 549480 43227 549536
rect 41492 549478 43227 549480
rect 43161 549475 43227 549478
rect 45369 549130 45435 549133
rect 41492 549128 45435 549130
rect 41492 549072 45374 549128
rect 45430 549072 45435 549128
rect 41492 549070 45435 549072
rect 45369 549067 45435 549070
rect 44173 548722 44239 548725
rect 41492 548720 44239 548722
rect 41492 548664 44178 548720
rect 44234 548664 44239 548720
rect 41492 548662 44239 548664
rect 44173 548659 44239 548662
rect 673177 548450 673243 548453
rect 675477 548450 675543 548453
rect 673177 548448 675543 548450
rect 673177 548392 673182 548448
rect 673238 548392 675482 548448
rect 675538 548392 675543 548448
rect 673177 548390 675543 548392
rect 673177 548387 673243 548390
rect 675477 548387 675543 548390
rect 41321 548314 41387 548317
rect 41308 548312 41387 548314
rect 41308 548256 41326 548312
rect 41382 548256 41387 548312
rect 41308 548254 41387 548256
rect 41321 548251 41387 548254
rect 675109 547908 675175 547909
rect 675109 547906 675156 547908
rect 675064 547904 675156 547906
rect 28766 547498 28826 547890
rect 675064 547848 675114 547904
rect 675064 547846 675156 547848
rect 675109 547844 675156 547846
rect 675220 547844 675226 547908
rect 675109 547843 675175 547844
rect 41689 547770 41755 547773
rect 43621 547770 43687 547773
rect 41689 547768 43687 547770
rect 41689 547712 41694 547768
rect 41750 547712 43626 547768
rect 43682 547712 43687 547768
rect 41689 547710 43687 547712
rect 41689 547707 41755 547710
rect 43621 547707 43687 547710
rect 675201 547634 675267 547637
rect 675518 547634 675524 547636
rect 675201 547632 675524 547634
rect 675201 547576 675206 547632
rect 675262 547576 675524 547632
rect 675201 547574 675524 547576
rect 675201 547571 675267 547574
rect 675518 547572 675524 547574
rect 675588 547572 675594 547636
rect 31753 547498 31819 547501
rect 28766 547496 31819 547498
rect 28766 547468 31758 547496
rect 28796 547440 31758 547468
rect 31814 547440 31819 547496
rect 28796 547438 31819 547440
rect 31753 547435 31819 547438
rect 674833 547362 674899 547365
rect 675845 547362 675911 547365
rect 674833 547360 675911 547362
rect 674833 547304 674838 547360
rect 674894 547304 675850 547360
rect 675906 547304 675911 547360
rect 674833 547302 675911 547304
rect 674833 547299 674899 547302
rect 675845 547299 675911 547302
rect 43805 547090 43871 547093
rect 41492 547088 43871 547090
rect 41492 547032 43810 547088
rect 43866 547032 43871 547088
rect 41492 547030 43871 547032
rect 43805 547027 43871 547030
rect 674373 547090 674439 547093
rect 683205 547090 683271 547093
rect 674373 547088 683271 547090
rect 674373 547032 674378 547088
rect 674434 547032 683210 547088
rect 683266 547032 683271 547088
rect 674373 547030 683271 547032
rect 674373 547027 674439 547030
rect 683205 547027 683271 547030
rect 676070 546484 676076 546548
rect 676140 546546 676146 546548
rect 679617 546546 679683 546549
rect 676140 546544 679683 546546
rect 676140 546488 679622 546544
rect 679678 546488 679683 546544
rect 676140 546486 679683 546488
rect 676140 546484 676146 546486
rect 679617 546483 679683 546486
rect 41321 546410 41387 546413
rect 41638 546410 41644 546412
rect 41321 546408 41644 546410
rect 41321 546352 41326 546408
rect 41382 546352 41644 546408
rect 41321 546350 41644 546352
rect 41321 546347 41387 546350
rect 41638 546348 41644 546350
rect 41708 546348 41714 546412
rect 672625 546274 672691 546277
rect 676397 546274 676463 546277
rect 672625 546272 676463 546274
rect 672625 546216 672630 546272
rect 672686 546216 676402 546272
rect 676458 546216 676463 546272
rect 672625 546214 676463 546216
rect 672625 546211 672691 546214
rect 676397 546211 676463 546214
rect 62113 545866 62179 545869
rect 62113 545864 64492 545866
rect 62113 545808 62118 545864
rect 62174 545808 64492 545864
rect 62113 545806 64492 545808
rect 62113 545803 62179 545806
rect 40534 545668 40540 545732
rect 40604 545730 40610 545732
rect 42057 545730 42123 545733
rect 40604 545728 42123 545730
rect 40604 545672 42062 545728
rect 42118 545672 42123 545728
rect 40604 545670 42123 545672
rect 40604 545668 40610 545670
rect 42057 545667 42123 545670
rect 674005 545730 674071 545733
rect 683389 545730 683455 545733
rect 674005 545728 683455 545730
rect 674005 545672 674010 545728
rect 674066 545672 683394 545728
rect 683450 545672 683455 545728
rect 674005 545670 683455 545672
rect 674005 545667 674071 545670
rect 683389 545667 683455 545670
rect 40718 545396 40724 545460
rect 40788 545458 40794 545460
rect 42006 545458 42012 545460
rect 40788 545398 42012 545458
rect 40788 545396 40794 545398
rect 42006 545396 42012 545398
rect 42076 545396 42082 545460
rect 674833 543828 674899 543829
rect 674782 543764 674788 543828
rect 674852 543826 674899 543828
rect 674852 543824 674944 543826
rect 674894 543768 674944 543824
rect 674852 543766 674944 543768
rect 674852 543764 674899 543766
rect 674833 543763 674899 543764
rect 41781 541106 41847 541109
rect 41781 541104 41890 541106
rect 41781 541048 41786 541104
rect 41842 541048 41890 541104
rect 41781 541043 41890 541048
rect 41830 540701 41890 541043
rect 41781 540696 41890 540701
rect 41781 540640 41786 540696
rect 41842 540640 41890 540696
rect 41781 540638 41890 540640
rect 41781 540635 41847 540638
rect 42609 540290 42675 540293
rect 56041 540290 56107 540293
rect 42609 540288 56107 540290
rect 42609 540232 42614 540288
rect 42670 540232 56046 540288
rect 56102 540232 56107 540288
rect 42609 540230 56107 540232
rect 42609 540227 42675 540230
rect 56041 540227 56107 540230
rect 40718 538596 40724 538660
rect 40788 538658 40794 538660
rect 42333 538658 42399 538661
rect 40788 538656 42399 538658
rect 40788 538600 42338 538656
rect 42394 538600 42399 538656
rect 40788 538598 42399 538600
rect 40788 538596 40794 538598
rect 42333 538595 42399 538598
rect 40534 538188 40540 538252
rect 40604 538250 40610 538252
rect 42241 538250 42307 538253
rect 40604 538248 42307 538250
rect 40604 538192 42246 538248
rect 42302 538192 42307 538248
rect 40604 538190 42307 538192
rect 40604 538188 40610 538190
rect 42241 538187 42307 538190
rect 42057 537978 42123 537981
rect 42609 537978 42675 537981
rect 42057 537976 42675 537978
rect 42057 537920 42062 537976
rect 42118 537920 42614 537976
rect 42670 537920 42675 537976
rect 42057 537918 42675 537920
rect 42057 537915 42123 537918
rect 42609 537915 42675 537918
rect 670141 537842 670207 537845
rect 676029 537842 676095 537845
rect 670141 537840 676095 537842
rect 670141 537784 670146 537840
rect 670202 537784 676034 537840
rect 676090 537784 676095 537840
rect 670141 537782 676095 537784
rect 670141 537779 670207 537782
rect 676029 537779 676095 537782
rect 651465 537570 651531 537573
rect 650164 537568 651531 537570
rect 650164 537512 651470 537568
rect 651526 537512 651531 537568
rect 650164 537510 651531 537512
rect 651465 537507 651531 537510
rect 42609 537162 42675 537165
rect 45369 537162 45435 537165
rect 42609 537160 45435 537162
rect 42609 537104 42614 537160
rect 42670 537104 45374 537160
rect 45430 537104 45435 537160
rect 42609 537102 45435 537104
rect 42609 537099 42675 537102
rect 45369 537099 45435 537102
rect 44173 536890 44239 536893
rect 42198 536888 44239 536890
rect 42198 536832 44178 536888
rect 44234 536832 44239 536888
rect 42198 536830 44239 536832
rect 42198 536349 42258 536830
rect 44173 536827 44239 536830
rect 42198 536344 42307 536349
rect 42198 536288 42246 536344
rect 42302 536288 42307 536344
rect 42198 536286 42307 536288
rect 42241 536283 42307 536286
rect 668577 535938 668643 535941
rect 676262 535938 676322 536112
rect 668577 535936 676322 535938
rect 668577 535880 668582 535936
rect 668638 535880 676322 535936
rect 668577 535878 676322 535880
rect 668577 535875 668643 535878
rect 676029 535734 676095 535737
rect 676029 535732 676292 535734
rect 676029 535676 676034 535732
rect 676090 535676 676292 535732
rect 676029 535674 676292 535676
rect 676029 535671 676095 535674
rect 674005 535394 674071 535397
rect 674005 535392 676322 535394
rect 674005 535336 674010 535392
rect 674066 535336 676322 535392
rect 674005 535334 676322 535336
rect 674005 535331 674071 535334
rect 676262 535296 676322 535334
rect 670785 535122 670851 535125
rect 674465 535122 674531 535125
rect 670785 535120 674531 535122
rect 670785 535064 670790 535120
rect 670846 535064 674470 535120
rect 674526 535064 674531 535120
rect 670785 535062 674531 535064
rect 670785 535059 670851 535062
rect 674465 535059 674531 535062
rect 671429 534714 671495 534717
rect 676262 534714 676322 534888
rect 671429 534712 676322 534714
rect 671429 534656 671434 534712
rect 671490 534656 676322 534712
rect 671429 534654 676322 534656
rect 671429 534651 671495 534654
rect 671429 534442 671495 534445
rect 676262 534442 676322 534480
rect 671429 534440 676322 534442
rect 671429 534384 671434 534440
rect 671490 534384 676322 534440
rect 671429 534382 676322 534384
rect 671429 534379 671495 534382
rect 667197 534170 667263 534173
rect 674005 534170 674071 534173
rect 667197 534168 674071 534170
rect 667197 534112 667202 534168
rect 667258 534112 674010 534168
rect 674066 534112 674071 534168
rect 667197 534110 674071 534112
rect 667197 534107 667263 534110
rect 674005 534107 674071 534110
rect 674465 534170 674531 534173
rect 674465 534168 676322 534170
rect 674465 534112 674470 534168
rect 674526 534112 676322 534168
rect 674465 534110 676322 534112
rect 674465 534107 674531 534110
rect 676262 534072 676322 534110
rect 42149 533898 42215 533901
rect 42977 533898 43043 533901
rect 42149 533896 43043 533898
rect 42149 533840 42154 533896
rect 42210 533840 42982 533896
rect 43038 533840 43043 533896
rect 42149 533838 43043 533840
rect 42149 533835 42215 533838
rect 42977 533835 43043 533838
rect 672533 533490 672599 533493
rect 676262 533490 676322 533664
rect 672533 533488 676322 533490
rect 672533 533432 672538 533488
rect 672594 533432 676322 533488
rect 672533 533430 676322 533432
rect 672533 533427 672599 533430
rect 42241 533218 42307 533221
rect 43161 533218 43227 533221
rect 42241 533216 43227 533218
rect 42241 533160 42246 533216
rect 42302 533160 43166 533216
rect 43222 533160 43227 533216
rect 42241 533158 43227 533160
rect 42241 533155 42307 533158
rect 43161 533155 43227 533158
rect 670877 533082 670943 533085
rect 676262 533082 676322 533256
rect 670877 533080 676322 533082
rect 670877 533024 670882 533080
rect 670938 533024 676322 533080
rect 670877 533022 676322 533024
rect 670877 533019 670943 533022
rect 42517 532810 42583 532813
rect 45185 532810 45251 532813
rect 42517 532808 45251 532810
rect 42517 532752 42522 532808
rect 42578 532752 45190 532808
rect 45246 532752 45251 532808
rect 42517 532750 45251 532752
rect 42517 532747 42583 532750
rect 45185 532747 45251 532750
rect 62113 532810 62179 532813
rect 671521 532810 671587 532813
rect 676262 532810 676322 532848
rect 62113 532808 64492 532810
rect 62113 532752 62118 532808
rect 62174 532752 64492 532808
rect 62113 532750 64492 532752
rect 671521 532808 676322 532810
rect 671521 532752 671526 532808
rect 671582 532752 676322 532808
rect 671521 532750 676322 532752
rect 62113 532747 62179 532750
rect 671521 532747 671587 532750
rect 673821 532538 673887 532541
rect 675845 532538 675911 532541
rect 673821 532536 675911 532538
rect 673821 532480 673826 532536
rect 673882 532480 675850 532536
rect 675906 532480 675911 532536
rect 673821 532478 675911 532480
rect 673821 532475 673887 532478
rect 675845 532475 675911 532478
rect 674465 532266 674531 532269
rect 676262 532266 676322 532440
rect 674465 532264 676322 532266
rect 674465 532208 674470 532264
rect 674526 532208 676322 532264
rect 674465 532206 676322 532208
rect 676581 532266 676647 532269
rect 683573 532266 683639 532269
rect 676581 532264 683639 532266
rect 676581 532208 676586 532264
rect 676642 532208 683578 532264
rect 683634 532208 683639 532264
rect 676581 532206 683639 532208
rect 674465 532203 674531 532206
rect 676581 532203 676647 532206
rect 683573 532203 683639 532206
rect 672717 531858 672783 531861
rect 676262 531858 676322 532032
rect 672717 531856 676322 531858
rect 672717 531800 672722 531856
rect 672778 531800 676322 531856
rect 672717 531798 676322 531800
rect 683205 531858 683271 531861
rect 683205 531856 683314 531858
rect 683205 531800 683210 531856
rect 683266 531800 683314 531856
rect 672717 531795 672783 531798
rect 683205 531795 683314 531800
rect 683254 531624 683314 531795
rect 672257 531450 672323 531453
rect 674465 531450 674531 531453
rect 672257 531448 674531 531450
rect 672257 531392 672262 531448
rect 672318 531392 674470 531448
rect 674526 531392 674531 531448
rect 672257 531390 674531 531392
rect 672257 531387 672323 531390
rect 674465 531387 674531 531390
rect 678237 531450 678303 531453
rect 678237 531448 678346 531450
rect 678237 531392 678242 531448
rect 678298 531392 678346 531448
rect 678237 531387 678346 531392
rect 678286 531216 678346 531387
rect 679617 531042 679683 531045
rect 679574 531040 679683 531042
rect 679574 530984 679622 531040
rect 679678 530984 679683 531040
rect 679574 530979 679683 530984
rect 679574 530808 679634 530979
rect 41454 530572 41460 530636
rect 41524 530634 41530 530636
rect 42517 530634 42583 530637
rect 41524 530632 42583 530634
rect 41524 530576 42522 530632
rect 42578 530576 42583 530632
rect 41524 530574 42583 530576
rect 41524 530572 41530 530574
rect 42517 530571 42583 530574
rect 672165 530226 672231 530229
rect 676262 530226 676322 530400
rect 672165 530224 676322 530226
rect 672165 530168 672170 530224
rect 672226 530168 676322 530224
rect 672165 530166 676322 530168
rect 672165 530163 672231 530166
rect 42149 530090 42215 530093
rect 42701 530090 42767 530093
rect 42149 530088 42767 530090
rect 42149 530032 42154 530088
rect 42210 530032 42706 530088
rect 42762 530032 42767 530088
rect 42149 530030 42767 530032
rect 42149 530027 42215 530030
rect 42701 530027 42767 530030
rect 666461 529954 666527 529957
rect 676262 529954 676322 529992
rect 666461 529952 676322 529954
rect 666461 529896 666466 529952
rect 666522 529896 676322 529952
rect 666461 529894 676322 529896
rect 666461 529891 666527 529894
rect 42609 529682 42675 529685
rect 45001 529682 45067 529685
rect 42609 529680 45067 529682
rect 42609 529624 42614 529680
rect 42670 529624 45006 529680
rect 45062 529624 45067 529680
rect 42609 529622 45067 529624
rect 42609 529619 42675 529622
rect 45001 529619 45067 529622
rect 41873 529412 41939 529413
rect 41822 529410 41828 529412
rect 41782 529350 41828 529410
rect 41892 529408 41939 529412
rect 41934 529352 41939 529408
rect 41822 529348 41828 529350
rect 41892 529348 41939 529352
rect 41873 529347 41939 529348
rect 672349 529410 672415 529413
rect 675753 529410 675819 529413
rect 672349 529408 675819 529410
rect 672349 529352 672354 529408
rect 672410 529352 675758 529408
rect 675814 529352 675819 529408
rect 672349 529350 675819 529352
rect 672349 529347 672415 529350
rect 675753 529347 675819 529350
rect 675937 529410 676003 529413
rect 676262 529410 676322 529584
rect 675937 529408 676322 529410
rect 675937 529352 675942 529408
rect 675998 529352 676322 529408
rect 675937 529350 676322 529352
rect 675937 529347 676003 529350
rect 41638 529076 41644 529140
rect 41708 529138 41714 529140
rect 42885 529138 42951 529141
rect 41708 529136 42951 529138
rect 41708 529080 42890 529136
rect 42946 529080 42951 529136
rect 41708 529078 42951 529080
rect 41708 529076 41714 529078
rect 42885 529075 42951 529078
rect 670601 529002 670667 529005
rect 676262 529002 676322 529176
rect 670601 529000 676322 529002
rect 670601 528944 670606 529000
rect 670662 528944 676322 529000
rect 670601 528942 676322 528944
rect 670601 528939 670667 528942
rect 675753 528798 675819 528801
rect 675753 528796 676292 528798
rect 675753 528740 675758 528796
rect 675814 528740 676292 528796
rect 675753 528738 676292 528740
rect 675753 528735 675819 528738
rect 668853 528594 668919 528597
rect 675937 528594 676003 528597
rect 668853 528592 676003 528594
rect 668853 528536 668858 528592
rect 668914 528536 675942 528592
rect 675998 528536 676003 528592
rect 668853 528534 676003 528536
rect 668853 528531 668919 528534
rect 675937 528531 676003 528534
rect 673637 528322 673703 528325
rect 676262 528322 676322 528360
rect 673637 528320 676322 528322
rect 673637 528264 673642 528320
rect 673698 528264 676322 528320
rect 673637 528262 676322 528264
rect 673637 528259 673703 528262
rect 670325 527778 670391 527781
rect 676262 527778 676322 527952
rect 670325 527776 676322 527778
rect 670325 527720 670330 527776
rect 670386 527720 676322 527776
rect 670325 527718 676322 527720
rect 683389 527778 683455 527781
rect 683389 527776 683498 527778
rect 683389 527720 683394 527776
rect 683450 527720 683498 527776
rect 670325 527715 670391 527718
rect 683389 527715 683498 527720
rect 683438 527544 683498 527715
rect 674414 527036 674420 527100
rect 674484 527098 674490 527100
rect 676262 527098 676322 527136
rect 674484 527038 676322 527098
rect 674484 527036 674490 527038
rect 668393 526554 668459 526557
rect 676262 526554 676322 526728
rect 668393 526552 676322 526554
rect 668393 526496 668398 526552
rect 668454 526496 676322 526552
rect 668393 526494 676322 526496
rect 683573 526554 683639 526557
rect 683573 526552 683682 526554
rect 683573 526496 683578 526552
rect 683634 526496 683682 526552
rect 668393 526491 668459 526494
rect 683573 526491 683682 526496
rect 683622 526320 683682 526491
rect 676814 525741 676874 525912
rect 676814 525736 676923 525741
rect 676814 525680 676862 525736
rect 676918 525680 676923 525736
rect 676814 525678 676923 525680
rect 676857 525675 676923 525678
rect 670877 524922 670943 524925
rect 676262 524922 676322 525504
rect 670877 524920 676322 524922
rect 670877 524864 670882 524920
rect 670938 524864 676322 524920
rect 670877 524862 676322 524864
rect 670877 524859 670943 524862
rect 677918 524517 677978 524688
rect 677869 524512 677978 524517
rect 677869 524456 677874 524512
rect 677930 524456 677978 524512
rect 677869 524454 677978 524456
rect 677869 524451 677935 524454
rect 651833 524242 651899 524245
rect 650164 524240 651899 524242
rect 650164 524184 651838 524240
rect 651894 524184 651899 524240
rect 650164 524182 651899 524184
rect 651833 524179 651899 524182
rect 62113 519754 62179 519757
rect 62113 519752 64492 519754
rect 62113 519696 62118 519752
rect 62174 519696 64492 519752
rect 62113 519694 64492 519696
rect 62113 519691 62179 519694
rect 651465 511050 651531 511053
rect 650164 511048 651531 511050
rect 650164 510992 651470 511048
rect 651526 510992 651531 511048
rect 650164 510990 651531 510992
rect 651465 510987 651531 510990
rect 62113 506698 62179 506701
rect 62113 506696 64492 506698
rect 62113 506640 62118 506696
rect 62174 506640 64492 506696
rect 62113 506638 64492 506640
rect 62113 506635 62179 506638
rect 674925 503842 674991 503845
rect 675845 503842 675911 503845
rect 674925 503840 675911 503842
rect 674925 503784 674930 503840
rect 674986 503784 675850 503840
rect 675906 503784 675911 503840
rect 674925 503782 675911 503784
rect 674925 503779 674991 503782
rect 675845 503779 675911 503782
rect 676806 503644 676812 503708
rect 676876 503706 676882 503708
rect 683205 503706 683271 503709
rect 676876 503704 683271 503706
rect 676876 503648 683210 503704
rect 683266 503648 683271 503704
rect 676876 503646 683271 503648
rect 676876 503644 676882 503646
rect 683205 503643 683271 503646
rect 675017 503570 675083 503573
rect 676029 503570 676095 503573
rect 675017 503568 676095 503570
rect 675017 503512 675022 503568
rect 675078 503512 676034 503568
rect 676090 503512 676095 503568
rect 675017 503510 676095 503512
rect 675017 503507 675083 503510
rect 676029 503507 676095 503510
rect 675017 503298 675083 503301
rect 676029 503298 676095 503301
rect 675017 503296 676095 503298
rect 675017 503240 675022 503296
rect 675078 503240 676034 503296
rect 676090 503240 676095 503296
rect 675017 503238 676095 503240
rect 675017 503235 675083 503238
rect 676029 503235 676095 503238
rect 669405 500986 669471 500989
rect 674925 500986 674991 500989
rect 669405 500984 674991 500986
rect 669405 500928 669410 500984
rect 669466 500928 674930 500984
rect 674986 500928 674991 500984
rect 669405 500926 674991 500928
rect 669405 500923 669471 500926
rect 674925 500923 674991 500926
rect 651465 497722 651531 497725
rect 650164 497720 651531 497722
rect 650164 497664 651470 497720
rect 651526 497664 651531 497720
rect 650164 497662 651531 497664
rect 651465 497659 651531 497662
rect 665817 494730 665883 494733
rect 683573 494730 683639 494733
rect 665817 494728 683639 494730
rect 665817 494672 665822 494728
rect 665878 494672 683578 494728
rect 683634 494672 683639 494728
rect 665817 494670 683639 494672
rect 665817 494667 665883 494670
rect 683573 494667 683639 494670
rect 664621 494050 664687 494053
rect 676029 494050 676095 494053
rect 664621 494048 676095 494050
rect 664621 493992 664626 494048
rect 664682 493992 676034 494048
rect 676090 493992 676095 494048
rect 664621 493990 676095 493992
rect 664621 493987 664687 493990
rect 676029 493987 676095 493990
rect 62113 493642 62179 493645
rect 62113 493640 64492 493642
rect 62113 493584 62118 493640
rect 62174 493584 64492 493640
rect 62113 493582 64492 493584
rect 62113 493579 62179 493582
rect 677317 492420 677383 492421
rect 677317 492416 677364 492420
rect 677428 492418 677434 492420
rect 677317 492360 677322 492416
rect 677317 492356 677364 492360
rect 677428 492358 677474 492418
rect 677428 492356 677434 492358
rect 677317 492355 677383 492356
rect 663750 492086 676292 492146
rect 662045 492010 662111 492013
rect 663750 492010 663810 492086
rect 662045 492008 663810 492010
rect 662045 491952 662050 492008
rect 662106 491952 663810 492008
rect 662045 491950 663810 491952
rect 662045 491947 662111 491950
rect 683389 491738 683455 491741
rect 683389 491736 683468 491738
rect 683389 491680 683394 491736
rect 683450 491680 683468 491736
rect 683389 491678 683468 491680
rect 683389 491675 683455 491678
rect 683573 491330 683639 491333
rect 683573 491328 683652 491330
rect 683573 491272 683578 491328
rect 683634 491272 683652 491328
rect 683573 491270 683652 491272
rect 683573 491267 683639 491270
rect 671337 490922 671403 490925
rect 671337 490920 676292 490922
rect 671337 490864 671342 490920
rect 671398 490864 676292 490920
rect 671337 490862 676292 490864
rect 671337 490859 671403 490862
rect 675886 490452 675892 490516
rect 675956 490514 675962 490516
rect 675956 490454 676292 490514
rect 675956 490452 675962 490454
rect 672717 490106 672783 490109
rect 672717 490104 676292 490106
rect 672717 490048 672722 490104
rect 672778 490048 676292 490104
rect 672717 490046 676292 490048
rect 672717 490043 672783 490046
rect 672441 489698 672507 489701
rect 672441 489696 676292 489698
rect 672441 489640 672446 489696
rect 672502 489640 676292 489696
rect 672441 489638 676292 489640
rect 672441 489635 672507 489638
rect 671521 489290 671587 489293
rect 671521 489288 676292 489290
rect 671521 489232 671526 489288
rect 671582 489232 676292 489288
rect 671521 489230 676292 489232
rect 671521 489227 671587 489230
rect 676949 488882 677015 488885
rect 676949 488880 677028 488882
rect 676949 488824 676954 488880
rect 677010 488824 677028 488880
rect 676949 488822 677028 488824
rect 676949 488819 677015 488822
rect 672901 488474 672967 488477
rect 672901 488472 676292 488474
rect 672901 488416 672906 488472
rect 672962 488416 676292 488472
rect 672901 488414 676292 488416
rect 672901 488411 672967 488414
rect 672625 488066 672691 488069
rect 672625 488064 676292 488066
rect 672625 488008 672630 488064
rect 672686 488008 676292 488064
rect 672625 488006 676292 488008
rect 672625 488003 672691 488006
rect 680997 487658 681063 487661
rect 680997 487656 681076 487658
rect 680997 487600 681002 487656
rect 681058 487600 681076 487656
rect 680997 487598 681076 487600
rect 680997 487595 681063 487598
rect 677317 487250 677383 487253
rect 677317 487248 677396 487250
rect 677317 487192 677322 487248
rect 677378 487192 677396 487248
rect 677317 487190 677396 487192
rect 677317 487187 677383 487190
rect 679617 486842 679683 486845
rect 679604 486840 679683 486842
rect 679604 486784 679622 486840
rect 679678 486784 679683 486840
rect 679604 486782 679683 486784
rect 679617 486779 679683 486782
rect 675293 486434 675359 486437
rect 675293 486432 676292 486434
rect 675293 486376 675298 486432
rect 675354 486376 676292 486432
rect 675293 486374 676292 486376
rect 675293 486371 675359 486374
rect 671705 486026 671771 486029
rect 671705 486024 676292 486026
rect 671705 485968 671710 486024
rect 671766 485968 676292 486024
rect 671705 485966 676292 485968
rect 671705 485963 671771 485966
rect 676949 485792 677015 485793
rect 676949 485788 676996 485792
rect 677060 485790 677066 485792
rect 676949 485732 676954 485788
rect 676949 485728 676996 485732
rect 677060 485730 677106 485790
rect 677060 485728 677066 485730
rect 676949 485727 677015 485728
rect 673177 485618 673243 485621
rect 673177 485616 676292 485618
rect 673177 485560 673182 485616
rect 673238 485560 676292 485616
rect 673177 485558 676292 485560
rect 673177 485555 673243 485558
rect 668209 485210 668275 485213
rect 668209 485208 676292 485210
rect 668209 485152 668214 485208
rect 668270 485152 676292 485208
rect 668209 485150 676292 485152
rect 668209 485147 668275 485150
rect 672993 484802 673059 484805
rect 672993 484800 676292 484802
rect 672993 484744 672998 484800
rect 673054 484744 676292 484800
rect 672993 484742 676292 484744
rect 672993 484739 673059 484742
rect 651465 484530 651531 484533
rect 650164 484528 651531 484530
rect 650164 484472 651470 484528
rect 651526 484472 651531 484528
rect 650164 484470 651531 484472
rect 651465 484467 651531 484470
rect 674649 484394 674715 484397
rect 674649 484392 676292 484394
rect 674649 484336 674654 484392
rect 674710 484336 676292 484392
rect 674649 484334 676292 484336
rect 674649 484331 674715 484334
rect 674189 483986 674255 483989
rect 674189 483984 676292 483986
rect 674189 483928 674194 483984
rect 674250 483928 676292 483984
rect 674189 483926 676292 483928
rect 674189 483923 674255 483926
rect 669773 483578 669839 483581
rect 669773 483576 676292 483578
rect 669773 483520 669778 483576
rect 669834 483520 676292 483576
rect 669773 483518 676292 483520
rect 669773 483515 669839 483518
rect 669037 483170 669103 483173
rect 669037 483168 676292 483170
rect 669037 483112 669042 483168
rect 669098 483112 676292 483168
rect 669037 483110 676292 483112
rect 669037 483107 669103 483110
rect 683205 482762 683271 482765
rect 683205 482760 683284 482762
rect 683205 482704 683210 482760
rect 683266 482704 683284 482760
rect 683205 482702 683284 482704
rect 683205 482699 683271 482702
rect 669589 482354 669655 482357
rect 669589 482352 676292 482354
rect 669589 482296 669594 482352
rect 669650 482296 676292 482352
rect 669589 482294 676292 482296
rect 669589 482291 669655 482294
rect 675845 481946 675911 481949
rect 675845 481944 676292 481946
rect 675845 481888 675850 481944
rect 675906 481888 676292 481944
rect 675845 481886 676292 481888
rect 675845 481883 675911 481886
rect 682377 481538 682443 481541
rect 682364 481536 682443 481538
rect 682364 481508 682382 481536
rect 682334 481480 682382 481508
rect 682438 481480 682443 481536
rect 682334 481475 682443 481480
rect 682334 481100 682394 481475
rect 676029 480722 676095 480725
rect 676029 480720 676292 480722
rect 676029 480664 676034 480720
rect 676090 480664 676292 480720
rect 676029 480662 676292 480664
rect 676029 480659 676095 480662
rect 62113 480586 62179 480589
rect 62113 480584 64492 480586
rect 62113 480528 62118 480584
rect 62174 480528 64492 480584
rect 62113 480526 64492 480528
rect 62113 480523 62179 480526
rect 673678 475356 673684 475420
rect 673748 475418 673754 475420
rect 674046 475418 674052 475420
rect 673748 475358 674052 475418
rect 673748 475356 673754 475358
rect 674046 475356 674052 475358
rect 674116 475356 674122 475420
rect 651465 471202 651531 471205
rect 650164 471200 651531 471202
rect 650164 471144 651470 471200
rect 651526 471144 651531 471200
rect 650164 471142 651531 471144
rect 651465 471139 651531 471142
rect 62113 467530 62179 467533
rect 62113 467528 64492 467530
rect 62113 467472 62118 467528
rect 62174 467472 64492 467528
rect 62113 467470 64492 467472
rect 62113 467467 62179 467470
rect 673678 464748 673684 464812
rect 673748 464810 673754 464812
rect 674741 464810 674807 464813
rect 673748 464808 674807 464810
rect 673748 464752 674746 464808
rect 674802 464752 674807 464808
rect 673748 464750 674807 464752
rect 673748 464748 673754 464750
rect 674741 464747 674807 464750
rect 652385 457874 652451 457877
rect 650164 457872 652451 457874
rect 650164 457816 652390 457872
rect 652446 457816 652451 457872
rect 650164 457814 652451 457816
rect 652385 457811 652451 457814
rect 673821 456922 673887 456925
rect 674741 456922 674807 456925
rect 673821 456920 674807 456922
rect 673821 456864 673826 456920
rect 673882 456864 674746 456920
rect 674802 456864 674807 456920
rect 673821 456862 674807 456864
rect 673821 456859 673887 456862
rect 674741 456859 674807 456862
rect 669221 456514 669287 456517
rect 673941 456514 674007 456517
rect 669221 456512 674007 456514
rect 669221 456456 669226 456512
rect 669282 456456 673946 456512
rect 674002 456456 674007 456512
rect 669221 456454 674007 456456
rect 669221 456451 669287 456454
rect 673941 456451 674007 456454
rect 673591 455698 673657 455701
rect 676765 455698 676831 455701
rect 673591 455696 676831 455698
rect 673591 455640 673596 455696
rect 673652 455640 676770 455696
rect 676826 455640 676831 455696
rect 673591 455638 676831 455640
rect 673591 455635 673657 455638
rect 676765 455635 676831 455638
rect 671981 455426 672047 455429
rect 673499 455426 673565 455429
rect 671981 455424 673565 455426
rect 671981 455368 671986 455424
rect 672042 455368 673504 455424
rect 673560 455368 673565 455424
rect 671981 455366 673565 455368
rect 671981 455363 672047 455366
rect 673499 455363 673565 455366
rect 673381 455154 673447 455157
rect 673862 455154 673868 455156
rect 673381 455152 673868 455154
rect 673381 455096 673386 455152
rect 673442 455096 673868 455152
rect 673381 455094 673868 455096
rect 673381 455091 673447 455094
rect 673862 455092 673868 455094
rect 673932 455092 673938 455156
rect 673157 454882 673223 454885
rect 674925 454882 674991 454885
rect 673157 454880 674991 454882
rect 673157 454824 673162 454880
rect 673218 454824 674930 454880
rect 674986 454824 674991 454880
rect 673157 454822 674991 454824
rect 673157 454819 673223 454822
rect 674925 454819 674991 454822
rect 62113 454610 62179 454613
rect 673039 454610 673105 454613
rect 675477 454610 675543 454613
rect 62113 454608 64492 454610
rect 62113 454552 62118 454608
rect 62174 454552 64492 454608
rect 62113 454550 64492 454552
rect 673039 454608 675543 454610
rect 673039 454552 673044 454608
rect 673100 454552 675482 454608
rect 675538 454552 675543 454608
rect 673039 454550 675543 454552
rect 62113 454547 62179 454550
rect 673039 454547 673105 454550
rect 675477 454547 675543 454550
rect 672947 454338 673013 454341
rect 675661 454338 675727 454341
rect 672947 454336 675727 454338
rect 672947 454280 672952 454336
rect 673008 454280 675666 454336
rect 675722 454280 675727 454336
rect 672947 454278 675727 454280
rect 672947 454275 673013 454278
rect 675661 454275 675727 454278
rect 672809 454066 672875 454069
rect 676029 454066 676095 454069
rect 672809 454064 676095 454066
rect 672809 454008 672814 454064
rect 672870 454008 676034 454064
rect 676090 454008 676095 454064
rect 672809 454006 676095 454008
rect 672809 454003 672875 454006
rect 676029 454003 676095 454006
rect 672257 453794 672323 453797
rect 675845 453794 675911 453797
rect 672257 453792 675911 453794
rect 672257 453736 672262 453792
rect 672318 453736 675850 453792
rect 675906 453736 675911 453792
rect 672257 453734 675911 453736
rect 672257 453731 672323 453734
rect 675845 453731 675911 453734
rect 651465 444546 651531 444549
rect 650164 444544 651531 444546
rect 650164 444488 651470 444544
rect 651526 444488 651531 444544
rect 650164 444486 651531 444488
rect 651465 444483 651531 444486
rect 62113 441554 62179 441557
rect 62113 441552 64492 441554
rect 62113 441496 62118 441552
rect 62174 441496 64492 441552
rect 62113 441494 64492 441496
rect 62113 441491 62179 441494
rect 651465 431354 651531 431357
rect 650164 431352 651531 431354
rect 650164 431296 651470 431352
rect 651526 431296 651531 431352
rect 650164 431294 651531 431296
rect 651465 431291 651531 431294
rect 50337 430946 50403 430949
rect 41492 430944 50403 430946
rect 41492 430888 50342 430944
rect 50398 430888 50403 430944
rect 41492 430886 50403 430888
rect 50337 430883 50403 430886
rect 54477 430538 54543 430541
rect 41492 430536 54543 430538
rect 41492 430480 54482 430536
rect 54538 430480 54543 430536
rect 41492 430478 54543 430480
rect 54477 430475 54543 430478
rect 47577 430130 47643 430133
rect 41492 430128 47643 430130
rect 41492 430072 47582 430128
rect 47638 430072 47643 430128
rect 41492 430070 47643 430072
rect 47577 430067 47643 430070
rect 45553 429722 45619 429725
rect 41492 429720 45619 429722
rect 41492 429664 45558 429720
rect 45614 429664 45619 429720
rect 41492 429662 45619 429664
rect 45553 429659 45619 429662
rect 45001 429314 45067 429317
rect 41492 429312 45067 429314
rect 41492 429256 45006 429312
rect 45062 429256 45067 429312
rect 41492 429254 45067 429256
rect 45001 429251 45067 429254
rect 44357 428906 44423 428909
rect 41492 428904 44423 428906
rect 41492 428848 44362 428904
rect 44418 428848 44423 428904
rect 41492 428846 44423 428848
rect 44357 428843 44423 428846
rect 44173 428498 44239 428501
rect 41492 428496 44239 428498
rect 41492 428440 44178 428496
rect 44234 428440 44239 428496
rect 41492 428438 44239 428440
rect 44173 428435 44239 428438
rect 62113 428498 62179 428501
rect 62113 428496 64492 428498
rect 62113 428440 62118 428496
rect 62174 428440 64492 428496
rect 62113 428438 64492 428440
rect 62113 428435 62179 428438
rect 44817 428090 44883 428093
rect 41492 428088 44883 428090
rect 41492 428032 44822 428088
rect 44878 428032 44883 428088
rect 41492 428030 44883 428032
rect 44817 428027 44883 428030
rect 44449 427682 44515 427685
rect 41492 427680 44515 427682
rect 41492 427624 44454 427680
rect 44510 427624 44515 427680
rect 41492 427622 44515 427624
rect 44449 427619 44515 427622
rect 44633 427274 44699 427277
rect 41492 427272 44699 427274
rect 41492 427216 44638 427272
rect 44694 427216 44699 427272
rect 41492 427214 44699 427216
rect 44633 427211 44699 427214
rect 45185 426866 45251 426869
rect 41492 426864 45251 426866
rect 41492 426808 45190 426864
rect 45246 426808 45251 426864
rect 41492 426806 45251 426808
rect 45185 426803 45251 426806
rect 45553 426458 45619 426461
rect 41492 426456 45619 426458
rect 41492 426400 45558 426456
rect 45614 426400 45619 426456
rect 41492 426398 45619 426400
rect 45553 426395 45619 426398
rect 41321 426050 41387 426053
rect 41308 426048 41387 426050
rect 41308 425992 41326 426048
rect 41382 425992 41387 426048
rect 41308 425990 41387 425992
rect 41321 425987 41387 425990
rect 40953 425642 41019 425645
rect 40940 425640 41019 425642
rect 40940 425584 40958 425640
rect 41014 425584 41019 425640
rect 40940 425582 41019 425584
rect 40953 425579 41019 425582
rect 41822 425234 41828 425236
rect 41492 425174 41828 425234
rect 41822 425172 41828 425174
rect 41892 425172 41898 425236
rect 42006 424826 42012 424828
rect 41492 424766 42012 424826
rect 42006 424764 42012 424766
rect 42076 424764 42082 424828
rect 36537 424418 36603 424421
rect 36524 424416 36603 424418
rect 36524 424360 36542 424416
rect 36598 424360 36603 424416
rect 36524 424358 36603 424360
rect 36537 424355 36603 424358
rect 41321 424010 41387 424013
rect 41308 424008 41387 424010
rect 41308 423952 41326 424008
rect 41382 423952 41387 424008
rect 41308 423950 41387 423952
rect 41321 423947 41387 423950
rect 46933 423602 46999 423605
rect 41492 423600 46999 423602
rect 41492 423544 46938 423600
rect 46994 423544 46999 423600
rect 41492 423542 46999 423544
rect 46933 423539 46999 423542
rect 43069 423194 43135 423197
rect 41492 423192 43135 423194
rect 41492 423136 43074 423192
rect 43130 423136 43135 423192
rect 41492 423134 43135 423136
rect 43069 423131 43135 423134
rect 41873 422786 41939 422789
rect 41492 422784 41939 422786
rect 41492 422728 41878 422784
rect 41934 422728 41939 422784
rect 41492 422726 41939 422728
rect 41873 422723 41939 422726
rect 45369 422378 45435 422381
rect 41492 422376 45435 422378
rect 41492 422320 45374 422376
rect 45430 422320 45435 422376
rect 41492 422318 45435 422320
rect 45369 422315 45435 422318
rect 42057 421970 42123 421973
rect 41492 421968 42123 421970
rect 41492 421912 42062 421968
rect 42118 421912 42123 421968
rect 41492 421910 42123 421912
rect 42057 421907 42123 421910
rect 44633 421562 44699 421565
rect 41492 421560 44699 421562
rect 41492 421504 44638 421560
rect 44694 421504 44699 421560
rect 41492 421502 44699 421504
rect 44633 421499 44699 421502
rect 43253 421154 43319 421157
rect 41492 421152 43319 421154
rect 41492 421096 43258 421152
rect 43314 421096 43319 421152
rect 41492 421094 43319 421096
rect 43253 421091 43319 421094
rect 44817 420746 44883 420749
rect 41492 420744 44883 420746
rect 41492 420688 44822 420744
rect 44878 420688 44883 420744
rect 41492 420686 44883 420688
rect 44817 420683 44883 420686
rect 41462 419930 41522 420308
rect 42425 419930 42491 419933
rect 41462 419928 42491 419930
rect 41462 419900 42430 419928
rect 41492 419872 42430 419900
rect 42486 419872 42491 419928
rect 41492 419870 42491 419872
rect 42425 419867 42491 419870
rect 43989 419522 44055 419525
rect 41492 419520 44055 419522
rect 41492 419464 43994 419520
rect 44050 419464 44055 419520
rect 41492 419462 44055 419464
rect 43989 419459 44055 419462
rect 41137 418842 41203 418845
rect 41454 418842 41460 418844
rect 41137 418840 41460 418842
rect 41137 418784 41142 418840
rect 41198 418784 41460 418840
rect 41137 418782 41460 418784
rect 41137 418779 41203 418782
rect 41454 418780 41460 418782
rect 41524 418780 41530 418844
rect 41505 418570 41571 418573
rect 42241 418570 42307 418573
rect 41505 418568 42307 418570
rect 41505 418512 41510 418568
rect 41566 418512 42246 418568
rect 42302 418512 42307 418568
rect 41505 418510 42307 418512
rect 41505 418507 41571 418510
rect 42241 418507 42307 418510
rect 651833 418026 651899 418029
rect 650164 418024 651899 418026
rect 650164 417968 651838 418024
rect 651894 417968 651899 418024
rect 650164 417966 651899 417968
rect 651833 417963 651899 417966
rect 40718 417828 40724 417892
rect 40788 417890 40794 417892
rect 41873 417890 41939 417893
rect 40788 417888 41939 417890
rect 40788 417832 41878 417888
rect 41934 417832 41939 417888
rect 40788 417830 41939 417832
rect 40788 417828 40794 417830
rect 41873 417827 41939 417830
rect 40534 417556 40540 417620
rect 40604 417618 40610 417620
rect 42057 417618 42123 417621
rect 40604 417616 42123 417618
rect 40604 417560 42062 417616
rect 42118 417560 42123 417616
rect 40604 417558 42123 417560
rect 40604 417556 40610 417558
rect 42057 417555 42123 417558
rect 62113 415442 62179 415445
rect 62113 415440 64492 415442
rect 62113 415384 62118 415440
rect 62174 415384 64492 415440
rect 62113 415382 64492 415384
rect 62113 415379 62179 415382
rect 42057 411906 42123 411909
rect 42517 411906 42583 411909
rect 42057 411904 42583 411906
rect 42057 411848 42062 411904
rect 42118 411848 42522 411904
rect 42578 411848 42583 411904
rect 42057 411846 42583 411848
rect 42057 411843 42123 411846
rect 42517 411843 42583 411846
rect 40718 409396 40724 409460
rect 40788 409458 40794 409460
rect 41781 409458 41847 409461
rect 40788 409456 41847 409458
rect 40788 409400 41786 409456
rect 41842 409400 41847 409456
rect 40788 409398 41847 409400
rect 40788 409396 40794 409398
rect 41781 409395 41847 409398
rect 42425 408506 42491 408509
rect 55857 408506 55923 408509
rect 42425 408504 55923 408506
rect 42425 408448 42430 408504
rect 42486 408448 55862 408504
rect 55918 408448 55923 408504
rect 42425 408446 55923 408448
rect 42425 408443 42491 408446
rect 55857 408443 55923 408446
rect 42425 407826 42491 407829
rect 43253 407826 43319 407829
rect 42425 407824 43319 407826
rect 42425 407768 42430 407824
rect 42486 407768 43258 407824
rect 43314 407768 43319 407824
rect 42425 407766 43319 407768
rect 42425 407763 42491 407766
rect 43253 407763 43319 407766
rect 42425 407010 42491 407013
rect 44633 407010 44699 407013
rect 42425 407008 44699 407010
rect 42425 406952 42430 407008
rect 42486 406952 44638 407008
rect 44694 406952 44699 407008
rect 42425 406950 44699 406952
rect 42425 406947 42491 406950
rect 44633 406947 44699 406950
rect 41781 406332 41847 406333
rect 41781 406328 41828 406332
rect 41892 406330 41898 406332
rect 661861 406330 661927 406333
rect 683113 406330 683179 406333
rect 41781 406272 41786 406328
rect 41781 406268 41828 406272
rect 41892 406270 41938 406330
rect 661861 406328 683179 406330
rect 661861 406272 661866 406328
rect 661922 406272 683118 406328
rect 683174 406272 683179 406328
rect 661861 406270 683179 406272
rect 41892 406268 41898 406270
rect 41781 406267 41847 406268
rect 661861 406267 661927 406270
rect 683113 406267 683179 406270
rect 42609 405650 42675 405653
rect 45369 405650 45435 405653
rect 42609 405648 45435 405650
rect 42609 405592 42614 405648
rect 42670 405592 45374 405648
rect 45430 405592 45435 405648
rect 42609 405590 45435 405592
rect 42609 405587 42675 405590
rect 45369 405587 45435 405590
rect 660297 405650 660363 405653
rect 676029 405650 676095 405653
rect 660297 405648 676095 405650
rect 660297 405592 660302 405648
rect 660358 405592 676034 405648
rect 676090 405592 676095 405648
rect 660297 405590 676095 405592
rect 660297 405587 660363 405590
rect 676029 405587 676095 405590
rect 651465 404698 651531 404701
rect 650164 404696 651531 404698
rect 650164 404640 651470 404696
rect 651526 404640 651531 404696
rect 650164 404638 651531 404640
rect 651465 404635 651531 404638
rect 40534 403820 40540 403884
rect 40604 403882 40610 403884
rect 41781 403882 41847 403885
rect 40604 403880 41847 403882
rect 40604 403824 41786 403880
rect 41842 403824 41847 403880
rect 40604 403822 41847 403824
rect 40604 403820 40610 403822
rect 41781 403819 41847 403822
rect 669957 403746 670023 403749
rect 676262 403746 676322 403852
rect 669957 403744 676322 403746
rect 669957 403688 669962 403744
rect 670018 403688 676322 403744
rect 669957 403686 676322 403688
rect 669957 403683 670023 403686
rect 676029 403474 676095 403477
rect 676029 403472 676292 403474
rect 676029 403416 676034 403472
rect 676090 403416 676292 403472
rect 676029 403414 676292 403416
rect 676029 403411 676095 403414
rect 683113 403338 683179 403341
rect 683070 403336 683179 403338
rect 683070 403280 683118 403336
rect 683174 403280 683179 403336
rect 683070 403275 683179 403280
rect 683070 403036 683130 403275
rect 42333 402930 42399 402933
rect 43069 402930 43135 402933
rect 42333 402928 43135 402930
rect 42333 402872 42338 402928
rect 42394 402872 43074 402928
rect 43130 402872 43135 402928
rect 42333 402870 43135 402872
rect 42333 402867 42399 402870
rect 43069 402867 43135 402870
rect 676806 402868 676812 402932
rect 676876 402868 676882 402932
rect 676814 402628 676874 402868
rect 62113 402386 62179 402389
rect 62113 402384 64492 402386
rect 62113 402328 62118 402384
rect 62174 402328 64492 402384
rect 62113 402326 64492 402328
rect 62113 402323 62179 402326
rect 674189 402250 674255 402253
rect 674189 402248 676292 402250
rect 674189 402192 674194 402248
rect 674250 402192 676292 402248
rect 674189 402190 676292 402192
rect 674189 402187 674255 402190
rect 41781 401844 41847 401845
rect 41781 401840 41828 401844
rect 41892 401842 41898 401844
rect 41781 401784 41786 401840
rect 41781 401780 41828 401784
rect 41892 401782 41938 401842
rect 41892 401780 41898 401782
rect 41781 401779 41847 401780
rect 672441 401706 672507 401709
rect 676262 401706 676322 401812
rect 672441 401704 676322 401706
rect 672441 401648 672446 401704
rect 672502 401648 676322 401704
rect 672441 401646 676322 401648
rect 672441 401643 672507 401646
rect 674649 401434 674715 401437
rect 674649 401432 676292 401434
rect 674649 401376 674654 401432
rect 674710 401376 676292 401432
rect 674649 401374 676292 401376
rect 674649 401371 674715 401374
rect 676990 401236 676996 401300
rect 677060 401236 677066 401300
rect 676998 400996 677058 401236
rect 672441 400482 672507 400485
rect 676262 400482 676322 400588
rect 672441 400480 676322 400482
rect 672441 400424 672446 400480
rect 672502 400424 676322 400480
rect 672441 400422 676322 400424
rect 672441 400419 672507 400422
rect 42425 400210 42491 400213
rect 46933 400210 46999 400213
rect 42425 400208 46999 400210
rect 42425 400152 42430 400208
rect 42486 400152 46938 400208
rect 46994 400152 46999 400208
rect 42425 400150 46999 400152
rect 42425 400147 42491 400150
rect 46933 400147 46999 400150
rect 672625 400074 672691 400077
rect 676262 400074 676322 400180
rect 672625 400072 676322 400074
rect 672625 400016 672630 400072
rect 672686 400016 676322 400072
rect 672625 400014 676322 400016
rect 672625 400011 672691 400014
rect 42425 399802 42491 399805
rect 45553 399802 45619 399805
rect 42425 399800 45619 399802
rect 42425 399744 42430 399800
rect 42486 399744 45558 399800
rect 45614 399744 45619 399800
rect 42425 399742 45619 399744
rect 42425 399739 42491 399742
rect 45553 399739 45619 399742
rect 676262 399666 676322 399772
rect 674790 399606 676322 399666
rect 41454 398788 41460 398852
rect 41524 398850 41530 398852
rect 41781 398850 41847 398853
rect 41524 398848 41847 398850
rect 41524 398792 41786 398848
rect 41842 398792 41847 398848
rect 41524 398790 41847 398792
rect 41524 398788 41530 398790
rect 41781 398787 41847 398790
rect 673177 398850 673243 398853
rect 674790 398850 674850 399606
rect 676029 399394 676095 399397
rect 676029 399392 676292 399394
rect 676029 399336 676034 399392
rect 676090 399336 676292 399392
rect 676029 399334 676292 399336
rect 676029 399331 676095 399334
rect 673177 398848 674850 398850
rect 673177 398792 673182 398848
rect 673238 398792 674850 398848
rect 673177 398790 674850 398792
rect 673177 398787 673243 398790
rect 675886 398788 675892 398852
rect 675956 398850 675962 398852
rect 676262 398850 676322 398956
rect 675956 398790 676322 398850
rect 675956 398788 675962 398790
rect 676262 398445 676322 398548
rect 676213 398440 676322 398445
rect 676213 398384 676218 398440
rect 676274 398384 676322 398440
rect 676213 398382 676322 398384
rect 676213 398379 676279 398382
rect 676446 398037 676506 398140
rect 676397 398032 676506 398037
rect 676397 397976 676402 398032
rect 676458 397976 676506 398032
rect 676397 397974 676506 397976
rect 676397 397971 676463 397974
rect 681046 397629 681106 397732
rect 680997 397624 681106 397629
rect 680997 397568 681002 397624
rect 681058 397568 681106 397624
rect 680997 397566 681106 397568
rect 680997 397563 681063 397566
rect 672993 397218 673059 397221
rect 676262 397218 676322 397324
rect 672993 397216 676322 397218
rect 672993 397160 672998 397216
rect 673054 397160 676322 397216
rect 672993 397158 676322 397160
rect 672993 397155 673059 397158
rect 676630 396812 676690 396916
rect 676622 396748 676628 396812
rect 676692 396748 676698 396812
rect 673361 396402 673427 396405
rect 676262 396402 676322 396508
rect 673361 396400 676322 396402
rect 673361 396344 673366 396400
rect 673422 396344 676322 396400
rect 673361 396342 676322 396344
rect 673361 396339 673427 396342
rect 673821 396130 673887 396133
rect 673821 396128 676292 396130
rect 673821 396072 673826 396128
rect 673882 396072 676292 396128
rect 673821 396070 676292 396072
rect 673821 396067 673887 396070
rect 674005 395722 674071 395725
rect 674005 395720 676292 395722
rect 674005 395664 674010 395720
rect 674066 395664 676292 395720
rect 674005 395662 676292 395664
rect 674005 395659 674071 395662
rect 676262 395180 676322 395284
rect 676254 395116 676260 395180
rect 676324 395116 676330 395180
rect 676446 394772 676506 394876
rect 676438 394708 676444 394772
rect 676508 394708 676514 394772
rect 674465 394498 674531 394501
rect 674465 394496 676292 394498
rect 674465 394440 674470 394496
rect 674526 394440 676292 394496
rect 674465 394438 676292 394440
rect 674465 394435 674531 394438
rect 672257 393954 672323 393957
rect 676262 393954 676322 394060
rect 672257 393952 676322 393954
rect 672257 393896 672262 393952
rect 672318 393896 676322 393952
rect 672257 393894 676322 393896
rect 672257 393891 672323 393894
rect 670601 393546 670667 393549
rect 676262 393546 676322 393652
rect 670601 393544 676322 393546
rect 670601 393488 670606 393544
rect 670662 393488 676322 393544
rect 670601 393486 676322 393488
rect 670601 393483 670667 393486
rect 676070 393076 676076 393140
rect 676140 393138 676146 393140
rect 676262 393138 676322 393244
rect 676140 393078 676322 393138
rect 676140 393076 676146 393078
rect 676262 392836 676322 393078
rect 672717 392594 672783 392597
rect 672717 392592 676322 392594
rect 672717 392536 672722 392592
rect 672778 392536 676322 392592
rect 672717 392534 676322 392536
rect 672717 392531 672783 392534
rect 676262 392428 676322 392534
rect 652569 391506 652635 391509
rect 650164 391504 652635 391506
rect 650164 391448 652574 391504
rect 652630 391448 652635 391504
rect 650164 391446 652635 391448
rect 652569 391443 652635 391446
rect 62113 389330 62179 389333
rect 62113 389328 64492 389330
rect 62113 389272 62118 389328
rect 62174 389272 64492 389328
rect 62113 389270 64492 389272
rect 62113 389267 62179 389270
rect 41492 387638 51090 387698
rect 41492 387230 49250 387290
rect 41137 387154 41203 387157
rect 41094 387152 41203 387154
rect 41094 387096 41142 387152
rect 41198 387096 41203 387152
rect 41094 387091 41203 387096
rect 41094 386852 41154 387091
rect 41873 387018 41939 387021
rect 48957 387018 49023 387021
rect 41873 387016 49023 387018
rect 41873 386960 41878 387016
rect 41934 386960 48962 387016
rect 49018 386960 49023 387016
rect 41873 386958 49023 386960
rect 41873 386955 41939 386958
rect 48957 386955 49023 386958
rect 41321 386746 41387 386749
rect 41278 386744 41387 386746
rect 41278 386688 41326 386744
rect 41382 386688 41387 386744
rect 41278 386683 41387 386688
rect 41505 386746 41571 386749
rect 45001 386746 45067 386749
rect 41505 386744 45067 386746
rect 41505 386688 41510 386744
rect 41566 386688 45006 386744
rect 45062 386688 45067 386744
rect 41505 386686 45067 386688
rect 41505 386683 41571 386686
rect 45001 386683 45067 386686
rect 41278 386444 41338 386683
rect 49190 386474 49250 387230
rect 51030 386746 51090 387638
rect 675702 387636 675708 387700
rect 675772 387698 675778 387700
rect 680997 387698 681063 387701
rect 675772 387696 681063 387698
rect 675772 387640 681002 387696
rect 681058 387640 681063 387696
rect 675772 387638 681063 387640
rect 675772 387636 675778 387638
rect 680997 387635 681063 387638
rect 51717 386746 51783 386749
rect 51030 386744 51783 386746
rect 51030 386688 51722 386744
rect 51778 386688 51783 386744
rect 51030 386686 51783 386688
rect 51717 386683 51783 386686
rect 51901 386474 51967 386477
rect 49190 386472 51967 386474
rect 49190 386416 51906 386472
rect 51962 386416 51967 386472
rect 49190 386414 51967 386416
rect 51901 386411 51967 386414
rect 45369 386066 45435 386069
rect 41492 386064 45435 386066
rect 41492 386008 45374 386064
rect 45430 386008 45435 386064
rect 41492 386006 45435 386008
rect 45369 386003 45435 386006
rect 44173 385658 44239 385661
rect 41492 385656 44239 385658
rect 41492 385600 44178 385656
rect 44234 385600 44239 385656
rect 41492 385598 44239 385600
rect 44173 385595 44239 385598
rect 44633 385250 44699 385253
rect 41492 385248 44699 385250
rect 41492 385192 44638 385248
rect 44694 385192 44699 385248
rect 41492 385190 44699 385192
rect 44633 385187 44699 385190
rect 675753 384978 675819 384981
rect 676622 384978 676628 384980
rect 675753 384976 676628 384978
rect 675753 384920 675758 384976
rect 675814 384920 676628 384976
rect 675753 384918 676628 384920
rect 675753 384915 675819 384918
rect 676622 384916 676628 384918
rect 676692 384916 676698 384980
rect 44449 384842 44515 384845
rect 41492 384840 44515 384842
rect 41492 384784 44454 384840
rect 44510 384784 44515 384840
rect 41492 384782 44515 384784
rect 44449 384779 44515 384782
rect 45001 384434 45067 384437
rect 41492 384432 45067 384434
rect 41492 384376 45006 384432
rect 45062 384376 45067 384432
rect 41492 384374 45067 384376
rect 45001 384371 45067 384374
rect 45185 384026 45251 384029
rect 41492 384024 45251 384026
rect 41492 383968 45190 384024
rect 45246 383968 45251 384024
rect 41492 383966 45251 383968
rect 45185 383963 45251 383966
rect 45185 383618 45251 383621
rect 41492 383616 45251 383618
rect 41492 383560 45190 383616
rect 45246 383560 45251 383616
rect 41492 383558 45251 383560
rect 45185 383555 45251 383558
rect 46933 383210 46999 383213
rect 41492 383208 46999 383210
rect 41492 383152 46938 383208
rect 46994 383152 46999 383208
rect 41492 383150 46999 383152
rect 46933 383147 46999 383150
rect 41278 382669 41338 382772
rect 41278 382664 41387 382669
rect 41278 382608 41326 382664
rect 41382 382608 41387 382664
rect 41278 382606 41387 382608
rect 41321 382603 41387 382606
rect 39990 382261 40050 382364
rect 39990 382256 40099 382261
rect 39990 382200 40038 382256
rect 40094 382200 40099 382256
rect 39990 382198 40099 382200
rect 40033 382195 40099 382198
rect 673361 382258 673427 382261
rect 675385 382258 675451 382261
rect 673361 382256 675451 382258
rect 673361 382200 673366 382256
rect 673422 382200 675390 382256
rect 675446 382200 675451 382256
rect 673361 382198 675451 382200
rect 673361 382195 673427 382198
rect 675385 382195 675451 382198
rect 41462 381852 41522 381956
rect 41454 381788 41460 381852
rect 41524 381788 41530 381852
rect 37966 381445 38026 381548
rect 37917 381440 38026 381445
rect 37917 381384 37922 381440
rect 37978 381384 38026 381440
rect 37917 381382 38026 381384
rect 673821 381442 673887 381445
rect 675109 381442 675175 381445
rect 673821 381440 675175 381442
rect 673821 381384 673826 381440
rect 673882 381384 675114 381440
rect 675170 381384 675175 381440
rect 673821 381382 675175 381384
rect 37917 381379 37983 381382
rect 673821 381379 673887 381382
rect 675109 381379 675175 381382
rect 40174 381037 40234 381140
rect 40174 381032 40283 381037
rect 40174 380976 40222 381032
rect 40278 380976 40283 381032
rect 40174 380974 40283 380976
rect 40217 380971 40283 380974
rect 45553 380762 45619 380765
rect 41492 380760 45619 380762
rect 41492 380704 45558 380760
rect 45614 380704 45619 380760
rect 41492 380702 45619 380704
rect 45553 380699 45619 380702
rect 675753 380626 675819 380629
rect 676438 380626 676444 380628
rect 675753 380624 676444 380626
rect 675753 380568 675758 380624
rect 675814 380568 676444 380624
rect 675753 380566 676444 380568
rect 675753 380563 675819 380566
rect 676438 380564 676444 380566
rect 676508 380564 676514 380628
rect 33734 380221 33794 380324
rect 33734 380216 33843 380221
rect 33734 380160 33782 380216
rect 33838 380160 33843 380216
rect 33734 380158 33843 380160
rect 33777 380155 33843 380158
rect 45737 379946 45803 379949
rect 41492 379944 45803 379946
rect 41492 379888 45742 379944
rect 45798 379888 45803 379944
rect 41492 379886 45803 379888
rect 45737 379883 45803 379886
rect 35758 379405 35818 379530
rect 35758 379400 35867 379405
rect 35758 379344 35806 379400
rect 35862 379344 35867 379400
rect 35758 379342 35867 379344
rect 35801 379339 35867 379342
rect 47117 379130 47183 379133
rect 41492 379128 47183 379130
rect 41492 379072 47122 379128
rect 47178 379072 47183 379128
rect 41492 379070 47183 379072
rect 47117 379067 47183 379070
rect 675753 378724 675819 378725
rect 675702 378722 675708 378724
rect 40542 378588 40602 378692
rect 675662 378662 675708 378722
rect 675772 378720 675819 378724
rect 675814 378664 675819 378720
rect 675702 378660 675708 378662
rect 675772 378660 675819 378664
rect 675753 378659 675819 378660
rect 40534 378524 40540 378588
rect 40604 378524 40610 378588
rect 40726 378180 40786 378284
rect 40718 378116 40724 378180
rect 40788 378116 40794 378180
rect 652017 378178 652083 378181
rect 650164 378176 652083 378178
rect 650164 378120 652022 378176
rect 652078 378120 652083 378176
rect 650164 378118 652083 378120
rect 652017 378115 652083 378118
rect 672993 378042 673059 378045
rect 674782 378042 674788 378044
rect 672993 378040 674788 378042
rect 672993 377984 672998 378040
rect 673054 377984 674788 378040
rect 672993 377982 674788 377984
rect 672993 377979 673059 377982
rect 674782 377980 674788 377982
rect 674852 377980 674858 378044
rect 44449 377906 44515 377909
rect 41492 377904 44515 377906
rect 41492 377848 44454 377904
rect 44510 377848 44515 377904
rect 41492 377846 44515 377848
rect 44449 377843 44515 377846
rect 674465 377770 674531 377773
rect 675109 377770 675175 377773
rect 674465 377768 675175 377770
rect 674465 377712 674470 377768
rect 674526 377712 675114 377768
rect 675170 377712 675175 377768
rect 674465 377710 675175 377712
rect 674465 377707 674531 377710
rect 675109 377707 675175 377710
rect 44265 377498 44331 377501
rect 41492 377496 44331 377498
rect 41492 377440 44270 377496
rect 44326 377440 44331 377496
rect 41492 377438 44331 377440
rect 44265 377435 44331 377438
rect 675753 377362 675819 377365
rect 676254 377362 676260 377364
rect 675753 377360 676260 377362
rect 675753 377304 675758 377360
rect 675814 377304 676260 377360
rect 675753 377302 676260 377304
rect 675753 377299 675819 377302
rect 676254 377300 676260 377302
rect 676324 377300 676330 377364
rect 27662 376546 27722 377060
rect 40033 376954 40099 376957
rect 41638 376954 41644 376956
rect 40033 376952 41644 376954
rect 40033 376896 40038 376952
rect 40094 376896 41644 376952
rect 40033 376894 41644 376896
rect 40033 376891 40099 376894
rect 41638 376892 41644 376894
rect 41708 376892 41714 376956
rect 675201 376954 675267 376957
rect 675886 376954 675892 376956
rect 675201 376952 675892 376954
rect 675201 376896 675206 376952
rect 675262 376896 675892 376952
rect 675201 376894 675892 376896
rect 675201 376891 675267 376894
rect 675886 376892 675892 376894
rect 675956 376892 675962 376956
rect 28533 376546 28599 376549
rect 27662 376544 28599 376546
rect 27662 376488 28538 376544
rect 28594 376488 28599 376544
rect 27662 376486 28599 376488
rect 28533 376483 28599 376486
rect 62113 376274 62179 376277
rect 672257 376274 672323 376277
rect 675385 376274 675451 376277
rect 62113 376272 64492 376274
rect 35758 376141 35818 376244
rect 62113 376216 62118 376272
rect 62174 376216 64492 376272
rect 62113 376214 64492 376216
rect 672257 376272 675451 376274
rect 672257 376216 672262 376272
rect 672318 376216 675390 376272
rect 675446 376216 675451 376272
rect 672257 376214 675451 376216
rect 62113 376211 62179 376214
rect 672257 376211 672323 376214
rect 675385 376211 675451 376214
rect 35758 376136 35867 376141
rect 35758 376080 35806 376136
rect 35862 376080 35867 376136
rect 35758 376078 35867 376080
rect 35801 376075 35867 376078
rect 41689 375458 41755 375461
rect 43345 375458 43411 375461
rect 41689 375456 43411 375458
rect 41689 375400 41694 375456
rect 41750 375400 43350 375456
rect 43406 375400 43411 375456
rect 41689 375398 43411 375400
rect 41689 375395 41755 375398
rect 43345 375395 43411 375398
rect 674005 375458 674071 375461
rect 675385 375458 675451 375461
rect 674005 375456 675451 375458
rect 674005 375400 674010 375456
rect 674066 375400 675390 375456
rect 675446 375400 675451 375456
rect 674005 375398 675451 375400
rect 674005 375395 674071 375398
rect 675385 375395 675451 375398
rect 28533 373282 28599 373285
rect 41270 373282 41276 373284
rect 28533 373280 41276 373282
rect 28533 373224 28538 373280
rect 28594 373224 41276 373280
rect 28533 373222 41276 373224
rect 28533 373219 28599 373222
rect 41270 373220 41276 373222
rect 41340 373220 41346 373284
rect 675753 373010 675819 373013
rect 676070 373010 676076 373012
rect 675753 373008 676076 373010
rect 675753 372952 675758 373008
rect 675814 372952 676076 373008
rect 675753 372950 676076 372952
rect 675753 372947 675819 372950
rect 676070 372948 676076 372950
rect 676140 372948 676146 373012
rect 41689 372602 41755 372605
rect 42609 372602 42675 372605
rect 41689 372600 42675 372602
rect 41689 372544 41694 372600
rect 41750 372544 42614 372600
rect 42670 372544 42675 372600
rect 41689 372542 42675 372544
rect 41689 372539 41755 372542
rect 42609 372539 42675 372542
rect 674782 372540 674788 372604
rect 674852 372602 674858 372604
rect 675109 372602 675175 372605
rect 674852 372600 675175 372602
rect 674852 372544 675114 372600
rect 675170 372544 675175 372600
rect 674852 372542 675175 372544
rect 674852 372540 674858 372542
rect 675109 372539 675175 372542
rect 33777 371922 33843 371925
rect 41822 371922 41828 371924
rect 33777 371920 41828 371922
rect 33777 371864 33782 371920
rect 33838 371864 41828 371920
rect 33777 371862 41828 371864
rect 33777 371859 33843 371862
rect 41822 371860 41828 371862
rect 41892 371860 41898 371924
rect 41270 368460 41276 368524
rect 41340 368522 41346 368524
rect 41781 368522 41847 368525
rect 41340 368520 41847 368522
rect 41340 368464 41786 368520
rect 41842 368464 41847 368520
rect 41340 368462 41847 368464
rect 41340 368460 41346 368462
rect 41781 368459 41847 368462
rect 42425 367026 42491 367029
rect 46197 367026 46263 367029
rect 42425 367024 46263 367026
rect 42425 366968 42430 367024
rect 42486 366968 46202 367024
rect 46258 366968 46263 367024
rect 42425 366966 46263 366968
rect 42425 366963 42491 366966
rect 46197 366963 46263 366966
rect 42333 365802 42399 365805
rect 42793 365802 42859 365805
rect 42333 365800 42859 365802
rect 42333 365744 42338 365800
rect 42394 365744 42798 365800
rect 42854 365744 42859 365800
rect 42333 365742 42859 365744
rect 42333 365739 42399 365742
rect 42793 365739 42859 365742
rect 42149 364986 42215 364989
rect 44449 364986 44515 364989
rect 42149 364984 44515 364986
rect 42149 364928 42154 364984
rect 42210 364928 44454 364984
rect 44510 364928 44515 364984
rect 42149 364926 44515 364928
rect 42149 364923 42215 364926
rect 44449 364923 44515 364926
rect 651649 364850 651715 364853
rect 650164 364848 651715 364850
rect 650164 364792 651654 364848
rect 651710 364792 651715 364848
rect 650164 364790 651715 364792
rect 651649 364787 651715 364790
rect 42425 364306 42491 364309
rect 47117 364306 47183 364309
rect 42425 364304 47183 364306
rect 42425 364248 42430 364304
rect 42486 364248 47122 364304
rect 47178 364248 47183 364304
rect 42425 364246 47183 364248
rect 42425 364243 42491 364246
rect 47117 364243 47183 364246
rect 40718 363564 40724 363628
rect 40788 363626 40794 363628
rect 41781 363626 41847 363629
rect 40788 363624 41847 363626
rect 40788 363568 41786 363624
rect 41842 363568 41847 363624
rect 40788 363566 41847 363568
rect 40788 363564 40794 363566
rect 41781 363563 41847 363566
rect 62113 363354 62179 363357
rect 62113 363352 64492 363354
rect 62113 363296 62118 363352
rect 62174 363296 64492 363352
rect 62113 363294 64492 363296
rect 62113 363291 62179 363294
rect 667197 360906 667263 360909
rect 675845 360906 675911 360909
rect 667197 360904 675911 360906
rect 667197 360848 667202 360904
rect 667258 360848 675850 360904
rect 675906 360848 675911 360904
rect 667197 360846 675911 360848
rect 667197 360843 667263 360846
rect 675845 360843 675911 360846
rect 40534 360028 40540 360092
rect 40604 360090 40610 360092
rect 41781 360090 41847 360093
rect 40604 360088 41847 360090
rect 40604 360032 41786 360088
rect 41842 360032 41847 360088
rect 40604 360030 41847 360032
rect 40604 360028 40610 360030
rect 41781 360027 41847 360030
rect 659101 360090 659167 360093
rect 676029 360090 676095 360093
rect 659101 360088 676095 360090
rect 659101 360032 659106 360088
rect 659162 360032 676034 360088
rect 676090 360032 676095 360088
rect 659101 360030 676095 360032
rect 659101 360027 659167 360030
rect 676029 360027 676095 360030
rect 42149 359954 42215 359957
rect 45737 359954 45803 359957
rect 42149 359952 45803 359954
rect 42149 359896 42154 359952
rect 42210 359896 45742 359952
rect 45798 359896 45803 359952
rect 42149 359894 45803 359896
rect 42149 359891 42215 359894
rect 45737 359891 45803 359894
rect 41781 359412 41847 359413
rect 41781 359408 41828 359412
rect 41892 359410 41898 359412
rect 41781 359352 41786 359408
rect 41781 359348 41828 359352
rect 41892 359350 41938 359410
rect 41892 359348 41898 359350
rect 41781 359347 41847 359348
rect 41454 358668 41460 358732
rect 41524 358730 41530 358732
rect 41781 358730 41847 358733
rect 41524 358728 41847 358730
rect 41524 358672 41786 358728
rect 41842 358672 41847 358728
rect 41524 358670 41847 358672
rect 41524 358668 41530 358670
rect 41781 358667 41847 358670
rect 663750 358670 676292 358730
rect 663241 358594 663307 358597
rect 663750 358594 663810 358670
rect 663241 358592 663810 358594
rect 663241 358536 663246 358592
rect 663302 358536 663810 358592
rect 663241 358534 663810 358536
rect 663241 358531 663307 358534
rect 676029 358322 676095 358325
rect 676029 358320 676292 358322
rect 676029 358264 676034 358320
rect 676090 358264 676292 358320
rect 676029 358262 676292 358264
rect 676029 358259 676095 358262
rect 675845 357914 675911 357917
rect 675845 357912 676292 357914
rect 675845 357856 675850 357912
rect 675906 357856 676292 357912
rect 675845 357854 676292 357856
rect 675845 357851 675911 357854
rect 674189 357506 674255 357509
rect 674189 357504 676292 357506
rect 674189 357448 674194 357504
rect 674250 357448 676292 357504
rect 674189 357446 676292 357448
rect 674189 357443 674255 357446
rect 674649 357098 674715 357101
rect 674649 357096 676292 357098
rect 674649 357040 674654 357096
rect 674710 357040 676292 357096
rect 674649 357038 676292 357040
rect 674649 357035 674715 357038
rect 42425 356962 42491 356965
rect 45553 356962 45619 356965
rect 42425 356960 45619 356962
rect 42425 356904 42430 356960
rect 42486 356904 45558 356960
rect 45614 356904 45619 356960
rect 42425 356902 45619 356904
rect 42425 356899 42491 356902
rect 45553 356899 45619 356902
rect 44265 356690 44331 356693
rect 45645 356690 45711 356693
rect 44265 356688 45711 356690
rect 44265 356632 44270 356688
rect 44326 356632 45650 356688
rect 45706 356632 45711 356688
rect 44265 356630 45711 356632
rect 44265 356627 44331 356630
rect 45645 356627 45711 356630
rect 674465 356690 674531 356693
rect 674465 356688 676292 356690
rect 674465 356632 674470 356688
rect 674526 356632 676292 356688
rect 674465 356630 676292 356632
rect 674465 356627 674531 356630
rect 42149 356418 42215 356421
rect 46933 356418 46999 356421
rect 42149 356416 46999 356418
rect 42149 356360 42154 356416
rect 42210 356360 46938 356416
rect 46994 356360 46999 356416
rect 42149 356358 46999 356360
rect 42149 356355 42215 356358
rect 46933 356355 46999 356358
rect 674097 356282 674163 356285
rect 674097 356280 676292 356282
rect 674097 356224 674102 356280
rect 674158 356224 676292 356280
rect 674097 356222 676292 356224
rect 674097 356219 674163 356222
rect 43345 355874 43411 355877
rect 45921 355874 45987 355877
rect 43345 355872 45987 355874
rect 43345 355816 43350 355872
rect 43406 355816 45926 355872
rect 45982 355816 45987 355872
rect 43345 355814 45987 355816
rect 43345 355811 43411 355814
rect 45921 355811 45987 355814
rect 672441 355874 672507 355877
rect 672441 355872 676292 355874
rect 672441 355816 672446 355872
rect 672502 355816 676292 355872
rect 672441 355814 676292 355816
rect 672441 355811 672507 355814
rect 41873 355740 41939 355741
rect 41822 355738 41828 355740
rect 41782 355678 41828 355738
rect 41892 355736 41939 355740
rect 41934 355680 41939 355736
rect 41822 355676 41828 355678
rect 41892 355676 41939 355680
rect 41873 355675 41939 355676
rect 673177 355466 673243 355469
rect 673177 355464 676292 355466
rect 673177 355408 673182 355464
rect 673238 355408 676292 355464
rect 673177 355406 676292 355408
rect 673177 355403 673243 355406
rect 673361 355058 673427 355061
rect 673361 355056 676292 355058
rect 673361 355000 673366 355056
rect 673422 355000 676292 355056
rect 673361 354998 676292 355000
rect 673361 354995 673427 354998
rect 672533 354650 672599 354653
rect 672533 354648 676292 354650
rect 672533 354592 672538 354648
rect 672594 354592 676292 354648
rect 672533 354590 676292 354592
rect 672533 354587 672599 354590
rect 43897 354244 43963 354245
rect 43846 354180 43852 354244
rect 43916 354242 43963 354244
rect 43916 354240 44008 354242
rect 43958 354184 44008 354240
rect 43916 354182 44008 354184
rect 43916 354180 43963 354182
rect 675334 354180 675340 354244
rect 675404 354242 675410 354244
rect 675404 354182 676292 354242
rect 675404 354180 675410 354182
rect 43897 354179 43963 354180
rect 44214 353772 44220 353836
rect 44284 353834 44290 353836
rect 44725 353834 44791 353837
rect 44284 353832 44791 353834
rect 44284 353776 44730 353832
rect 44786 353776 44791 353832
rect 44284 353774 44791 353776
rect 44284 353772 44290 353774
rect 44725 353771 44791 353774
rect 676029 353834 676095 353837
rect 676029 353832 676292 353834
rect 676029 353776 676034 353832
rect 676090 353776 676292 353832
rect 676029 353774 676292 353776
rect 676029 353771 676095 353774
rect 672165 353426 672231 353429
rect 672165 353424 676292 353426
rect 672165 353368 672170 353424
rect 672226 353368 676292 353424
rect 672165 353366 676292 353368
rect 672165 353363 672231 353366
rect 675702 352956 675708 353020
rect 675772 353018 675778 353020
rect 675772 352958 676292 353018
rect 675772 352956 675778 352958
rect 673913 352610 673979 352613
rect 673913 352608 676292 352610
rect 673913 352552 673918 352608
rect 673974 352552 676292 352608
rect 673913 352550 676292 352552
rect 673913 352547 673979 352550
rect 673545 352202 673611 352205
rect 673545 352200 676292 352202
rect 673545 352144 673550 352200
rect 673606 352144 676292 352200
rect 673545 352142 676292 352144
rect 673545 352139 673611 352142
rect 675886 351732 675892 351796
rect 675956 351794 675962 351796
rect 675956 351734 676292 351794
rect 675956 351732 675962 351734
rect 651465 351658 651531 351661
rect 650164 351656 651531 351658
rect 650164 351600 651470 351656
rect 651526 351600 651531 351656
rect 650164 351598 651531 351600
rect 651465 351595 651531 351598
rect 672993 351386 673059 351389
rect 672993 351384 676292 351386
rect 672993 351328 672998 351384
rect 673054 351328 676292 351384
rect 672993 351326 676292 351328
rect 672993 351323 673059 351326
rect 28533 351250 28599 351253
rect 50521 351250 50587 351253
rect 28533 351248 50587 351250
rect 28533 351192 28538 351248
rect 28594 351192 50526 351248
rect 50582 351192 50587 351248
rect 28533 351190 50587 351192
rect 28533 351187 28599 351190
rect 50521 351187 50587 351190
rect 675886 350916 675892 350980
rect 675956 350978 675962 350980
rect 675956 350918 676292 350978
rect 675956 350916 675962 350918
rect 673729 350570 673795 350573
rect 673729 350568 676292 350570
rect 673729 350512 673734 350568
rect 673790 350512 676292 350568
rect 673729 350510 676292 350512
rect 673729 350507 673795 350510
rect 62757 350298 62823 350301
rect 62757 350296 64492 350298
rect 62757 350240 62762 350296
rect 62818 350240 64492 350296
rect 62757 350238 64492 350240
rect 62757 350235 62823 350238
rect 675886 350100 675892 350164
rect 675956 350162 675962 350164
rect 675956 350102 676292 350162
rect 675956 350100 675962 350102
rect 673361 349754 673427 349757
rect 673361 349752 676292 349754
rect 673361 349696 673366 349752
rect 673422 349696 676292 349752
rect 673361 349694 676292 349696
rect 673361 349691 673427 349694
rect 674465 349482 674531 349485
rect 674465 349480 676230 349482
rect 674465 349424 674470 349480
rect 674526 349424 676230 349480
rect 674465 349422 676230 349424
rect 674465 349419 674531 349422
rect 676170 349346 676230 349422
rect 676170 349286 676292 349346
rect 675937 349212 676003 349213
rect 675886 349210 675892 349212
rect 675846 349150 675892 349210
rect 675956 349208 676003 349212
rect 675998 349152 676003 349208
rect 675886 349148 675892 349150
rect 675956 349148 676003 349152
rect 675937 349147 676003 349148
rect 671981 348938 672047 348941
rect 671981 348936 676292 348938
rect 671981 348880 671986 348936
rect 672042 348880 676292 348936
rect 671981 348878 676292 348880
rect 671981 348875 672047 348878
rect 672349 348530 672415 348533
rect 672349 348528 676292 348530
rect 672349 348472 672354 348528
rect 672410 348472 676292 348528
rect 672349 348470 676292 348472
rect 672349 348467 672415 348470
rect 674281 347714 674347 347717
rect 683070 347714 683130 348092
rect 674281 347712 683130 347714
rect 674281 347656 674286 347712
rect 674342 347684 683130 347712
rect 674342 347656 683100 347684
rect 674281 347654 683100 347656
rect 674281 347651 674347 347654
rect 669957 347306 670023 347309
rect 669957 347304 676292 347306
rect 669957 347248 669962 347304
rect 670018 347248 676292 347304
rect 669957 347246 676292 347248
rect 669957 347243 670023 347246
rect 40217 345402 40283 345405
rect 47577 345402 47643 345405
rect 40217 345400 47643 345402
rect 40217 345344 40222 345400
rect 40278 345344 47582 345400
rect 47638 345344 47643 345400
rect 40217 345342 47643 345344
rect 40217 345339 40283 345342
rect 47577 345339 47643 345342
rect 28901 344314 28967 344317
rect 41462 344314 41522 344556
rect 54477 344314 54543 344317
rect 28901 344312 29010 344314
rect 28901 344256 28906 344312
rect 28962 344256 29010 344312
rect 28901 344251 29010 344256
rect 41462 344312 54543 344314
rect 41462 344256 54482 344312
rect 54538 344256 54543 344312
rect 41462 344254 54543 344256
rect 54477 344251 54543 344254
rect 28950 344148 29010 344251
rect 28533 343906 28599 343909
rect 28533 343904 28642 343906
rect 28533 343848 28538 343904
rect 28594 343848 28642 343904
rect 28533 343843 28642 343848
rect 28582 343740 28642 343843
rect 45369 343362 45435 343365
rect 41492 343360 45435 343362
rect 41492 343304 45374 343360
rect 45430 343304 45435 343360
rect 41492 343302 45435 343304
rect 45369 343299 45435 343302
rect 44398 342954 44404 342956
rect 41492 342894 44404 342954
rect 44398 342892 44404 342894
rect 44468 342892 44474 342956
rect 44214 342682 44220 342684
rect 41462 342622 44220 342682
rect 41462 342516 41522 342622
rect 44214 342620 44220 342622
rect 44284 342620 44290 342684
rect 44398 342138 44404 342140
rect 41492 342078 44404 342138
rect 44398 342076 44404 342078
rect 44468 342076 44474 342140
rect 45001 341730 45067 341733
rect 41492 341728 45067 341730
rect 41492 341672 45006 341728
rect 45062 341672 45067 341728
rect 41492 341670 45067 341672
rect 45001 341667 45067 341670
rect 44582 341322 44588 341324
rect 41492 341262 44588 341322
rect 44582 341260 44588 341262
rect 44652 341260 44658 341324
rect 45185 340914 45251 340917
rect 41492 340912 45251 340914
rect 41492 340856 45190 340912
rect 45246 340856 45251 340912
rect 41492 340854 45251 340856
rect 45185 340851 45251 340854
rect 672165 340778 672231 340781
rect 675109 340778 675175 340781
rect 672165 340776 675175 340778
rect 672165 340720 672170 340776
rect 672226 340720 675114 340776
rect 675170 340720 675175 340776
rect 672165 340718 675175 340720
rect 672165 340715 672231 340718
rect 675109 340715 675175 340718
rect 43662 340506 43668 340508
rect 41492 340446 43668 340506
rect 43662 340444 43668 340446
rect 43732 340444 43738 340508
rect 675753 340370 675819 340373
rect 676622 340370 676628 340372
rect 675753 340368 676628 340370
rect 675753 340312 675758 340368
rect 675814 340312 676628 340368
rect 675753 340310 676628 340312
rect 675753 340307 675819 340310
rect 676622 340308 676628 340310
rect 676692 340308 676698 340372
rect 45553 340098 45619 340101
rect 41492 340096 45619 340098
rect 41492 340040 45558 340096
rect 45614 340040 45619 340096
rect 41492 340038 45619 340040
rect 45553 340035 45619 340038
rect 35801 339826 35867 339829
rect 35758 339824 35867 339826
rect 35758 339768 35806 339824
rect 35862 339768 35867 339824
rect 35758 339763 35867 339768
rect 35758 339660 35818 339763
rect 35758 339013 35818 339252
rect 35758 339008 35867 339013
rect 675385 339012 675451 339013
rect 675334 339010 675340 339012
rect 35758 338952 35806 339008
rect 35862 338952 35867 339008
rect 35758 338950 35867 338952
rect 675294 338950 675340 339010
rect 675404 339008 675451 339012
rect 675446 338952 675451 339008
rect 35801 338947 35867 338950
rect 675334 338948 675340 338950
rect 675404 338948 675451 338952
rect 675385 338947 675451 338948
rect 30974 338605 31034 338844
rect 30974 338600 31083 338605
rect 30974 338544 31022 338600
rect 31078 338544 31083 338600
rect 30974 338542 31083 338544
rect 31017 338539 31083 338542
rect 46933 338466 46999 338469
rect 41492 338464 46999 338466
rect 41492 338408 46938 338464
rect 46994 338408 46999 338464
rect 41492 338406 46999 338408
rect 46933 338403 46999 338406
rect 651465 338330 651531 338333
rect 650164 338328 651531 338330
rect 650164 338272 651470 338328
rect 651526 338272 651531 338328
rect 650164 338270 651531 338272
rect 651465 338267 651531 338270
rect 672993 338058 673059 338061
rect 675109 338058 675175 338061
rect 672993 338056 675175 338058
rect 40726 337788 40786 338028
rect 672993 338000 672998 338056
rect 673054 338000 675114 338056
rect 675170 338000 675175 338056
rect 672993 337998 675175 338000
rect 672993 337995 673059 337998
rect 675109 337995 675175 337998
rect 675569 337788 675635 337789
rect 40718 337724 40724 337788
rect 40788 337724 40794 337788
rect 675518 337786 675524 337788
rect 675478 337726 675524 337786
rect 675588 337784 675635 337788
rect 675630 337728 675635 337784
rect 675518 337724 675524 337726
rect 675588 337724 675635 337728
rect 675569 337723 675635 337724
rect 42926 337650 42932 337652
rect 41492 337590 42932 337650
rect 42926 337588 42932 337590
rect 42996 337588 43002 337652
rect 45369 337242 45435 337245
rect 41492 337240 45435 337242
rect 41492 337184 45374 337240
rect 45430 337184 45435 337240
rect 41492 337182 45435 337184
rect 45369 337179 45435 337182
rect 62113 337242 62179 337245
rect 62113 337240 64492 337242
rect 62113 337184 62118 337240
rect 62174 337184 64492 337240
rect 62113 337182 64492 337184
rect 62113 337179 62179 337182
rect 43110 336834 43116 336836
rect 41492 336774 43116 336834
rect 43110 336772 43116 336774
rect 43180 336772 43186 336836
rect 673913 336698 673979 336701
rect 675109 336698 675175 336701
rect 673913 336696 675175 336698
rect 673913 336640 673918 336696
rect 673974 336640 675114 336696
rect 675170 336640 675175 336696
rect 673913 336638 675175 336640
rect 673913 336635 673979 336638
rect 675109 336635 675175 336638
rect 675753 336698 675819 336701
rect 676438 336698 676444 336700
rect 675753 336696 676444 336698
rect 675753 336640 675758 336696
rect 675814 336640 676444 336696
rect 675753 336638 676444 336640
rect 675753 336635 675819 336638
rect 676438 336636 676444 336638
rect 676508 336636 676514 336700
rect 41462 336154 41522 336396
rect 43294 336154 43300 336156
rect 41462 336094 43300 336154
rect 43294 336092 43300 336094
rect 43364 336092 43370 336156
rect 40542 335748 40602 335988
rect 673361 335882 673427 335885
rect 675477 335882 675543 335885
rect 673361 335880 675543 335882
rect 673361 335824 673366 335880
rect 673422 335824 675482 335880
rect 675538 335824 675543 335880
rect 673361 335822 675543 335824
rect 673361 335819 673427 335822
rect 675477 335819 675543 335822
rect 40534 335684 40540 335748
rect 40604 335684 40610 335748
rect 41462 335474 41522 335580
rect 41462 335414 44098 335474
rect 44038 335202 44098 335414
rect 41462 335066 41522 335172
rect 44038 335142 44282 335202
rect 42190 335066 42196 335068
rect 41462 335006 42196 335066
rect 42190 335004 42196 335006
rect 42260 335004 42266 335068
rect 41492 334734 42074 334794
rect 42014 334658 42074 334734
rect 44222 334661 44282 335142
rect 42885 334658 42951 334661
rect 43253 334660 43319 334661
rect 43253 334658 43300 334660
rect 42014 334656 42951 334658
rect 42014 334600 42890 334656
rect 42946 334600 42951 334656
rect 42014 334598 42951 334600
rect 43208 334656 43300 334658
rect 43208 334600 43258 334656
rect 43208 334598 43300 334600
rect 42885 334595 42951 334598
rect 43253 334596 43300 334598
rect 43364 334596 43370 334660
rect 44173 334656 44282 334661
rect 44173 334600 44178 334656
rect 44234 334600 44282 334656
rect 44173 334598 44282 334600
rect 43253 334595 43319 334596
rect 44173 334595 44239 334598
rect 37917 334522 37983 334525
rect 41822 334522 41828 334524
rect 37917 334520 41828 334522
rect 37917 334464 37922 334520
rect 37978 334464 41828 334520
rect 37917 334462 41828 334464
rect 37917 334459 37983 334462
rect 41822 334460 41828 334462
rect 41892 334460 41898 334524
rect 41462 334114 41522 334356
rect 42190 334324 42196 334388
rect 42260 334386 42266 334388
rect 42609 334386 42675 334389
rect 42260 334384 42675 334386
rect 42260 334328 42614 334384
rect 42670 334328 42675 334384
rect 42260 334326 42675 334328
rect 42260 334324 42266 334326
rect 42609 334323 42675 334326
rect 48957 334114 49023 334117
rect 41462 334112 49023 334114
rect 41462 334056 48962 334112
rect 49018 334056 49023 334112
rect 41462 334054 49023 334056
rect 48957 334051 49023 334054
rect 27662 333540 27722 333948
rect 40910 333708 40970 333948
rect 40902 333644 40908 333708
rect 40972 333644 40978 333708
rect 47577 333162 47643 333165
rect 41492 333160 47643 333162
rect 41492 333104 47582 333160
rect 47638 333104 47643 333160
rect 41492 333102 47643 333104
rect 47577 333099 47643 333102
rect 674465 332890 674531 332893
rect 675385 332890 675451 332893
rect 674465 332888 675451 332890
rect 674465 332832 674470 332888
rect 674526 332832 675390 332888
rect 675446 332832 675451 332888
rect 674465 332830 675451 332832
rect 674465 332827 674531 332830
rect 675385 332827 675451 332830
rect 671981 332346 672047 332349
rect 675109 332346 675175 332349
rect 671981 332344 675175 332346
rect 671981 332288 671986 332344
rect 672042 332288 675114 332344
rect 675170 332288 675175 332344
rect 671981 332286 675175 332288
rect 671981 332283 672047 332286
rect 675109 332283 675175 332286
rect 675753 332210 675819 332213
rect 676254 332210 676260 332212
rect 675753 332208 676260 332210
rect 675753 332152 675758 332208
rect 675814 332152 676260 332208
rect 675753 332150 676260 332152
rect 675753 332147 675819 332150
rect 676254 332148 676260 332150
rect 676324 332148 676330 332212
rect 673729 331122 673795 331125
rect 675109 331122 675175 331125
rect 673729 331120 675175 331122
rect 673729 331064 673734 331120
rect 673790 331064 675114 331120
rect 675170 331064 675175 331120
rect 673729 331062 675175 331064
rect 673729 331059 673795 331062
rect 675109 331059 675175 331062
rect 31017 329082 31083 329085
rect 41638 329082 41644 329084
rect 31017 329080 41644 329082
rect 31017 329024 31022 329080
rect 31078 329024 41644 329080
rect 31017 329022 41644 329024
rect 31017 329019 31083 329022
rect 41638 329020 41644 329022
rect 41708 329020 41714 329084
rect 36537 328402 36603 328405
rect 41454 328402 41460 328404
rect 36537 328400 41460 328402
rect 36537 328344 36542 328400
rect 36598 328344 41460 328400
rect 36537 328342 41460 328344
rect 36537 328339 36603 328342
rect 41454 328340 41460 328342
rect 41524 328340 41530 328404
rect 675753 328402 675819 328405
rect 676070 328402 676076 328404
rect 675753 328400 676076 328402
rect 675753 328344 675758 328400
rect 675814 328344 676076 328400
rect 675753 328342 676076 328344
rect 675753 328339 675819 328342
rect 676070 328340 676076 328342
rect 676140 328340 676146 328404
rect 674281 327586 674347 327589
rect 675109 327586 675175 327589
rect 674281 327584 675175 327586
rect 674281 327528 674286 327584
rect 674342 327528 675114 327584
rect 675170 327528 675175 327584
rect 674281 327526 675175 327528
rect 674281 327523 674347 327526
rect 675109 327523 675175 327526
rect 40718 326708 40724 326772
rect 40788 326770 40794 326772
rect 41781 326770 41847 326773
rect 40788 326768 41847 326770
rect 40788 326712 41786 326768
rect 41842 326712 41847 326768
rect 40788 326710 41847 326712
rect 40788 326708 40794 326710
rect 41781 326707 41847 326710
rect 42609 326498 42675 326501
rect 42977 326498 43043 326501
rect 42609 326496 43043 326498
rect 42609 326440 42614 326496
rect 42670 326440 42982 326496
rect 43038 326440 43043 326496
rect 42609 326438 43043 326440
rect 42609 326435 42675 326438
rect 42977 326435 43043 326438
rect 673545 325682 673611 325685
rect 675109 325682 675175 325685
rect 673545 325680 675175 325682
rect 673545 325624 673550 325680
rect 673606 325624 675114 325680
rect 675170 325624 675175 325680
rect 673545 325622 675175 325624
rect 673545 325619 673611 325622
rect 675109 325619 675175 325622
rect 40902 325348 40908 325412
rect 40972 325410 40978 325412
rect 41781 325410 41847 325413
rect 40972 325408 41847 325410
rect 40972 325352 41786 325408
rect 41842 325352 41847 325408
rect 40972 325350 41847 325352
rect 40972 325348 40978 325350
rect 41781 325347 41847 325350
rect 651465 325002 651531 325005
rect 650164 325000 651531 325002
rect 650164 324944 651470 325000
rect 651526 324944 651531 325000
rect 650164 324942 651531 324944
rect 651465 324939 651531 324942
rect 41873 324732 41939 324733
rect 41822 324730 41828 324732
rect 41782 324670 41828 324730
rect 41892 324728 41939 324732
rect 41934 324672 41939 324728
rect 41822 324668 41828 324670
rect 41892 324668 41939 324672
rect 41873 324667 41939 324668
rect 62113 324186 62179 324189
rect 62113 324184 64492 324186
rect 62113 324128 62118 324184
rect 62174 324128 64492 324184
rect 62113 324126 64492 324128
rect 62113 324123 62179 324126
rect 42057 322826 42123 322829
rect 43253 322826 43319 322829
rect 42057 322824 43319 322826
rect 42057 322768 42062 322824
rect 42118 322768 43258 322824
rect 43314 322768 43319 322824
rect 42057 322766 43319 322768
rect 42057 322763 42123 322766
rect 43253 322763 43319 322766
rect 42425 321466 42491 321469
rect 53097 321466 53163 321469
rect 42425 321464 53163 321466
rect 42425 321408 42430 321464
rect 42486 321408 53102 321464
rect 53158 321408 53163 321464
rect 42425 321406 53163 321408
rect 42425 321403 42491 321406
rect 53097 321403 53163 321406
rect 40534 320996 40540 321060
rect 40604 321058 40610 321060
rect 41781 321058 41847 321061
rect 40604 321056 41847 321058
rect 40604 321000 41786 321056
rect 41842 321000 41847 321056
rect 40604 320998 41847 321000
rect 40604 320996 40610 320998
rect 41781 320995 41847 320998
rect 42425 319018 42491 319021
rect 46933 319018 46999 319021
rect 42425 319016 46999 319018
rect 42425 318960 42430 319016
rect 42486 318960 46938 319016
rect 46994 318960 46999 319016
rect 42425 318958 46999 318960
rect 42425 318955 42491 318958
rect 46933 318955 46999 318958
rect 42425 317386 42491 317389
rect 44173 317386 44239 317389
rect 42425 317384 44239 317386
rect 42425 317328 42430 317384
rect 42486 317328 44178 317384
rect 44234 317328 44239 317384
rect 42425 317326 44239 317328
rect 42425 317323 42491 317326
rect 44173 317323 44239 317326
rect 42425 316434 42491 316437
rect 43110 316434 43116 316436
rect 42425 316432 43116 316434
rect 42425 316376 42430 316432
rect 42486 316376 43116 316432
rect 42425 316374 43116 316376
rect 42425 316371 42491 316374
rect 43110 316372 43116 316374
rect 43180 316372 43186 316436
rect 42149 316026 42215 316029
rect 45461 316026 45527 316029
rect 42149 316024 45527 316026
rect 42149 315968 42154 316024
rect 42210 315968 45466 316024
rect 45522 315968 45527 316024
rect 42149 315966 45527 315968
rect 42149 315963 42215 315966
rect 45461 315963 45527 315966
rect 41781 315620 41847 315621
rect 41781 315616 41828 315620
rect 41892 315618 41898 315620
rect 41781 315560 41786 315616
rect 41781 315556 41828 315560
rect 41892 315558 41938 315618
rect 41892 315556 41898 315558
rect 41781 315555 41847 315556
rect 665817 315482 665883 315485
rect 676029 315482 676095 315485
rect 665817 315480 676095 315482
rect 665817 315424 665822 315480
rect 665878 315424 676034 315480
rect 676090 315424 676095 315480
rect 665817 315422 676095 315424
rect 665817 315419 665883 315422
rect 676029 315419 676095 315422
rect 42149 313714 42215 313717
rect 45645 313714 45711 313717
rect 42149 313712 45711 313714
rect 42149 313656 42154 313712
rect 42210 313656 45650 313712
rect 45706 313656 45711 313712
rect 42149 313654 45711 313656
rect 42149 313651 42215 313654
rect 45645 313651 45711 313654
rect 663750 313654 676292 313714
rect 661677 313578 661743 313581
rect 663750 313578 663810 313654
rect 661677 313576 663810 313578
rect 661677 313520 661682 313576
rect 661738 313520 663810 313576
rect 661677 313518 663810 313520
rect 661677 313515 661743 313518
rect 676029 313306 676095 313309
rect 676029 313304 676292 313306
rect 676029 313248 676034 313304
rect 676090 313248 676292 313304
rect 676029 313246 676292 313248
rect 676029 313243 676095 313246
rect 668577 312898 668643 312901
rect 668577 312896 676292 312898
rect 668577 312840 668582 312896
rect 668638 312840 676292 312896
rect 668577 312838 676292 312840
rect 668577 312835 668643 312838
rect 42425 312762 42491 312765
rect 42926 312762 42932 312764
rect 42425 312760 42932 312762
rect 42425 312704 42430 312760
rect 42486 312704 42932 312760
rect 42425 312702 42932 312704
rect 42425 312699 42491 312702
rect 42926 312700 42932 312702
rect 42996 312700 43002 312764
rect 41454 312564 41460 312628
rect 41524 312626 41530 312628
rect 41781 312626 41847 312629
rect 41524 312624 41847 312626
rect 41524 312568 41786 312624
rect 41842 312568 41847 312624
rect 41524 312566 41847 312568
rect 41524 312564 41530 312566
rect 41781 312563 41847 312566
rect 674649 312490 674715 312493
rect 674649 312488 676292 312490
rect 674649 312432 674654 312488
rect 674710 312432 676292 312488
rect 674649 312430 676292 312432
rect 674649 312427 674715 312430
rect 673913 312082 673979 312085
rect 673913 312080 676292 312082
rect 673913 312024 673918 312080
rect 673974 312024 676292 312080
rect 673913 312022 676292 312024
rect 673913 312019 673979 312022
rect 44214 311748 44220 311812
rect 44284 311810 44290 311812
rect 44725 311810 44791 311813
rect 651465 311810 651531 311813
rect 44284 311808 44791 311810
rect 44284 311752 44730 311808
rect 44786 311752 44791 311808
rect 44284 311750 44791 311752
rect 650164 311808 651531 311810
rect 650164 311752 651470 311808
rect 651526 311752 651531 311808
rect 650164 311750 651531 311752
rect 44284 311748 44290 311750
rect 44725 311747 44791 311750
rect 651465 311747 651531 311750
rect 674097 311674 674163 311677
rect 674097 311672 676292 311674
rect 674097 311616 674102 311672
rect 674158 311616 676292 311672
rect 674097 311614 676292 311616
rect 674097 311611 674163 311614
rect 44173 311538 44239 311541
rect 44398 311538 44404 311540
rect 44173 311536 44404 311538
rect 44173 311480 44178 311536
rect 44234 311480 44404 311536
rect 44173 311478 44404 311480
rect 44173 311475 44239 311478
rect 44398 311476 44404 311478
rect 44468 311476 44474 311540
rect 44541 311268 44607 311269
rect 44541 311266 44588 311268
rect 44496 311264 44588 311266
rect 44496 311208 44546 311264
rect 44496 311206 44588 311208
rect 44541 311204 44588 311206
rect 44652 311204 44658 311268
rect 672165 311266 672231 311269
rect 672165 311264 676292 311266
rect 672165 311208 672170 311264
rect 672226 311208 676292 311264
rect 672165 311206 676292 311208
rect 44541 311203 44607 311204
rect 672165 311203 672231 311206
rect 62113 311130 62179 311133
rect 62113 311128 64492 311130
rect 62113 311072 62118 311128
rect 62174 311072 64492 311128
rect 62113 311070 64492 311072
rect 62113 311067 62179 311070
rect 673177 310858 673243 310861
rect 673177 310856 676292 310858
rect 673177 310800 673182 310856
rect 673238 310800 676292 310856
rect 673177 310798 676292 310800
rect 673177 310795 673243 310798
rect 674189 310450 674255 310453
rect 674189 310448 676292 310450
rect 674189 310392 674194 310448
rect 674250 310392 676292 310448
rect 674189 310390 676292 310392
rect 674189 310387 674255 310390
rect 672533 310042 672599 310045
rect 672533 310040 676292 310042
rect 672533 309984 672538 310040
rect 672594 309984 676292 310040
rect 672533 309982 676292 309984
rect 672533 309979 672599 309982
rect 674557 309634 674623 309637
rect 674557 309632 676292 309634
rect 674557 309576 674562 309632
rect 674618 309576 676292 309632
rect 674557 309574 676292 309576
rect 674557 309571 674623 309574
rect 674833 309226 674899 309229
rect 674833 309224 676292 309226
rect 674833 309168 674838 309224
rect 674894 309168 676292 309224
rect 674833 309166 676292 309168
rect 674833 309163 674899 309166
rect 675702 308756 675708 308820
rect 675772 308818 675778 308820
rect 675772 308758 676292 308818
rect 675772 308756 675778 308758
rect 676029 308410 676095 308413
rect 676029 308408 676292 308410
rect 676029 308352 676034 308408
rect 676090 308352 676292 308408
rect 676029 308350 676292 308352
rect 676029 308347 676095 308350
rect 675150 307940 675156 308004
rect 675220 308002 675226 308004
rect 675220 307942 676292 308002
rect 675220 307940 675226 307942
rect 680997 307594 681063 307597
rect 680997 307592 681076 307594
rect 680997 307536 681002 307592
rect 681058 307536 681076 307592
rect 680997 307534 681076 307536
rect 680997 307531 681063 307534
rect 678237 307186 678303 307189
rect 678237 307184 678316 307186
rect 678237 307128 678242 307184
rect 678298 307128 678316 307184
rect 678237 307126 678316 307128
rect 678237 307123 678303 307126
rect 675886 306716 675892 306780
rect 675956 306778 675962 306780
rect 675956 306718 676292 306778
rect 675956 306716 675962 306718
rect 678973 306370 679039 306373
rect 678973 306368 679052 306370
rect 678973 306312 678978 306368
rect 679034 306312 679052 306368
rect 678973 306310 679052 306312
rect 678973 306307 679039 306310
rect 676397 305962 676463 305965
rect 676397 305960 676476 305962
rect 676397 305904 676402 305960
rect 676458 305904 676476 305960
rect 676397 305902 676476 305904
rect 676397 305899 676463 305902
rect 674373 305554 674439 305557
rect 674373 305552 676292 305554
rect 674373 305496 674378 305552
rect 674434 305496 676292 305552
rect 674373 305494 676292 305496
rect 674373 305491 674439 305494
rect 676581 305146 676647 305149
rect 676581 305144 676660 305146
rect 676581 305088 676586 305144
rect 676642 305088 676660 305144
rect 676581 305086 676660 305088
rect 676581 305083 676647 305086
rect 673361 304738 673427 304741
rect 673361 304736 676292 304738
rect 673361 304680 673366 304736
rect 673422 304680 676292 304736
rect 673361 304678 676292 304680
rect 673361 304675 673427 304678
rect 672993 304330 673059 304333
rect 672993 304328 676292 304330
rect 672993 304272 672998 304328
rect 673054 304272 676292 304328
rect 672993 304270 676292 304272
rect 672993 304267 673059 304270
rect 673729 303922 673795 303925
rect 673729 303920 676292 303922
rect 673729 303864 673734 303920
rect 673790 303864 676292 303920
rect 673729 303862 676292 303864
rect 673729 303859 673795 303862
rect 674833 303650 674899 303653
rect 675385 303650 675451 303653
rect 674833 303648 675451 303650
rect 674833 303592 674838 303648
rect 674894 303592 675390 303648
rect 675446 303592 675451 303648
rect 674833 303590 675451 303592
rect 674833 303587 674899 303590
rect 675385 303587 675451 303590
rect 676029 303514 676095 303517
rect 676029 303512 676292 303514
rect 676029 303456 676034 303512
rect 676090 303456 676292 303512
rect 676029 303454 676292 303456
rect 676029 303451 676095 303454
rect 41781 303106 41847 303109
rect 46381 303106 46447 303109
rect 41781 303104 46447 303106
rect 41781 303048 41786 303104
rect 41842 303048 46386 303104
rect 46442 303048 46447 303104
rect 41781 303046 46447 303048
rect 41781 303043 41847 303046
rect 46381 303043 46447 303046
rect 675886 302636 675892 302700
rect 675956 302698 675962 302700
rect 676262 302698 676322 303076
rect 675956 302668 676322 302698
rect 675956 302638 676292 302668
rect 675956 302636 675962 302638
rect 668301 302290 668367 302293
rect 668301 302288 676292 302290
rect 668301 302232 668306 302288
rect 668362 302232 676292 302288
rect 668301 302230 676292 302232
rect 668301 302227 668367 302230
rect 671981 302018 672047 302021
rect 676029 302018 676095 302021
rect 671981 302016 676095 302018
rect 671981 301960 671986 302016
rect 672042 301960 676034 302016
rect 676090 301960 676095 302016
rect 671981 301958 676095 301960
rect 671981 301955 672047 301958
rect 676029 301955 676095 301958
rect 675109 301748 675175 301749
rect 675109 301746 675156 301748
rect 675064 301744 675156 301746
rect 675064 301688 675114 301744
rect 675064 301686 675156 301688
rect 675109 301684 675156 301686
rect 675220 301684 675226 301748
rect 675109 301683 675175 301684
rect 676581 301612 676647 301613
rect 676581 301608 676628 301612
rect 676692 301610 676698 301612
rect 676581 301552 676586 301608
rect 676581 301548 676628 301552
rect 676692 301550 676738 301610
rect 676692 301548 676698 301550
rect 676581 301547 676647 301548
rect 676397 301476 676463 301477
rect 676397 301474 676444 301476
rect 676352 301472 676444 301474
rect 676352 301416 676402 301472
rect 676352 301414 676444 301416
rect 676397 301412 676444 301414
rect 676508 301412 676514 301476
rect 676397 301411 676463 301412
rect 51717 301338 51783 301341
rect 41492 301336 51783 301338
rect 41492 301280 51722 301336
rect 51778 301280 51783 301336
rect 41492 301278 51783 301280
rect 51717 301275 51783 301278
rect 41781 300930 41847 300933
rect 41492 300928 41847 300930
rect 41492 300872 41786 300928
rect 41842 300872 41847 300928
rect 41492 300870 41847 300872
rect 41781 300867 41847 300870
rect 47761 300522 47827 300525
rect 41492 300520 47827 300522
rect 41492 300464 47766 300520
rect 47822 300464 47827 300520
rect 41492 300462 47827 300464
rect 47761 300459 47827 300462
rect 44725 300114 44791 300117
rect 41492 300112 44791 300114
rect 41492 300056 44730 300112
rect 44786 300056 44791 300112
rect 41492 300054 44791 300056
rect 44725 300051 44791 300054
rect 44725 299706 44791 299709
rect 41492 299704 44791 299706
rect 41492 299648 44730 299704
rect 44786 299648 44791 299704
rect 41492 299646 44791 299648
rect 44725 299643 44791 299646
rect 44173 299298 44239 299301
rect 41492 299296 44239 299298
rect 41492 299240 44178 299296
rect 44234 299240 44239 299296
rect 41492 299238 44239 299240
rect 44173 299235 44239 299238
rect 44265 298890 44331 298893
rect 41492 298888 44331 298890
rect 41492 298832 44270 298888
rect 44326 298832 44331 298888
rect 41492 298830 44331 298832
rect 44265 298827 44331 298830
rect 44541 298482 44607 298485
rect 652201 298482 652267 298485
rect 41492 298480 44607 298482
rect 41492 298424 44546 298480
rect 44602 298424 44607 298480
rect 41492 298422 44607 298424
rect 650164 298480 652267 298482
rect 650164 298424 652206 298480
rect 652262 298424 652267 298480
rect 650164 298422 652267 298424
rect 44541 298419 44607 298422
rect 652201 298419 652267 298422
rect 62113 298210 62179 298213
rect 62113 298208 64492 298210
rect 62113 298152 62118 298208
rect 62174 298152 64492 298208
rect 62113 298150 64492 298152
rect 62113 298147 62179 298150
rect 43253 298074 43319 298077
rect 41492 298072 43319 298074
rect 41492 298016 43258 298072
rect 43314 298016 43319 298072
rect 41492 298014 43319 298016
rect 43253 298011 43319 298014
rect 43662 297666 43668 297668
rect 41492 297606 43668 297666
rect 43662 297604 43668 297606
rect 43732 297604 43738 297668
rect 675702 297332 675708 297396
rect 675772 297394 675778 297396
rect 678237 297394 678303 297397
rect 675772 297392 678303 297394
rect 675772 297336 678242 297392
rect 678298 297336 678303 297392
rect 675772 297334 678303 297336
rect 675772 297332 675778 297334
rect 678237 297331 678303 297334
rect 42885 297258 42951 297261
rect 41492 297256 42951 297258
rect 41492 297200 42890 297256
rect 42946 297200 42951 297256
rect 41492 297198 42951 297200
rect 42885 297195 42951 297198
rect 41781 296850 41847 296853
rect 41492 296848 41847 296850
rect 41492 296792 41786 296848
rect 41842 296792 41847 296848
rect 41492 296790 41847 296792
rect 41781 296787 41847 296790
rect 674833 296850 674899 296853
rect 676121 296850 676187 296853
rect 674833 296848 676187 296850
rect 674833 296792 674838 296848
rect 674894 296792 676126 296848
rect 676182 296792 676187 296848
rect 674833 296790 676187 296792
rect 674833 296787 674899 296790
rect 676121 296787 676187 296790
rect 675017 296578 675083 296581
rect 675845 296578 675911 296581
rect 675017 296576 675911 296578
rect 675017 296520 675022 296576
rect 675078 296520 675850 296576
rect 675906 296520 675911 296576
rect 675017 296518 675911 296520
rect 675017 296515 675083 296518
rect 675845 296515 675911 296518
rect 42006 296442 42012 296444
rect 41492 296382 42012 296442
rect 42006 296380 42012 296382
rect 42076 296380 42082 296444
rect 675569 296306 675635 296309
rect 675526 296304 675635 296306
rect 675526 296248 675574 296304
rect 675630 296248 675635 296304
rect 675526 296243 675635 296248
rect 42057 296034 42123 296037
rect 41492 296032 42123 296034
rect 41492 295976 42062 296032
rect 42118 295976 42123 296032
rect 41492 295974 42123 295976
rect 42057 295971 42123 295974
rect 675526 295901 675586 296243
rect 675477 295896 675586 295901
rect 675477 295840 675482 295896
rect 675538 295840 675586 295896
rect 675477 295838 675586 295840
rect 675477 295835 675543 295838
rect 41822 295626 41828 295628
rect 41492 295566 41828 295626
rect 41822 295564 41828 295566
rect 41892 295564 41898 295628
rect 45001 295218 45067 295221
rect 41492 295216 45067 295218
rect 41492 295160 45006 295216
rect 45062 295160 45067 295216
rect 41492 295158 45067 295160
rect 45001 295155 45067 295158
rect 675753 295218 675819 295221
rect 676254 295218 676260 295220
rect 675753 295216 676260 295218
rect 675753 295160 675758 295216
rect 675814 295160 676260 295216
rect 675753 295158 676260 295160
rect 675753 295155 675819 295158
rect 676254 295156 676260 295158
rect 676324 295156 676330 295220
rect 32397 294810 32463 294813
rect 32397 294808 32476 294810
rect 32397 294752 32402 294808
rect 32458 294752 32476 294808
rect 32397 294750 32476 294752
rect 32397 294747 32463 294750
rect 43437 294402 43503 294405
rect 41492 294400 43503 294402
rect 41492 294344 43442 294400
rect 43498 294344 43503 294400
rect 41492 294342 43503 294344
rect 43437 294339 43503 294342
rect 45185 293994 45251 293997
rect 41492 293992 45251 293994
rect 41492 293936 45190 293992
rect 45246 293936 45251 293992
rect 41492 293934 45251 293936
rect 45185 293931 45251 293934
rect 43069 293586 43135 293589
rect 41492 293584 43135 293586
rect 41492 293528 43074 293584
rect 43130 293528 43135 293584
rect 41492 293526 43135 293528
rect 43069 293523 43135 293526
rect 43621 293178 43687 293181
rect 41492 293176 43687 293178
rect 41492 293120 43626 293176
rect 43682 293120 43687 293176
rect 41492 293118 43687 293120
rect 43621 293115 43687 293118
rect 41781 292772 41847 292773
rect 41781 292768 41828 292772
rect 41892 292770 41898 292772
rect 40726 292592 40786 292740
rect 41781 292712 41786 292768
rect 41781 292708 41828 292712
rect 41892 292710 41938 292770
rect 41892 292708 41898 292710
rect 41781 292707 41847 292708
rect 674373 292634 674439 292637
rect 674373 292632 674482 292634
rect 40534 292528 40540 292592
rect 40604 292528 40610 292592
rect 40718 292528 40724 292592
rect 40788 292528 40794 292592
rect 674373 292576 674378 292632
rect 674434 292576 674482 292632
rect 674373 292571 674482 292576
rect 40542 292332 40602 292528
rect 41822 292300 41828 292364
rect 41892 292362 41898 292364
rect 42057 292362 42123 292365
rect 41892 292360 42123 292362
rect 41892 292304 42062 292360
rect 42118 292304 42123 292360
rect 41892 292302 42123 292304
rect 674422 292362 674482 292571
rect 674649 292362 674715 292365
rect 674422 292360 674715 292362
rect 674422 292304 674654 292360
rect 674710 292304 674715 292360
rect 674422 292302 674715 292304
rect 41892 292300 41898 292302
rect 42057 292299 42123 292302
rect 674649 292299 674715 292302
rect 43805 291954 43871 291957
rect 41492 291952 43871 291954
rect 41492 291896 43810 291952
rect 43866 291896 43871 291952
rect 41492 291894 43871 291896
rect 43805 291891 43871 291894
rect 44449 291546 44515 291549
rect 41492 291544 44515 291546
rect 41492 291488 44454 291544
rect 44510 291488 44515 291544
rect 41492 291486 44515 291488
rect 44449 291483 44515 291486
rect 675753 291546 675819 291549
rect 676438 291546 676444 291548
rect 675753 291544 676444 291546
rect 675753 291488 675758 291544
rect 675814 291488 676444 291544
rect 675753 291486 676444 291488
rect 675753 291483 675819 291486
rect 676438 291484 676444 291486
rect 676508 291484 676514 291548
rect 42241 291138 42307 291141
rect 41492 291136 42307 291138
rect 41492 291080 42246 291136
rect 42302 291080 42307 291136
rect 41492 291078 42307 291080
rect 42241 291075 42307 291078
rect 41492 290670 41890 290730
rect 41321 290322 41387 290325
rect 41308 290320 41387 290322
rect 41308 290264 41326 290320
rect 41382 290264 41387 290320
rect 41308 290262 41387 290264
rect 41321 290259 41387 290262
rect 41830 290186 41890 290670
rect 673361 290594 673427 290597
rect 675109 290594 675175 290597
rect 673361 290592 675175 290594
rect 673361 290536 673366 290592
rect 673422 290536 675114 290592
rect 675170 290536 675175 290592
rect 673361 290534 675175 290536
rect 673361 290531 673427 290534
rect 675109 290531 675175 290534
rect 42057 290458 42123 290461
rect 49141 290458 49207 290461
rect 42057 290456 49207 290458
rect 42057 290400 42062 290456
rect 42118 290400 49146 290456
rect 49202 290400 49207 290456
rect 42057 290398 49207 290400
rect 42057 290395 42123 290398
rect 49141 290395 49207 290398
rect 50337 290186 50403 290189
rect 41830 290184 50403 290186
rect 41830 290128 50342 290184
rect 50398 290128 50403 290184
rect 41830 290126 50403 290128
rect 50337 290123 50403 290126
rect 42057 289914 42123 289917
rect 41492 289912 42123 289914
rect 41492 289856 42062 289912
rect 42118 289856 42123 289912
rect 41492 289854 42123 289856
rect 42057 289851 42123 289854
rect 42241 289914 42307 289917
rect 51717 289914 51783 289917
rect 42241 289912 51783 289914
rect 42241 289856 42246 289912
rect 42302 289856 51722 289912
rect 51778 289856 51783 289912
rect 42241 289854 51783 289856
rect 42241 289851 42307 289854
rect 51717 289851 51783 289854
rect 672993 287874 673059 287877
rect 675109 287874 675175 287877
rect 672993 287872 675175 287874
rect 672993 287816 672998 287872
rect 673054 287816 675114 287872
rect 675170 287816 675175 287872
rect 672993 287814 675175 287816
rect 672993 287811 673059 287814
rect 675109 287811 675175 287814
rect 675753 287058 675819 287061
rect 676622 287058 676628 287060
rect 675753 287056 676628 287058
rect 675753 287000 675758 287056
rect 675814 287000 676628 287056
rect 675753 286998 676628 287000
rect 675753 286995 675819 286998
rect 676622 286996 676628 286998
rect 676692 286996 676698 287060
rect 673729 286514 673795 286517
rect 675385 286514 675451 286517
rect 673729 286512 675451 286514
rect 673729 286456 673734 286512
rect 673790 286456 675390 286512
rect 675446 286456 675451 286512
rect 673729 286454 675451 286456
rect 673729 286451 673795 286454
rect 675385 286451 675451 286454
rect 651465 285290 651531 285293
rect 650164 285288 651531 285290
rect 650164 285232 651470 285288
rect 651526 285232 651531 285288
rect 650164 285230 651531 285232
rect 651465 285227 651531 285230
rect 62941 285154 63007 285157
rect 62941 285152 64492 285154
rect 62941 285096 62946 285152
rect 63002 285096 64492 285152
rect 62941 285094 64492 285096
rect 62941 285091 63007 285094
rect 675753 283658 675819 283661
rect 676070 283658 676076 283660
rect 675753 283656 676076 283658
rect 675753 283600 675758 283656
rect 675814 283600 676076 283656
rect 675753 283598 676076 283600
rect 675753 283595 675819 283598
rect 676070 283596 676076 283598
rect 676140 283596 676146 283660
rect 675661 282842 675727 282845
rect 675886 282842 675892 282844
rect 675661 282840 675892 282842
rect 675661 282784 675666 282840
rect 675722 282784 675892 282840
rect 675661 282782 675892 282784
rect 675661 282779 675727 282782
rect 675886 282780 675892 282782
rect 675956 282780 675962 282844
rect 675661 281620 675727 281621
rect 675661 281616 675708 281620
rect 675772 281618 675778 281620
rect 675661 281560 675666 281616
rect 675661 281556 675708 281560
rect 675772 281558 675818 281618
rect 675772 281556 675778 281558
rect 675661 281555 675727 281556
rect 41965 281484 42031 281485
rect 41965 281480 42012 281484
rect 42076 281482 42082 281484
rect 41965 281424 41970 281480
rect 41965 281420 42012 281424
rect 42076 281422 42122 281482
rect 42076 281420 42082 281422
rect 41965 281419 42031 281420
rect 42149 279850 42215 279853
rect 43621 279850 43687 279853
rect 42149 279848 43687 279850
rect 42149 279792 42154 279848
rect 42210 279792 43626 279848
rect 43682 279792 43687 279848
rect 42149 279790 43687 279792
rect 42149 279787 42215 279790
rect 43621 279787 43687 279790
rect 42425 278762 42491 278765
rect 55857 278762 55923 278765
rect 42425 278760 55923 278762
rect 42425 278704 42430 278760
rect 42486 278704 55862 278760
rect 55918 278704 55923 278760
rect 42425 278702 55923 278704
rect 42425 278699 42491 278702
rect 55857 278699 55923 278702
rect 42425 278218 42491 278221
rect 44449 278218 44515 278221
rect 42425 278216 44515 278218
rect 42425 278160 42430 278216
rect 42486 278160 44454 278216
rect 44510 278160 44515 278216
rect 42425 278158 44515 278160
rect 42425 278155 42491 278158
rect 44449 278155 44515 278158
rect 40718 277884 40724 277948
rect 40788 277946 40794 277948
rect 41781 277946 41847 277949
rect 40788 277944 41847 277946
rect 40788 277888 41786 277944
rect 41842 277888 41847 277944
rect 40788 277886 41847 277888
rect 40788 277884 40794 277886
rect 41781 277883 41847 277886
rect 40902 277612 40908 277676
rect 40972 277674 40978 277676
rect 42333 277674 42399 277677
rect 40972 277672 42399 277674
rect 40972 277616 42338 277672
rect 42394 277616 42399 277672
rect 40972 277614 42399 277616
rect 40972 277612 40978 277614
rect 42333 277611 42399 277614
rect 42057 277130 42123 277133
rect 43805 277130 43871 277133
rect 42057 277128 43871 277130
rect 42057 277072 42062 277128
rect 42118 277072 43810 277128
rect 43866 277072 43871 277128
rect 42057 277070 43871 277072
rect 42057 277067 42123 277070
rect 43805 277067 43871 277070
rect 42057 276586 42123 276589
rect 45001 276586 45067 276589
rect 42057 276584 45067 276586
rect 42057 276528 42062 276584
rect 42118 276528 45006 276584
rect 45062 276528 45067 276584
rect 42057 276526 45067 276528
rect 42057 276523 42123 276526
rect 45001 276523 45067 276526
rect 525793 275770 525859 275773
rect 530853 275770 530919 275773
rect 525793 275768 530919 275770
rect 525793 275712 525798 275768
rect 525854 275712 530858 275768
rect 530914 275712 530919 275768
rect 525793 275710 530919 275712
rect 525793 275707 525859 275710
rect 530853 275707 530919 275710
rect 536833 275634 536899 275637
rect 537937 275634 538003 275637
rect 536833 275632 538003 275634
rect 536833 275576 536838 275632
rect 536894 275576 537942 275632
rect 537998 275576 538003 275632
rect 536833 275574 538003 275576
rect 536833 275571 536899 275574
rect 537937 275571 538003 275574
rect 535085 275362 535151 275365
rect 538673 275362 538739 275365
rect 535085 275360 538739 275362
rect 535085 275304 535090 275360
rect 535146 275304 538678 275360
rect 538734 275304 538739 275360
rect 535085 275302 538739 275304
rect 535085 275299 535151 275302
rect 538673 275299 538739 275302
rect 538673 274954 538739 274957
rect 541157 274954 541223 274957
rect 538673 274952 541223 274954
rect 538673 274896 538678 274952
rect 538734 274896 541162 274952
rect 541218 274896 541223 274952
rect 538673 274894 541223 274896
rect 538673 274891 538739 274894
rect 541157 274891 541223 274894
rect 527817 274682 527883 274685
rect 543181 274682 543247 274685
rect 527817 274680 543247 274682
rect 527817 274624 527822 274680
rect 527878 274624 543186 274680
rect 543242 274624 543247 274680
rect 527817 274622 543247 274624
rect 527817 274619 527883 274622
rect 543181 274619 543247 274622
rect 40534 274212 40540 274276
rect 40604 274274 40610 274276
rect 41781 274274 41847 274277
rect 40604 274272 41847 274274
rect 40604 274216 41786 274272
rect 41842 274216 41847 274272
rect 40604 274214 41847 274216
rect 40604 274212 40610 274214
rect 41781 274211 41847 274214
rect 516593 274138 516659 274141
rect 519721 274138 519787 274141
rect 516593 274136 519787 274138
rect 516593 274080 516598 274136
rect 516654 274080 519726 274136
rect 519782 274080 519787 274136
rect 516593 274078 519787 274080
rect 516593 274075 516659 274078
rect 519721 274075 519787 274078
rect 536741 273866 536807 273869
rect 635641 273866 635707 273869
rect 536741 273864 635707 273866
rect 536741 273808 536746 273864
rect 536802 273808 635646 273864
rect 635702 273808 635707 273864
rect 536741 273806 635707 273808
rect 536741 273803 536807 273806
rect 635641 273803 635707 273806
rect 521101 273730 521167 273733
rect 524229 273730 524295 273733
rect 521101 273728 524295 273730
rect 521101 273672 521106 273728
rect 521162 273672 524234 273728
rect 524290 273672 524295 273728
rect 521101 273670 524295 273672
rect 521101 273667 521167 273670
rect 524229 273667 524295 273670
rect 42057 273458 42123 273461
rect 43069 273458 43135 273461
rect 42057 273456 43135 273458
rect 42057 273400 42062 273456
rect 42118 273400 43074 273456
rect 43130 273400 43135 273456
rect 42057 273398 43135 273400
rect 42057 273395 42123 273398
rect 43069 273395 43135 273398
rect 42057 272914 42123 272917
rect 45185 272914 45251 272917
rect 42057 272912 45251 272914
rect 42057 272856 42062 272912
rect 42118 272856 45190 272912
rect 45246 272856 45251 272912
rect 42057 272854 45251 272856
rect 42057 272851 42123 272854
rect 45185 272851 45251 272854
rect 534073 272778 534139 272781
rect 544837 272778 544903 272781
rect 534073 272776 544903 272778
rect 534073 272720 534078 272776
rect 534134 272720 544842 272776
rect 544898 272720 544903 272776
rect 534073 272718 544903 272720
rect 534073 272715 534139 272718
rect 544837 272715 544903 272718
rect 521469 272506 521535 272509
rect 524873 272506 524939 272509
rect 521469 272504 524939 272506
rect 521469 272448 521474 272504
rect 521530 272448 524878 272504
rect 524934 272448 524939 272504
rect 521469 272446 524939 272448
rect 521469 272443 521535 272446
rect 524873 272443 524939 272446
rect 533521 272506 533587 272509
rect 534165 272506 534231 272509
rect 533521 272504 534231 272506
rect 533521 272448 533526 272504
rect 533582 272448 534170 272504
rect 534226 272448 534231 272504
rect 533521 272446 534231 272448
rect 533521 272443 533587 272446
rect 534165 272443 534231 272446
rect 542997 272506 543063 272509
rect 645117 272506 645183 272509
rect 542997 272504 645183 272506
rect 542997 272448 543002 272504
rect 543058 272448 645122 272504
rect 645178 272448 645183 272504
rect 542997 272446 645183 272448
rect 542997 272443 543063 272446
rect 645117 272443 645183 272446
rect 513189 272370 513255 272373
rect 518433 272370 518499 272373
rect 513189 272368 518499 272370
rect 513189 272312 513194 272368
rect 513250 272312 518438 272368
rect 518494 272312 518499 272368
rect 513189 272310 518499 272312
rect 513189 272307 513255 272310
rect 518433 272307 518499 272310
rect 524597 272234 524663 272237
rect 531497 272234 531563 272237
rect 524597 272232 531563 272234
rect 524597 272176 524602 272232
rect 524658 272176 531502 272232
rect 531558 272176 531563 272232
rect 524597 272174 531563 272176
rect 524597 272171 524663 272174
rect 531497 272171 531563 272174
rect 523953 271690 524019 271693
rect 524781 271690 524847 271693
rect 523953 271688 524847 271690
rect 523953 271632 523958 271688
rect 524014 271632 524786 271688
rect 524842 271632 524847 271688
rect 523953 271630 524847 271632
rect 523953 271627 524019 271630
rect 524781 271627 524847 271630
rect 543549 271554 543615 271557
rect 546217 271554 546283 271557
rect 543549 271552 546283 271554
rect 543549 271496 543554 271552
rect 543610 271496 546222 271552
rect 546278 271496 546283 271552
rect 543549 271494 546283 271496
rect 543549 271491 543615 271494
rect 546217 271491 546283 271494
rect 511717 271418 511783 271421
rect 515305 271418 515371 271421
rect 511717 271416 515371 271418
rect 511717 271360 511722 271416
rect 511778 271360 515310 271416
rect 515366 271360 515371 271416
rect 511717 271358 515371 271360
rect 511717 271355 511783 271358
rect 515305 271355 515371 271358
rect 526253 271146 526319 271149
rect 529565 271146 529631 271149
rect 526253 271144 529631 271146
rect 526253 271088 526258 271144
rect 526314 271088 529570 271144
rect 529626 271088 529631 271144
rect 526253 271086 529631 271088
rect 526253 271083 526319 271086
rect 529565 271083 529631 271086
rect 529749 271146 529815 271149
rect 625061 271146 625127 271149
rect 529749 271144 625127 271146
rect 529749 271088 529754 271144
rect 529810 271088 625066 271144
rect 625122 271088 625127 271144
rect 529749 271086 625127 271088
rect 529749 271083 529815 271086
rect 625061 271083 625127 271086
rect 664437 271146 664503 271149
rect 683113 271146 683179 271149
rect 664437 271144 683179 271146
rect 664437 271088 664442 271144
rect 664498 271088 683118 271144
rect 683174 271088 683179 271144
rect 664437 271086 683179 271088
rect 664437 271083 664503 271086
rect 683113 271083 683179 271086
rect 523953 270874 524019 270877
rect 524873 270874 524939 270877
rect 523953 270872 524939 270874
rect 523953 270816 523958 270872
rect 524014 270816 524878 270872
rect 524934 270816 524939 270872
rect 523953 270814 524939 270816
rect 523953 270811 524019 270814
rect 524873 270811 524939 270814
rect 533889 270874 533955 270877
rect 534349 270874 534415 270877
rect 533889 270872 534415 270874
rect 533889 270816 533894 270872
rect 533950 270816 534354 270872
rect 534410 270816 534415 270872
rect 533889 270814 534415 270816
rect 533889 270811 533955 270814
rect 534349 270811 534415 270814
rect 528645 270738 528711 270741
rect 533153 270738 533219 270741
rect 528645 270736 533219 270738
rect 528645 270680 528650 270736
rect 528706 270680 533158 270736
rect 533214 270680 533219 270736
rect 528645 270678 533219 270680
rect 528645 270675 528711 270678
rect 533153 270675 533219 270678
rect 552197 270738 552263 270741
rect 553393 270738 553459 270741
rect 552197 270736 553459 270738
rect 552197 270680 552202 270736
rect 552258 270680 553398 270736
rect 553454 270680 553459 270736
rect 552197 270678 553459 270680
rect 552197 270675 552263 270678
rect 553393 270675 553459 270678
rect 504173 270602 504239 270605
rect 507853 270602 507919 270605
rect 504173 270600 507919 270602
rect 504173 270544 504178 270600
rect 504234 270544 507858 270600
rect 507914 270544 507919 270600
rect 504173 270542 507919 270544
rect 504173 270539 504239 270542
rect 507853 270539 507919 270542
rect 539501 270602 539567 270605
rect 543549 270602 543615 270605
rect 539501 270600 543615 270602
rect 539501 270544 539506 270600
rect 539562 270544 543554 270600
rect 543610 270544 543615 270600
rect 539501 270542 543615 270544
rect 539501 270539 539567 270542
rect 543549 270539 543615 270542
rect 41454 270404 41460 270468
rect 41524 270466 41530 270468
rect 41781 270466 41847 270469
rect 41524 270464 41847 270466
rect 41524 270408 41786 270464
rect 41842 270408 41847 270464
rect 41524 270406 41847 270408
rect 41524 270404 41530 270406
rect 41781 270403 41847 270406
rect 42425 270466 42491 270469
rect 43437 270466 43503 270469
rect 42425 270464 43503 270466
rect 42425 270408 42430 270464
rect 42486 270408 43442 270464
rect 43498 270408 43503 270464
rect 42425 270406 43503 270408
rect 42425 270403 42491 270406
rect 43437 270403 43503 270406
rect 494329 270330 494395 270333
rect 494881 270330 494947 270333
rect 574461 270330 574527 270333
rect 494329 270328 494947 270330
rect 494329 270272 494334 270328
rect 494390 270272 494886 270328
rect 494942 270272 494947 270328
rect 494329 270270 494947 270272
rect 494329 270267 494395 270270
rect 494881 270267 494947 270270
rect 499530 270328 574527 270330
rect 499530 270272 574466 270328
rect 574522 270272 574527 270328
rect 499530 270270 574527 270272
rect 494145 270058 494211 270061
rect 499530 270058 499590 270270
rect 574461 270267 574527 270270
rect 494145 270056 499590 270058
rect 494145 270000 494150 270056
rect 494206 270000 499590 270056
rect 494145 269998 499590 270000
rect 531405 270058 531471 270061
rect 627913 270058 627979 270061
rect 531405 270056 627979 270058
rect 531405 270000 531410 270056
rect 531466 270000 627918 270056
rect 627974 270000 627979 270056
rect 531405 269998 627979 270000
rect 494145 269995 494211 269998
rect 531405 269995 531471 269998
rect 627913 269995 627979 269998
rect 136541 269786 136607 269789
rect 139945 269786 140011 269789
rect 136541 269784 140011 269786
rect 136541 269728 136546 269784
rect 136602 269728 139950 269784
rect 140006 269728 140011 269784
rect 136541 269726 140011 269728
rect 136541 269723 136607 269726
rect 139945 269723 140011 269726
rect 509877 269786 509943 269789
rect 523309 269786 523375 269789
rect 509877 269784 523375 269786
rect 509877 269728 509882 269784
rect 509938 269728 523314 269784
rect 523370 269728 523375 269784
rect 509877 269726 523375 269728
rect 509877 269723 509943 269726
rect 523309 269723 523375 269726
rect 532877 269786 532943 269789
rect 533889 269786 533955 269789
rect 532877 269784 533955 269786
rect 532877 269728 532882 269784
rect 532938 269728 533894 269784
rect 533950 269728 533955 269784
rect 532877 269726 533955 269728
rect 532877 269723 532943 269726
rect 533889 269723 533955 269726
rect 538121 269786 538187 269789
rect 637573 269786 637639 269789
rect 538121 269784 637639 269786
rect 538121 269728 538126 269784
rect 538182 269728 637578 269784
rect 637634 269728 637639 269784
rect 538121 269726 637639 269728
rect 538121 269723 538187 269726
rect 637573 269723 637639 269726
rect 671337 269786 671403 269789
rect 676029 269786 676095 269789
rect 671337 269784 676095 269786
rect 671337 269728 671342 269784
rect 671398 269728 676034 269784
rect 676090 269728 676095 269784
rect 671337 269726 676095 269728
rect 671337 269723 671403 269726
rect 676029 269723 676095 269726
rect 502333 269650 502399 269653
rect 504541 269650 504607 269653
rect 502333 269648 504607 269650
rect 502333 269592 502338 269648
rect 502394 269592 504546 269648
rect 504602 269592 504607 269648
rect 502333 269590 504607 269592
rect 502333 269587 502399 269590
rect 504541 269587 504607 269590
rect 521653 269514 521719 269517
rect 532693 269514 532759 269517
rect 521653 269512 532759 269514
rect 521653 269456 521658 269512
rect 521714 269456 532698 269512
rect 532754 269456 532759 269512
rect 521653 269454 532759 269456
rect 521653 269451 521719 269454
rect 532693 269451 532759 269454
rect 535913 269514 535979 269517
rect 541985 269514 542051 269517
rect 535913 269512 542051 269514
rect 535913 269456 535918 269512
rect 535974 269456 541990 269512
rect 542046 269456 542051 269512
rect 535913 269454 542051 269456
rect 535913 269451 535979 269454
rect 541985 269451 542051 269454
rect 537017 269242 537083 269245
rect 538673 269242 538739 269245
rect 537017 269240 538739 269242
rect 537017 269184 537022 269240
rect 537078 269184 538678 269240
rect 538734 269184 538739 269240
rect 537017 269182 538739 269184
rect 537017 269179 537083 269182
rect 538673 269179 538739 269182
rect 41781 269108 41847 269109
rect 41781 269104 41828 269108
rect 41892 269106 41898 269108
rect 41781 269048 41786 269104
rect 41781 269044 41828 269048
rect 41892 269046 41938 269106
rect 41892 269044 41898 269046
rect 41781 269043 41847 269044
rect 525517 268698 525583 268701
rect 533889 268698 533955 268701
rect 525517 268696 533955 268698
rect 525517 268640 525522 268696
rect 525578 268640 533894 268696
rect 533950 268640 533955 268696
rect 525517 268638 533955 268640
rect 525517 268635 525583 268638
rect 533889 268635 533955 268638
rect 518433 268562 518499 268565
rect 518985 268562 519051 268565
rect 676262 268562 676322 268668
rect 518433 268560 519051 268562
rect 518433 268504 518438 268560
rect 518494 268504 518990 268560
rect 519046 268504 519051 268560
rect 518433 268502 519051 268504
rect 518433 268499 518499 268502
rect 518985 268499 519051 268502
rect 663750 268502 676322 268562
rect 519169 268426 519235 268429
rect 520457 268426 520523 268429
rect 519169 268424 520523 268426
rect 519169 268368 519174 268424
rect 519230 268368 520462 268424
rect 520518 268368 520523 268424
rect 519169 268366 520523 268368
rect 519169 268363 519235 268366
rect 520457 268363 520523 268366
rect 547505 268426 547571 268429
rect 549253 268426 549319 268429
rect 547505 268424 549319 268426
rect 547505 268368 547510 268424
rect 547566 268368 549258 268424
rect 549314 268368 549319 268424
rect 547505 268366 549319 268368
rect 547505 268363 547571 268366
rect 549253 268363 549319 268366
rect 539225 268154 539291 268157
rect 547689 268154 547755 268157
rect 539225 268152 547755 268154
rect 539225 268096 539230 268152
rect 539286 268096 547694 268152
rect 547750 268096 547755 268152
rect 539225 268094 547755 268096
rect 539225 268091 539291 268094
rect 547689 268091 547755 268094
rect 663057 268154 663123 268157
rect 663750 268154 663810 268502
rect 676029 268290 676095 268293
rect 676029 268288 676292 268290
rect 676029 268232 676034 268288
rect 676090 268232 676292 268288
rect 676029 268230 676292 268232
rect 676029 268227 676095 268230
rect 683113 268154 683179 268157
rect 663057 268152 663810 268154
rect 663057 268096 663062 268152
rect 663118 268096 663810 268152
rect 663057 268094 663810 268096
rect 683070 268152 683179 268154
rect 683070 268096 683118 268152
rect 683174 268096 683179 268152
rect 663057 268091 663123 268094
rect 683070 268091 683179 268096
rect 683070 267852 683130 268091
rect 533889 267746 533955 267749
rect 535453 267746 535519 267749
rect 533889 267744 535519 267746
rect 533889 267688 533894 267744
rect 533950 267688 535458 267744
rect 535514 267688 535519 267744
rect 533889 267686 535519 267688
rect 533889 267683 533955 267686
rect 535453 267683 535519 267686
rect 537569 267610 537635 267613
rect 543549 267610 543615 267613
rect 537569 267608 543615 267610
rect 537569 267552 537574 267608
rect 537630 267552 543554 267608
rect 543610 267552 543615 267608
rect 537569 267550 543615 267552
rect 537569 267547 537635 267550
rect 543549 267547 543615 267550
rect 673913 267474 673979 267477
rect 673913 267472 676292 267474
rect 673913 267416 673918 267472
rect 673974 267416 676292 267472
rect 673913 267414 676292 267416
rect 673913 267411 673979 267414
rect 518893 267338 518959 267341
rect 527173 267338 527239 267341
rect 518893 267336 527239 267338
rect 518893 267280 518898 267336
rect 518954 267280 527178 267336
rect 527234 267280 527239 267336
rect 518893 267278 527239 267280
rect 518893 267275 518959 267278
rect 527173 267275 527239 267278
rect 527633 267338 527699 267341
rect 533705 267338 533771 267341
rect 527633 267336 533771 267338
rect 527633 267280 527638 267336
rect 527694 267280 533710 267336
rect 533766 267280 533771 267336
rect 527633 267278 533771 267280
rect 527633 267275 527699 267278
rect 533705 267275 533771 267278
rect 542169 267338 542235 267341
rect 607857 267338 607923 267341
rect 542169 267336 607923 267338
rect 542169 267280 542174 267336
rect 542230 267280 607862 267336
rect 607918 267280 607923 267336
rect 542169 267278 607923 267280
rect 542169 267275 542235 267278
rect 607857 267275 607923 267278
rect 499757 267202 499823 267205
rect 501045 267202 501111 267205
rect 499757 267200 501111 267202
rect 499757 267144 499762 267200
rect 499818 267144 501050 267200
rect 501106 267144 501111 267200
rect 499757 267142 501111 267144
rect 499757 267139 499823 267142
rect 501045 267139 501111 267142
rect 506197 267202 506263 267205
rect 507853 267202 507919 267205
rect 506197 267200 507919 267202
rect 506197 267144 506202 267200
rect 506258 267144 507858 267200
rect 507914 267144 507919 267200
rect 506197 267142 507919 267144
rect 506197 267139 506263 267142
rect 507853 267139 507919 267142
rect 533889 267202 533955 267205
rect 534165 267202 534231 267205
rect 533889 267200 534231 267202
rect 533889 267144 533894 267200
rect 533950 267144 534170 267200
rect 534226 267144 534231 267200
rect 533889 267142 534231 267144
rect 533889 267139 533955 267142
rect 534165 267139 534231 267142
rect 40677 267066 40743 267069
rect 62757 267066 62823 267069
rect 40677 267064 62823 267066
rect 40677 267008 40682 267064
rect 40738 267008 62762 267064
rect 62818 267008 62823 267064
rect 40677 267006 62823 267008
rect 40677 267003 40743 267006
rect 62757 267003 62823 267006
rect 524505 267066 524571 267069
rect 525885 267066 525951 267069
rect 629293 267066 629359 267069
rect 524505 267064 525951 267066
rect 524505 267008 524510 267064
rect 524566 267008 525890 267064
rect 525946 267008 525951 267064
rect 524505 267006 525951 267008
rect 524505 267003 524571 267006
rect 525885 267003 525951 267006
rect 547830 267064 629359 267066
rect 547830 267008 629298 267064
rect 629354 267008 629359 267064
rect 547830 267006 629359 267008
rect 532233 266930 532299 266933
rect 547830 266930 547890 267006
rect 629293 267003 629359 267006
rect 674649 267066 674715 267069
rect 674649 267064 676292 267066
rect 674649 267008 674654 267064
rect 674710 267008 676292 267064
rect 674649 267006 676292 267008
rect 674649 267003 674715 267006
rect 532233 266928 547890 266930
rect 532233 266872 532238 266928
rect 532294 266872 547890 266928
rect 532233 266870 547890 266872
rect 532233 266867 532299 266870
rect 518709 266794 518775 266797
rect 518893 266794 518959 266797
rect 518709 266792 518994 266794
rect 518709 266736 518714 266792
rect 518770 266736 518898 266792
rect 518954 266736 518994 266792
rect 518709 266734 518994 266736
rect 518709 266731 518775 266734
rect 518893 266731 518959 266734
rect 473261 266658 473327 266661
rect 474825 266658 474891 266661
rect 473261 266656 474891 266658
rect 473261 266600 473266 266656
rect 473322 266600 474830 266656
rect 474886 266600 474891 266656
rect 473261 266598 474891 266600
rect 473261 266595 473327 266598
rect 474825 266595 474891 266598
rect 534073 266658 534139 266661
rect 537385 266658 537451 266661
rect 534073 266656 537451 266658
rect 534073 266600 534078 266656
rect 534134 266600 537390 266656
rect 537446 266600 537451 266656
rect 534073 266598 537451 266600
rect 534073 266595 534139 266598
rect 537385 266595 537451 266598
rect 672165 266522 672231 266525
rect 676262 266522 676322 266628
rect 672165 266520 676322 266522
rect 672165 266464 672170 266520
rect 672226 266464 676322 266520
rect 672165 266462 676322 266464
rect 672165 266459 672231 266462
rect 674005 266250 674071 266253
rect 674005 266248 676292 266250
rect 674005 266192 674010 266248
rect 674066 266192 676292 266248
rect 674005 266190 676292 266192
rect 674005 266187 674071 266190
rect 674189 265842 674255 265845
rect 674189 265840 676292 265842
rect 674189 265784 674194 265840
rect 674250 265784 676292 265840
rect 674189 265782 676292 265784
rect 674189 265779 674255 265782
rect 674281 265434 674347 265437
rect 674281 265432 676292 265434
rect 674281 265376 674286 265432
rect 674342 265376 676292 265432
rect 674281 265374 676292 265376
rect 674281 265371 674347 265374
rect 674465 265026 674531 265029
rect 674465 265024 676292 265026
rect 674465 264968 674470 265024
rect 674526 264968 676292 265024
rect 674465 264966 676292 264968
rect 674465 264963 674531 264966
rect 674833 264482 674899 264485
rect 676262 264482 676322 264588
rect 674833 264480 676322 264482
rect 674833 264424 674838 264480
rect 674894 264424 676322 264480
rect 674833 264422 676322 264424
rect 674833 264419 674899 264422
rect 676446 264077 676506 264180
rect 671337 264074 671403 264077
rect 671337 264072 676322 264074
rect 671337 264016 671342 264072
rect 671398 264016 676322 264072
rect 671337 264014 676322 264016
rect 676446 264072 676555 264077
rect 676446 264016 676494 264072
rect 676550 264016 676555 264072
rect 676446 264014 676555 264016
rect 671337 264011 671403 264014
rect 673085 263802 673151 263805
rect 674833 263802 674899 263805
rect 673085 263800 674899 263802
rect 673085 263744 673090 263800
rect 673146 263744 674838 263800
rect 674894 263744 674899 263800
rect 676262 263772 676322 264014
rect 676489 264011 676555 264014
rect 673085 263742 674899 263744
rect 673085 263739 673151 263742
rect 674833 263739 674899 263742
rect 674966 263604 674972 263668
rect 675036 263666 675042 263668
rect 676489 263666 676555 263669
rect 675036 263664 676555 263666
rect 675036 263608 676494 263664
rect 676550 263608 676555 263664
rect 675036 263606 676555 263608
rect 675036 263604 675042 263606
rect 676489 263603 676555 263606
rect 678286 263261 678346 263364
rect 678237 263256 678346 263261
rect 678237 263200 678242 263256
rect 678298 263200 678346 263256
rect 678237 263198 678346 263200
rect 678237 263195 678303 263198
rect 676262 262853 676322 262956
rect 676213 262848 676322 262853
rect 676213 262792 676218 262848
rect 676274 262792 676322 262848
rect 676213 262790 676322 262792
rect 676213 262787 676279 262790
rect 676070 262380 676076 262444
rect 676140 262442 676146 262444
rect 676262 262442 676322 262548
rect 676140 262382 676322 262442
rect 676140 262380 676146 262382
rect 554405 262170 554471 262173
rect 552460 262168 554471 262170
rect 552460 262112 554410 262168
rect 554466 262112 554471 262168
rect 552460 262110 554471 262112
rect 554405 262107 554471 262110
rect 671705 262034 671771 262037
rect 676262 262034 676322 262140
rect 671705 262032 676322 262034
rect 671705 261976 671710 262032
rect 671766 261976 676322 262032
rect 671705 261974 676322 261976
rect 671705 261971 671771 261974
rect 676998 261628 677058 261732
rect 676990 261564 676996 261628
rect 677060 261564 677066 261628
rect 678470 261221 678530 261324
rect 678421 261216 678530 261221
rect 678421 261160 678426 261216
rect 678482 261160 678530 261216
rect 678421 261158 678530 261160
rect 678421 261155 678487 261158
rect 674189 260946 674255 260949
rect 674189 260944 676292 260946
rect 674189 260888 674194 260944
rect 674250 260888 676292 260944
rect 674189 260886 676292 260888
rect 674189 260883 674255 260886
rect 673361 260402 673427 260405
rect 676262 260402 676322 260508
rect 673361 260400 676322 260402
rect 673361 260344 673366 260400
rect 673422 260344 676322 260400
rect 673361 260342 676322 260344
rect 673361 260339 673427 260342
rect 554313 259994 554379 259997
rect 676814 259996 676874 260100
rect 552460 259992 554379 259994
rect 552460 259936 554318 259992
rect 554374 259936 554379 259992
rect 552460 259934 554379 259936
rect 554313 259931 554379 259934
rect 676806 259932 676812 259996
rect 676876 259932 676882 259996
rect 673729 259722 673795 259725
rect 673729 259720 676292 259722
rect 673729 259664 673734 259720
rect 673790 259664 676292 259720
rect 673729 259662 676292 259664
rect 673729 259659 673795 259662
rect 672901 259178 672967 259181
rect 676262 259178 676322 259284
rect 672901 259176 676322 259178
rect 672901 259120 672906 259176
rect 672962 259120 676322 259176
rect 672901 259118 676322 259120
rect 672901 259115 672967 259118
rect 675937 258770 676003 258773
rect 676262 258770 676322 258876
rect 675937 258768 676322 258770
rect 675937 258712 675942 258768
rect 675998 258712 676322 258768
rect 675937 258710 676322 258712
rect 675937 258707 676003 258710
rect 673913 258498 673979 258501
rect 673913 258496 676292 258498
rect 673913 258440 673918 258496
rect 673974 258440 676292 258496
rect 673913 258438 676292 258440
rect 673913 258435 673979 258438
rect 675937 258226 676003 258229
rect 675894 258224 676003 258226
rect 675894 258168 675942 258224
rect 675998 258168 676003 258224
rect 675894 258163 676003 258168
rect 41492 258030 42074 258090
rect 42014 257954 42074 258030
rect 46197 257954 46263 257957
rect 42014 257952 46263 257954
rect 42014 257896 46202 257952
rect 46258 257896 46263 257952
rect 42014 257894 46263 257896
rect 46197 257891 46263 257894
rect 671521 257954 671587 257957
rect 675894 257954 675954 258163
rect 671521 257952 675954 257954
rect 671521 257896 671526 257952
rect 671582 257896 675954 257952
rect 671521 257894 675954 257896
rect 671521 257891 671587 257894
rect 553945 257818 554011 257821
rect 552460 257816 554011 257818
rect 552460 257760 553950 257816
rect 554006 257760 554011 257816
rect 552460 257758 554011 257760
rect 553945 257755 554011 257758
rect 41462 257546 41522 257652
rect 53281 257546 53347 257549
rect 41462 257544 53347 257546
rect 41462 257488 53286 257544
rect 53342 257488 53347 257544
rect 41462 257486 53347 257488
rect 53281 257483 53347 257486
rect 675293 257546 675359 257549
rect 676262 257546 676322 258060
rect 675293 257544 676322 257546
rect 675293 257488 675298 257544
rect 675354 257488 676322 257544
rect 675293 257486 676322 257488
rect 675293 257483 675359 257486
rect 35758 257141 35818 257244
rect 35758 257136 35867 257141
rect 35758 257080 35806 257136
rect 35862 257080 35867 257136
rect 35758 257078 35867 257080
rect 35801 257075 35867 257078
rect 673177 257138 673243 257141
rect 676262 257138 676322 257244
rect 673177 257136 676322 257138
rect 673177 257080 673182 257136
rect 673238 257080 676322 257136
rect 673177 257078 676322 257080
rect 673177 257075 673243 257078
rect 44633 256866 44699 256869
rect 41492 256864 44699 256866
rect 41492 256808 44638 256864
rect 44694 256808 44699 256864
rect 41492 256806 44699 256808
rect 44633 256803 44699 256806
rect 670417 256730 670483 256733
rect 675293 256730 675359 256733
rect 670417 256728 675359 256730
rect 670417 256672 670422 256728
rect 670478 256672 675298 256728
rect 675354 256672 675359 256728
rect 670417 256670 675359 256672
rect 670417 256667 670483 256670
rect 675293 256667 675359 256670
rect 43713 256458 43779 256461
rect 41492 256456 43779 256458
rect 41492 256400 43718 256456
rect 43774 256400 43779 256456
rect 41492 256398 43779 256400
rect 43713 256395 43779 256398
rect 44265 256050 44331 256053
rect 41492 256048 44331 256050
rect 41492 255992 44270 256048
rect 44326 255992 44331 256048
rect 41492 255990 44331 255992
rect 44265 255987 44331 255990
rect 43437 255642 43503 255645
rect 553669 255642 553735 255645
rect 41492 255640 43503 255642
rect 41492 255584 43442 255640
rect 43498 255584 43503 255640
rect 41492 255582 43503 255584
rect 552460 255640 553735 255642
rect 552460 255584 553674 255640
rect 553730 255584 553735 255640
rect 552460 255582 553735 255584
rect 43437 255579 43503 255582
rect 553669 255579 553735 255582
rect 43253 255234 43319 255237
rect 41492 255232 43319 255234
rect 41492 255176 43258 255232
rect 43314 255176 43319 255232
rect 41492 255174 43319 255176
rect 43253 255171 43319 255174
rect 42885 254826 42951 254829
rect 41492 254824 42951 254826
rect 41492 254768 42890 254824
rect 42946 254768 42951 254824
rect 41492 254766 42951 254768
rect 42885 254763 42951 254766
rect 43069 254418 43135 254421
rect 41492 254416 43135 254418
rect 41492 254360 43074 254416
rect 43130 254360 43135 254416
rect 41492 254358 43135 254360
rect 43069 254355 43135 254358
rect 44173 254010 44239 254013
rect 41492 254008 44239 254010
rect 41492 253952 44178 254008
rect 44234 253952 44239 254008
rect 41492 253950 44239 253952
rect 44173 253947 44239 253950
rect 35574 253469 35634 253572
rect 35574 253464 35683 253469
rect 554497 253466 554563 253469
rect 35574 253408 35622 253464
rect 35678 253408 35683 253464
rect 35574 253406 35683 253408
rect 552460 253464 554563 253466
rect 552460 253408 554502 253464
rect 554558 253408 554563 253464
rect 552460 253406 554563 253408
rect 35617 253403 35683 253406
rect 554497 253403 554563 253406
rect 35390 253061 35450 253164
rect 35390 253056 35499 253061
rect 35801 253058 35867 253061
rect 35390 253000 35438 253056
rect 35494 253000 35499 253056
rect 35390 252998 35499 253000
rect 35433 252995 35499 252998
rect 35758 253056 35867 253058
rect 35758 253000 35806 253056
rect 35862 253000 35867 253056
rect 35758 252995 35867 253000
rect 35758 252756 35818 252995
rect 35758 252245 35818 252348
rect 35758 252240 35867 252245
rect 35758 252184 35806 252240
rect 35862 252184 35867 252240
rect 35758 252182 35867 252184
rect 35801 252179 35867 252182
rect 44633 251970 44699 251973
rect 41492 251968 44699 251970
rect 41492 251912 44638 251968
rect 44694 251912 44699 251968
rect 41492 251910 44699 251912
rect 44633 251907 44699 251910
rect 674925 251562 674991 251565
rect 675845 251562 675911 251565
rect 674925 251560 675911 251562
rect 40542 251428 40602 251532
rect 674925 251504 674930 251560
rect 674986 251504 675850 251560
rect 675906 251504 675911 251560
rect 674925 251502 675911 251504
rect 674925 251499 674991 251502
rect 675845 251499 675911 251502
rect 40534 251364 40540 251428
rect 40604 251364 40610 251428
rect 553485 251290 553551 251293
rect 552460 251288 553551 251290
rect 552460 251232 553490 251288
rect 553546 251232 553551 251288
rect 552460 251230 553551 251232
rect 553485 251227 553551 251230
rect 43529 251154 43595 251157
rect 41492 251152 43595 251154
rect 41492 251096 43534 251152
rect 43590 251096 43595 251152
rect 41492 251094 43595 251096
rect 43529 251091 43595 251094
rect 45829 250746 45895 250749
rect 41492 250744 45895 250746
rect 41492 250688 45834 250744
rect 45890 250688 45895 250744
rect 41492 250686 45895 250688
rect 45829 250683 45895 250686
rect 45553 250338 45619 250341
rect 41492 250336 45619 250338
rect 41492 250280 45558 250336
rect 45614 250280 45619 250336
rect 41492 250278 45619 250280
rect 45553 250275 45619 250278
rect 675753 250338 675819 250341
rect 676990 250338 676996 250340
rect 675753 250336 676996 250338
rect 675753 250280 675758 250336
rect 675814 250280 676996 250336
rect 675753 250278 676996 250280
rect 675753 250275 675819 250278
rect 676990 250276 676996 250278
rect 677060 250276 677066 250340
rect 40726 249796 40786 249900
rect 40718 249732 40724 249796
rect 40788 249732 40794 249796
rect 674782 249596 674788 249660
rect 674852 249658 674858 249660
rect 675385 249658 675451 249661
rect 674852 249656 675451 249658
rect 674852 249600 675390 249656
rect 675446 249600 675451 249656
rect 674852 249598 675451 249600
rect 674852 249596 674858 249598
rect 675385 249595 675451 249598
rect 676070 249596 676076 249660
rect 676140 249596 676146 249660
rect 46013 249522 46079 249525
rect 41492 249520 46079 249522
rect 41492 249464 46018 249520
rect 46074 249464 46079 249520
rect 41492 249462 46079 249464
rect 46013 249459 46079 249462
rect 674925 249386 674991 249389
rect 676078 249386 676138 249596
rect 674925 249384 676138 249386
rect 674925 249328 674930 249384
rect 674986 249328 676138 249384
rect 674925 249326 676138 249328
rect 674925 249323 674991 249326
rect 43069 249114 43135 249117
rect 553853 249114 553919 249117
rect 41492 249112 43135 249114
rect 41492 249056 43074 249112
rect 43130 249056 43135 249112
rect 41492 249054 43135 249056
rect 552460 249112 553919 249114
rect 552460 249056 553858 249112
rect 553914 249056 553919 249112
rect 552460 249054 553919 249056
rect 43069 249051 43135 249054
rect 553853 249051 553919 249054
rect 44541 248706 44607 248709
rect 41492 248704 44607 248706
rect 41492 248648 44546 248704
rect 44602 248648 44607 248704
rect 41492 248646 44607 248648
rect 44541 248643 44607 248646
rect 44357 248298 44423 248301
rect 41492 248296 44423 248298
rect 41492 248240 44362 248296
rect 44418 248240 44423 248296
rect 41492 248238 44423 248240
rect 44357 248235 44423 248238
rect 46197 247890 46263 247893
rect 41492 247888 46263 247890
rect 41492 247832 46202 247888
rect 46258 247832 46263 247888
rect 41492 247830 46263 247832
rect 46197 247827 46263 247830
rect 47761 247482 47827 247485
rect 41492 247480 47827 247482
rect 41492 247424 47766 247480
rect 47822 247424 47827 247480
rect 41492 247422 47827 247424
rect 47761 247419 47827 247422
rect 46933 247074 46999 247077
rect 41492 247072 46999 247074
rect 41492 247016 46938 247072
rect 46994 247016 46999 247072
rect 41492 247014 46999 247016
rect 46933 247011 46999 247014
rect 554405 246938 554471 246941
rect 552460 246936 554471 246938
rect 552460 246880 554410 246936
rect 554466 246880 554471 246936
rect 552460 246878 554471 246880
rect 554405 246875 554471 246878
rect 674281 246938 674347 246941
rect 675109 246938 675175 246941
rect 674281 246936 675175 246938
rect 674281 246880 674286 246936
rect 674342 246880 675114 246936
rect 675170 246880 675175 246936
rect 674281 246878 675175 246880
rect 674281 246875 674347 246878
rect 675109 246875 675175 246878
rect 41462 246530 41522 246636
rect 50521 246530 50587 246533
rect 41462 246528 50587 246530
rect 41462 246472 50526 246528
rect 50582 246472 50587 246528
rect 41462 246470 50587 246472
rect 50521 246467 50587 246470
rect 673729 245578 673795 245581
rect 675109 245578 675175 245581
rect 673729 245576 675175 245578
rect 673729 245520 673734 245576
rect 673790 245520 675114 245576
rect 675170 245520 675175 245576
rect 673729 245518 675175 245520
rect 673729 245515 673795 245518
rect 675109 245515 675175 245518
rect 674833 245306 674899 245309
rect 676806 245306 676812 245308
rect 674833 245304 676812 245306
rect 674833 245248 674838 245304
rect 674894 245248 676812 245304
rect 674833 245246 676812 245248
rect 674833 245243 674899 245246
rect 676806 245244 676812 245246
rect 676876 245244 676882 245308
rect 673361 245034 673427 245037
rect 675150 245034 675156 245036
rect 673361 245032 675156 245034
rect 673361 244976 673366 245032
rect 673422 244976 675156 245032
rect 673361 244974 675156 244976
rect 673361 244971 673427 244974
rect 675150 244972 675156 244974
rect 675220 244972 675226 245036
rect 554497 244762 554563 244765
rect 552460 244760 554563 244762
rect 552460 244704 554502 244760
rect 554558 244704 554563 244760
rect 552460 244702 554563 244704
rect 554497 244699 554563 244702
rect 671705 244762 671771 244765
rect 675334 244762 675340 244764
rect 671705 244760 675340 244762
rect 671705 244704 671710 244760
rect 671766 244704 675340 244760
rect 671705 244702 675340 244704
rect 671705 244699 671771 244702
rect 675334 244700 675340 244702
rect 675404 244700 675410 244764
rect 41689 242858 41755 242861
rect 42701 242858 42767 242861
rect 41689 242856 42767 242858
rect 41689 242800 41694 242856
rect 41750 242800 42706 242856
rect 42762 242800 42767 242856
rect 41689 242798 42767 242800
rect 41689 242795 41755 242798
rect 42701 242795 42767 242798
rect 672809 242858 672875 242861
rect 675385 242858 675451 242861
rect 672809 242856 675451 242858
rect 672809 242800 672814 242856
rect 672870 242800 675390 242856
rect 675446 242800 675451 242856
rect 672809 242798 675451 242800
rect 672809 242795 672875 242798
rect 675385 242795 675451 242798
rect 40677 242586 40743 242589
rect 43253 242586 43319 242589
rect 553945 242586 554011 242589
rect 40677 242584 43319 242586
rect 40677 242528 40682 242584
rect 40738 242528 43258 242584
rect 43314 242528 43319 242584
rect 40677 242526 43319 242528
rect 552460 242584 554011 242586
rect 552460 242528 553950 242584
rect 554006 242528 554011 242584
rect 552460 242526 554011 242528
rect 40677 242523 40743 242526
rect 43253 242523 43319 242526
rect 553945 242523 554011 242526
rect 671521 241498 671587 241501
rect 675109 241498 675175 241501
rect 671521 241496 675175 241498
rect 671521 241440 671526 241496
rect 671582 241440 675114 241496
rect 675170 241440 675175 241496
rect 671521 241438 675175 241440
rect 671521 241435 671587 241438
rect 675109 241435 675175 241438
rect 553853 240410 553919 240413
rect 552460 240408 553919 240410
rect 552460 240352 553858 240408
rect 553914 240352 553919 240408
rect 552460 240350 553919 240352
rect 553853 240347 553919 240350
rect 675201 240276 675267 240277
rect 675150 240274 675156 240276
rect 675110 240214 675156 240274
rect 675220 240272 675267 240276
rect 675262 240216 675267 240272
rect 675150 240212 675156 240214
rect 675220 240212 675267 240216
rect 675201 240211 675267 240212
rect 40534 240076 40540 240140
rect 40604 240138 40610 240140
rect 41781 240138 41847 240141
rect 40604 240136 41847 240138
rect 40604 240080 41786 240136
rect 41842 240080 41847 240136
rect 40604 240078 41847 240080
rect 40604 240076 40610 240078
rect 41781 240075 41847 240078
rect 42057 238506 42123 238509
rect 46933 238506 46999 238509
rect 42057 238504 46999 238506
rect 42057 238448 42062 238504
rect 42118 238448 46938 238504
rect 46994 238448 46999 238504
rect 42057 238446 46999 238448
rect 42057 238443 42123 238446
rect 46933 238443 46999 238446
rect 554313 238234 554379 238237
rect 552460 238232 554379 238234
rect 552460 238176 554318 238232
rect 554374 238176 554379 238232
rect 552460 238174 554379 238176
rect 554313 238171 554379 238174
rect 671337 238234 671403 238237
rect 675109 238234 675175 238237
rect 671337 238232 675175 238234
rect 671337 238176 671342 238232
rect 671398 238176 675114 238232
rect 675170 238176 675175 238232
rect 671337 238174 675175 238176
rect 671337 238171 671403 238174
rect 675109 238171 675175 238174
rect 42006 237356 42012 237420
rect 42076 237418 42082 237420
rect 42517 237418 42583 237421
rect 42076 237416 42583 237418
rect 42076 237360 42522 237416
rect 42578 237360 42583 237416
rect 42076 237358 42583 237360
rect 42076 237356 42082 237358
rect 42517 237355 42583 237358
rect 672993 237418 673059 237421
rect 674833 237418 674899 237421
rect 672993 237416 674899 237418
rect 672993 237360 672998 237416
rect 673054 237360 674838 237416
rect 674894 237360 674899 237416
rect 672993 237358 674899 237360
rect 672993 237355 673059 237358
rect 674833 237355 674899 237358
rect 673297 237146 673363 237149
rect 674230 237146 674236 237148
rect 673297 237144 674236 237146
rect 673297 237088 673302 237144
rect 673358 237088 674236 237144
rect 673297 237086 674236 237088
rect 673297 237083 673363 237086
rect 674230 237084 674236 237086
rect 674300 237084 674306 237148
rect 675385 236876 675451 236877
rect 675334 236874 675340 236876
rect 675294 236814 675340 236874
rect 675404 236872 675451 236876
rect 675446 236816 675451 236872
rect 675334 236812 675340 236814
rect 675404 236812 675451 236816
rect 675385 236811 675451 236812
rect 668945 236738 669011 236741
rect 673521 236738 673587 236741
rect 668945 236736 673587 236738
rect 668945 236680 668950 236736
rect 669006 236680 673526 236736
rect 673582 236680 673587 236736
rect 668945 236678 673587 236680
rect 668945 236675 669011 236678
rect 673521 236675 673587 236678
rect 554497 236058 554563 236061
rect 552460 236056 554563 236058
rect 552460 236000 554502 236056
rect 554558 236000 554563 236056
rect 552460 235998 554563 236000
rect 554497 235995 554563 235998
rect 40718 235860 40724 235924
rect 40788 235922 40794 235924
rect 41781 235922 41847 235925
rect 40788 235920 41847 235922
rect 40788 235864 41786 235920
rect 41842 235864 41847 235920
rect 40788 235862 41847 235864
rect 40788 235860 40794 235862
rect 41781 235859 41847 235862
rect 42425 235922 42491 235925
rect 44357 235922 44423 235925
rect 42425 235920 44423 235922
rect 42425 235864 42430 235920
rect 42486 235864 44362 235920
rect 44418 235864 44423 235920
rect 42425 235862 44423 235864
rect 42425 235859 42491 235862
rect 44357 235859 44423 235862
rect 670417 235922 670483 235925
rect 675109 235922 675175 235925
rect 670417 235920 675175 235922
rect 670417 235864 670422 235920
rect 670478 235864 675114 235920
rect 675170 235864 675175 235920
rect 670417 235862 675175 235864
rect 670417 235859 670483 235862
rect 675109 235859 675175 235862
rect 674189 235650 674255 235653
rect 674189 235648 674298 235650
rect 674189 235592 674194 235648
rect 674250 235592 674298 235648
rect 674189 235587 674298 235592
rect 674238 235514 674298 235587
rect 675661 235514 675727 235517
rect 674238 235512 675727 235514
rect 674238 235456 675666 235512
rect 675722 235456 675727 235512
rect 674238 235454 675727 235456
rect 675661 235451 675727 235454
rect 674833 235242 674899 235245
rect 676029 235242 676095 235245
rect 674833 235240 676095 235242
rect 674833 235184 674838 235240
rect 674894 235184 676034 235240
rect 676090 235184 676095 235240
rect 674833 235182 676095 235184
rect 674833 235179 674899 235182
rect 676029 235179 676095 235182
rect 674465 234970 674531 234973
rect 675845 234970 675911 234973
rect 674465 234968 675911 234970
rect 674465 234912 674470 234968
rect 674526 234912 675850 234968
rect 675906 234912 675911 234968
rect 674465 234910 675911 234912
rect 674465 234907 674531 234910
rect 675845 234907 675911 234910
rect 42241 234562 42307 234565
rect 46013 234562 46079 234565
rect 42241 234560 46079 234562
rect 42241 234504 42246 234560
rect 42302 234504 46018 234560
rect 46074 234504 46079 234560
rect 42241 234502 46079 234504
rect 42241 234499 42307 234502
rect 46013 234499 46079 234502
rect 668485 234562 668551 234565
rect 672165 234562 672231 234565
rect 668485 234560 672231 234562
rect 668485 234504 668490 234560
rect 668546 234504 672170 234560
rect 672226 234504 672231 234560
rect 668485 234502 672231 234504
rect 668485 234499 668551 234502
rect 672165 234499 672231 234502
rect 674649 234426 674715 234429
rect 675845 234426 675911 234429
rect 674649 234424 675911 234426
rect 674649 234368 674654 234424
rect 674710 234368 675850 234424
rect 675906 234368 675911 234424
rect 674649 234366 675911 234368
rect 674649 234363 674715 234366
rect 675845 234363 675911 234366
rect 42333 234154 42399 234157
rect 44541 234154 44607 234157
rect 42333 234152 44607 234154
rect 42333 234096 42338 234152
rect 42394 234096 44546 234152
rect 44602 234096 44607 234152
rect 42333 234094 44607 234096
rect 42333 234091 42399 234094
rect 44541 234091 44607 234094
rect 661861 234154 661927 234157
rect 683849 234154 683915 234157
rect 661861 234152 683915 234154
rect 661861 234096 661866 234152
rect 661922 234096 683854 234152
rect 683910 234096 683915 234152
rect 661861 234094 683915 234096
rect 661861 234091 661927 234094
rect 683849 234091 683915 234094
rect 554405 233882 554471 233885
rect 552460 233880 554471 233882
rect 552460 233824 554410 233880
rect 554466 233824 554471 233880
rect 552460 233822 554471 233824
rect 554405 233819 554471 233822
rect 658917 233882 658983 233885
rect 683297 233882 683363 233885
rect 658917 233880 683363 233882
rect 658917 233824 658922 233880
rect 658978 233824 683302 233880
rect 683358 233824 683363 233880
rect 658917 233822 683363 233824
rect 658917 233819 658983 233822
rect 683297 233819 683363 233822
rect 42333 233202 42399 233205
rect 44541 233202 44607 233205
rect 42333 233200 44607 233202
rect 42333 233144 42338 233200
rect 42394 233144 44546 233200
rect 44602 233144 44607 233200
rect 42333 233142 44607 233144
rect 42333 233139 42399 233142
rect 44541 233139 44607 233142
rect 670325 233202 670391 233205
rect 671153 233202 671219 233205
rect 670325 233200 671219 233202
rect 670325 233144 670330 233200
rect 670386 233144 671158 233200
rect 671214 233144 671219 233200
rect 670325 233142 671219 233144
rect 670325 233139 670391 233142
rect 671153 233139 671219 233142
rect 670141 232930 670207 232933
rect 673913 232930 673979 232933
rect 670141 232928 673979 232930
rect 670141 232872 670146 232928
rect 670202 232872 673918 232928
rect 673974 232872 673979 232928
rect 670141 232870 673979 232872
rect 670141 232867 670207 232870
rect 673913 232867 673979 232870
rect 42333 231842 42399 231845
rect 43069 231842 43135 231845
rect 675173 231842 675239 231845
rect 42333 231840 43135 231842
rect 42333 231784 42338 231840
rect 42394 231784 43074 231840
rect 43130 231784 43135 231840
rect 42333 231782 43135 231784
rect 42333 231779 42399 231782
rect 43069 231779 43135 231782
rect 663750 231840 675239 231842
rect 663750 231784 675178 231840
rect 675234 231784 675239 231840
rect 663750 231782 675239 231784
rect 663057 231706 663123 231709
rect 663750 231706 663810 231782
rect 675173 231779 675239 231782
rect 663057 231704 663810 231706
rect 663057 231648 663062 231704
rect 663118 231648 663810 231704
rect 663057 231646 663810 231648
rect 663057 231643 663123 231646
rect 672390 231508 672396 231572
rect 672460 231570 672466 231572
rect 675063 231570 675129 231573
rect 672460 231568 675129 231570
rect 672460 231512 675068 231568
rect 675124 231512 675129 231568
rect 672460 231510 675129 231512
rect 672460 231508 672466 231510
rect 675063 231507 675129 231510
rect 640241 231434 640307 231437
rect 671797 231434 671863 231437
rect 640241 231432 671863 231434
rect 640241 231376 640246 231432
rect 640302 231376 671802 231432
rect 671858 231376 671863 231432
rect 640241 231374 671863 231376
rect 640241 231371 640307 231374
rect 671797 231371 671863 231374
rect 665817 231162 665883 231165
rect 674833 231162 674899 231165
rect 665817 231160 674899 231162
rect 665817 231104 665822 231160
rect 665878 231104 674838 231160
rect 674894 231104 674899 231160
rect 665817 231102 674899 231104
rect 665817 231099 665883 231102
rect 674833 231099 674899 231102
rect 664437 230890 664503 230893
rect 674725 230890 674791 230893
rect 664437 230888 674791 230890
rect 664437 230832 664442 230888
rect 664498 230832 674730 230888
rect 674786 230832 674791 230888
rect 664437 230830 674791 230832
rect 664437 230827 664503 230830
rect 674725 230827 674791 230830
rect 674833 230754 674899 230757
rect 675845 230754 675911 230757
rect 674833 230752 675911 230754
rect 674833 230696 674838 230752
rect 674894 230696 675850 230752
rect 675906 230696 675911 230752
rect 674833 230694 675911 230696
rect 674833 230691 674899 230694
rect 675845 230691 675911 230694
rect 663701 230618 663767 230621
rect 672390 230618 672396 230620
rect 663701 230616 672396 230618
rect 663701 230560 663706 230616
rect 663762 230560 672396 230616
rect 663701 230558 672396 230560
rect 663701 230555 663767 230558
rect 672390 230556 672396 230558
rect 672460 230556 672466 230620
rect 674005 230618 674071 230621
rect 674005 230616 674114 230618
rect 674005 230560 674010 230616
rect 674066 230560 674114 230616
rect 674005 230555 674114 230560
rect 42149 230346 42215 230349
rect 45553 230346 45619 230349
rect 42149 230344 45619 230346
rect 42149 230288 42154 230344
rect 42210 230288 45558 230344
rect 45614 230288 45619 230344
rect 42149 230286 45619 230288
rect 42149 230283 42215 230286
rect 45553 230283 45619 230286
rect 661677 230346 661743 230349
rect 674054 230346 674114 230555
rect 674741 230482 674807 230485
rect 676765 230482 676831 230485
rect 674741 230480 676831 230482
rect 674741 230424 674746 230480
rect 674802 230424 676770 230480
rect 676826 230424 676831 230480
rect 674741 230422 676831 230424
rect 674741 230419 674807 230422
rect 676765 230419 676831 230422
rect 661677 230344 674114 230346
rect 661677 230288 661682 230344
rect 661738 230288 674114 230344
rect 661677 230286 674114 230288
rect 661677 230283 661743 230286
rect 674165 230210 674231 230213
rect 674414 230210 674420 230212
rect 674165 230208 674420 230210
rect 674165 230152 674170 230208
rect 674226 230152 674420 230208
rect 674165 230150 674420 230152
rect 674165 230147 674231 230150
rect 674414 230148 674420 230150
rect 674484 230148 674490 230212
rect 676581 230210 676647 230213
rect 674974 230208 676647 230210
rect 674974 230152 676586 230208
rect 676642 230152 676647 230208
rect 674974 230150 676647 230152
rect 639597 230074 639663 230077
rect 673821 230074 673887 230077
rect 639597 230072 673887 230074
rect 639597 230016 639602 230072
rect 639658 230016 673826 230072
rect 673882 230016 673887 230072
rect 639597 230014 673887 230016
rect 639597 230011 639663 230014
rect 673821 230011 673887 230014
rect 673941 229938 674007 229941
rect 674974 229938 675034 230150
rect 676581 230147 676647 230150
rect 673941 229936 675034 229938
rect 673941 229880 673946 229936
rect 674002 229880 675034 229936
rect 673941 229878 675034 229880
rect 673941 229875 674007 229878
rect 103605 229802 103671 229805
rect 145649 229802 145715 229805
rect 103605 229800 145715 229802
rect 103605 229744 103610 229800
rect 103666 229744 145654 229800
rect 145710 229744 145715 229800
rect 103605 229742 145715 229744
rect 103605 229739 103671 229742
rect 145649 229739 145715 229742
rect 660941 229802 661007 229805
rect 673453 229802 673519 229805
rect 660941 229800 673519 229802
rect 660941 229744 660946 229800
rect 661002 229744 673458 229800
rect 673514 229744 673519 229800
rect 660941 229742 673519 229744
rect 660941 229739 661007 229742
rect 673453 229739 673519 229742
rect 674189 229666 674255 229669
rect 675109 229666 675175 229669
rect 674189 229664 675175 229666
rect 674189 229608 674194 229664
rect 674250 229608 675114 229664
rect 675170 229608 675175 229664
rect 674189 229606 675175 229608
rect 674189 229603 674255 229606
rect 675109 229603 675175 229606
rect 667974 229468 667980 229532
rect 668044 229530 668050 229532
rect 668301 229530 668367 229533
rect 668044 229528 668367 229530
rect 668044 229472 668306 229528
rect 668362 229472 668367 229528
rect 668044 229470 668367 229472
rect 668044 229468 668050 229470
rect 668301 229467 668367 229470
rect 42333 229394 42399 229397
rect 45829 229394 45895 229397
rect 42333 229392 45895 229394
rect 42333 229336 42338 229392
rect 42394 229336 45834 229392
rect 45890 229336 45895 229392
rect 42333 229334 45895 229336
rect 42333 229331 42399 229334
rect 45829 229331 45895 229334
rect 673453 229394 673519 229397
rect 675109 229394 675175 229397
rect 673453 229392 675175 229394
rect 673453 229336 673458 229392
rect 673514 229336 675114 229392
rect 675170 229336 675175 229392
rect 673453 229334 675175 229336
rect 673453 229331 673519 229334
rect 675109 229331 675175 229334
rect 146293 229258 146359 229261
rect 147949 229258 148015 229261
rect 146293 229256 148015 229258
rect 146293 229200 146298 229256
rect 146354 229200 147954 229256
rect 148010 229200 148015 229256
rect 146293 229198 148015 229200
rect 146293 229195 146359 229198
rect 147949 229195 148015 229198
rect 167637 229258 167703 229261
rect 172421 229258 172487 229261
rect 167637 229256 172487 229258
rect 167637 229200 167642 229256
rect 167698 229200 172426 229256
rect 172482 229200 172487 229256
rect 167637 229198 172487 229200
rect 167637 229195 167703 229198
rect 172421 229195 172487 229198
rect 673591 229122 673657 229125
rect 675109 229122 675175 229125
rect 673591 229120 675175 229122
rect 673591 229064 673596 229120
rect 673652 229064 675114 229120
rect 675170 229064 675175 229120
rect 673591 229062 675175 229064
rect 673591 229059 673657 229062
rect 675109 229059 675175 229062
rect 157977 228986 158043 228989
rect 163865 228986 163931 228989
rect 157977 228984 163931 228986
rect 157977 228928 157982 228984
rect 158038 228928 163870 228984
rect 163926 228928 163931 228984
rect 157977 228926 163931 228928
rect 157977 228923 158043 228926
rect 163865 228923 163931 228926
rect 172421 228986 172487 228989
rect 175641 228986 175707 228989
rect 172421 228984 175707 228986
rect 172421 228928 172426 228984
rect 172482 228928 175646 228984
rect 175702 228928 175707 228984
rect 172421 228926 175707 228928
rect 172421 228923 172487 228926
rect 175641 228923 175707 228926
rect 180609 228986 180675 228989
rect 181897 228986 181963 228989
rect 180609 228984 181963 228986
rect 180609 228928 180614 228984
rect 180670 228928 181902 228984
rect 181958 228928 181963 228984
rect 180609 228926 181963 228928
rect 180609 228923 180675 228926
rect 181897 228923 181963 228926
rect 166441 228850 166507 228853
rect 168189 228850 168255 228853
rect 166441 228848 168255 228850
rect 166441 228792 166446 228848
rect 166502 228792 168194 228848
rect 168250 228792 168255 228848
rect 166441 228790 168255 228792
rect 166441 228787 166507 228790
rect 168189 228787 168255 228790
rect 190545 228850 190611 228853
rect 192845 228850 192911 228853
rect 190545 228848 192911 228850
rect 190545 228792 190550 228848
rect 190606 228792 192850 228848
rect 192906 228792 192911 228848
rect 190545 228790 192911 228792
rect 190545 228787 190611 228790
rect 192845 228787 192911 228790
rect 672257 228850 672323 228853
rect 673126 228850 673132 228852
rect 672257 228848 673132 228850
rect 672257 228792 672262 228848
rect 672318 228792 673132 228848
rect 672257 228790 673132 228792
rect 672257 228787 672323 228790
rect 673126 228788 673132 228790
rect 673196 228788 673202 228852
rect 673499 228850 673565 228853
rect 675109 228850 675175 228853
rect 673499 228848 675175 228850
rect 673499 228792 673504 228848
rect 673560 228792 675114 228848
rect 675170 228792 675175 228848
rect 673499 228790 675175 228792
rect 673499 228787 673565 228790
rect 675109 228787 675175 228790
rect 181253 228714 181319 228717
rect 181897 228714 181963 228717
rect 181253 228712 181963 228714
rect 181253 228656 181258 228712
rect 181314 228656 181902 228712
rect 181958 228656 181963 228712
rect 181253 228654 181963 228656
rect 181253 228651 181319 228654
rect 181897 228651 181963 228654
rect 147673 228578 147739 228581
rect 149789 228578 149855 228581
rect 147673 228576 149855 228578
rect 147673 228520 147678 228576
rect 147734 228520 149794 228576
rect 149850 228520 149855 228576
rect 147673 228518 149855 228520
rect 147673 228515 147739 228518
rect 149789 228515 149855 228518
rect 157425 228578 157491 228581
rect 158805 228578 158871 228581
rect 672901 228580 672967 228581
rect 672901 228578 672948 228580
rect 157425 228576 158871 228578
rect 157425 228520 157430 228576
rect 157486 228520 158810 228576
rect 158866 228520 158871 228576
rect 157425 228518 158871 228520
rect 672856 228576 672948 228578
rect 672856 228520 672906 228576
rect 672856 228518 672948 228520
rect 157425 228515 157491 228518
rect 158805 228515 158871 228518
rect 672901 228516 672948 228518
rect 673012 228516 673018 228580
rect 673381 228578 673447 228581
rect 675150 228578 675156 228580
rect 673381 228576 675156 228578
rect 673381 228520 673386 228576
rect 673442 228520 675156 228576
rect 673381 228518 675156 228520
rect 672901 228515 672967 228516
rect 673381 228515 673447 228518
rect 675150 228516 675156 228518
rect 675220 228516 675226 228580
rect 166441 228442 166507 228445
rect 168005 228442 168071 228445
rect 166441 228440 168071 228442
rect 166441 228384 166446 228440
rect 166502 228384 168010 228440
rect 168066 228384 168071 228440
rect 166441 228382 168071 228384
rect 166441 228379 166507 228382
rect 168005 228379 168071 228382
rect 79961 228306 80027 228309
rect 160461 228306 160527 228309
rect 79961 228304 160527 228306
rect 79961 228248 79966 228304
rect 80022 228248 160466 228304
rect 160522 228248 160527 228304
rect 79961 228246 160527 228248
rect 79961 228243 80027 228246
rect 160461 228243 160527 228246
rect 135161 228034 135227 228037
rect 141141 228034 141207 228037
rect 135161 228032 141207 228034
rect 135161 227976 135166 228032
rect 135222 227976 141146 228032
rect 141202 227976 141207 228032
rect 135161 227974 141207 227976
rect 135161 227971 135227 227974
rect 141141 227971 141207 227974
rect 155861 228034 155927 228037
rect 157793 228034 157859 228037
rect 155861 228032 157859 228034
rect 155861 227976 155866 228032
rect 155922 227976 157798 228032
rect 157854 227976 157859 228032
rect 155861 227974 157859 227976
rect 155861 227971 155927 227974
rect 157793 227971 157859 227974
rect 181069 228034 181135 228037
rect 181713 228034 181779 228037
rect 181069 228032 181779 228034
rect 181069 227976 181074 228032
rect 181130 227976 181718 228032
rect 181774 227976 181779 228032
rect 181069 227974 181779 227976
rect 181069 227971 181135 227974
rect 181713 227971 181779 227974
rect 42425 227626 42491 227629
rect 43529 227626 43595 227629
rect 42425 227624 43595 227626
rect 42425 227568 42430 227624
rect 42486 227568 43534 227624
rect 43590 227568 43595 227624
rect 42425 227566 43595 227568
rect 42425 227563 42491 227566
rect 43529 227563 43595 227566
rect 151905 227490 151971 227493
rect 152917 227490 152983 227493
rect 151905 227488 152983 227490
rect 151905 227432 151910 227488
rect 151966 227432 152922 227488
rect 152978 227432 152983 227488
rect 151905 227430 152983 227432
rect 151905 227427 151971 227430
rect 152917 227427 152983 227430
rect 159633 227490 159699 227493
rect 166625 227490 166691 227493
rect 159633 227488 166691 227490
rect 159633 227432 159638 227488
rect 159694 227432 166630 227488
rect 166686 227432 166691 227488
rect 159633 227430 166691 227432
rect 159633 227427 159699 227430
rect 166625 227427 166691 227430
rect 41965 227356 42031 227357
rect 41965 227352 42012 227356
rect 42076 227354 42082 227356
rect 41965 227296 41970 227352
rect 41965 227292 42012 227296
rect 42076 227294 42122 227354
rect 42076 227292 42082 227294
rect 41965 227291 42031 227292
rect 142153 227218 142219 227221
rect 143073 227218 143139 227221
rect 142153 227216 143139 227218
rect 142153 227160 142158 227216
rect 142214 227160 143078 227216
rect 143134 227160 143139 227216
rect 142153 227158 143139 227160
rect 142153 227155 142219 227158
rect 143073 227155 143139 227158
rect 150157 227218 150223 227221
rect 154573 227218 154639 227221
rect 150157 227216 154639 227218
rect 150157 227160 150162 227216
rect 150218 227160 154578 227216
rect 154634 227160 154639 227216
rect 150157 227158 154639 227160
rect 150157 227155 150223 227158
rect 154573 227155 154639 227158
rect 672441 227084 672507 227085
rect 672390 227082 672396 227084
rect 672350 227022 672396 227082
rect 672460 227080 672507 227084
rect 672502 227024 672507 227080
rect 672390 227020 672396 227022
rect 672460 227020 672507 227024
rect 672441 227019 672507 227020
rect 672597 227082 672663 227085
rect 672758 227082 672764 227084
rect 672597 227080 672764 227082
rect 672597 227024 672602 227080
rect 672658 227024 672764 227080
rect 672597 227022 672764 227024
rect 672597 227019 672663 227022
rect 672758 227020 672764 227022
rect 672828 227020 672834 227084
rect 673453 227082 673519 227085
rect 673913 227082 673979 227085
rect 673453 227080 673979 227082
rect 673453 227024 673458 227080
rect 673514 227024 673918 227080
rect 673974 227024 673979 227080
rect 673453 227022 673979 227024
rect 673453 227019 673519 227022
rect 673913 227019 673979 227022
rect 73061 226946 73127 226949
rect 155309 226946 155375 226949
rect 73061 226944 155375 226946
rect 73061 226888 73066 226944
rect 73122 226888 155314 226944
rect 155370 226888 155375 226944
rect 73061 226886 155375 226888
rect 73061 226883 73127 226886
rect 155309 226883 155375 226886
rect 672373 226810 672439 226813
rect 675385 226810 675451 226813
rect 672373 226808 675451 226810
rect 672373 226752 672378 226808
rect 672434 226752 675390 226808
rect 675446 226752 675451 226808
rect 672373 226750 675451 226752
rect 672373 226747 672439 226750
rect 675385 226747 675451 226750
rect 134977 226674 135043 226677
rect 135621 226674 135687 226677
rect 134977 226672 135687 226674
rect 134977 226616 134982 226672
rect 135038 226616 135626 226672
rect 135682 226616 135687 226672
rect 134977 226614 135687 226616
rect 134977 226611 135043 226614
rect 135621 226611 135687 226614
rect 139301 226538 139367 226541
rect 142245 226538 142311 226541
rect 139301 226536 142311 226538
rect 139301 226480 139306 226536
rect 139362 226480 142250 226536
rect 142306 226480 142311 226536
rect 139301 226478 142311 226480
rect 139301 226475 139367 226478
rect 142245 226475 142311 226478
rect 672809 226538 672875 226541
rect 675017 226538 675083 226541
rect 672809 226536 675083 226538
rect 672809 226480 672814 226536
rect 672870 226480 675022 226536
rect 675078 226480 675083 226536
rect 672809 226478 675083 226480
rect 672809 226475 672875 226478
rect 675017 226475 675083 226478
rect 652753 226402 652819 226405
rect 668301 226402 668367 226405
rect 652753 226400 668367 226402
rect 652753 226344 652758 226400
rect 652814 226344 668306 226400
rect 668362 226344 668367 226400
rect 652753 226342 668367 226344
rect 652753 226339 652819 226342
rect 668301 226339 668367 226342
rect 672027 226266 672093 226269
rect 674097 226266 674163 226269
rect 672027 226264 674163 226266
rect 672027 226208 672032 226264
rect 672088 226208 674102 226264
rect 674158 226208 674163 226264
rect 672027 226206 674163 226208
rect 672027 226203 672093 226206
rect 674097 226203 674163 226206
rect 136541 226130 136607 226133
rect 141693 226130 141759 226133
rect 136541 226128 141759 226130
rect 136541 226072 136546 226128
rect 136602 226072 141698 226128
rect 141754 226072 141759 226128
rect 136541 226070 141759 226072
rect 136541 226067 136607 226070
rect 141693 226067 141759 226070
rect 153101 226130 153167 226133
rect 157609 226130 157675 226133
rect 153101 226128 157675 226130
rect 153101 226072 153106 226128
rect 153162 226072 157614 226128
rect 157670 226072 157675 226128
rect 153101 226070 157675 226072
rect 153101 226067 153167 226070
rect 157609 226067 157675 226070
rect 161197 226130 161263 226133
rect 162301 226130 162367 226133
rect 161197 226128 162367 226130
rect 161197 226072 161202 226128
rect 161258 226072 162306 226128
rect 162362 226072 162367 226128
rect 161197 226070 162367 226072
rect 161197 226067 161263 226070
rect 162301 226067 162367 226070
rect 169201 226130 169267 226133
rect 169201 226128 173910 226130
rect 169201 226072 169206 226128
rect 169262 226072 173910 226128
rect 169201 226070 173910 226072
rect 169201 226067 169267 226070
rect 146937 225994 147003 225997
rect 152825 225994 152891 225997
rect 146937 225992 152891 225994
rect 146937 225936 146942 225992
rect 146998 225936 152830 225992
rect 152886 225936 152891 225992
rect 146937 225934 152891 225936
rect 146937 225931 147003 225934
rect 152825 225931 152891 225934
rect 166809 225994 166875 225997
rect 169017 225994 169083 225997
rect 166809 225992 169083 225994
rect 166809 225936 166814 225992
rect 166870 225936 169022 225992
rect 169078 225936 169083 225992
rect 166809 225934 169083 225936
rect 173850 225994 173910 226070
rect 178677 225994 178743 225997
rect 173850 225992 178743 225994
rect 173850 225936 178682 225992
rect 178738 225936 178743 225992
rect 173850 225934 178743 225936
rect 166809 225931 166875 225934
rect 169017 225931 169083 225934
rect 178677 225931 178743 225934
rect 185669 225994 185735 225997
rect 195421 225994 195487 225997
rect 185669 225992 195487 225994
rect 185669 225936 185674 225992
rect 185730 225936 195426 225992
rect 195482 225936 195487 225992
rect 185669 225934 195487 225936
rect 185669 225931 185735 225934
rect 195421 225931 195487 225934
rect 671797 225994 671863 225997
rect 675334 225994 675340 225996
rect 671797 225992 675340 225994
rect 671797 225936 671802 225992
rect 671858 225936 675340 225992
rect 671797 225934 675340 225936
rect 671797 225931 671863 225934
rect 675334 225932 675340 225934
rect 675404 225932 675410 225996
rect 42425 225722 42491 225725
rect 43161 225722 43227 225725
rect 42425 225720 43227 225722
rect 42425 225664 42430 225720
rect 42486 225664 43166 225720
rect 43222 225664 43227 225720
rect 42425 225662 43227 225664
rect 42425 225659 42491 225662
rect 43161 225659 43227 225662
rect 184841 225722 184907 225725
rect 187325 225722 187391 225725
rect 671061 225722 671127 225725
rect 184841 225720 187391 225722
rect 184841 225664 184846 225720
rect 184902 225664 187330 225720
rect 187386 225664 187391 225720
rect 184841 225662 187391 225664
rect 184841 225659 184907 225662
rect 187325 225659 187391 225662
rect 663750 225720 671127 225722
rect 663750 225664 671066 225720
rect 671122 225664 671127 225720
rect 663750 225662 671127 225664
rect 143165 225586 143231 225589
rect 147121 225586 147187 225589
rect 143165 225584 147187 225586
rect 143165 225528 143170 225584
rect 143226 225528 147126 225584
rect 147182 225528 147187 225584
rect 143165 225526 147187 225528
rect 143165 225523 143231 225526
rect 147121 225523 147187 225526
rect 162301 225586 162367 225589
rect 166901 225586 166967 225589
rect 162301 225584 166967 225586
rect 162301 225528 162306 225584
rect 162362 225528 166906 225584
rect 166962 225528 166967 225584
rect 162301 225526 166967 225528
rect 162301 225523 162367 225526
rect 166901 225523 166967 225526
rect 176469 225586 176535 225589
rect 177021 225586 177087 225589
rect 176469 225584 177087 225586
rect 176469 225528 176474 225584
rect 176530 225528 177026 225584
rect 177082 225528 177087 225584
rect 176469 225526 177087 225528
rect 176469 225523 176535 225526
rect 177021 225523 177087 225526
rect 658917 225586 658983 225589
rect 663750 225586 663810 225662
rect 671061 225659 671127 225662
rect 671813 225722 671879 225725
rect 672022 225722 672028 225724
rect 671813 225720 672028 225722
rect 671813 225664 671818 225720
rect 671874 225664 672028 225720
rect 671813 225662 672028 225664
rect 671813 225659 671879 225662
rect 672022 225660 672028 225662
rect 672092 225660 672098 225724
rect 658917 225584 663810 225586
rect 658917 225528 658922 225584
rect 658978 225528 663810 225584
rect 658917 225526 663810 225528
rect 672533 225586 672599 225589
rect 675201 225586 675267 225589
rect 672533 225584 675267 225586
rect 672533 225528 672538 225584
rect 672594 225528 675206 225584
rect 675262 225528 675267 225584
rect 672533 225526 675267 225528
rect 658917 225523 658983 225526
rect 672533 225523 672599 225526
rect 675201 225523 675267 225526
rect 185669 225450 185735 225453
rect 194869 225450 194935 225453
rect 185669 225448 194935 225450
rect 185669 225392 185674 225448
rect 185730 225392 194874 225448
rect 194930 225392 194935 225448
rect 185669 225390 194935 225392
rect 185669 225387 185735 225390
rect 194869 225387 194935 225390
rect 145925 225314 145991 225317
rect 153285 225314 153351 225317
rect 145925 225312 153351 225314
rect 145925 225256 145930 225312
rect 145986 225256 153290 225312
rect 153346 225256 153351 225312
rect 145925 225254 153351 225256
rect 145925 225251 145991 225254
rect 153285 225251 153351 225254
rect 166993 225314 167059 225317
rect 169845 225314 169911 225317
rect 166993 225312 169911 225314
rect 166993 225256 166998 225312
rect 167054 225256 169850 225312
rect 169906 225256 169911 225312
rect 166993 225254 169911 225256
rect 166993 225251 167059 225254
rect 169845 225251 169911 225254
rect 176469 225314 176535 225317
rect 177205 225314 177271 225317
rect 176469 225312 177271 225314
rect 176469 225256 176474 225312
rect 176530 225256 177210 225312
rect 177266 225256 177271 225312
rect 176469 225254 177271 225256
rect 176469 225251 176535 225254
rect 177205 225251 177271 225254
rect 655513 225314 655579 225317
rect 668301 225314 668367 225317
rect 655513 225312 668367 225314
rect 655513 225256 655518 225312
rect 655574 225256 668306 225312
rect 668362 225256 668367 225312
rect 655513 225254 668367 225256
rect 655513 225251 655579 225254
rect 668301 225251 668367 225254
rect 671061 225314 671127 225317
rect 673545 225314 673611 225317
rect 671061 225312 673611 225314
rect 671061 225256 671066 225312
rect 671122 225256 673550 225312
rect 673606 225256 673611 225312
rect 671061 225254 673611 225256
rect 671061 225251 671127 225254
rect 673545 225251 673611 225254
rect 183277 225178 183343 225181
rect 187509 225178 187575 225181
rect 183277 225176 187575 225178
rect 183277 225120 183282 225176
rect 183338 225120 187514 225176
rect 187570 225120 187575 225176
rect 183277 225118 187575 225120
rect 183277 225115 183343 225118
rect 187509 225115 187575 225118
rect 166441 225042 166507 225045
rect 167361 225042 167427 225045
rect 166441 225040 167427 225042
rect 166441 224984 166446 225040
rect 166502 224984 167366 225040
rect 167422 224984 167427 225040
rect 166441 224982 167427 224984
rect 166441 224979 166507 224982
rect 167361 224979 167427 224982
rect 654777 225042 654843 225045
rect 669405 225042 669471 225045
rect 654777 225040 669471 225042
rect 654777 224984 654782 225040
rect 654838 224984 669410 225040
rect 669466 224984 669471 225040
rect 654777 224982 669471 224984
rect 654777 224979 654843 224982
rect 669405 224979 669471 224982
rect 673494 224980 673500 225044
rect 673564 225042 673570 225044
rect 674414 225042 674420 225044
rect 673564 224982 674420 225042
rect 673564 224980 673570 224982
rect 674414 224980 674420 224982
rect 674484 224980 674490 225044
rect 185669 224906 185735 224909
rect 187049 224906 187115 224909
rect 185669 224904 187115 224906
rect 185669 224848 185674 224904
rect 185730 224848 187054 224904
rect 187110 224848 187115 224904
rect 185669 224846 187115 224848
rect 185669 224843 185735 224846
rect 187049 224843 187115 224846
rect 671061 224906 671127 224909
rect 672717 224906 672783 224909
rect 671061 224904 672783 224906
rect 671061 224848 671066 224904
rect 671122 224848 672722 224904
rect 672778 224848 672783 224904
rect 671061 224846 672783 224848
rect 671061 224843 671127 224846
rect 672717 224843 672783 224846
rect 142153 224634 142219 224637
rect 147305 224634 147371 224637
rect 142153 224632 147371 224634
rect 142153 224576 142158 224632
rect 142214 224576 147310 224632
rect 147366 224576 147371 224632
rect 142153 224574 147371 224576
rect 142153 224571 142219 224574
rect 147305 224571 147371 224574
rect 157333 224634 157399 224637
rect 162945 224634 163011 224637
rect 157333 224632 163011 224634
rect 157333 224576 157338 224632
rect 157394 224576 162950 224632
rect 163006 224576 163011 224632
rect 157333 224574 163011 224576
rect 157333 224571 157399 224574
rect 162945 224571 163011 224574
rect 672533 224634 672599 224637
rect 673126 224634 673132 224636
rect 672533 224632 673132 224634
rect 672533 224576 672538 224632
rect 672594 224576 673132 224632
rect 672533 224574 673132 224576
rect 672533 224571 672599 224574
rect 673126 224572 673132 224574
rect 673196 224572 673202 224636
rect 163957 224498 164023 224501
rect 170765 224498 170831 224501
rect 163957 224496 170831 224498
rect 163957 224440 163962 224496
rect 164018 224440 170770 224496
rect 170826 224440 170831 224496
rect 163957 224438 170831 224440
rect 163957 224435 164023 224438
rect 170765 224435 170831 224438
rect 659285 224498 659351 224501
rect 671015 224498 671081 224501
rect 659285 224496 671081 224498
rect 659285 224440 659290 224496
rect 659346 224440 671020 224496
rect 671076 224440 671081 224496
rect 659285 224438 671081 224440
rect 659285 224435 659351 224438
rect 671015 224435 671081 224438
rect 152549 224362 152615 224365
rect 142110 224360 152615 224362
rect 142110 224304 152554 224360
rect 152610 224304 152615 224360
rect 142110 224302 152615 224304
rect 68921 224226 68987 224229
rect 142110 224226 142170 224302
rect 152549 224299 152615 224302
rect 672758 224300 672764 224364
rect 672828 224362 672834 224364
rect 674833 224362 674899 224365
rect 672828 224360 674899 224362
rect 672828 224304 674838 224360
rect 674894 224304 674899 224360
rect 672828 224302 674899 224304
rect 672828 224300 672834 224302
rect 674833 224299 674899 224302
rect 68921 224224 142170 224226
rect 68921 224168 68926 224224
rect 68982 224168 142170 224224
rect 68921 224166 142170 224168
rect 154573 224226 154639 224229
rect 157425 224226 157491 224229
rect 154573 224224 157491 224226
rect 154573 224168 154578 224224
rect 154634 224168 157430 224224
rect 157486 224168 157491 224224
rect 154573 224166 157491 224168
rect 68921 224163 68987 224166
rect 154573 224163 154639 224166
rect 157425 224163 157491 224166
rect 170949 224226 171015 224229
rect 171409 224226 171475 224229
rect 170949 224224 171475 224226
rect 170949 224168 170954 224224
rect 171010 224168 171414 224224
rect 171470 224168 171475 224224
rect 170949 224166 171475 224168
rect 170949 224163 171015 224166
rect 171409 224163 171475 224166
rect 145557 224090 145623 224093
rect 145557 224088 147690 224090
rect 145557 224032 145562 224088
rect 145618 224032 147690 224088
rect 145557 224030 147690 224032
rect 145557 224027 145623 224030
rect 147630 223957 147690 224030
rect 141785 223954 141851 223957
rect 142613 223954 142679 223957
rect 141785 223952 142679 223954
rect 141785 223896 141790 223952
rect 141846 223896 142618 223952
rect 142674 223896 142679 223952
rect 141785 223894 142679 223896
rect 147630 223952 147739 223957
rect 147630 223896 147678 223952
rect 147734 223896 147739 223952
rect 147630 223894 147739 223896
rect 141785 223891 141851 223894
rect 142613 223891 142679 223894
rect 147673 223891 147739 223894
rect 656617 223954 656683 223957
rect 667933 223954 667999 223957
rect 656617 223952 667999 223954
rect 656617 223896 656622 223952
rect 656678 223896 667938 223952
rect 667994 223896 667999 223952
rect 656617 223894 667999 223896
rect 656617 223891 656683 223894
rect 667933 223891 667999 223894
rect 151721 223818 151787 223821
rect 156873 223818 156939 223821
rect 679249 223818 679315 223821
rect 151721 223816 156939 223818
rect 151721 223760 151726 223816
rect 151782 223760 156878 223816
rect 156934 223760 156939 223816
rect 151721 223758 156939 223760
rect 151721 223755 151787 223758
rect 156873 223755 156939 223758
rect 679206 223816 679315 223818
rect 679206 223760 679254 223816
rect 679310 223760 679315 223816
rect 679206 223755 679315 223760
rect 658181 223682 658247 223685
rect 669405 223682 669471 223685
rect 658181 223680 669471 223682
rect 658181 223624 658186 223680
rect 658242 223624 669410 223680
rect 669466 223624 669471 223680
rect 658181 223622 669471 223624
rect 658181 223619 658247 223622
rect 669405 223619 669471 223622
rect 679206 223516 679266 223755
rect 156873 223274 156939 223277
rect 157425 223274 157491 223277
rect 666645 223274 666711 223277
rect 156873 223272 157491 223274
rect 156873 223216 156878 223272
rect 156934 223216 157430 223272
rect 157486 223216 157491 223272
rect 156873 223214 157491 223216
rect 156873 223211 156939 223214
rect 157425 223211 157491 223214
rect 659610 223272 666711 223274
rect 659610 223216 666650 223272
rect 666706 223216 666711 223272
rect 659610 223214 666711 223216
rect 158345 223138 158411 223141
rect 165061 223138 165127 223141
rect 158345 223136 165127 223138
rect 158345 223080 158350 223136
rect 158406 223080 165066 223136
rect 165122 223080 165127 223136
rect 158345 223078 165127 223080
rect 158345 223075 158411 223078
rect 165061 223075 165127 223078
rect 166441 223138 166507 223141
rect 170397 223138 170463 223141
rect 166441 223136 170463 223138
rect 166441 223080 166446 223136
rect 166502 223080 170402 223136
rect 170458 223080 170463 223136
rect 166441 223078 170463 223080
rect 166441 223075 166507 223078
rect 170397 223075 170463 223078
rect 650637 223138 650703 223141
rect 659610 223138 659670 223214
rect 666645 223211 666711 223214
rect 683297 223138 683363 223141
rect 650637 223136 659670 223138
rect 650637 223080 650642 223136
rect 650698 223080 659670 223136
rect 650637 223078 659670 223080
rect 683284 223136 683363 223138
rect 683284 223080 683302 223136
rect 683358 223080 683363 223136
rect 683284 223078 683363 223080
rect 650637 223075 650703 223078
rect 683297 223075 683363 223078
rect 672073 223004 672139 223005
rect 672022 222940 672028 223004
rect 672092 223002 672139 223004
rect 672092 223000 672184 223002
rect 672134 222944 672184 223000
rect 672092 222942 672184 222944
rect 672092 222940 672139 222942
rect 672073 222939 672139 222940
rect 40677 222866 40743 222869
rect 62941 222866 63007 222869
rect 40677 222864 63007 222866
rect 40677 222808 40682 222864
rect 40738 222808 62946 222864
rect 63002 222808 63007 222864
rect 40677 222806 63007 222808
rect 40677 222803 40743 222806
rect 62941 222803 63007 222806
rect 123477 222866 123543 222869
rect 165613 222866 165679 222869
rect 123477 222864 165679 222866
rect 123477 222808 123482 222864
rect 123538 222808 165618 222864
rect 165674 222808 165679 222864
rect 123477 222806 165679 222808
rect 123477 222803 123543 222806
rect 165613 222803 165679 222806
rect 652017 222866 652083 222869
rect 666829 222866 666895 222869
rect 652017 222864 666895 222866
rect 652017 222808 652022 222864
rect 652078 222808 666834 222864
rect 666890 222808 666895 222864
rect 652017 222806 666895 222808
rect 652017 222803 652083 222806
rect 666829 222803 666895 222806
rect 683849 222730 683915 222733
rect 683836 222728 683915 222730
rect 683836 222672 683854 222728
rect 683910 222672 683915 222728
rect 683836 222670 683915 222672
rect 683849 222667 683915 222670
rect 155033 222594 155099 222597
rect 157241 222594 157307 222597
rect 155033 222592 157307 222594
rect 155033 222536 155038 222592
rect 155094 222536 157246 222592
rect 157302 222536 157307 222592
rect 155033 222534 157307 222536
rect 155033 222531 155099 222534
rect 157241 222531 157307 222534
rect 565629 222594 565695 222597
rect 572478 222594 572484 222596
rect 565629 222592 572484 222594
rect 565629 222536 565634 222592
rect 565690 222536 572484 222592
rect 565629 222534 572484 222536
rect 565629 222531 565695 222534
rect 572478 222532 572484 222534
rect 572548 222532 572554 222596
rect 142981 222458 143047 222461
rect 145005 222458 145071 222461
rect 142981 222456 145071 222458
rect 142981 222400 142986 222456
rect 143042 222400 145010 222456
rect 145066 222400 145071 222456
rect 142981 222398 145071 222400
rect 142981 222395 143047 222398
rect 145005 222395 145071 222398
rect 171225 222322 171291 222325
rect 179965 222322 180031 222325
rect 171225 222320 180031 222322
rect 171225 222264 171230 222320
rect 171286 222264 179970 222320
rect 180026 222264 180031 222320
rect 171225 222262 180031 222264
rect 171225 222259 171291 222262
rect 179965 222259 180031 222262
rect 560661 222322 560727 222325
rect 561254 222322 561260 222324
rect 560661 222320 561260 222322
rect 560661 222264 560666 222320
rect 560722 222264 561260 222320
rect 560661 222262 561260 222264
rect 560661 222259 560727 222262
rect 561254 222260 561260 222262
rect 561324 222260 561330 222324
rect 561949 222322 562015 222325
rect 562685 222322 562751 222325
rect 582189 222322 582255 222325
rect 679985 222322 680051 222325
rect 561949 222320 582255 222322
rect 561949 222264 561954 222320
rect 562010 222264 562690 222320
rect 562746 222264 582194 222320
rect 582250 222264 582255 222320
rect 561949 222262 582255 222264
rect 679972 222320 680051 222322
rect 679972 222264 679990 222320
rect 680046 222264 680051 222320
rect 679972 222262 680051 222264
rect 561949 222259 562015 222262
rect 562685 222259 562751 222262
rect 582189 222259 582255 222262
rect 679985 222259 680051 222262
rect 674833 222186 674899 222189
rect 669270 222184 674899 222186
rect 669270 222128 674838 222184
rect 674894 222128 674899 222184
rect 669270 222126 674899 222128
rect 176101 222050 176167 222053
rect 177021 222050 177087 222053
rect 176101 222048 177087 222050
rect 176101 221992 176106 222048
rect 176162 221992 177026 222048
rect 177082 221992 177087 222048
rect 176101 221990 177087 221992
rect 176101 221987 176167 221990
rect 177021 221987 177087 221990
rect 555785 222050 555851 222053
rect 562910 222050 562916 222052
rect 555785 222048 562916 222050
rect 555785 221992 555790 222048
rect 555846 221992 562916 222048
rect 555785 221990 562916 221992
rect 555785 221987 555851 221990
rect 562910 221988 562916 221990
rect 562980 221988 562986 222052
rect 563094 221988 563100 222052
rect 563164 222050 563170 222052
rect 563421 222050 563487 222053
rect 563164 222048 563487 222050
rect 563164 221992 563426 222048
rect 563482 221992 563487 222048
rect 563164 221990 563487 221992
rect 563164 221988 563170 221990
rect 563421 221987 563487 221990
rect 563646 221988 563652 222052
rect 563716 222050 563722 222052
rect 572110 222050 572116 222052
rect 563716 221990 572116 222050
rect 563716 221988 563722 221990
rect 572110 221988 572116 221990
rect 572180 221988 572186 222052
rect 572299 222050 572365 222053
rect 576577 222050 576643 222053
rect 572299 222048 576643 222050
rect 572299 221992 572304 222048
rect 572360 221992 576582 222048
rect 576638 221992 576643 222048
rect 572299 221990 576643 221992
rect 572299 221987 572365 221990
rect 576577 221987 576643 221990
rect 142153 221914 142219 221917
rect 149053 221914 149119 221917
rect 142153 221912 149119 221914
rect 142153 221856 142158 221912
rect 142214 221856 149058 221912
rect 149114 221856 149119 221912
rect 142153 221854 149119 221856
rect 142153 221851 142219 221854
rect 149053 221851 149119 221854
rect 171041 221914 171107 221917
rect 171501 221914 171567 221917
rect 171041 221912 171567 221914
rect 171041 221856 171046 221912
rect 171102 221856 171506 221912
rect 171562 221856 171567 221912
rect 171041 221854 171567 221856
rect 171041 221851 171107 221854
rect 171501 221851 171567 221854
rect 513373 221914 513439 221917
rect 513373 221912 514770 221914
rect 513373 221856 513378 221912
rect 513434 221856 514770 221912
rect 513373 221854 514770 221856
rect 513373 221851 513439 221854
rect 514710 221778 514770 221854
rect 599485 221778 599551 221781
rect 514710 221776 599551 221778
rect 514710 221720 599490 221776
rect 599546 221720 599551 221776
rect 514710 221718 599551 221720
rect 599485 221715 599551 221718
rect 601509 221778 601575 221781
rect 602245 221778 602311 221781
rect 601509 221776 602311 221778
rect 601509 221720 601514 221776
rect 601570 221720 602250 221776
rect 602306 221720 602311 221776
rect 601509 221718 602311 221720
rect 601509 221715 601575 221718
rect 602245 221715 602311 221718
rect 659469 221778 659535 221781
rect 669270 221778 669330 222126
rect 674833 222123 674899 222126
rect 674649 221914 674715 221917
rect 674649 221912 676292 221914
rect 674649 221856 674654 221912
rect 674710 221856 676292 221912
rect 674649 221854 676292 221856
rect 674649 221851 674715 221854
rect 659469 221776 669330 221778
rect 659469 221720 659474 221776
rect 659530 221720 669330 221776
rect 659469 221718 669330 221720
rect 659469 221715 659535 221718
rect 101857 221506 101923 221509
rect 178033 221506 178099 221509
rect 101857 221504 178099 221506
rect 101857 221448 101862 221504
rect 101918 221448 178038 221504
rect 178094 221448 178099 221504
rect 101857 221446 178099 221448
rect 101857 221443 101923 221446
rect 178033 221443 178099 221446
rect 517789 221506 517855 221509
rect 616873 221506 616939 221509
rect 517789 221504 616939 221506
rect 517789 221448 517794 221504
rect 517850 221448 616878 221504
rect 616934 221448 616939 221504
rect 517789 221446 616939 221448
rect 517789 221443 517855 221446
rect 616873 221443 616939 221446
rect 657997 221506 658063 221509
rect 671797 221506 671863 221509
rect 679801 221506 679867 221509
rect 657997 221504 671863 221506
rect 657997 221448 658002 221504
rect 658058 221448 671802 221504
rect 671858 221448 671863 221504
rect 657997 221446 671863 221448
rect 679788 221504 679867 221506
rect 679788 221448 679806 221504
rect 679862 221448 679867 221504
rect 679788 221446 679867 221448
rect 657997 221443 658063 221446
rect 671797 221443 671863 221446
rect 679801 221443 679867 221446
rect 138473 221234 138539 221237
rect 142245 221234 142311 221237
rect 138473 221232 142311 221234
rect 138473 221176 138478 221232
rect 138534 221176 142250 221232
rect 142306 221176 142311 221232
rect 138473 221174 142311 221176
rect 138473 221171 138539 221174
rect 142245 221171 142311 221174
rect 180609 221234 180675 221237
rect 180885 221234 180951 221237
rect 180609 221232 180951 221234
rect 180609 221176 180614 221232
rect 180670 221176 180890 221232
rect 180946 221176 180951 221232
rect 180609 221174 180951 221176
rect 180609 221171 180675 221174
rect 180885 221171 180951 221174
rect 515949 221234 516015 221237
rect 600589 221234 600655 221237
rect 515949 221232 600655 221234
rect 515949 221176 515954 221232
rect 516010 221176 600594 221232
rect 600650 221176 600655 221232
rect 515949 221174 600655 221176
rect 515949 221171 516015 221174
rect 600589 221171 600655 221174
rect 666645 221098 666711 221101
rect 666645 221096 676292 221098
rect 666645 221040 666650 221096
rect 666706 221040 676292 221096
rect 666645 221038 676292 221040
rect 666645 221035 666711 221038
rect 486601 220962 486667 220965
rect 611629 220962 611695 220965
rect 486601 220960 611695 220962
rect 486601 220904 486606 220960
rect 486662 220904 611634 220960
rect 611690 220904 611695 220960
rect 486601 220902 611695 220904
rect 486601 220899 486667 220902
rect 611629 220899 611695 220902
rect 142153 220826 142219 220829
rect 148409 220826 148475 220829
rect 142153 220824 148475 220826
rect 142153 220768 142158 220824
rect 142214 220768 148414 220824
rect 148470 220768 148475 220824
rect 142153 220766 148475 220768
rect 142153 220763 142219 220766
rect 148409 220763 148475 220766
rect 150709 220826 150775 220829
rect 156137 220826 156203 220829
rect 150709 220824 156203 220826
rect 150709 220768 150714 220824
rect 150770 220768 156142 220824
rect 156198 220768 156203 220824
rect 150709 220766 156203 220768
rect 150709 220763 150775 220766
rect 156137 220763 156203 220766
rect 180793 220826 180859 220829
rect 185945 220826 186011 220829
rect 180793 220824 186011 220826
rect 180793 220768 180798 220824
rect 180854 220768 185950 220824
rect 186006 220768 186011 220824
rect 180793 220766 186011 220768
rect 180793 220763 180859 220766
rect 185945 220763 186011 220766
rect 194777 220826 194843 220829
rect 196065 220826 196131 220829
rect 194777 220824 196131 220826
rect 194777 220768 194782 220824
rect 194838 220768 196070 220824
rect 196126 220768 196131 220824
rect 194777 220766 196131 220768
rect 194777 220763 194843 220766
rect 196065 220763 196131 220766
rect 582373 220690 582439 220693
rect 591849 220690 591915 220693
rect 582373 220688 591915 220690
rect 582373 220632 582378 220688
rect 582434 220632 591854 220688
rect 591910 220632 591915 220688
rect 582373 220630 591915 220632
rect 582373 220627 582439 220630
rect 591849 220627 591915 220630
rect 592309 220690 592375 220693
rect 600405 220690 600471 220693
rect 592309 220688 600471 220690
rect 592309 220632 592314 220688
rect 592370 220632 600410 220688
rect 600466 220632 600471 220688
rect 592309 220630 600471 220632
rect 592309 220627 592375 220630
rect 600405 220627 600471 220630
rect 653029 220690 653095 220693
rect 673545 220690 673611 220693
rect 676029 220690 676095 220693
rect 679617 220690 679683 220693
rect 653029 220688 673611 220690
rect 653029 220632 653034 220688
rect 653090 220632 673550 220688
rect 673606 220632 673611 220688
rect 653029 220630 673611 220632
rect 653029 220627 653095 220630
rect 673545 220627 673611 220630
rect 674422 220688 676095 220690
rect 674422 220632 676034 220688
rect 676090 220632 676095 220688
rect 674422 220630 676095 220632
rect 679604 220688 679683 220690
rect 679604 220632 679622 220688
rect 679678 220632 679683 220688
rect 679604 220630 679683 220632
rect 153653 220554 153719 220557
rect 142110 220552 153719 220554
rect 142110 220496 153658 220552
rect 153714 220496 153719 220552
rect 142110 220494 153719 220496
rect 72877 220418 72943 220421
rect 142110 220418 142170 220494
rect 153653 220491 153719 220494
rect 157333 220554 157399 220557
rect 161749 220554 161815 220557
rect 157333 220552 161815 220554
rect 157333 220496 157338 220552
rect 157394 220496 161754 220552
rect 161810 220496 161815 220552
rect 157333 220494 161815 220496
rect 157333 220491 157399 220494
rect 161749 220491 161815 220494
rect 161933 220554 161999 220557
rect 162853 220554 162919 220557
rect 545021 220556 545087 220557
rect 545021 220554 545068 220556
rect 161933 220552 162919 220554
rect 161933 220496 161938 220552
rect 161994 220496 162858 220552
rect 162914 220496 162919 220552
rect 161933 220494 162919 220496
rect 544976 220552 545068 220554
rect 544976 220496 545026 220552
rect 544976 220494 545068 220496
rect 161933 220491 161999 220494
rect 162853 220491 162919 220494
rect 545021 220492 545068 220494
rect 545132 220492 545138 220556
rect 545297 220554 545363 220557
rect 545297 220552 553410 220554
rect 545297 220496 545302 220552
rect 545358 220496 553410 220552
rect 545297 220494 553410 220496
rect 545021 220491 545087 220492
rect 545297 220491 545363 220494
rect 72877 220416 142170 220418
rect 72877 220360 72882 220416
rect 72938 220360 142170 220416
rect 72877 220358 142170 220360
rect 72877 220355 72943 220358
rect 519537 220282 519603 220285
rect 542537 220282 542603 220285
rect 543365 220282 543431 220285
rect 519537 220280 534090 220282
rect 519537 220224 519542 220280
rect 519598 220224 534090 220280
rect 519537 220222 534090 220224
rect 519537 220219 519603 220222
rect 69749 220146 69815 220149
rect 151077 220146 151143 220149
rect 69749 220144 151143 220146
rect 69749 220088 69754 220144
rect 69810 220088 151082 220144
rect 151138 220088 151143 220144
rect 69749 220086 151143 220088
rect 69749 220083 69815 220086
rect 151077 220083 151143 220086
rect 510981 220012 511047 220013
rect 510981 220008 511028 220012
rect 511092 220010 511098 220012
rect 512637 220010 512703 220013
rect 530025 220012 530091 220013
rect 529974 220010 529980 220012
rect 510981 219952 510986 220008
rect 510981 219948 511028 219952
rect 511092 219950 511138 220010
rect 512637 220008 524430 220010
rect 512637 219952 512642 220008
rect 512698 219952 524430 220008
rect 512637 219950 524430 219952
rect 529934 219950 529980 220010
rect 530044 220008 530091 220012
rect 530301 220012 530367 220013
rect 530301 220010 530348 220012
rect 530086 219952 530091 220008
rect 511092 219948 511098 219950
rect 510981 219947 511047 219948
rect 512637 219947 512703 219950
rect 141969 219874 142035 219877
rect 142245 219874 142311 219877
rect 141969 219872 142311 219874
rect 141969 219816 141974 219872
rect 142030 219816 142250 219872
rect 142306 219816 142311 219872
rect 141969 219814 142311 219816
rect 141969 219811 142035 219814
rect 142245 219811 142311 219814
rect 494789 219738 494855 219741
rect 519537 219738 519603 219741
rect 519813 219740 519879 219741
rect 522573 219740 522639 219741
rect 519813 219738 519860 219740
rect 494789 219736 519603 219738
rect 494789 219680 494794 219736
rect 494850 219680 519542 219736
rect 519598 219680 519603 219736
rect 494789 219678 519603 219680
rect 519768 219736 519860 219738
rect 519768 219680 519818 219736
rect 519768 219678 519860 219680
rect 494789 219675 494855 219678
rect 519537 219675 519603 219678
rect 519813 219676 519860 219678
rect 519924 219676 519930 219740
rect 522573 219736 522620 219740
rect 522684 219738 522690 219740
rect 524370 219738 524430 219950
rect 529974 219948 529980 219950
rect 530044 219948 530091 219952
rect 530256 220008 530348 220010
rect 530256 219952 530306 220008
rect 530256 219950 530348 219952
rect 530025 219947 530091 219948
rect 530301 219948 530348 219950
rect 530412 219948 530418 220012
rect 534030 220010 534090 220222
rect 542537 220280 543431 220282
rect 542537 220224 542542 220280
rect 542598 220224 543370 220280
rect 543426 220224 543431 220280
rect 542537 220222 543431 220224
rect 542537 220219 542603 220222
rect 543365 220219 543431 220222
rect 543774 220220 543780 220284
rect 543844 220282 543850 220284
rect 553025 220282 553091 220285
rect 543844 220280 553091 220282
rect 543844 220224 553030 220280
rect 553086 220224 553091 220280
rect 543844 220222 553091 220224
rect 553350 220282 553410 220494
rect 553894 220492 553900 220556
rect 553964 220554 553970 220556
rect 563278 220554 563284 220556
rect 553964 220494 563284 220554
rect 553964 220492 553970 220494
rect 563278 220492 563284 220494
rect 563348 220492 563354 220556
rect 566825 220554 566891 220557
rect 563470 220552 566891 220554
rect 563470 220496 566830 220552
rect 566886 220496 566891 220552
rect 563470 220494 566891 220496
rect 556470 220282 556476 220284
rect 553350 220222 556476 220282
rect 543844 220220 543850 220222
rect 553025 220219 553091 220222
rect 556470 220220 556476 220222
rect 556540 220220 556546 220284
rect 556705 220282 556771 220285
rect 562501 220282 562567 220285
rect 556705 220280 562567 220282
rect 556705 220224 556710 220280
rect 556766 220224 562506 220280
rect 562562 220224 562567 220280
rect 556705 220222 562567 220224
rect 556705 220219 556771 220222
rect 562501 220219 562567 220222
rect 562869 220282 562935 220285
rect 563470 220282 563530 220494
rect 566825 220491 566891 220494
rect 567009 220554 567075 220557
rect 577681 220554 577747 220557
rect 567009 220552 577747 220554
rect 567009 220496 567014 220552
rect 567070 220496 577686 220552
rect 577742 220496 577747 220552
rect 567009 220494 577747 220496
rect 567009 220491 567075 220494
rect 577681 220491 577747 220494
rect 582189 220418 582255 220421
rect 582373 220418 582439 220421
rect 582189 220416 582439 220418
rect 582189 220360 582194 220416
rect 582250 220360 582378 220416
rect 582434 220360 582439 220416
rect 582189 220358 582439 220360
rect 582189 220355 582255 220358
rect 582373 220355 582439 220358
rect 591849 220418 591915 220421
rect 592125 220418 592191 220421
rect 591849 220416 592191 220418
rect 591849 220360 591854 220416
rect 591910 220360 592130 220416
rect 592186 220360 592191 220416
rect 591849 220358 592191 220360
rect 591849 220355 591915 220358
rect 592125 220355 592191 220358
rect 643185 220418 643251 220421
rect 664253 220418 664319 220421
rect 643185 220416 664319 220418
rect 643185 220360 643190 220416
rect 643246 220360 664258 220416
rect 664314 220360 664319 220416
rect 643185 220358 664319 220360
rect 643185 220355 643251 220358
rect 664253 220355 664319 220358
rect 669270 220358 673378 220418
rect 562869 220280 563530 220282
rect 562869 220224 562874 220280
rect 562930 220224 563530 220280
rect 562869 220222 563530 220224
rect 562869 220219 562935 220222
rect 563830 220220 563836 220284
rect 563900 220282 563906 220284
rect 572989 220282 573055 220285
rect 563900 220280 573055 220282
rect 563900 220224 572994 220280
rect 573050 220224 573055 220280
rect 563900 220222 573055 220224
rect 563900 220220 563906 220222
rect 572989 220219 573055 220222
rect 573214 220220 573220 220284
rect 573284 220282 573290 220284
rect 575841 220282 575907 220285
rect 610801 220282 610867 220285
rect 573284 220280 575907 220282
rect 573284 220224 575846 220280
rect 575902 220224 575907 220280
rect 573284 220222 575907 220224
rect 573284 220220 573290 220222
rect 575841 220219 575907 220222
rect 605790 220280 610867 220282
rect 605790 220224 610806 220280
rect 610862 220224 610867 220280
rect 605790 220222 610867 220224
rect 605790 220010 605850 220222
rect 610801 220219 610867 220222
rect 641437 220146 641503 220149
rect 669270 220146 669330 220358
rect 641437 220144 669330 220146
rect 641437 220088 641442 220144
rect 641498 220088 669330 220144
rect 641437 220086 669330 220088
rect 641437 220083 641503 220086
rect 670734 220084 670740 220148
rect 670804 220146 670810 220148
rect 671981 220146 672047 220149
rect 670804 220144 672047 220146
rect 670804 220088 671986 220144
rect 672042 220088 672047 220144
rect 670804 220086 672047 220088
rect 670804 220084 670810 220086
rect 671981 220083 672047 220086
rect 617057 220010 617123 220013
rect 534030 219950 605850 220010
rect 610574 220008 617123 220010
rect 610574 219952 617062 220008
rect 617118 219952 617123 220008
rect 610574 219950 617123 219952
rect 673318 220010 673378 220358
rect 673545 220282 673611 220285
rect 674097 220282 674163 220285
rect 673545 220280 674163 220282
rect 673545 220224 673550 220280
rect 673606 220224 674102 220280
rect 674158 220224 674163 220280
rect 673545 220222 674163 220224
rect 673545 220219 673611 220222
rect 674097 220219 674163 220222
rect 674422 220146 674482 220630
rect 676029 220627 676095 220630
rect 679617 220627 679683 220630
rect 674598 220356 674604 220420
rect 674668 220418 674674 220420
rect 676029 220418 676095 220421
rect 674668 220416 676095 220418
rect 674668 220360 676034 220416
rect 676090 220360 676095 220416
rect 674668 220358 676095 220360
rect 674668 220356 674674 220358
rect 676029 220355 676095 220358
rect 676170 220222 676292 220282
rect 674238 220086 674482 220146
rect 674238 220010 674298 220086
rect 674782 220084 674788 220148
rect 674852 220146 674858 220148
rect 676170 220146 676230 220222
rect 674852 220086 676230 220146
rect 674852 220084 674858 220086
rect 673318 219950 674298 220010
rect 530301 219947 530367 219948
rect 610574 219738 610634 219950
rect 617057 219947 617123 219950
rect 683481 219874 683547 219877
rect 683468 219872 683547 219874
rect 683468 219816 683486 219872
rect 683542 219816 683547 219872
rect 683468 219814 683547 219816
rect 683481 219811 683547 219814
rect 522573 219680 522578 219736
rect 522573 219676 522620 219680
rect 522684 219678 522730 219738
rect 524370 219678 610634 219738
rect 610801 219738 610867 219741
rect 630949 219738 631015 219741
rect 610801 219736 631015 219738
rect 610801 219680 610806 219736
rect 610862 219680 630954 219736
rect 631010 219680 631015 219736
rect 610801 219678 631015 219680
rect 522684 219676 522690 219678
rect 519813 219675 519879 219676
rect 522573 219675 522639 219676
rect 610801 219675 610867 219678
rect 630949 219675 631015 219678
rect 664253 219738 664319 219741
rect 675017 219738 675083 219741
rect 664253 219736 675083 219738
rect 664253 219680 664258 219736
rect 664314 219680 675022 219736
rect 675078 219680 675083 219736
rect 664253 219678 675083 219680
rect 664253 219675 664319 219678
rect 675017 219675 675083 219678
rect 140773 219602 140839 219605
rect 142153 219602 142219 219605
rect 140773 219600 142219 219602
rect 140773 219544 140778 219600
rect 140834 219544 142158 219600
rect 142214 219544 142219 219600
rect 140773 219542 142219 219544
rect 140773 219539 140839 219542
rect 142153 219539 142219 219542
rect 484577 219466 484643 219469
rect 630765 219466 630831 219469
rect 484577 219464 630831 219466
rect 484577 219408 484582 219464
rect 484638 219408 630770 219464
rect 630826 219408 630831 219464
rect 484577 219406 630831 219408
rect 484577 219403 484643 219406
rect 630765 219403 630831 219406
rect 671889 219466 671955 219469
rect 671889 219464 676292 219466
rect 671889 219408 671894 219464
rect 671950 219408 676292 219464
rect 671889 219406 676292 219408
rect 671889 219403 671955 219406
rect 148409 219330 148475 219333
rect 152917 219330 152983 219333
rect 148409 219328 152983 219330
rect 148409 219272 148414 219328
rect 148470 219272 152922 219328
rect 152978 219272 152983 219328
rect 148409 219270 152983 219272
rect 148409 219267 148475 219270
rect 152917 219267 152983 219270
rect 166257 219330 166323 219333
rect 169109 219330 169175 219333
rect 166257 219328 169175 219330
rect 166257 219272 166262 219328
rect 166318 219272 169114 219328
rect 169170 219272 169175 219328
rect 166257 219270 169175 219272
rect 166257 219267 166323 219270
rect 169109 219267 169175 219270
rect 195053 219330 195119 219333
rect 196065 219330 196131 219333
rect 195053 219328 196131 219330
rect 195053 219272 195058 219328
rect 195114 219272 196070 219328
rect 196126 219272 196131 219328
rect 195053 219270 196131 219272
rect 195053 219267 195119 219270
rect 196065 219267 196131 219270
rect 490557 219194 490623 219197
rect 491109 219194 491175 219197
rect 490557 219192 491175 219194
rect 490557 219136 490562 219192
rect 490618 219136 491114 219192
rect 491170 219136 491175 219192
rect 490557 219134 491175 219136
rect 490557 219131 490623 219134
rect 491109 219131 491175 219134
rect 492949 219194 493015 219197
rect 493593 219194 493659 219197
rect 492949 219192 493659 219194
rect 492949 219136 492954 219192
rect 493010 219136 493598 219192
rect 493654 219136 493659 219192
rect 492949 219134 493659 219136
rect 492949 219131 493015 219134
rect 493593 219131 493659 219134
rect 497733 219194 497799 219197
rect 502517 219194 502583 219197
rect 497733 219192 502583 219194
rect 497733 219136 497738 219192
rect 497794 219136 502522 219192
rect 502578 219136 502583 219192
rect 497733 219134 502583 219136
rect 497733 219131 497799 219134
rect 502517 219131 502583 219134
rect 502701 219194 502767 219197
rect 505093 219194 505159 219197
rect 502701 219192 505159 219194
rect 502701 219136 502706 219192
rect 502762 219136 505098 219192
rect 505154 219136 505159 219192
rect 502701 219134 505159 219136
rect 502701 219131 502767 219134
rect 505093 219131 505159 219134
rect 505277 219194 505343 219197
rect 514477 219194 514543 219197
rect 514753 219196 514819 219197
rect 514702 219194 514708 219196
rect 505277 219192 514543 219194
rect 505277 219136 505282 219192
rect 505338 219136 514482 219192
rect 514538 219136 514543 219192
rect 505277 219134 514543 219136
rect 514626 219134 514708 219194
rect 514772 219192 514819 219196
rect 514814 219136 514819 219192
rect 505277 219131 505343 219134
rect 514477 219131 514543 219134
rect 514702 219132 514708 219134
rect 514772 219132 514819 219136
rect 514753 219131 514819 219132
rect 516593 219194 516659 219197
rect 524413 219194 524479 219197
rect 516593 219192 524479 219194
rect 516593 219136 516598 219192
rect 516654 219136 524418 219192
rect 524474 219136 524479 219192
rect 516593 219134 524479 219136
rect 516593 219131 516659 219134
rect 524413 219131 524479 219134
rect 524597 219194 524663 219197
rect 534165 219194 534231 219197
rect 524597 219192 534231 219194
rect 524597 219136 524602 219192
rect 524658 219136 534170 219192
rect 534226 219136 534231 219192
rect 524597 219134 534231 219136
rect 524597 219131 524663 219134
rect 534165 219131 534231 219134
rect 534625 219194 534691 219197
rect 542353 219194 542419 219197
rect 534625 219192 542419 219194
rect 534625 219136 534630 219192
rect 534686 219136 542358 219192
rect 542414 219136 542419 219192
rect 534625 219134 542419 219136
rect 534625 219131 534691 219134
rect 542353 219131 542419 219134
rect 543365 219194 543431 219197
rect 553158 219194 553164 219196
rect 543365 219192 553164 219194
rect 543365 219136 543370 219192
rect 543426 219136 553164 219192
rect 543365 219134 553164 219136
rect 543365 219131 543431 219134
rect 553158 219132 553164 219134
rect 553228 219132 553234 219196
rect 553526 219132 553532 219196
rect 553596 219194 553602 219196
rect 567653 219194 567719 219197
rect 553596 219192 567719 219194
rect 553596 219136 567658 219192
rect 567714 219136 567719 219192
rect 553596 219134 567719 219136
rect 553596 219132 553602 219134
rect 567653 219131 567719 219134
rect 567878 219132 567884 219196
rect 567948 219194 567954 219196
rect 592125 219194 592191 219197
rect 567948 219192 592191 219194
rect 567948 219136 592130 219192
rect 592186 219136 592191 219192
rect 567948 219134 592191 219136
rect 567948 219132 567954 219134
rect 592125 219131 592191 219134
rect 592309 219194 592375 219197
rect 596541 219194 596607 219197
rect 603073 219194 603139 219197
rect 592309 219192 596607 219194
rect 592309 219136 592314 219192
rect 592370 219136 596546 219192
rect 596602 219136 596607 219192
rect 592309 219134 596607 219136
rect 592309 219131 592375 219134
rect 596541 219131 596607 219134
rect 596774 219192 603139 219194
rect 596774 219136 603078 219192
rect 603134 219136 603139 219192
rect 596774 219134 603139 219136
rect 152089 218922 152155 218925
rect 153837 218922 153903 218925
rect 152089 218920 153903 218922
rect 152089 218864 152094 218920
rect 152150 218864 153842 218920
rect 153898 218864 153903 218920
rect 152089 218862 153903 218864
rect 152089 218859 152155 218862
rect 153837 218859 153903 218862
rect 166073 218922 166139 218925
rect 167085 218922 167151 218925
rect 166073 218920 167151 218922
rect 166073 218864 166078 218920
rect 166134 218864 167090 218920
rect 167146 218864 167151 218920
rect 166073 218862 167151 218864
rect 166073 218859 166139 218862
rect 167085 218859 167151 218862
rect 490281 218922 490347 218925
rect 596774 218922 596834 219134
rect 603073 219131 603139 219134
rect 638861 219194 638927 219197
rect 674598 219194 674604 219196
rect 638861 219192 674604 219194
rect 638861 219136 638866 219192
rect 638922 219136 674604 219192
rect 638861 219134 674604 219136
rect 638861 219131 638927 219134
rect 674598 219132 674604 219134
rect 674668 219132 674674 219196
rect 674833 219058 674899 219061
rect 674833 219056 676292 219058
rect 674833 219000 674838 219056
rect 674894 219000 676292 219056
rect 674833 218998 676292 219000
rect 674833 218995 674899 218998
rect 490281 218920 596834 218922
rect 490281 218864 490286 218920
rect 490342 218864 596834 218920
rect 490281 218862 596834 218864
rect 597001 218922 597067 218925
rect 640057 218922 640123 218925
rect 597001 218920 615510 218922
rect 597001 218864 597006 218920
rect 597062 218864 615510 218920
rect 597001 218862 615510 218864
rect 490281 218859 490347 218862
rect 597001 218859 597067 218862
rect 142245 218786 142311 218789
rect 148593 218786 148659 218789
rect 142245 218784 148659 218786
rect 142245 218728 142250 218784
rect 142306 218728 148598 218784
rect 148654 218728 148659 218784
rect 142245 218726 148659 218728
rect 142245 218723 142311 218726
rect 148593 218723 148659 218726
rect 505277 218684 505343 218687
rect 505277 218682 505570 218684
rect 157241 218650 157307 218653
rect 491109 218650 491175 218653
rect 504817 218650 504883 218653
rect 157241 218648 157350 218650
rect 157241 218592 157246 218648
rect 157302 218592 157350 218648
rect 157241 218587 157350 218592
rect 491109 218648 504883 218650
rect 491109 218592 491114 218648
rect 491170 218592 504822 218648
rect 504878 218592 504883 218648
rect 505277 218626 505282 218682
rect 505338 218650 505570 218682
rect 614481 218650 614547 218653
rect 505338 218648 614547 218650
rect 505338 218626 614486 218648
rect 505277 218624 614486 218626
rect 505277 218621 505343 218624
rect 491109 218590 504883 218592
rect 505510 218592 614486 218624
rect 614542 218592 614547 218648
rect 505510 218590 614547 218592
rect 615450 218650 615510 218862
rect 640057 218920 673930 218922
rect 640057 218864 640062 218920
rect 640118 218864 673930 218920
rect 640057 218862 673930 218864
rect 640057 218859 640123 218862
rect 631133 218650 631199 218653
rect 615450 218648 631199 218650
rect 615450 218592 631138 218648
rect 631194 218592 631199 218648
rect 615450 218590 631199 218592
rect 491109 218587 491175 218590
rect 504817 218587 504883 218590
rect 614481 218587 614547 218590
rect 631133 218587 631199 218590
rect 649901 218650 649967 218653
rect 673545 218650 673611 218653
rect 649901 218648 673611 218650
rect 649901 218592 649906 218648
rect 649962 218592 673550 218648
rect 673606 218592 673611 218648
rect 649901 218590 673611 218592
rect 649901 218587 649967 218590
rect 673545 218587 673611 218590
rect 157290 218514 157350 218587
rect 157701 218514 157767 218517
rect 157290 218512 157767 218514
rect 157290 218456 157706 218512
rect 157762 218456 157767 218512
rect 157290 218454 157767 218456
rect 157701 218451 157767 218454
rect 496905 218378 496971 218381
rect 500033 218378 500099 218381
rect 496905 218376 500099 218378
rect 496905 218320 496910 218376
rect 496966 218320 500038 218376
rect 500094 218320 500099 218376
rect 496905 218318 500099 218320
rect 496905 218315 496971 218318
rect 500033 218315 500099 218318
rect 500217 218378 500283 218381
rect 504633 218378 504699 218381
rect 500217 218376 504699 218378
rect 500217 218320 500222 218376
rect 500278 218320 504638 218376
rect 504694 218320 504699 218376
rect 500217 218318 504699 218320
rect 500217 218315 500283 218318
rect 504633 218315 504699 218318
rect 507301 218378 507367 218381
rect 514334 218378 514340 218380
rect 507301 218376 514340 218378
rect 507301 218320 507306 218376
rect 507362 218320 514340 218376
rect 507301 218318 514340 218320
rect 507301 218315 507367 218318
rect 514334 218316 514340 218318
rect 514404 218316 514410 218380
rect 524137 218378 524203 218381
rect 514710 218376 524203 218378
rect 514710 218347 524142 218376
rect 514661 218342 524142 218347
rect 514661 218286 514666 218342
rect 514722 218320 524142 218342
rect 524198 218320 524203 218376
rect 514722 218318 524203 218320
rect 514722 218286 514770 218318
rect 524137 218315 524203 218318
rect 524597 218378 524663 218381
rect 533705 218378 533771 218381
rect 524597 218376 533771 218378
rect 524597 218320 524602 218376
rect 524658 218320 533710 218376
rect 533766 218320 533771 218376
rect 524597 218318 533771 218320
rect 524597 218315 524663 218318
rect 533705 218315 533771 218318
rect 533889 218378 533955 218381
rect 543774 218378 543780 218380
rect 533889 218376 543780 218378
rect 533889 218320 533894 218376
rect 533950 218320 543780 218376
rect 533889 218318 543780 218320
rect 533889 218315 533955 218318
rect 543774 218316 543780 218318
rect 543844 218316 543850 218380
rect 544009 218378 544075 218381
rect 553894 218378 553900 218380
rect 544009 218376 553900 218378
rect 544009 218320 544014 218376
rect 544070 218320 553900 218376
rect 544009 218318 553900 218320
rect 544009 218315 544075 218318
rect 553894 218316 553900 218318
rect 553964 218316 553970 218380
rect 554078 218316 554084 218380
rect 554148 218378 554154 218380
rect 558361 218378 558427 218381
rect 554148 218376 558427 218378
rect 554148 218320 558366 218376
rect 558422 218320 558427 218376
rect 554148 218318 558427 218320
rect 554148 218316 554154 218318
rect 558361 218315 558427 218318
rect 558545 218378 558611 218381
rect 567878 218378 567884 218380
rect 558545 218376 567884 218378
rect 558545 218320 558550 218376
rect 558606 218320 567884 218376
rect 558545 218318 567884 218320
rect 558545 218315 558611 218318
rect 567878 218316 567884 218318
rect 567948 218316 567954 218380
rect 568113 218378 568179 218381
rect 571609 218378 571675 218381
rect 568113 218376 571675 218378
rect 568113 218320 568118 218376
rect 568174 218320 571614 218376
rect 571670 218320 571675 218376
rect 568113 218318 571675 218320
rect 568113 218315 568179 218318
rect 571609 218315 571675 218318
rect 572110 218316 572116 218380
rect 572180 218378 572186 218380
rect 582097 218378 582163 218381
rect 572180 218376 582163 218378
rect 572180 218320 582102 218376
rect 582158 218320 582163 218376
rect 572180 218318 582163 218320
rect 572180 218316 572186 218318
rect 582097 218315 582163 218318
rect 582281 218378 582347 218381
rect 582741 218378 582807 218381
rect 582281 218376 582807 218378
rect 582281 218320 582286 218376
rect 582342 218320 582746 218376
rect 582802 218320 582807 218376
rect 582281 218318 582807 218320
rect 582281 218315 582347 218318
rect 582741 218315 582807 218318
rect 582925 218378 582991 218381
rect 591941 218378 592007 218381
rect 582925 218376 592007 218378
rect 582925 218320 582930 218376
rect 582986 218320 591946 218376
rect 592002 218320 592007 218376
rect 582925 218318 592007 218320
rect 582925 218315 582991 218318
rect 591941 218315 592007 218318
rect 592125 218378 592191 218381
rect 629937 218378 630003 218381
rect 592125 218376 630003 218378
rect 592125 218320 592130 218376
rect 592186 218320 629942 218376
rect 629998 218320 630003 218376
rect 592125 218318 630003 218320
rect 673870 218378 673930 218862
rect 674966 218588 674972 218652
rect 675036 218650 675042 218652
rect 675036 218590 676292 218650
rect 675036 218588 675042 218590
rect 675661 218378 675727 218381
rect 673870 218376 675727 218378
rect 673870 218320 675666 218376
rect 675722 218320 675727 218376
rect 673870 218318 675727 218320
rect 592125 218315 592191 218318
rect 629937 218315 630003 218318
rect 675661 218315 675727 218318
rect 514661 218284 514770 218286
rect 514661 218281 514727 218284
rect 159633 218242 159699 218245
rect 162853 218242 162919 218245
rect 159633 218240 162919 218242
rect 159633 218184 159638 218240
rect 159694 218184 162858 218240
rect 162914 218184 162919 218240
rect 159633 218182 162919 218184
rect 159633 218179 159699 218182
rect 162853 218179 162919 218182
rect 675886 218180 675892 218244
rect 675956 218242 675962 218244
rect 675956 218182 676292 218242
rect 675956 218180 675962 218182
rect 487797 218106 487863 218109
rect 534073 218106 534139 218109
rect 487797 218104 534139 218106
rect 487797 218048 487802 218104
rect 487858 218048 534078 218104
rect 534134 218048 534139 218104
rect 487797 218046 534139 218048
rect 487797 218043 487863 218046
rect 534073 218043 534139 218046
rect 534257 218106 534323 218109
rect 543457 218106 543523 218109
rect 534257 218104 543523 218106
rect 534257 218048 534262 218104
rect 534318 218048 543462 218104
rect 543518 218048 543523 218104
rect 534257 218046 543523 218048
rect 534257 218043 534323 218046
rect 543457 218043 543523 218046
rect 543641 218106 543707 218109
rect 582925 218106 582991 218109
rect 591849 218106 591915 218109
rect 626441 218106 626507 218109
rect 543641 218104 582666 218106
rect 543641 218048 543646 218104
rect 543702 218048 582666 218104
rect 543641 218046 582666 218048
rect 543641 218043 543707 218046
rect 35525 217970 35591 217973
rect 54477 217970 54543 217973
rect 35525 217968 54543 217970
rect 35525 217912 35530 217968
rect 35586 217912 54482 217968
rect 54538 217912 54543 217968
rect 35525 217910 54543 217912
rect 582606 217970 582666 218046
rect 582925 218104 591915 218106
rect 582925 218048 582930 218104
rect 582986 218048 591854 218104
rect 591910 218048 591915 218104
rect 582925 218046 591915 218048
rect 582925 218043 582991 218046
rect 591849 218043 591915 218046
rect 598890 218104 626507 218106
rect 598890 218048 626446 218104
rect 626502 218048 626507 218104
rect 598890 218046 626507 218048
rect 592125 217970 592191 217973
rect 598890 217970 598950 218046
rect 626441 218043 626507 218046
rect 582606 217910 582850 217970
rect 35525 217907 35591 217910
rect 54477 217907 54543 217910
rect 504817 217834 504883 217837
rect 505461 217834 505527 217837
rect 504817 217832 505527 217834
rect 504817 217776 504822 217832
rect 504878 217776 505466 217832
rect 505522 217776 505527 217832
rect 504817 217774 505527 217776
rect 504817 217771 504883 217774
rect 505461 217771 505527 217774
rect 508497 217834 508563 217837
rect 524413 217834 524479 217837
rect 508497 217832 524479 217834
rect 508497 217776 508502 217832
rect 508558 217776 524418 217832
rect 524474 217776 524479 217832
rect 508497 217774 524479 217776
rect 508497 217771 508563 217774
rect 524413 217771 524479 217774
rect 524597 217834 524663 217837
rect 563053 217834 563119 217837
rect 524597 217832 563119 217834
rect 524597 217776 524602 217832
rect 524658 217776 563058 217832
rect 563114 217776 563119 217832
rect 524597 217774 563119 217776
rect 524597 217771 524663 217774
rect 563053 217771 563119 217774
rect 563237 217834 563303 217837
rect 563830 217834 563836 217836
rect 563237 217832 563836 217834
rect 563237 217776 563242 217832
rect 563298 217776 563836 217832
rect 563237 217774 563836 217776
rect 563237 217771 563303 217774
rect 563830 217772 563836 217774
rect 563900 217772 563906 217836
rect 564014 217772 564020 217836
rect 564084 217834 564090 217836
rect 564341 217834 564407 217837
rect 564084 217832 564407 217834
rect 564084 217776 564346 217832
rect 564402 217776 564407 217832
rect 564084 217774 564407 217776
rect 564084 217772 564090 217774
rect 564341 217771 564407 217774
rect 564525 217834 564591 217837
rect 571149 217834 571215 217837
rect 564525 217832 571215 217834
rect 564525 217776 564530 217832
rect 564586 217776 571154 217832
rect 571210 217776 571215 217832
rect 564525 217774 571215 217776
rect 564525 217771 564591 217774
rect 571149 217771 571215 217774
rect 572110 217772 572116 217836
rect 572180 217834 572186 217836
rect 574369 217834 574435 217837
rect 572180 217832 574435 217834
rect 572180 217776 574374 217832
rect 574430 217776 574435 217832
rect 572180 217774 574435 217776
rect 572180 217772 572186 217774
rect 574369 217771 574435 217774
rect 574553 217834 574619 217837
rect 582373 217834 582439 217837
rect 574553 217832 582439 217834
rect 574553 217776 574558 217832
rect 574614 217776 582378 217832
rect 582434 217776 582439 217832
rect 574553 217774 582439 217776
rect 582790 217834 582850 217910
rect 592125 217968 598950 217970
rect 592125 217912 592130 217968
rect 592186 217912 598950 217968
rect 592125 217910 598950 217912
rect 592125 217907 592191 217910
rect 591665 217834 591731 217837
rect 582790 217832 591731 217834
rect 582790 217776 591670 217832
rect 591726 217776 591731 217832
rect 582790 217774 591731 217776
rect 574553 217771 574619 217774
rect 582373 217771 582439 217774
rect 591665 217771 591731 217774
rect 675017 217834 675083 217837
rect 675017 217832 676292 217834
rect 675017 217776 675022 217832
rect 675078 217776 676292 217832
rect 675017 217774 676292 217776
rect 675017 217771 675083 217774
rect 498653 217562 498719 217565
rect 500718 217562 500724 217564
rect 498653 217560 500724 217562
rect 498653 217504 498658 217560
rect 498714 217504 500724 217560
rect 498653 217502 500724 217504
rect 498653 217499 498719 217502
rect 500718 217500 500724 217502
rect 500788 217500 500794 217564
rect 503529 217562 503595 217565
rect 504766 217562 504772 217564
rect 503529 217560 504772 217562
rect 503529 217504 503534 217560
rect 503590 217504 504772 217560
rect 503529 217502 504772 217504
rect 503529 217499 503595 217502
rect 504766 217500 504772 217502
rect 504836 217500 504842 217564
rect 506013 217562 506079 217565
rect 590101 217562 590167 217565
rect 506013 217560 590167 217562
rect 506013 217504 506018 217560
rect 506074 217504 590106 217560
rect 590162 217504 590167 217560
rect 506013 217502 590167 217504
rect 506013 217499 506079 217502
rect 590101 217499 590167 217502
rect 644933 217562 644999 217565
rect 672206 217562 672212 217564
rect 644933 217560 672212 217562
rect 644933 217504 644938 217560
rect 644994 217504 672212 217560
rect 644933 217502 672212 217504
rect 644933 217499 644999 217502
rect 672206 217500 672212 217502
rect 672276 217500 672282 217564
rect 675518 217364 675524 217428
rect 675588 217426 675594 217428
rect 675588 217366 676292 217426
rect 675588 217364 675594 217366
rect 493593 217292 493659 217293
rect 493542 217290 493548 217292
rect 493502 217230 493548 217290
rect 493612 217288 493659 217292
rect 493654 217232 493659 217288
rect 493542 217228 493548 217230
rect 493612 217228 493659 217232
rect 493593 217227 493659 217228
rect 497549 217290 497615 217293
rect 541750 217290 541756 217292
rect 497549 217288 541756 217290
rect 497549 217232 497554 217288
rect 497610 217232 541756 217288
rect 497549 217230 541756 217232
rect 497549 217227 497615 217230
rect 541750 217228 541756 217230
rect 541820 217228 541826 217292
rect 541985 217290 542051 217293
rect 543825 217290 543891 217293
rect 541985 217288 543891 217290
rect 541985 217232 541990 217288
rect 542046 217232 543830 217288
rect 543886 217232 543891 217288
rect 541985 217230 543891 217232
rect 541985 217227 542051 217230
rect 543825 217227 543891 217230
rect 544142 217228 544148 217292
rect 544212 217290 544218 217292
rect 572118 217290 572730 217324
rect 591757 217290 591823 217293
rect 544212 217288 591823 217290
rect 544212 217264 591762 217288
rect 544212 217230 572178 217264
rect 572670 217232 591762 217264
rect 591818 217232 591823 217288
rect 572670 217230 591823 217232
rect 544212 217228 544218 217230
rect 591757 217227 591823 217230
rect 592217 217290 592283 217293
rect 594793 217290 594859 217293
rect 592217 217288 594859 217290
rect 592217 217232 592222 217288
rect 592278 217232 594798 217288
rect 594854 217232 594859 217288
rect 592217 217230 594859 217232
rect 592217 217227 592283 217230
rect 594793 217227 594859 217230
rect 642081 217290 642147 217293
rect 675150 217290 675156 217292
rect 642081 217288 675156 217290
rect 642081 217232 642086 217288
rect 642142 217232 675156 217288
rect 642081 217230 675156 217232
rect 642081 217227 642147 217230
rect 675150 217228 675156 217230
rect 675220 217228 675226 217292
rect 492121 217154 492187 217157
rect 492121 217152 492506 217154
rect 492121 217096 492126 217152
rect 492182 217096 492506 217152
rect 492121 217094 492506 217096
rect 492121 217091 492187 217094
rect 492446 216746 492506 217094
rect 500718 216956 500724 217020
rect 500788 217018 500794 217020
rect 582327 217018 582393 217021
rect 500788 217016 582393 217018
rect 500788 216960 582332 217016
rect 582388 216960 582393 217016
rect 500788 216958 582393 216960
rect 500788 216956 500794 216958
rect 582327 216955 582393 216958
rect 582598 216956 582604 217020
rect 582668 217018 582674 217020
rect 591614 217018 591620 217020
rect 582668 216958 591620 217018
rect 582668 216956 582674 216958
rect 591614 216956 591620 216958
rect 591684 216956 591690 217020
rect 592166 216956 592172 217020
rect 592236 217018 592242 217020
rect 592236 216958 595546 217018
rect 592236 216956 592242 216958
rect 595161 216746 595227 216749
rect 492446 216744 595227 216746
rect 492446 216688 595166 216744
rect 595222 216688 595227 216744
rect 492446 216686 595227 216688
rect 595161 216683 595227 216686
rect 595486 216610 595546 216958
rect 675702 216956 675708 217020
rect 675772 217018 675778 217020
rect 675772 216958 676292 217018
rect 675772 216956 675778 216958
rect 675201 216882 675267 216885
rect 674422 216880 675267 216882
rect 674422 216824 675206 216880
rect 675262 216824 675267 216880
rect 674422 216822 675267 216824
rect 664253 216746 664319 216749
rect 664253 216744 664730 216746
rect 664253 216688 664258 216744
rect 664314 216688 664730 216744
rect 664253 216686 664730 216688
rect 664253 216683 664319 216686
rect 597553 216610 597619 216613
rect 595486 216608 597619 216610
rect 595486 216552 597558 216608
rect 597614 216552 597619 216608
rect 595486 216550 597619 216552
rect 664670 216610 664730 216686
rect 674422 216610 674482 216822
rect 675201 216819 675267 216822
rect 664670 216550 674482 216610
rect 674741 216610 674807 216613
rect 674741 216608 676292 216610
rect 674741 216552 674746 216608
rect 674802 216552 676292 216608
rect 674741 216550 676292 216552
rect 597553 216547 597619 216550
rect 674741 216547 674807 216550
rect 511022 216412 511028 216476
rect 511092 216474 511098 216476
rect 519302 216474 519308 216476
rect 511092 216414 519308 216474
rect 511092 216412 511098 216414
rect 519302 216412 519308 216414
rect 519372 216412 519378 216476
rect 519854 216412 519860 216476
rect 519924 216474 519930 216476
rect 566590 216474 566596 216476
rect 519924 216414 566596 216474
rect 519924 216412 519930 216414
rect 566590 216412 566596 216414
rect 566660 216412 566666 216476
rect 566774 216412 566780 216476
rect 566844 216474 566850 216476
rect 572110 216474 572116 216476
rect 566844 216414 572116 216474
rect 566844 216412 566850 216414
rect 572110 216412 572116 216414
rect 572180 216412 572186 216476
rect 572478 216412 572484 216476
rect 572548 216474 572554 216476
rect 577313 216474 577379 216477
rect 572548 216472 577379 216474
rect 572548 216416 577318 216472
rect 577374 216416 577379 216472
rect 572548 216414 577379 216416
rect 572548 216412 572554 216414
rect 577313 216411 577379 216414
rect 577630 216412 577636 216476
rect 577700 216474 577706 216476
rect 582373 216474 582439 216477
rect 577700 216472 582439 216474
rect 577700 216416 582378 216472
rect 582434 216416 582439 216472
rect 577700 216414 582439 216416
rect 577700 216412 577706 216414
rect 582373 216411 582439 216414
rect 582557 216474 582623 216477
rect 591757 216474 591823 216477
rect 592033 216474 592099 216477
rect 582557 216472 591823 216474
rect 582557 216416 582562 216472
rect 582618 216416 591762 216472
rect 591818 216416 591823 216472
rect 582557 216414 591823 216416
rect 582557 216411 582623 216414
rect 591757 216411 591823 216414
rect 591990 216472 592099 216474
rect 591990 216416 592038 216472
rect 592094 216416 592099 216472
rect 591990 216411 592099 216416
rect 654041 216474 654107 216477
rect 654041 216472 664546 216474
rect 654041 216416 654046 216472
rect 654102 216416 664546 216472
rect 654041 216414 664546 216416
rect 654041 216411 654107 216414
rect 504766 216140 504772 216204
rect 504836 216202 504842 216204
rect 582414 216202 582420 216204
rect 504836 216142 582420 216202
rect 504836 216140 504842 216142
rect 582414 216140 582420 216142
rect 582484 216140 582490 216204
rect 582741 216202 582807 216205
rect 591990 216202 592050 216411
rect 592217 216338 592283 216341
rect 595713 216338 595779 216341
rect 592217 216336 595779 216338
rect 592217 216280 592222 216336
rect 592278 216280 595718 216336
rect 595774 216280 595779 216336
rect 592217 216278 595779 216280
rect 592217 216275 592283 216278
rect 595713 216275 595779 216278
rect 595897 216338 595963 216341
rect 599025 216338 599091 216341
rect 595897 216336 599091 216338
rect 595897 216280 595902 216336
rect 595958 216280 599030 216336
rect 599086 216280 599091 216336
rect 595897 216278 599091 216280
rect 664486 216338 664546 216414
rect 672717 216338 672783 216341
rect 664486 216336 672783 216338
rect 664486 216280 672722 216336
rect 672778 216280 672783 216336
rect 664486 216278 672783 216280
rect 595897 216275 595963 216278
rect 599025 216275 599091 216278
rect 672717 216275 672783 216278
rect 582741 216200 592050 216202
rect 582741 216144 582746 216200
rect 582802 216144 592050 216200
rect 582741 216142 592050 216144
rect 646589 216202 646655 216205
rect 664253 216202 664319 216205
rect 646589 216200 664319 216202
rect 646589 216144 646594 216200
rect 646650 216144 664258 216200
rect 664314 216144 664319 216200
rect 646589 216142 664319 216144
rect 582741 216139 582807 216142
rect 646589 216139 646655 216142
rect 664253 216139 664319 216142
rect 673453 216202 673519 216205
rect 673453 216200 676292 216202
rect 673453 216144 673458 216200
rect 673514 216144 676292 216200
rect 673453 216142 676292 216144
rect 673453 216139 673519 216142
rect 519302 215868 519308 215932
rect 519372 215930 519378 215932
rect 529238 215930 529244 215932
rect 519372 215870 529244 215930
rect 519372 215868 519378 215870
rect 529238 215868 529244 215870
rect 529308 215868 529314 215932
rect 530342 215868 530348 215932
rect 530412 215930 530418 215932
rect 546902 215930 546908 215932
rect 530412 215870 546908 215930
rect 530412 215868 530418 215870
rect 546902 215868 546908 215870
rect 546972 215868 546978 215932
rect 548558 215868 548564 215932
rect 548628 215930 548634 215932
rect 577078 215930 577084 215932
rect 548628 215870 577084 215930
rect 548628 215868 548634 215870
rect 577078 215868 577084 215870
rect 577148 215868 577154 215932
rect 577313 215930 577379 215933
rect 611353 215930 611419 215933
rect 577313 215928 611419 215930
rect 577313 215872 577318 215928
rect 577374 215872 611358 215928
rect 611414 215872 611419 215928
rect 577313 215870 611419 215872
rect 577313 215867 577379 215870
rect 611353 215867 611419 215870
rect 643001 215930 643067 215933
rect 675334 215930 675340 215932
rect 643001 215928 675340 215930
rect 643001 215872 643006 215928
rect 643062 215872 675340 215928
rect 643001 215870 675340 215872
rect 643001 215867 643067 215870
rect 675334 215868 675340 215870
rect 675404 215868 675410 215932
rect 547278 215734 548442 215794
rect 547278 215658 547338 215734
rect 524370 215598 547338 215658
rect 548382 215658 548442 215734
rect 676170 215734 676292 215794
rect 556470 215658 556476 215660
rect 548382 215598 556476 215658
rect 522614 215324 522620 215388
rect 522684 215386 522690 215388
rect 524370 215386 524430 215598
rect 556470 215596 556476 215598
rect 556540 215596 556546 215660
rect 556846 215598 558010 215658
rect 556846 215522 556906 215598
rect 547462 215462 548258 215522
rect 522684 215326 524430 215386
rect 522684 215324 522690 215326
rect 529238 215324 529244 215388
rect 529308 215386 529314 215388
rect 536966 215386 536972 215388
rect 529308 215326 536972 215386
rect 529308 215324 529314 215326
rect 536966 215324 536972 215326
rect 537036 215324 537042 215388
rect 538622 215324 538628 215388
rect 538692 215386 538698 215388
rect 547462 215386 547522 215462
rect 538692 215326 547522 215386
rect 548198 215386 548258 215462
rect 556708 215462 556906 215522
rect 557950 215522 558010 215598
rect 558310 215596 558316 215660
rect 558380 215658 558386 215660
rect 618897 215658 618963 215661
rect 558380 215656 618963 215658
rect 558380 215600 618902 215656
rect 618958 215600 618963 215656
rect 558380 215598 618963 215600
rect 558380 215596 558386 215598
rect 618897 215595 618963 215598
rect 666318 215596 666324 215660
rect 666388 215658 666394 215660
rect 676170 215658 676230 215734
rect 666388 215598 676230 215658
rect 666388 215596 666394 215598
rect 557950 215462 558194 215522
rect 556708 215386 556768 215462
rect 548198 215326 556768 215386
rect 558134 215386 558194 215462
rect 566774 215386 566780 215388
rect 558134 215326 566780 215386
rect 538692 215324 538698 215326
rect 566774 215324 566780 215326
rect 566844 215324 566850 215388
rect 620553 215386 620619 215389
rect 566966 215384 620619 215386
rect 566966 215328 620558 215384
rect 620614 215328 620619 215384
rect 566966 215326 620619 215328
rect 547646 215250 548074 215310
rect 529974 215052 529980 215116
rect 530044 215114 530050 215116
rect 547646 215114 547706 215250
rect 530044 215054 547706 215114
rect 548014 215114 548074 215250
rect 566966 215114 567026 215326
rect 620553 215323 620619 215326
rect 674557 215386 674623 215389
rect 674782 215386 674788 215388
rect 674557 215384 674788 215386
rect 674557 215328 674562 215384
rect 674618 215328 674788 215384
rect 674557 215326 674788 215328
rect 674557 215323 674623 215326
rect 674782 215324 674788 215326
rect 674852 215324 674858 215388
rect 675201 215386 675267 215389
rect 675201 215384 676292 215386
rect 675201 215328 675206 215384
rect 675262 215328 676292 215384
rect 675201 215326 676292 215328
rect 675201 215323 675267 215326
rect 548014 215054 567026 215114
rect 530044 215052 530050 215054
rect 568246 215052 568252 215116
rect 568316 215114 568322 215116
rect 577037 215114 577103 215117
rect 568316 215112 577103 215114
rect 568316 215056 577042 215112
rect 577098 215056 577103 215112
rect 568316 215054 577103 215056
rect 568316 215052 568322 215054
rect 577037 215051 577103 215054
rect 659653 215114 659719 215117
rect 675937 215114 676003 215117
rect 659653 215112 676003 215114
rect 659653 215056 659658 215112
rect 659714 215056 675942 215112
rect 675998 215056 676003 215112
rect 676254 215086 676260 215150
rect 676324 215086 676330 215150
rect 659653 215054 676003 215056
rect 659653 215051 659719 215054
rect 675937 215051 676003 215054
rect 44817 214978 44883 214981
rect 41492 214976 44883 214978
rect 41492 214920 44822 214976
rect 44878 214920 44883 214976
rect 676262 214948 676322 215086
rect 41492 214918 44883 214920
rect 44817 214915 44883 214918
rect 651281 214842 651347 214845
rect 672073 214842 672139 214845
rect 651281 214840 672139 214842
rect 651281 214784 651286 214840
rect 651342 214784 672078 214840
rect 672134 214784 672139 214840
rect 651281 214782 672139 214784
rect 651281 214779 651347 214782
rect 672073 214779 672139 214782
rect 672533 214842 672599 214845
rect 673126 214842 673132 214844
rect 672533 214840 673132 214842
rect 672533 214784 672538 214840
rect 672594 214784 673132 214840
rect 672533 214782 673132 214784
rect 672533 214779 672599 214782
rect 673126 214780 673132 214782
rect 673196 214780 673202 214844
rect 647141 214570 647207 214573
rect 675661 214570 675727 214573
rect 647141 214568 675727 214570
rect 35758 214301 35818 214540
rect 647141 214512 647146 214568
rect 647202 214512 675666 214568
rect 675722 214512 675727 214568
rect 647141 214510 675727 214512
rect 647141 214507 647207 214510
rect 675661 214507 675727 214510
rect 675886 214508 675892 214572
rect 675956 214570 675962 214572
rect 675956 214510 676292 214570
rect 675956 214508 675962 214510
rect 35525 214298 35591 214301
rect 35525 214296 35634 214298
rect 35525 214240 35530 214296
rect 35586 214240 35634 214296
rect 35525 214235 35634 214240
rect 35758 214296 35867 214301
rect 35758 214240 35806 214296
rect 35862 214240 35867 214296
rect 35758 214238 35867 214240
rect 35801 214235 35867 214238
rect 35574 214132 35634 214235
rect 575982 214026 576042 214404
rect 669405 214162 669471 214165
rect 669405 214160 676292 214162
rect 669405 214104 669410 214160
rect 669466 214104 676292 214160
rect 669405 214102 676292 214104
rect 669405 214099 669471 214102
rect 578877 214026 578943 214029
rect 575982 214024 578943 214026
rect 575982 213968 578882 214024
rect 578938 213968 578943 214024
rect 575982 213966 578943 213968
rect 578877 213963 578943 213966
rect 43713 213754 43779 213757
rect 41492 213752 43779 213754
rect 41492 213696 43718 213752
rect 43774 213696 43779 213752
rect 41492 213694 43779 213696
rect 43713 213691 43779 213694
rect 664805 213754 664871 213757
rect 672165 213754 672231 213757
rect 664805 213752 671906 213754
rect 664805 213696 664810 213752
rect 664866 213696 671906 213752
rect 664805 213694 671906 213696
rect 664805 213691 664871 213694
rect 575657 213620 575723 213621
rect 575606 213618 575612 213620
rect 575566 213558 575612 213618
rect 575676 213616 575723 213620
rect 575718 213560 575723 213616
rect 575606 213556 575612 213558
rect 575676 213556 575723 213560
rect 575657 213555 575723 213556
rect 661493 213482 661559 213485
rect 671846 213482 671906 213694
rect 672165 213752 676292 213754
rect 672165 213696 672170 213752
rect 672226 213696 676292 213752
rect 672165 213694 676292 213696
rect 672165 213691 672231 213694
rect 676029 213482 676095 213485
rect 661493 213480 669330 213482
rect 661493 213424 661498 213480
rect 661554 213424 669330 213480
rect 661493 213422 669330 213424
rect 671846 213480 676095 213482
rect 671846 213424 676034 213480
rect 676090 213424 676095 213480
rect 671846 213422 676095 213424
rect 661493 213419 661559 213422
rect 47945 213346 48011 213349
rect 41492 213344 48011 213346
rect 41492 213288 47950 213344
rect 48006 213288 48011 213344
rect 41492 213286 48011 213288
rect 47945 213283 48011 213286
rect 642173 213210 642239 213213
rect 669270 213210 669330 213422
rect 676029 213419 676095 213422
rect 683297 213346 683363 213349
rect 683284 213344 683363 213346
rect 683284 213288 683302 213344
rect 683358 213288 683363 213344
rect 683284 213286 683363 213288
rect 683297 213283 683363 213286
rect 676029 213210 676095 213213
rect 642173 213208 663810 213210
rect 642173 213152 642178 213208
rect 642234 213152 663810 213208
rect 642173 213150 663810 213152
rect 669270 213208 676095 213210
rect 669270 213152 676034 213208
rect 676090 213152 676095 213208
rect 669270 213150 676095 213152
rect 642173 213147 642239 213150
rect 43437 212938 43503 212941
rect 41492 212936 43503 212938
rect 41492 212880 43442 212936
rect 43498 212880 43503 212936
rect 41492 212878 43503 212880
rect 663750 212938 663810 213150
rect 676029 213147 676095 213150
rect 673913 212938 673979 212941
rect 663750 212936 673979 212938
rect 663750 212880 673918 212936
rect 673974 212880 673979 212936
rect 663750 212878 673979 212880
rect 43437 212875 43503 212878
rect 673913 212875 673979 212878
rect 683070 212533 683130 212908
rect 43437 212530 43503 212533
rect 41492 212528 43503 212530
rect 41492 212472 43442 212528
rect 43498 212472 43503 212528
rect 683070 212528 683179 212533
rect 683070 212500 683118 212528
rect 41492 212470 43503 212472
rect 683100 212472 683118 212500
rect 683174 212472 683179 212528
rect 683100 212470 683179 212472
rect 43437 212467 43503 212470
rect 683113 212467 683179 212470
rect 42885 212122 42951 212125
rect 41492 212120 42951 212122
rect 41492 212064 42890 212120
rect 42946 212064 42951 212120
rect 41492 212062 42951 212064
rect 42885 212059 42951 212062
rect 575982 211714 576042 212228
rect 674046 212060 674052 212124
rect 674116 212122 674122 212124
rect 674116 212062 676292 212122
rect 674116 212060 674122 212062
rect 578509 211714 578575 211717
rect 575982 211712 578575 211714
rect 35758 211445 35818 211684
rect 575982 211656 578514 211712
rect 578570 211656 578575 211712
rect 575982 211654 578575 211656
rect 578509 211651 578575 211654
rect 35758 211440 35867 211445
rect 35758 211384 35806 211440
rect 35862 211384 35867 211440
rect 35758 211382 35867 211384
rect 35801 211379 35867 211382
rect 675886 211380 675892 211444
rect 675956 211442 675962 211444
rect 676438 211442 676444 211444
rect 675956 211382 676444 211442
rect 675956 211380 675962 211382
rect 676438 211380 676444 211382
rect 676508 211380 676514 211444
rect 44173 211306 44239 211309
rect 41492 211304 44239 211306
rect 41492 211248 44178 211304
rect 44234 211248 44239 211304
rect 41492 211246 44239 211248
rect 44173 211243 44239 211246
rect 669446 211108 669452 211172
rect 669516 211170 669522 211172
rect 670601 211170 670667 211173
rect 683113 211170 683179 211173
rect 669516 211168 670667 211170
rect 669516 211112 670606 211168
rect 670662 211112 670667 211168
rect 669516 211110 670667 211112
rect 669516 211108 669522 211110
rect 670601 211107 670667 211110
rect 670926 211168 683179 211170
rect 670926 211112 683118 211168
rect 683174 211112 683179 211168
rect 670926 211110 683179 211112
rect 48129 210898 48195 210901
rect 41492 210896 48195 210898
rect 41492 210840 48134 210896
rect 48190 210840 48195 210896
rect 41492 210838 48195 210840
rect 48129 210835 48195 210838
rect 670601 210898 670667 210901
rect 670926 210898 670986 211110
rect 683113 211107 683179 211110
rect 670601 210896 670986 210898
rect 670601 210840 670606 210896
rect 670662 210840 670986 210896
rect 670601 210838 670986 210840
rect 670601 210835 670667 210838
rect 44173 210490 44239 210493
rect 41492 210488 44239 210490
rect 41492 210432 44178 210488
rect 44234 210432 44239 210488
rect 41492 210430 44239 210432
rect 44173 210427 44239 210430
rect 674966 210428 674972 210492
rect 675036 210490 675042 210492
rect 675886 210490 675892 210492
rect 675036 210430 675892 210490
rect 675036 210428 675042 210430
rect 675886 210428 675892 210430
rect 675956 210428 675962 210492
rect 683297 210354 683363 210357
rect 678930 210352 683363 210354
rect 678930 210296 683302 210352
rect 683358 210296 683363 210352
rect 678930 210294 683363 210296
rect 672717 210218 672783 210221
rect 678930 210218 678990 210294
rect 683297 210291 683363 210294
rect 672717 210216 678990 210218
rect 672717 210160 672722 210216
rect 672778 210160 678990 210216
rect 672717 210158 678990 210160
rect 672717 210155 672783 210158
rect 41462 209812 41522 210052
rect 41454 209748 41460 209812
rect 41524 209748 41530 209812
rect 575982 209810 576042 210052
rect 579245 209810 579311 209813
rect 575982 209808 579311 209810
rect 575982 209752 579250 209808
rect 579306 209752 579311 209808
rect 575982 209750 579311 209752
rect 579245 209747 579311 209750
rect 673913 209674 673979 209677
rect 676857 209674 676923 209677
rect 673913 209672 676923 209674
rect 41278 209402 41338 209644
rect 673913 209616 673918 209672
rect 673974 209616 676862 209672
rect 676918 209616 676923 209672
rect 673913 209614 676923 209616
rect 673913 209611 673979 209614
rect 676857 209611 676923 209614
rect 42793 209402 42859 209405
rect 41278 209400 42859 209402
rect 41278 209344 42798 209400
rect 42854 209344 42859 209400
rect 41278 209342 42859 209344
rect 42793 209339 42859 209342
rect 35758 208997 35818 209236
rect 35758 208992 35867 208997
rect 35758 208936 35806 208992
rect 35862 208936 35867 208992
rect 35758 208934 35867 208936
rect 35801 208931 35867 208934
rect 41689 208994 41755 208997
rect 49509 208994 49575 208997
rect 41689 208992 49575 208994
rect 41689 208936 41694 208992
rect 41750 208936 49514 208992
rect 49570 208936 49575 208992
rect 41689 208934 49575 208936
rect 41689 208931 41755 208934
rect 49509 208931 49575 208934
rect 41462 208586 41522 208828
rect 44541 208586 44607 208589
rect 41462 208584 44607 208586
rect 41462 208528 44546 208584
rect 44602 208528 44607 208584
rect 41462 208526 44607 208528
rect 44541 208523 44607 208526
rect 40542 208180 40602 208420
rect 669221 208314 669287 208317
rect 675845 208314 675911 208317
rect 669221 208312 675911 208314
rect 669221 208256 669226 208312
rect 669282 208256 675850 208312
rect 675906 208256 675911 208312
rect 669221 208254 675911 208256
rect 669221 208251 669287 208254
rect 675845 208251 675911 208254
rect 40534 208116 40540 208180
rect 40604 208116 40610 208180
rect 43253 208042 43319 208045
rect 41492 208040 43319 208042
rect 41492 207984 43258 208040
rect 43314 207984 43319 208040
rect 41492 207982 43319 207984
rect 43253 207979 43319 207982
rect 589457 208042 589523 208045
rect 589457 208040 592572 208042
rect 589457 207984 589462 208040
rect 589518 207984 592572 208040
rect 589457 207982 592572 207984
rect 589457 207979 589523 207982
rect 40033 207770 40099 207773
rect 42374 207770 42380 207772
rect 40033 207768 42380 207770
rect 40033 207712 40038 207768
rect 40094 207712 42380 207768
rect 40033 207710 42380 207712
rect 40033 207707 40099 207710
rect 42374 207708 42380 207710
rect 42444 207708 42450 207772
rect 40910 207364 40970 207604
rect 575982 207498 576042 207876
rect 579521 207498 579587 207501
rect 575982 207496 579587 207498
rect 575982 207440 579526 207496
rect 579582 207440 579587 207496
rect 575982 207438 579587 207440
rect 579521 207435 579587 207438
rect 40902 207300 40908 207364
rect 40972 207300 40978 207364
rect 669221 207362 669287 207365
rect 666694 207360 669287 207362
rect 666694 207304 669226 207360
rect 669282 207304 669287 207360
rect 666694 207302 669287 207304
rect 666694 207294 666754 207302
rect 669221 207299 669287 207302
rect 666356 207234 666754 207294
rect 40726 206956 40786 207196
rect 40718 206892 40724 206956
rect 40788 206892 40794 206956
rect 673545 206954 673611 206957
rect 677777 206954 677843 206957
rect 673545 206952 677843 206954
rect 673545 206896 673550 206952
rect 673606 206896 677782 206952
rect 677838 206896 677843 206952
rect 673545 206894 677843 206896
rect 673545 206891 673611 206894
rect 677777 206891 677843 206894
rect 43805 206818 43871 206821
rect 41492 206816 43871 206818
rect 41492 206760 43810 206816
rect 43866 206760 43871 206816
rect 41492 206758 43871 206760
rect 43805 206755 43871 206758
rect 42977 206410 43043 206413
rect 41492 206408 43043 206410
rect 41492 206352 42982 206408
rect 43038 206352 43043 206408
rect 41492 206350 43043 206352
rect 42977 206347 43043 206350
rect 589457 206410 589523 206413
rect 589457 206408 592572 206410
rect 589457 206352 589462 206408
rect 589518 206352 592572 206408
rect 589457 206350 592572 206352
rect 589457 206347 589523 206350
rect 43437 206274 43503 206277
rect 48773 206274 48839 206277
rect 43437 206272 48839 206274
rect 43437 206216 43442 206272
rect 43498 206216 48778 206272
rect 48834 206216 48839 206272
rect 43437 206214 48839 206216
rect 43437 206211 43503 206214
rect 48773 206211 48839 206214
rect 44357 206002 44423 206005
rect 41492 206000 44423 206002
rect 41492 205944 44362 206000
rect 44418 205944 44423 206000
rect 41492 205942 44423 205944
rect 44357 205939 44423 205942
rect 579521 205866 579587 205869
rect 575798 205864 579587 205866
rect 575798 205808 579526 205864
rect 579582 205808 579587 205864
rect 575798 205806 579587 205808
rect 575798 205700 575858 205806
rect 579521 205803 579587 205806
rect 43621 205594 43687 205597
rect 41492 205592 43687 205594
rect 41492 205536 43626 205592
rect 43682 205536 43687 205592
rect 41492 205534 43687 205536
rect 43621 205531 43687 205534
rect 675753 205594 675819 205597
rect 676622 205594 676628 205596
rect 675753 205592 676628 205594
rect 675753 205536 675758 205592
rect 675814 205536 676628 205592
rect 675753 205534 676628 205536
rect 675753 205531 675819 205534
rect 676622 205532 676628 205534
rect 676692 205532 676698 205596
rect 43989 205186 44055 205189
rect 41492 205184 44055 205186
rect 41492 205128 43994 205184
rect 44050 205128 44055 205184
rect 41492 205126 44055 205128
rect 43989 205123 44055 205126
rect 674741 205050 674807 205053
rect 675477 205050 675543 205053
rect 674741 205048 675543 205050
rect 674741 204992 674746 205048
rect 674802 204992 675482 205048
rect 675538 204992 675543 205048
rect 674741 204990 675543 204992
rect 674741 204987 674807 204990
rect 675477 204987 675543 204990
rect 44817 204778 44883 204781
rect 41492 204776 44883 204778
rect 41492 204720 44822 204776
rect 44878 204720 44883 204776
rect 41492 204718 44883 204720
rect 44817 204715 44883 204718
rect 589641 204778 589707 204781
rect 589641 204776 592572 204778
rect 589641 204720 589646 204776
rect 589702 204720 592572 204776
rect 589641 204718 592572 204720
rect 589641 204715 589707 204718
rect 674925 204506 674991 204509
rect 675477 204506 675543 204509
rect 674925 204504 675543 204506
rect 674925 204448 674930 204504
rect 674986 204448 675482 204504
rect 675538 204448 675543 204504
rect 674925 204446 675543 204448
rect 674925 204443 674991 204446
rect 675477 204443 675543 204446
rect 35574 204101 35634 204340
rect 674833 204234 674899 204237
rect 675293 204234 675359 204237
rect 674833 204232 675359 204234
rect 674833 204176 674838 204232
rect 674894 204176 675298 204232
rect 675354 204176 675359 204232
rect 674833 204174 675359 204176
rect 674833 204171 674899 204174
rect 675293 204171 675359 204174
rect 35574 204096 35683 204101
rect 35574 204040 35622 204096
rect 35678 204040 35683 204096
rect 35574 204038 35683 204040
rect 35617 204035 35683 204038
rect 666356 203970 666938 204030
rect 666878 203962 666938 203970
rect 35758 203693 35818 203932
rect 666878 203902 667122 203962
rect 35758 203688 35867 203693
rect 35758 203632 35806 203688
rect 35862 203632 35867 203688
rect 35758 203630 35867 203632
rect 35801 203627 35867 203630
rect 46381 203554 46447 203557
rect 41492 203552 46447 203554
rect 41492 203496 46386 203552
rect 46442 203496 46447 203552
rect 667062 203554 667122 203902
rect 673913 203554 673979 203557
rect 667062 203552 673979 203554
rect 41492 203494 46447 203496
rect 46381 203491 46447 203494
rect 575982 203282 576042 203524
rect 667062 203496 673918 203552
rect 673974 203496 673979 203552
rect 667062 203494 673979 203496
rect 673913 203491 673979 203494
rect 578325 203282 578391 203285
rect 575982 203280 578391 203282
rect 575982 203224 578330 203280
rect 578386 203224 578391 203280
rect 575982 203222 578391 203224
rect 578325 203219 578391 203222
rect 589457 203146 589523 203149
rect 589457 203144 592572 203146
rect 589457 203088 589462 203144
rect 589518 203088 592572 203144
rect 589457 203086 592572 203088
rect 589457 203083 589523 203086
rect 669221 202466 669287 202469
rect 666694 202464 669287 202466
rect 666694 202408 669226 202464
rect 669282 202408 669287 202464
rect 666694 202406 669287 202408
rect 666694 202398 666754 202406
rect 669221 202403 669287 202406
rect 666356 202338 666754 202398
rect 35617 202194 35683 202197
rect 43437 202194 43503 202197
rect 35617 202192 43503 202194
rect 35617 202136 35622 202192
rect 35678 202136 43442 202192
rect 43498 202136 43503 202192
rect 35617 202134 43503 202136
rect 35617 202131 35683 202134
rect 43437 202131 43503 202134
rect 673361 201922 673427 201925
rect 675477 201922 675543 201925
rect 673361 201920 675543 201922
rect 673361 201864 673366 201920
rect 673422 201864 675482 201920
rect 675538 201864 675543 201920
rect 673361 201862 675543 201864
rect 673361 201859 673427 201862
rect 675477 201859 675543 201862
rect 673269 201652 673335 201653
rect 673269 201650 673316 201652
rect 673224 201648 673316 201650
rect 673224 201592 673274 201648
rect 673224 201590 673316 201592
rect 673269 201588 673316 201590
rect 673380 201588 673386 201652
rect 673269 201587 673335 201588
rect 589457 201514 589523 201517
rect 589457 201512 592572 201514
rect 589457 201456 589462 201512
rect 589518 201456 592572 201512
rect 589457 201454 592572 201456
rect 589457 201451 589523 201454
rect 575982 200834 576042 201348
rect 578785 200834 578851 200837
rect 575982 200832 578851 200834
rect 575982 200776 578790 200832
rect 578846 200776 578851 200832
rect 575982 200774 578851 200776
rect 578785 200771 578851 200774
rect 672165 200834 672231 200837
rect 675293 200834 675359 200837
rect 672165 200832 675359 200834
rect 672165 200776 672170 200832
rect 672226 200776 675298 200832
rect 675354 200776 675359 200832
rect 672165 200774 675359 200776
rect 672165 200771 672231 200774
rect 675293 200771 675359 200774
rect 675753 200698 675819 200701
rect 676438 200698 676444 200700
rect 675753 200696 676444 200698
rect 675753 200640 675758 200696
rect 675814 200640 676444 200696
rect 675753 200638 676444 200640
rect 675753 200635 675819 200638
rect 676438 200636 676444 200638
rect 676508 200636 676514 200700
rect 589457 199882 589523 199885
rect 589457 199880 592572 199882
rect 589457 199824 589462 199880
rect 589518 199824 592572 199880
rect 589457 199822 592572 199824
rect 589457 199819 589523 199822
rect 669129 199338 669195 199341
rect 666878 199336 669195 199338
rect 666878 199280 669134 199336
rect 669190 199280 669195 199336
rect 666878 199278 669195 199280
rect 575982 198930 576042 199172
rect 666878 199134 666938 199278
rect 669129 199275 669195 199278
rect 666356 199074 666938 199134
rect 579521 198930 579587 198933
rect 575982 198928 579587 198930
rect 575982 198872 579526 198928
rect 579582 198872 579587 198928
rect 575982 198870 579587 198872
rect 579521 198867 579587 198870
rect 669221 198794 669287 198797
rect 672533 198794 672599 198797
rect 669221 198792 672599 198794
rect 669221 198736 669226 198792
rect 669282 198736 672538 198792
rect 672594 198736 672599 198792
rect 669221 198734 672599 198736
rect 669221 198731 669287 198734
rect 672533 198731 672599 198734
rect 590377 198250 590443 198253
rect 675569 198252 675635 198253
rect 675518 198250 675524 198252
rect 590377 198248 592572 198250
rect 590377 198192 590382 198248
rect 590438 198192 592572 198248
rect 590377 198190 592572 198192
rect 675478 198190 675524 198250
rect 675588 198248 675635 198252
rect 675630 198192 675635 198248
rect 590377 198187 590443 198190
rect 675518 198188 675524 198190
rect 675588 198188 675635 198192
rect 675569 198187 675635 198188
rect 666502 197916 666508 197980
rect 666572 197978 666578 197980
rect 675109 197978 675175 197981
rect 666572 197976 675175 197978
rect 666572 197920 675114 197976
rect 675170 197920 675175 197976
rect 666572 197918 675175 197920
rect 666572 197916 666578 197918
rect 675109 197915 675175 197918
rect 37917 197842 37983 197845
rect 41822 197842 41828 197844
rect 37917 197840 41828 197842
rect 37917 197784 37922 197840
rect 37978 197784 41828 197840
rect 37917 197782 41828 197784
rect 37917 197779 37983 197782
rect 41822 197780 41828 197782
rect 41892 197780 41898 197844
rect 673545 197706 673611 197709
rect 666878 197704 673611 197706
rect 666878 197648 673550 197704
rect 673606 197648 673611 197704
rect 666878 197646 673611 197648
rect 666878 197502 666938 197646
rect 673545 197643 673611 197646
rect 666356 197442 666938 197502
rect 40534 197100 40540 197164
rect 40604 197162 40610 197164
rect 41781 197162 41847 197165
rect 40604 197160 41847 197162
rect 40604 197104 41786 197160
rect 41842 197104 41847 197160
rect 40604 197102 41847 197104
rect 40604 197100 40610 197102
rect 41781 197099 41847 197102
rect 669405 197162 669471 197165
rect 675477 197162 675543 197165
rect 669405 197160 675543 197162
rect 669405 197104 669410 197160
rect 669466 197104 675482 197160
rect 675538 197104 675543 197160
rect 669405 197102 675543 197104
rect 669405 197099 669471 197102
rect 675477 197099 675543 197102
rect 675753 197162 675819 197165
rect 676254 197162 676260 197164
rect 675753 197160 676260 197162
rect 675753 197104 675758 197160
rect 675814 197104 676260 197160
rect 675753 197102 676260 197104
rect 675753 197099 675819 197102
rect 676254 197100 676260 197102
rect 676324 197100 676330 197164
rect 49509 196482 49575 196485
rect 575982 196482 576042 196996
rect 589457 196618 589523 196621
rect 589457 196616 592572 196618
rect 589457 196560 589462 196616
rect 589518 196560 592572 196616
rect 589457 196558 592572 196560
rect 589457 196555 589523 196558
rect 578509 196482 578575 196485
rect 49509 196480 52164 196482
rect 49509 196424 49514 196480
rect 49570 196424 52164 196480
rect 49509 196422 52164 196424
rect 575982 196480 578575 196482
rect 575982 196424 578514 196480
rect 578570 196424 578575 196480
rect 575982 196422 578575 196424
rect 49509 196419 49575 196422
rect 578509 196419 578575 196422
rect 41873 195804 41939 195805
rect 41822 195802 41828 195804
rect 41782 195742 41828 195802
rect 41892 195800 41939 195804
rect 41934 195744 41939 195800
rect 41822 195740 41828 195742
rect 41892 195740 41939 195744
rect 41873 195739 41939 195740
rect 41454 195196 41460 195260
rect 41524 195258 41530 195260
rect 41781 195258 41847 195261
rect 41524 195256 41847 195258
rect 41524 195200 41786 195256
rect 41842 195200 41847 195256
rect 41524 195198 41847 195200
rect 41524 195196 41530 195198
rect 41781 195195 41847 195198
rect 40902 194924 40908 194988
rect 40972 194986 40978 194988
rect 42241 194986 42307 194989
rect 579521 194986 579587 194989
rect 40972 194984 42307 194986
rect 40972 194928 42246 194984
rect 42302 194928 42307 194984
rect 40972 194926 42307 194928
rect 40972 194924 40978 194926
rect 42241 194923 42307 194926
rect 575798 194984 579587 194986
rect 575798 194928 579526 194984
rect 579582 194928 579587 194984
rect 575798 194926 579587 194928
rect 575798 194820 575858 194926
rect 579521 194923 579587 194926
rect 589273 194986 589339 194989
rect 589273 194984 592572 194986
rect 589273 194928 589278 194984
rect 589334 194928 592572 194984
rect 589273 194926 592572 194928
rect 589273 194923 589339 194926
rect 40718 194516 40724 194580
rect 40788 194578 40794 194580
rect 41638 194578 41644 194580
rect 40788 194518 41644 194578
rect 40788 194516 40794 194518
rect 41638 194516 41644 194518
rect 41708 194516 41714 194580
rect 48129 194442 48195 194445
rect 48129 194440 52164 194442
rect 48129 194384 48134 194440
rect 48190 194384 52164 194440
rect 48129 194382 52164 194384
rect 48129 194379 48195 194382
rect 669129 194306 669195 194309
rect 666694 194304 669195 194306
rect 666694 194248 669134 194304
rect 669190 194248 669195 194304
rect 666694 194246 669195 194248
rect 666694 194238 666754 194246
rect 669129 194243 669195 194246
rect 666356 194178 666754 194238
rect 589457 193354 589523 193357
rect 589457 193352 592572 193354
rect 589457 193296 589462 193352
rect 589518 193296 592572 193352
rect 589457 193294 592572 193296
rect 589457 193291 589523 193294
rect 42241 193220 42307 193221
rect 42190 193156 42196 193220
rect 42260 193218 42307 193220
rect 675661 193218 675727 193221
rect 675886 193218 675892 193220
rect 42260 193216 42352 193218
rect 42302 193160 42352 193216
rect 42260 193158 42352 193160
rect 675661 193216 675892 193218
rect 675661 193160 675666 193216
rect 675722 193160 675892 193216
rect 675661 193158 675892 193160
rect 42260 193156 42307 193158
rect 42241 193155 42307 193156
rect 675661 193155 675727 193158
rect 675886 193156 675892 193158
rect 675956 193156 675962 193220
rect 42333 192946 42399 192949
rect 43805 192946 43871 192949
rect 42333 192944 43871 192946
rect 42333 192888 42338 192944
rect 42394 192888 43810 192944
rect 43866 192888 43871 192944
rect 42333 192886 43871 192888
rect 42333 192883 42399 192886
rect 43805 192883 43871 192886
rect 667933 192674 667999 192677
rect 666694 192672 667999 192674
rect 48773 192402 48839 192405
rect 48773 192400 52164 192402
rect 48773 192344 48778 192400
rect 48834 192344 52164 192400
rect 48773 192342 52164 192344
rect 48773 192339 48839 192342
rect 575982 192266 576042 192644
rect 666694 192616 667938 192672
rect 667994 192616 667999 192672
rect 666694 192614 667999 192616
rect 666694 192606 666754 192614
rect 667933 192611 667999 192614
rect 666356 192546 666754 192606
rect 579521 192266 579587 192269
rect 575982 192264 579587 192266
rect 575982 192208 579526 192264
rect 579582 192208 579587 192264
rect 575982 192206 579587 192208
rect 579521 192203 579587 192206
rect 42333 191722 42399 191725
rect 43989 191722 44055 191725
rect 42333 191720 44055 191722
rect 42333 191664 42338 191720
rect 42394 191664 43994 191720
rect 44050 191664 44055 191720
rect 42333 191662 44055 191664
rect 42333 191659 42399 191662
rect 43989 191659 44055 191662
rect 589457 191722 589523 191725
rect 589457 191720 592572 191722
rect 589457 191664 589462 191720
rect 589518 191664 592572 191720
rect 589457 191662 592572 191664
rect 589457 191659 589523 191662
rect 675753 191586 675819 191589
rect 676070 191586 676076 191588
rect 675753 191584 676076 191586
rect 675753 191528 675758 191584
rect 675814 191528 676076 191584
rect 675753 191526 676076 191528
rect 675753 191523 675819 191526
rect 676070 191524 676076 191526
rect 676140 191524 676146 191588
rect 42425 191178 42491 191181
rect 42977 191178 43043 191181
rect 42425 191176 43043 191178
rect 42425 191120 42430 191176
rect 42486 191120 42982 191176
rect 43038 191120 43043 191176
rect 42425 191118 43043 191120
rect 42425 191115 42491 191118
rect 42977 191115 43043 191118
rect 579521 190770 579587 190773
rect 575798 190768 579587 190770
rect 575798 190712 579526 190768
rect 579582 190712 579587 190768
rect 575798 190710 579587 190712
rect 42425 190498 42491 190501
rect 43621 190498 43687 190501
rect 42425 190496 43687 190498
rect 42425 190440 42430 190496
rect 42486 190440 43626 190496
rect 43682 190440 43687 190496
rect 42425 190438 43687 190440
rect 42425 190435 42491 190438
rect 43621 190435 43687 190438
rect 47945 190498 48011 190501
rect 47945 190496 52164 190498
rect 47945 190440 47950 190496
rect 48006 190440 52164 190496
rect 575798 190468 575858 190710
rect 579521 190707 579587 190710
rect 47945 190438 52164 190440
rect 47945 190435 48011 190438
rect 670601 190362 670667 190365
rect 675293 190362 675359 190365
rect 670601 190360 675359 190362
rect 670601 190304 670606 190360
rect 670662 190304 675298 190360
rect 675354 190304 675359 190360
rect 670601 190302 675359 190304
rect 670601 190299 670667 190302
rect 675293 190299 675359 190302
rect 590561 190090 590627 190093
rect 590561 190088 592572 190090
rect 590561 190032 590566 190088
rect 590622 190032 592572 190088
rect 590561 190030 592572 190032
rect 590561 190027 590627 190030
rect 42425 189954 42491 189957
rect 44541 189954 44607 189957
rect 42425 189952 44607 189954
rect 42425 189896 42430 189952
rect 42486 189896 44546 189952
rect 44602 189896 44607 189952
rect 42425 189894 44607 189896
rect 42425 189891 42491 189894
rect 44541 189891 44607 189894
rect 667933 189410 667999 189413
rect 666694 189408 667999 189410
rect 666694 189352 667938 189408
rect 667994 189352 667999 189408
rect 666694 189350 667999 189352
rect 666694 189342 666754 189350
rect 667933 189347 667999 189350
rect 666356 189282 666754 189342
rect 589641 188458 589707 188461
rect 589641 188456 592572 188458
rect 589641 188400 589646 188456
rect 589702 188400 592572 188456
rect 589641 188398 592572 188400
rect 589641 188395 589707 188398
rect 575982 188050 576042 188292
rect 579521 188050 579587 188053
rect 575982 188048 579587 188050
rect 575982 187992 579526 188048
rect 579582 187992 579587 188048
rect 575982 187990 579587 187992
rect 579521 187987 579587 187990
rect 666356 187650 666754 187710
rect 42425 187642 42491 187645
rect 44357 187642 44423 187645
rect 42425 187640 44423 187642
rect 42425 187584 42430 187640
rect 42486 187584 44362 187640
rect 44418 187584 44423 187640
rect 42425 187582 44423 187584
rect 666694 187642 666754 187650
rect 669129 187642 669195 187645
rect 666694 187640 669195 187642
rect 666694 187584 669134 187640
rect 669190 187584 669195 187640
rect 666694 187582 669195 187584
rect 42425 187579 42491 187582
rect 44357 187579 44423 187582
rect 669129 187579 669195 187582
rect 41781 187236 41847 187237
rect 41781 187232 41828 187236
rect 41892 187234 41898 187236
rect 41781 187176 41786 187232
rect 41781 187172 41828 187176
rect 41892 187174 41938 187234
rect 41892 187172 41898 187174
rect 41781 187171 41847 187172
rect 667565 186962 667631 186965
rect 683113 186962 683179 186965
rect 667565 186960 683179 186962
rect 667565 186904 667570 186960
rect 667626 186904 683118 186960
rect 683174 186904 683179 186960
rect 667565 186902 683179 186904
rect 667565 186899 667631 186902
rect 683113 186899 683179 186902
rect 589457 186826 589523 186829
rect 589457 186824 592572 186826
rect 589457 186768 589462 186824
rect 589518 186768 592572 186824
rect 589457 186766 592572 186768
rect 589457 186763 589523 186766
rect 42333 186284 42399 186285
rect 42333 186282 42380 186284
rect 42288 186280 42380 186282
rect 42288 186224 42338 186280
rect 42288 186222 42380 186224
rect 42333 186220 42380 186222
rect 42444 186220 42450 186284
rect 579521 186282 579587 186285
rect 575798 186280 579587 186282
rect 575798 186224 579526 186280
rect 579582 186224 579587 186280
rect 575798 186222 579587 186224
rect 42333 186219 42399 186220
rect 575798 186116 575858 186222
rect 579521 186219 579587 186222
rect 42149 186012 42215 186013
rect 42149 186010 42196 186012
rect 42104 186008 42196 186010
rect 42104 185952 42154 186008
rect 42104 185950 42196 185952
rect 42149 185948 42196 185950
rect 42260 185948 42266 186012
rect 42149 185947 42215 185948
rect 589457 185194 589523 185197
rect 589457 185192 592572 185194
rect 589457 185136 589462 185192
rect 589518 185136 592572 185192
rect 589457 185134 592572 185136
rect 589457 185131 589523 185134
rect 42425 184922 42491 184925
rect 44173 184922 44239 184925
rect 42425 184920 44239 184922
rect 42425 184864 42430 184920
rect 42486 184864 44178 184920
rect 44234 184864 44239 184920
rect 42425 184862 44239 184864
rect 42425 184859 42491 184862
rect 44173 184859 44239 184862
rect 669221 184514 669287 184517
rect 666694 184512 669287 184514
rect 666694 184456 669226 184512
rect 669282 184456 669287 184512
rect 666694 184454 669287 184456
rect 666694 184446 666754 184454
rect 669221 184451 669287 184454
rect 666356 184386 666754 184446
rect 579521 184378 579587 184381
rect 575798 184376 579587 184378
rect 575798 184320 579526 184376
rect 579582 184320 579587 184376
rect 575798 184318 579587 184320
rect 575798 183940 575858 184318
rect 579521 184315 579587 184318
rect 589457 183562 589523 183565
rect 672073 183562 672139 183565
rect 672942 183562 672948 183564
rect 589457 183560 592572 183562
rect 589457 183504 589462 183560
rect 589518 183504 592572 183560
rect 589457 183502 592572 183504
rect 672073 183560 672948 183562
rect 672073 183504 672078 183560
rect 672134 183504 672948 183560
rect 672073 183502 672948 183504
rect 589457 183499 589523 183502
rect 672073 183499 672139 183502
rect 672942 183500 672948 183502
rect 673012 183500 673018 183564
rect 42425 183154 42491 183157
rect 43253 183154 43319 183157
rect 42425 183152 43319 183154
rect 42425 183096 42430 183152
rect 42486 183096 43258 183152
rect 43314 183096 43319 183152
rect 42425 183094 43319 183096
rect 42425 183091 42491 183094
rect 43253 183091 43319 183094
rect 668117 182882 668183 182885
rect 666694 182880 668183 182882
rect 666694 182824 668122 182880
rect 668178 182824 668183 182880
rect 666694 182822 668183 182824
rect 666694 182814 666754 182822
rect 668117 182819 668183 182822
rect 666356 182754 666754 182814
rect 672257 182066 672323 182069
rect 673126 182066 673132 182068
rect 672257 182064 673132 182066
rect 672257 182008 672262 182064
rect 672318 182008 673132 182064
rect 672257 182006 673132 182008
rect 672257 182003 672323 182006
rect 673126 182004 673132 182006
rect 673196 182004 673202 182068
rect 579521 181930 579587 181933
rect 575798 181928 579587 181930
rect 575798 181872 579526 181928
rect 579582 181872 579587 181928
rect 575798 181870 579587 181872
rect 575798 181764 575858 181870
rect 579521 181867 579587 181870
rect 590561 181930 590627 181933
rect 590561 181928 592572 181930
rect 590561 181872 590566 181928
rect 590622 181872 592572 181928
rect 590561 181870 592572 181872
rect 590561 181867 590627 181870
rect 667381 181386 667447 181389
rect 676489 181386 676555 181389
rect 667381 181384 676555 181386
rect 667381 181328 667386 181384
rect 667442 181328 676494 181384
rect 676550 181328 676555 181384
rect 667381 181326 676555 181328
rect 667381 181323 667447 181326
rect 676489 181323 676555 181326
rect 589641 180298 589707 180301
rect 589641 180296 592572 180298
rect 589641 180240 589646 180296
rect 589702 180240 592572 180296
rect 589641 180238 592572 180240
rect 589641 180235 589707 180238
rect 578785 180162 578851 180165
rect 575798 180160 578851 180162
rect 575798 180104 578790 180160
rect 578846 180104 578851 180160
rect 575798 180102 578851 180104
rect 575798 179588 575858 180102
rect 578785 180099 578851 180102
rect 666356 179490 666938 179550
rect 666878 179482 666938 179490
rect 674097 179482 674163 179485
rect 666878 179480 674163 179482
rect 666878 179424 674102 179480
rect 674158 179424 674163 179480
rect 666878 179422 674163 179424
rect 674097 179419 674163 179422
rect 667013 178802 667079 178805
rect 683113 178802 683179 178805
rect 667013 178800 675770 178802
rect 667013 178744 667018 178800
rect 667074 178744 675770 178800
rect 667013 178742 675770 178744
rect 667013 178739 667079 178742
rect 589457 178666 589523 178669
rect 589457 178664 592572 178666
rect 589457 178608 589462 178664
rect 589518 178608 592572 178664
rect 589457 178606 592572 178608
rect 589457 178603 589523 178606
rect 672993 177986 673059 177989
rect 666694 177984 673059 177986
rect 666694 177928 672998 177984
rect 673054 177928 673059 177984
rect 666694 177926 673059 177928
rect 675710 177986 675770 178742
rect 683070 178800 683179 178802
rect 683070 178744 683118 178800
rect 683174 178744 683179 178800
rect 683070 178739 683179 178744
rect 683070 178500 683130 178739
rect 676029 178122 676095 178125
rect 676029 178120 676292 178122
rect 676029 178064 676034 178120
rect 676090 178064 676292 178120
rect 676029 178062 676292 178064
rect 676029 178059 676095 178062
rect 675710 177926 675954 177986
rect 666694 177918 666754 177926
rect 672993 177923 673059 177926
rect 666356 177858 666754 177918
rect 579521 177714 579587 177717
rect 575798 177712 579587 177714
rect 575798 177656 579526 177712
rect 579582 177656 579587 177712
rect 575798 177654 579587 177656
rect 675894 177714 675954 177926
rect 675894 177654 676292 177714
rect 575798 177412 575858 177654
rect 579521 177651 579587 177654
rect 674373 177306 674439 177309
rect 674373 177304 676292 177306
rect 674373 177248 674378 177304
rect 674434 177248 676292 177304
rect 674373 177246 676292 177248
rect 674373 177243 674439 177246
rect 589641 177034 589707 177037
rect 589641 177032 592572 177034
rect 589641 176976 589646 177032
rect 589702 176976 592572 177032
rect 589641 176974 592572 176976
rect 589641 176971 589707 176974
rect 674281 176898 674347 176901
rect 674281 176896 676292 176898
rect 674281 176840 674286 176896
rect 674342 176840 676292 176896
rect 674281 176838 676292 176840
rect 674281 176835 674347 176838
rect 666645 176490 666711 176493
rect 666645 176488 676292 176490
rect 666645 176432 666650 176488
rect 666706 176432 676292 176488
rect 666645 176430 676292 176432
rect 666645 176427 666711 176430
rect 673913 176082 673979 176085
rect 673913 176080 676292 176082
rect 673913 176024 673918 176080
rect 673974 176024 676292 176080
rect 673913 176022 676292 176024
rect 673913 176019 673979 176022
rect 674557 175674 674623 175677
rect 674557 175672 676292 175674
rect 674557 175616 674562 175672
rect 674618 175616 676292 175672
rect 674557 175614 676292 175616
rect 674557 175611 674623 175614
rect 589457 175402 589523 175405
rect 589457 175400 592572 175402
rect 589457 175344 589462 175400
rect 589518 175344 592572 175400
rect 589457 175342 592572 175344
rect 589457 175339 589523 175342
rect 672533 175266 672599 175269
rect 672533 175264 676292 175266
rect 575982 175130 576042 175236
rect 672533 175208 672538 175264
rect 672594 175208 676292 175264
rect 672533 175206 676292 175208
rect 672533 175203 672599 175206
rect 578785 175130 578851 175133
rect 575982 175128 578851 175130
rect 575982 175072 578790 175128
rect 578846 175072 578851 175128
rect 575982 175070 578851 175072
rect 578785 175067 578851 175070
rect 671889 174858 671955 174861
rect 671889 174856 676292 174858
rect 671889 174800 671894 174856
rect 671950 174800 676292 174856
rect 671889 174798 676292 174800
rect 671889 174795 671955 174798
rect 667933 174722 667999 174725
rect 666694 174720 667999 174722
rect 666694 174664 667938 174720
rect 667994 174664 667999 174720
rect 666694 174662 667999 174664
rect 666694 174654 666754 174662
rect 667933 174659 667999 174662
rect 666356 174594 666754 174654
rect 673361 174450 673427 174453
rect 673361 174448 676292 174450
rect 673361 174392 673366 174448
rect 673422 174392 676292 174448
rect 673361 174390 676292 174392
rect 673361 174387 673427 174390
rect 675886 173980 675892 174044
rect 675956 174042 675962 174044
rect 675956 173982 676292 174042
rect 675956 173980 675962 173982
rect 589457 173770 589523 173773
rect 589457 173768 592572 173770
rect 589457 173712 589462 173768
rect 589518 173712 592572 173768
rect 589457 173710 592572 173712
rect 589457 173707 589523 173710
rect 675702 173572 675708 173636
rect 675772 173634 675778 173636
rect 675772 173574 676292 173634
rect 675772 173572 675778 173574
rect 578417 173498 578483 173501
rect 575798 173496 578483 173498
rect 575798 173440 578422 173496
rect 578478 173440 578483 173496
rect 575798 173438 578483 173440
rect 575798 173060 575858 173438
rect 578417 173435 578483 173438
rect 678237 173226 678303 173229
rect 678237 173224 678316 173226
rect 678237 173168 678242 173224
rect 678298 173168 678316 173224
rect 678237 173166 678316 173168
rect 678237 173163 678303 173166
rect 672901 173090 672967 173093
rect 666694 173088 672967 173090
rect 666694 173032 672906 173088
rect 672962 173032 672967 173088
rect 666694 173030 672967 173032
rect 666694 173022 666754 173030
rect 672901 173027 672967 173030
rect 666356 172962 666754 173022
rect 674833 172818 674899 172821
rect 674833 172816 676292 172818
rect 674833 172760 674838 172816
rect 674894 172760 676292 172816
rect 674833 172758 676292 172760
rect 674833 172755 674899 172758
rect 675886 172348 675892 172412
rect 675956 172410 675962 172412
rect 675956 172350 676292 172410
rect 675956 172348 675962 172350
rect 589457 172138 589523 172141
rect 589457 172136 592572 172138
rect 589457 172080 589462 172136
rect 589518 172080 592572 172136
rect 589457 172078 592572 172080
rect 589457 172075 589523 172078
rect 675886 171940 675892 172004
rect 675956 172002 675962 172004
rect 675956 171942 676292 172002
rect 675956 171940 675962 171942
rect 680997 171594 681063 171597
rect 680997 171592 681076 171594
rect 680997 171536 681002 171592
rect 681058 171536 681076 171592
rect 680997 171534 681076 171536
rect 680997 171531 681063 171534
rect 679617 171186 679683 171189
rect 679604 171184 679683 171186
rect 679604 171128 679622 171184
rect 679678 171128 679683 171184
rect 679604 171126 679683 171128
rect 679617 171123 679683 171126
rect 578233 171050 578299 171053
rect 575798 171048 578299 171050
rect 575798 170992 578238 171048
rect 578294 170992 578299 171048
rect 575798 170990 578299 170992
rect 575798 170884 575858 170990
rect 578233 170987 578299 170990
rect 676581 170778 676647 170781
rect 676581 170776 676660 170778
rect 676581 170720 676586 170776
rect 676642 170720 676660 170776
rect 676581 170718 676660 170720
rect 676581 170715 676647 170718
rect 589457 170506 589523 170509
rect 589457 170504 592572 170506
rect 589457 170448 589462 170504
rect 589518 170448 592572 170504
rect 589457 170446 592572 170448
rect 589457 170443 589523 170446
rect 670601 170370 670667 170373
rect 670601 170368 676292 170370
rect 670601 170312 670606 170368
rect 670662 170312 676292 170368
rect 670601 170310 676292 170312
rect 670601 170307 670667 170310
rect 673177 169962 673243 169965
rect 673177 169960 676292 169962
rect 673177 169904 673182 169960
rect 673238 169904 676292 169960
rect 673177 169902 676292 169904
rect 673177 169899 673243 169902
rect 666356 169698 666754 169758
rect 666694 169690 666754 169698
rect 668025 169690 668091 169693
rect 666694 169688 668091 169690
rect 666694 169632 668030 169688
rect 668086 169632 668091 169688
rect 666694 169630 668091 169632
rect 668025 169627 668091 169630
rect 674097 169554 674163 169557
rect 674097 169552 676292 169554
rect 674097 169496 674102 169552
rect 674158 169496 676292 169552
rect 674097 169494 676292 169496
rect 674097 169491 674163 169494
rect 578693 169282 578759 169285
rect 575798 169280 578759 169282
rect 575798 169224 578698 169280
rect 578754 169224 578759 169280
rect 575798 169222 578759 169224
rect 575798 168708 575858 169222
rect 578693 169219 578759 169222
rect 672993 169146 673059 169149
rect 672993 169144 676292 169146
rect 672993 169088 672998 169144
rect 673054 169088 676292 169144
rect 672993 169086 676292 169088
rect 672993 169083 673059 169086
rect 589457 168874 589523 168877
rect 589457 168872 592572 168874
rect 589457 168816 589462 168872
rect 589518 168816 592572 168872
rect 589457 168814 592572 168816
rect 589457 168811 589523 168814
rect 674465 168738 674531 168741
rect 674465 168736 676292 168738
rect 674465 168680 674470 168736
rect 674526 168680 676292 168736
rect 674465 168678 676292 168680
rect 674465 168675 674531 168678
rect 673729 168466 673795 168469
rect 667982 168464 673795 168466
rect 667982 168408 673734 168464
rect 673790 168408 673795 168464
rect 667982 168406 673795 168408
rect 667982 168194 668042 168406
rect 673729 168403 673795 168406
rect 673870 168270 676292 168330
rect 666878 168134 668042 168194
rect 669773 168194 669839 168197
rect 673870 168194 673930 168270
rect 669773 168192 673930 168194
rect 669773 168136 669778 168192
rect 669834 168136 673930 168192
rect 669773 168134 673930 168136
rect 666878 168126 666938 168134
rect 669773 168131 669839 168134
rect 666356 168066 666938 168126
rect 676029 167922 676095 167925
rect 676029 167920 676292 167922
rect 676029 167864 676034 167920
rect 676090 167864 676292 167920
rect 676029 167862 676292 167864
rect 676029 167859 676095 167862
rect 675518 167452 675524 167516
rect 675588 167514 675594 167516
rect 675588 167454 676292 167514
rect 675588 167452 675594 167454
rect 589457 167242 589523 167245
rect 589457 167240 592572 167242
rect 589457 167184 589462 167240
rect 589518 167184 592572 167240
rect 589457 167182 592572 167184
rect 589457 167179 589523 167182
rect 676170 167046 676292 167106
rect 579521 166970 579587 166973
rect 575798 166968 579587 166970
rect 575798 166912 579526 166968
rect 579582 166912 579587 166968
rect 575798 166910 579587 166912
rect 575798 166532 575858 166910
rect 579521 166907 579587 166910
rect 671889 166970 671955 166973
rect 676170 166970 676230 167046
rect 671889 166968 676230 166970
rect 671889 166912 671894 166968
rect 671950 166912 676230 166968
rect 671889 166910 676230 166912
rect 671889 166907 671955 166910
rect 676581 166428 676647 166429
rect 676581 166424 676628 166428
rect 676692 166426 676698 166428
rect 676581 166368 676586 166424
rect 676581 166364 676628 166368
rect 676692 166366 676738 166426
rect 676692 166364 676698 166366
rect 676581 166363 676647 166364
rect 589457 165610 589523 165613
rect 670325 165610 670391 165613
rect 676029 165610 676095 165613
rect 589457 165608 592572 165610
rect 589457 165552 589462 165608
rect 589518 165552 592572 165608
rect 589457 165550 592572 165552
rect 670325 165608 676095 165610
rect 670325 165552 670330 165608
rect 670386 165552 676034 165608
rect 676090 165552 676095 165608
rect 670325 165550 676095 165552
rect 589457 165547 589523 165550
rect 670325 165547 670391 165550
rect 676029 165547 676095 165550
rect 667933 164930 667999 164933
rect 666694 164928 667999 164930
rect 666694 164872 667938 164928
rect 667994 164872 667999 164928
rect 666694 164870 667999 164872
rect 666694 164862 666754 164870
rect 667933 164867 667999 164870
rect 666356 164802 666754 164862
rect 578877 164522 578943 164525
rect 575798 164520 578943 164522
rect 575798 164464 578882 164520
rect 578938 164464 578943 164520
rect 575798 164462 578943 164464
rect 575798 164356 575858 164462
rect 578877 164459 578943 164462
rect 669129 164250 669195 164253
rect 672257 164250 672323 164253
rect 669129 164248 672323 164250
rect 669129 164192 669134 164248
rect 669190 164192 672262 164248
rect 672318 164192 672323 164248
rect 669129 164190 672323 164192
rect 669129 164187 669195 164190
rect 672257 164187 672323 164190
rect 589457 163978 589523 163981
rect 589457 163976 592572 163978
rect 589457 163920 589462 163976
rect 589518 163920 592572 163976
rect 589457 163918 592572 163920
rect 589457 163915 589523 163918
rect 668301 163298 668367 163301
rect 666694 163296 668367 163298
rect 666694 163240 668306 163296
rect 668362 163240 668367 163296
rect 666694 163238 668367 163240
rect 666694 163230 666754 163238
rect 668301 163235 668367 163238
rect 666356 163170 666754 163230
rect 579521 162754 579587 162757
rect 575798 162752 579587 162754
rect 575798 162696 579526 162752
rect 579582 162696 579587 162752
rect 575798 162694 579587 162696
rect 575798 162180 575858 162694
rect 579521 162691 579587 162694
rect 589457 162346 589523 162349
rect 589457 162344 592572 162346
rect 589457 162288 589462 162344
rect 589518 162288 592572 162344
rect 589457 162286 592572 162288
rect 589457 162283 589523 162286
rect 675334 161876 675340 161940
rect 675404 161938 675410 161940
rect 675937 161938 676003 161941
rect 675404 161936 676003 161938
rect 675404 161880 675942 161936
rect 675998 161880 676003 161936
rect 675404 161878 676003 161880
rect 675404 161876 675410 161878
rect 675937 161875 676003 161878
rect 676121 161394 676187 161397
rect 676078 161392 676187 161394
rect 676078 161336 676126 161392
rect 676182 161336 676187 161392
rect 676078 161331 676187 161336
rect 589457 160714 589523 160717
rect 675753 160714 675819 160717
rect 676078 160714 676138 161331
rect 589457 160712 592572 160714
rect 589457 160656 589462 160712
rect 589518 160656 592572 160712
rect 589457 160654 592572 160656
rect 675753 160712 676138 160714
rect 675753 160656 675758 160712
rect 675814 160656 676138 160712
rect 675753 160654 676138 160656
rect 589457 160651 589523 160654
rect 675753 160651 675819 160654
rect 668945 160034 669011 160037
rect 666694 160032 669011 160034
rect 575982 159898 576042 160004
rect 666694 159976 668950 160032
rect 669006 159976 669011 160032
rect 666694 159974 669011 159976
rect 666694 159966 666754 159974
rect 668945 159971 669011 159974
rect 666356 159906 666754 159966
rect 578233 159898 578299 159901
rect 575982 159896 578299 159898
rect 575982 159840 578238 159896
rect 578294 159840 578299 159896
rect 575982 159838 578299 159840
rect 578233 159835 578299 159838
rect 675753 159354 675819 159357
rect 676438 159354 676444 159356
rect 675753 159352 676444 159354
rect 675753 159296 675758 159352
rect 675814 159296 676444 159352
rect 675753 159294 676444 159296
rect 675753 159291 675819 159294
rect 676438 159292 676444 159294
rect 676508 159292 676514 159356
rect 589825 159082 589891 159085
rect 589825 159080 592572 159082
rect 589825 159024 589830 159080
rect 589886 159024 592572 159080
rect 589825 159022 592572 159024
rect 589825 159019 589891 159022
rect 578417 158402 578483 158405
rect 671705 158402 671771 158405
rect 575798 158400 578483 158402
rect 575798 158344 578422 158400
rect 578478 158344 578483 158400
rect 575798 158342 578483 158344
rect 575798 157828 575858 158342
rect 578417 158339 578483 158342
rect 666694 158400 671771 158402
rect 666694 158344 671710 158400
rect 671766 158344 671771 158400
rect 666694 158342 671771 158344
rect 666694 158334 666754 158342
rect 671705 158339 671771 158342
rect 666356 158274 666754 158334
rect 674833 157586 674899 157589
rect 675477 157586 675543 157589
rect 674833 157584 675543 157586
rect 674833 157528 674838 157584
rect 674894 157528 675482 157584
rect 675538 157528 675543 157584
rect 674833 157526 675543 157528
rect 674833 157523 674899 157526
rect 675477 157523 675543 157526
rect 589457 157450 589523 157453
rect 589457 157448 592572 157450
rect 589457 157392 589462 157448
rect 589518 157392 592572 157448
rect 589457 157390 592572 157392
rect 589457 157387 589523 157390
rect 675385 157044 675451 157045
rect 675334 156980 675340 157044
rect 675404 157042 675451 157044
rect 675404 157040 675496 157042
rect 675446 156984 675496 157040
rect 675404 156982 675496 156984
rect 675404 156980 675451 156982
rect 675385 156979 675451 156980
rect 675753 156362 675819 156365
rect 676622 156362 676628 156364
rect 675753 156360 676628 156362
rect 675753 156304 675758 156360
rect 675814 156304 676628 156360
rect 675753 156302 676628 156304
rect 675753 156299 675819 156302
rect 676622 156300 676628 156302
rect 676692 156300 676698 156364
rect 578877 155954 578943 155957
rect 575798 155952 578943 155954
rect 575798 155896 578882 155952
rect 578938 155896 578943 155952
rect 575798 155894 578943 155896
rect 575798 155652 575858 155894
rect 578877 155891 578943 155894
rect 589457 155818 589523 155821
rect 589457 155816 592572 155818
rect 589457 155760 589462 155816
rect 589518 155760 592572 155816
rect 589457 155758 592572 155760
rect 589457 155755 589523 155758
rect 674097 155410 674163 155413
rect 675109 155410 675175 155413
rect 674097 155408 675175 155410
rect 674097 155352 674102 155408
rect 674158 155352 675114 155408
rect 675170 155352 675175 155408
rect 674097 155350 675175 155352
rect 674097 155347 674163 155350
rect 675109 155347 675175 155350
rect 666356 155010 666938 155070
rect 666878 155002 666938 155010
rect 674230 155002 674236 155004
rect 666878 154942 674236 155002
rect 674230 154940 674236 154942
rect 674300 154940 674306 155004
rect 589457 154186 589523 154189
rect 589457 154184 592572 154186
rect 589457 154128 589462 154184
rect 589518 154128 592572 154184
rect 589457 154126 592572 154128
rect 589457 154123 589523 154126
rect 578325 154050 578391 154053
rect 575798 154048 578391 154050
rect 575798 153992 578330 154048
rect 578386 153992 578391 154048
rect 575798 153990 578391 153992
rect 575798 153476 575858 153990
rect 578325 153987 578391 153990
rect 668761 153506 668827 153509
rect 666694 153504 668827 153506
rect 666694 153448 668766 153504
rect 668822 153448 668827 153504
rect 666694 153446 668827 153448
rect 666694 153438 666754 153446
rect 668761 153443 668827 153446
rect 666356 153378 666754 153438
rect 672993 153098 673059 153101
rect 675109 153098 675175 153101
rect 672993 153096 675175 153098
rect 672993 153040 672998 153096
rect 673054 153040 675114 153096
rect 675170 153040 675175 153096
rect 672993 153038 675175 153040
rect 672993 153035 673059 153038
rect 675109 153035 675175 153038
rect 675753 153098 675819 153101
rect 676254 153098 676260 153100
rect 675753 153096 676260 153098
rect 675753 153040 675758 153096
rect 675814 153040 676260 153096
rect 675753 153038 676260 153040
rect 675753 153035 675819 153038
rect 676254 153036 676260 153038
rect 676324 153036 676330 153100
rect 589457 152554 589523 152557
rect 589457 152552 592572 152554
rect 589457 152496 589462 152552
rect 589518 152496 592572 152552
rect 589457 152494 592572 152496
rect 589457 152491 589523 152494
rect 578233 151738 578299 151741
rect 575798 151736 578299 151738
rect 575798 151680 578238 151736
rect 578294 151680 578299 151736
rect 575798 151678 578299 151680
rect 575798 151300 575858 151678
rect 578233 151675 578299 151678
rect 673177 151738 673243 151741
rect 675109 151738 675175 151741
rect 673177 151736 675175 151738
rect 673177 151680 673182 151736
rect 673238 151680 675114 151736
rect 675170 151680 675175 151736
rect 673177 151678 675175 151680
rect 673177 151675 673243 151678
rect 675109 151675 675175 151678
rect 590009 150922 590075 150925
rect 590009 150920 592572 150922
rect 590009 150864 590014 150920
rect 590070 150864 592572 150920
rect 590009 150862 592572 150864
rect 590009 150859 590075 150862
rect 671521 150242 671587 150245
rect 666694 150240 671587 150242
rect 666694 150184 671526 150240
rect 671582 150184 671587 150240
rect 666694 150182 671587 150184
rect 666694 150174 666754 150182
rect 671521 150179 671587 150182
rect 666356 150114 666754 150174
rect 578325 149698 578391 149701
rect 575798 149696 578391 149698
rect 575798 149640 578330 149696
rect 578386 149640 578391 149696
rect 575798 149638 578391 149640
rect 575798 149124 575858 149638
rect 578325 149635 578391 149638
rect 589457 149290 589523 149293
rect 589457 149288 592572 149290
rect 589457 149232 589462 149288
rect 589518 149232 592572 149288
rect 589457 149230 592572 149232
rect 589457 149227 589523 149230
rect 668761 149154 668827 149157
rect 673310 149154 673316 149156
rect 668761 149152 673316 149154
rect 668761 149096 668766 149152
rect 668822 149096 673316 149152
rect 668761 149094 673316 149096
rect 668761 149091 668827 149094
rect 673310 149092 673316 149094
rect 673380 149092 673386 149156
rect 668485 148610 668551 148613
rect 666694 148608 668551 148610
rect 666694 148552 668490 148608
rect 668546 148552 668551 148608
rect 666694 148550 668551 148552
rect 666694 148542 666754 148550
rect 668485 148547 668551 148550
rect 666356 148482 666754 148542
rect 675661 148474 675727 148477
rect 675886 148474 675892 148476
rect 675661 148472 675892 148474
rect 675661 148416 675666 148472
rect 675722 148416 675892 148472
rect 675661 148414 675892 148416
rect 675661 148411 675727 148414
rect 675886 148412 675892 148414
rect 675956 148412 675962 148476
rect 588537 147658 588603 147661
rect 670601 147658 670667 147661
rect 675109 147658 675175 147661
rect 588537 147656 592572 147658
rect 588537 147600 588542 147656
rect 588598 147600 592572 147656
rect 588537 147598 592572 147600
rect 670601 147656 675175 147658
rect 670601 147600 670606 147656
rect 670662 147600 675114 147656
rect 675170 147600 675175 147656
rect 670601 147598 675175 147600
rect 588537 147595 588603 147598
rect 670601 147595 670667 147598
rect 675109 147595 675175 147598
rect 675661 147660 675727 147661
rect 675661 147656 675708 147660
rect 675772 147658 675778 147660
rect 675661 147600 675666 147656
rect 675661 147596 675708 147600
rect 675772 147598 675818 147658
rect 675772 147596 675778 147598
rect 675661 147595 675727 147596
rect 578693 147250 578759 147253
rect 575798 147248 578759 147250
rect 575798 147192 578698 147248
rect 578754 147192 578759 147248
rect 575798 147190 578759 147192
rect 575798 146948 575858 147190
rect 578693 147187 578759 147190
rect 589457 146026 589523 146029
rect 675753 146026 675819 146029
rect 676070 146026 676076 146028
rect 589457 146024 592572 146026
rect 589457 145968 589462 146024
rect 589518 145968 592572 146024
rect 589457 145966 592572 145968
rect 675753 146024 676076 146026
rect 675753 145968 675758 146024
rect 675814 145968 676076 146024
rect 675753 145966 676076 145968
rect 589457 145963 589523 145966
rect 675753 145963 675819 145966
rect 676070 145964 676076 145966
rect 676140 145964 676146 146028
rect 668577 145346 668643 145349
rect 666694 145344 668643 145346
rect 666694 145288 668582 145344
rect 668638 145288 668643 145344
rect 666694 145286 668643 145288
rect 666694 145278 666754 145286
rect 668577 145283 668643 145286
rect 666356 145218 666754 145278
rect 575982 144666 576042 144772
rect 579245 144666 579311 144669
rect 575982 144664 579311 144666
rect 575982 144608 579250 144664
rect 579306 144608 579311 144664
rect 575982 144606 579311 144608
rect 579245 144603 579311 144606
rect 589457 144394 589523 144397
rect 589457 144392 592572 144394
rect 589457 144336 589462 144392
rect 589518 144336 592572 144392
rect 589457 144334 592572 144336
rect 589457 144331 589523 144334
rect 669262 143714 669268 143716
rect 666694 143654 669268 143714
rect 666694 143646 666754 143654
rect 669262 143652 669268 143654
rect 669332 143652 669338 143716
rect 666356 143586 666754 143646
rect 579521 143034 579587 143037
rect 575798 143032 579587 143034
rect 575798 142976 579526 143032
rect 579582 142976 579587 143032
rect 575798 142974 579587 142976
rect 575798 142596 575858 142974
rect 579521 142971 579587 142974
rect 589825 142762 589891 142765
rect 589825 142760 592572 142762
rect 589825 142704 589830 142760
rect 589886 142704 592572 142760
rect 589825 142702 592572 142704
rect 589825 142699 589891 142702
rect 589457 141130 589523 141133
rect 589457 141128 592572 141130
rect 589457 141072 589462 141128
rect 589518 141072 592572 141128
rect 589457 141070 592572 141072
rect 589457 141067 589523 141070
rect 578601 140586 578667 140589
rect 575798 140584 578667 140586
rect 575798 140528 578606 140584
rect 578662 140528 578667 140584
rect 575798 140526 578667 140528
rect 575798 140420 575858 140526
rect 578601 140523 578667 140526
rect 672073 140450 672139 140453
rect 666694 140448 672139 140450
rect 666694 140392 672078 140448
rect 672134 140392 672139 140448
rect 666694 140390 672139 140392
rect 666694 140382 666754 140390
rect 672073 140387 672139 140390
rect 666356 140322 666754 140382
rect 589457 139498 589523 139501
rect 589457 139496 592572 139498
rect 589457 139440 589462 139496
rect 589518 139440 592572 139496
rect 589457 139438 592572 139440
rect 589457 139435 589523 139438
rect 578601 138818 578667 138821
rect 669129 138818 669195 138821
rect 575798 138816 578667 138818
rect 575798 138760 578606 138816
rect 578662 138760 578667 138816
rect 575798 138758 578667 138760
rect 575798 138244 575858 138758
rect 578601 138755 578667 138758
rect 666694 138816 669195 138818
rect 666694 138760 669134 138816
rect 669190 138760 669195 138816
rect 666694 138758 669195 138760
rect 666694 138750 666754 138758
rect 669129 138755 669195 138758
rect 666356 138690 666754 138750
rect 589457 137866 589523 137869
rect 589457 137864 592572 137866
rect 589457 137808 589462 137864
rect 589518 137808 592572 137864
rect 589457 137806 592572 137808
rect 589457 137803 589523 137806
rect 578877 136642 578943 136645
rect 575798 136640 578943 136642
rect 575798 136584 578882 136640
rect 578938 136584 578943 136640
rect 575798 136582 578943 136584
rect 575798 136068 575858 136582
rect 578877 136579 578943 136582
rect 589457 136234 589523 136237
rect 589457 136232 592572 136234
rect 589457 136176 589462 136232
rect 589518 136176 592572 136232
rect 589457 136174 592572 136176
rect 589457 136171 589523 136174
rect 667749 135962 667815 135965
rect 683113 135962 683179 135965
rect 667749 135960 683179 135962
rect 667749 135904 667754 135960
rect 667810 135904 683118 135960
rect 683174 135904 683179 135960
rect 667749 135902 683179 135904
rect 667749 135899 667815 135902
rect 683113 135899 683179 135902
rect 667933 135554 667999 135557
rect 666694 135552 667999 135554
rect 666694 135496 667938 135552
rect 667994 135496 667999 135552
rect 666694 135494 667999 135496
rect 666694 135486 666754 135494
rect 667933 135491 667999 135494
rect 666356 135426 666754 135486
rect 590285 134602 590351 134605
rect 667197 134602 667263 134605
rect 675845 134602 675911 134605
rect 590285 134600 592572 134602
rect 590285 134544 590290 134600
rect 590346 134544 592572 134600
rect 590285 134542 592572 134544
rect 667197 134600 675911 134602
rect 667197 134544 667202 134600
rect 667258 134544 675850 134600
rect 675906 134544 675911 134600
rect 667197 134542 675911 134544
rect 590285 134539 590351 134542
rect 667197 134539 667263 134542
rect 675845 134539 675911 134542
rect 578693 134466 578759 134469
rect 575798 134464 578759 134466
rect 575798 134408 578698 134464
rect 578754 134408 578759 134464
rect 575798 134406 578759 134408
rect 575798 133892 575858 134406
rect 578693 134403 578759 134406
rect 666356 133794 666754 133854
rect 666694 133786 666754 133794
rect 670734 133786 670740 133788
rect 666694 133726 670740 133786
rect 670734 133724 670740 133726
rect 670804 133724 670810 133788
rect 666829 133106 666895 133109
rect 676262 133106 676322 133348
rect 676489 133106 676555 133109
rect 666829 133104 676322 133106
rect 666829 133048 666834 133104
rect 666890 133048 676322 133104
rect 666829 133046 676322 133048
rect 676446 133104 676555 133106
rect 676446 133048 676494 133104
rect 676550 133048 676555 133104
rect 666829 133043 666895 133046
rect 676446 133043 676555 133048
rect 588721 132970 588787 132973
rect 588721 132968 592572 132970
rect 588721 132912 588726 132968
rect 588782 132912 592572 132968
rect 676446 132940 676506 133043
rect 588721 132910 592572 132912
rect 588721 132907 588787 132910
rect 683113 132698 683179 132701
rect 683070 132696 683179 132698
rect 683070 132640 683118 132696
rect 683174 132640 683179 132696
rect 683070 132635 683179 132640
rect 683070 132532 683130 132635
rect 579061 132290 579127 132293
rect 575798 132288 579127 132290
rect 575798 132232 579066 132288
rect 579122 132232 579127 132288
rect 575798 132230 579127 132232
rect 575798 131716 575858 132230
rect 579061 132227 579127 132230
rect 674281 132154 674347 132157
rect 674281 132152 676292 132154
rect 674281 132096 674286 132152
rect 674342 132096 676292 132152
rect 674281 132094 676292 132096
rect 674281 132091 674347 132094
rect 671337 131746 671403 131749
rect 671337 131744 676292 131746
rect 671337 131688 671342 131744
rect 671398 131688 676292 131744
rect 671337 131686 676292 131688
rect 671337 131683 671403 131686
rect 589457 131338 589523 131341
rect 673913 131338 673979 131341
rect 589457 131336 592572 131338
rect 589457 131280 589462 131336
rect 589518 131280 592572 131336
rect 589457 131278 592572 131280
rect 673913 131336 676292 131338
rect 673913 131280 673918 131336
rect 673974 131280 676292 131336
rect 673913 131278 676292 131280
rect 589457 131275 589523 131278
rect 673913 131275 673979 131278
rect 671521 130930 671587 130933
rect 671521 130928 676292 130930
rect 671521 130872 671526 130928
rect 671582 130872 676292 130928
rect 671521 130870 676292 130872
rect 671521 130867 671587 130870
rect 667974 130658 667980 130660
rect 666694 130598 667980 130658
rect 666694 130590 666754 130598
rect 667974 130596 667980 130598
rect 668044 130596 668050 130660
rect 666356 130530 666754 130590
rect 672533 130522 672599 130525
rect 672533 130520 676292 130522
rect 672533 130464 672538 130520
rect 672594 130464 676292 130520
rect 672533 130462 676292 130464
rect 672533 130459 672599 130462
rect 675937 130114 676003 130117
rect 675937 130112 676292 130114
rect 675937 130056 675942 130112
rect 675998 130056 676292 130112
rect 675937 130054 676292 130056
rect 675937 130051 676003 130054
rect 579061 129706 579127 129709
rect 575798 129704 579127 129706
rect 575798 129648 579066 129704
rect 579122 129648 579127 129704
rect 575798 129646 579127 129648
rect 575798 129540 575858 129646
rect 579061 129643 579127 129646
rect 589641 129706 589707 129709
rect 673361 129706 673427 129709
rect 589641 129704 592572 129706
rect 589641 129648 589646 129704
rect 589702 129648 592572 129704
rect 589641 129646 592572 129648
rect 673361 129704 676292 129706
rect 673361 129648 673366 129704
rect 673422 129648 676292 129704
rect 673361 129646 676292 129648
rect 589641 129643 589707 129646
rect 673361 129643 673427 129646
rect 674097 129298 674163 129301
rect 674097 129296 676292 129298
rect 674097 129240 674102 129296
rect 674158 129240 676292 129296
rect 674097 129238 676292 129240
rect 674097 129235 674163 129238
rect 666356 128898 666938 128958
rect 666878 128890 666938 128898
rect 673494 128890 673500 128892
rect 666878 128830 673500 128890
rect 673494 128828 673500 128830
rect 673564 128828 673570 128892
rect 676630 128620 676690 128860
rect 676622 128556 676628 128620
rect 676692 128556 676698 128620
rect 668577 128346 668643 128349
rect 674046 128346 674052 128348
rect 668577 128344 674052 128346
rect 668577 128288 668582 128344
rect 668638 128288 674052 128344
rect 668577 128286 674052 128288
rect 668577 128283 668643 128286
rect 674046 128284 674052 128286
rect 674116 128284 674122 128348
rect 674281 128346 674347 128349
rect 675937 128346 676003 128349
rect 674281 128344 676003 128346
rect 674281 128288 674286 128344
rect 674342 128288 675942 128344
rect 675998 128288 676003 128344
rect 674281 128286 676003 128288
rect 674281 128283 674347 128286
rect 675937 128283 676003 128286
rect 676070 128148 676076 128212
rect 676140 128210 676146 128212
rect 676262 128210 676322 128452
rect 676140 128150 676322 128210
rect 676140 128148 676146 128150
rect 589457 128074 589523 128077
rect 589457 128072 592572 128074
rect 589457 128016 589462 128072
rect 589518 128016 592572 128072
rect 589457 128014 592572 128016
rect 589457 128011 589523 128014
rect 682334 127805 682394 128044
rect 579153 127802 579219 127805
rect 575798 127800 579219 127802
rect 575798 127744 579158 127800
rect 579214 127744 579219 127800
rect 575798 127742 579219 127744
rect 682334 127800 682443 127805
rect 682334 127744 682382 127800
rect 682438 127744 682443 127800
rect 682334 127742 682443 127744
rect 575798 127364 575858 127742
rect 579153 127739 579219 127742
rect 682377 127739 682443 127742
rect 674833 127666 674899 127669
rect 674833 127664 676292 127666
rect 674833 127608 674838 127664
rect 674894 127608 676292 127664
rect 674833 127606 676292 127608
rect 674833 127603 674899 127606
rect 675886 127196 675892 127260
rect 675956 127258 675962 127260
rect 675956 127198 676292 127258
rect 675956 127196 675962 127198
rect 676254 126924 676260 126988
rect 676324 126924 676330 126988
rect 676262 126820 676322 126924
rect 590101 126442 590167 126445
rect 675017 126442 675083 126445
rect 590101 126440 592572 126442
rect 590101 126384 590106 126440
rect 590162 126384 592572 126440
rect 590101 126382 592572 126384
rect 675017 126440 676292 126442
rect 675017 126384 675022 126440
rect 675078 126384 676292 126440
rect 675017 126382 676292 126384
rect 590101 126379 590167 126382
rect 675017 126379 675083 126382
rect 673085 126034 673151 126037
rect 673085 126032 676292 126034
rect 673085 125976 673090 126032
rect 673146 125976 676292 126032
rect 673085 125974 676292 125976
rect 673085 125971 673151 125974
rect 668761 125762 668827 125765
rect 666694 125760 668827 125762
rect 666694 125704 668766 125760
rect 668822 125704 668827 125760
rect 666694 125702 668827 125704
rect 666694 125694 666754 125702
rect 668761 125699 668827 125702
rect 666356 125634 666754 125694
rect 674649 125626 674715 125629
rect 674649 125624 676292 125626
rect 674649 125568 674654 125624
rect 674710 125568 676292 125624
rect 674649 125566 676292 125568
rect 674649 125563 674715 125566
rect 579521 125354 579587 125357
rect 575798 125352 579587 125354
rect 575798 125296 579526 125352
rect 579582 125296 579587 125352
rect 575798 125294 579587 125296
rect 575798 125188 575858 125294
rect 579521 125291 579587 125294
rect 674465 125218 674531 125221
rect 674465 125216 676292 125218
rect 674465 125160 674470 125216
rect 674526 125160 676292 125216
rect 674465 125158 676292 125160
rect 674465 125155 674531 125158
rect 589917 124810 589983 124813
rect 589917 124808 592572 124810
rect 589917 124752 589922 124808
rect 589978 124752 592572 124808
rect 589917 124750 592572 124752
rect 589917 124747 589983 124750
rect 676446 124540 676506 124780
rect 676438 124476 676444 124540
rect 676508 124476 676514 124540
rect 672901 124402 672967 124405
rect 672901 124400 676292 124402
rect 672901 124344 672906 124400
rect 672962 124344 676292 124400
rect 672901 124342 676292 124344
rect 672901 124339 672967 124342
rect 672717 124130 672783 124133
rect 666694 124128 672783 124130
rect 666694 124072 672722 124128
rect 672778 124072 672783 124128
rect 666694 124070 672783 124072
rect 666694 124062 666754 124070
rect 672717 124067 672783 124070
rect 666356 124002 666754 124062
rect 672950 123934 676292 123994
rect 672533 123858 672599 123861
rect 672950 123858 673010 123934
rect 672533 123856 673010 123858
rect 672533 123800 672538 123856
rect 672594 123800 673010 123856
rect 672533 123798 673010 123800
rect 672533 123795 672599 123798
rect 578325 123586 578391 123589
rect 575798 123584 578391 123586
rect 575798 123528 578330 123584
rect 578386 123528 578391 123584
rect 575798 123526 578391 123528
rect 575798 123012 575858 123526
rect 578325 123523 578391 123526
rect 673361 123586 673427 123589
rect 673361 123584 676292 123586
rect 673361 123528 673366 123584
rect 673422 123528 676292 123584
rect 673361 123526 676292 123528
rect 673361 123523 673427 123526
rect 589457 123178 589523 123181
rect 672349 123178 672415 123181
rect 589457 123176 592572 123178
rect 589457 123120 589462 123176
rect 589518 123120 592572 123176
rect 589457 123118 592572 123120
rect 672349 123176 676292 123178
rect 672349 123120 672354 123176
rect 672410 123120 676292 123176
rect 672349 123118 676292 123120
rect 589457 123115 589523 123118
rect 672349 123115 672415 123118
rect 669957 122770 670023 122773
rect 669957 122768 676292 122770
rect 669957 122712 669962 122768
rect 670018 122712 676292 122768
rect 669957 122710 676292 122712
rect 669957 122707 670023 122710
rect 675702 122300 675708 122364
rect 675772 122362 675778 122364
rect 675772 122302 676292 122362
rect 675772 122300 675778 122302
rect 673913 121682 673979 121685
rect 676262 121682 676322 121924
rect 673913 121680 676322 121682
rect 673913 121624 673918 121680
rect 673974 121624 676322 121680
rect 673913 121622 676322 121624
rect 673913 121619 673979 121622
rect 589273 121546 589339 121549
rect 589273 121544 592572 121546
rect 589273 121488 589278 121544
rect 589334 121488 592572 121544
rect 589273 121486 592572 121488
rect 589273 121483 589339 121486
rect 579521 121138 579587 121141
rect 575798 121136 579587 121138
rect 575798 121080 579526 121136
rect 579582 121080 579587 121136
rect 575798 121078 579587 121080
rect 575798 120836 575858 121078
rect 579521 121075 579587 121078
rect 668577 120866 668643 120869
rect 666694 120864 668643 120866
rect 666694 120808 668582 120864
rect 668638 120808 668643 120864
rect 666694 120806 668643 120808
rect 666694 120798 666754 120806
rect 668577 120803 668643 120806
rect 666356 120738 666754 120798
rect 668945 120186 669011 120189
rect 672349 120186 672415 120189
rect 668945 120184 672415 120186
rect 668945 120128 668950 120184
rect 669006 120128 672354 120184
rect 672410 120128 672415 120184
rect 668945 120126 672415 120128
rect 668945 120123 669011 120126
rect 672349 120123 672415 120126
rect 589457 119914 589523 119917
rect 589457 119912 592572 119914
rect 589457 119856 589462 119912
rect 589518 119856 592572 119912
rect 589457 119854 592572 119856
rect 589457 119851 589523 119854
rect 667933 119234 667999 119237
rect 666694 119232 667999 119234
rect 666694 119176 667938 119232
rect 667994 119176 667999 119232
rect 666694 119174 667999 119176
rect 666694 119166 666754 119174
rect 667933 119171 667999 119174
rect 666356 119106 666754 119166
rect 575982 118418 576042 118660
rect 578693 118418 578759 118421
rect 575982 118416 578759 118418
rect 575982 118360 578698 118416
rect 578754 118360 578759 118416
rect 575982 118358 578759 118360
rect 578693 118355 578759 118358
rect 589457 118282 589523 118285
rect 589457 118280 592572 118282
rect 589457 118224 589462 118280
rect 589518 118224 592572 118280
rect 589457 118222 592572 118224
rect 589457 118219 589523 118222
rect 672717 117874 672783 117877
rect 673913 117874 673979 117877
rect 672717 117872 673979 117874
rect 672717 117816 672722 117872
rect 672778 117816 673918 117872
rect 673974 117816 673979 117872
rect 672717 117814 673979 117816
rect 672717 117811 672783 117814
rect 673913 117811 673979 117814
rect 668025 117602 668091 117605
rect 666694 117600 668091 117602
rect 666694 117544 668030 117600
rect 668086 117544 668091 117600
rect 666694 117542 668091 117544
rect 666694 117534 666754 117542
rect 668025 117539 668091 117542
rect 666356 117474 666754 117534
rect 578693 116922 578759 116925
rect 575798 116920 578759 116922
rect 575798 116864 578698 116920
rect 578754 116864 578759 116920
rect 575798 116862 578759 116864
rect 575798 116484 575858 116862
rect 578693 116859 578759 116862
rect 589457 116650 589523 116653
rect 589457 116648 592572 116650
rect 589457 116592 589462 116648
rect 589518 116592 592572 116648
rect 589457 116590 592572 116592
rect 589457 116587 589523 116590
rect 666356 115842 666754 115902
rect 666694 115834 666754 115842
rect 671889 115834 671955 115837
rect 666694 115832 671955 115834
rect 666694 115776 671894 115832
rect 671950 115776 671955 115832
rect 666694 115774 671955 115776
rect 671889 115771 671955 115774
rect 588537 115018 588603 115021
rect 588537 115016 592572 115018
rect 588537 114960 588542 115016
rect 588598 114960 592572 115016
rect 588537 114958 592572 114960
rect 588537 114955 588603 114958
rect 579245 114474 579311 114477
rect 575798 114472 579311 114474
rect 575798 114416 579250 114472
rect 579306 114416 579311 114472
rect 575798 114414 579311 114416
rect 575798 114308 575858 114414
rect 579245 114411 579311 114414
rect 668945 114338 669011 114341
rect 666694 114336 669011 114338
rect 666694 114280 668950 114336
rect 669006 114280 669011 114336
rect 666694 114278 669011 114280
rect 666694 114270 666754 114278
rect 668945 114275 669011 114278
rect 666356 114210 666754 114270
rect 589457 113386 589523 113389
rect 589457 113384 592572 113386
rect 589457 113328 589462 113384
rect 589518 113328 592572 113384
rect 589457 113326 592572 113328
rect 589457 113323 589523 113326
rect 675293 113114 675359 113117
rect 676622 113114 676628 113116
rect 675293 113112 676628 113114
rect 675293 113056 675298 113112
rect 675354 113056 676628 113112
rect 675293 113054 676628 113056
rect 675293 113051 675359 113054
rect 676622 113052 676628 113054
rect 676692 113052 676698 113116
rect 668117 112706 668183 112709
rect 666694 112704 668183 112706
rect 666694 112648 668122 112704
rect 668178 112648 668183 112704
rect 666694 112646 668183 112648
rect 666694 112638 666754 112646
rect 668117 112643 668183 112646
rect 666356 112578 666754 112638
rect 579153 112570 579219 112573
rect 575798 112568 579219 112570
rect 575798 112512 579158 112568
rect 579214 112512 579219 112568
rect 575798 112510 579219 112512
rect 575798 112132 575858 112510
rect 579153 112507 579219 112510
rect 668577 111890 668643 111893
rect 674097 111890 674163 111893
rect 668577 111888 674163 111890
rect 668577 111832 668582 111888
rect 668638 111832 674102 111888
rect 674158 111832 674163 111888
rect 668577 111830 674163 111832
rect 668577 111827 668643 111830
rect 674097 111827 674163 111830
rect 589365 111754 589431 111757
rect 589365 111752 592572 111754
rect 589365 111696 589370 111752
rect 589426 111696 592572 111752
rect 589365 111694 592572 111696
rect 589365 111691 589431 111694
rect 673085 111482 673151 111485
rect 675109 111482 675175 111485
rect 673085 111480 675175 111482
rect 673085 111424 673090 111480
rect 673146 111424 675114 111480
rect 675170 111424 675175 111480
rect 673085 111422 675175 111424
rect 673085 111419 673151 111422
rect 675109 111419 675175 111422
rect 672717 111074 672783 111077
rect 666694 111072 672783 111074
rect 666694 111016 672722 111072
rect 672778 111016 672783 111072
rect 666694 111014 672783 111016
rect 666694 111006 666754 111014
rect 672717 111011 672783 111014
rect 666356 110946 666754 111006
rect 578877 110394 578943 110397
rect 575798 110392 578943 110394
rect 575798 110336 578882 110392
rect 578938 110336 578943 110392
rect 575798 110334 578943 110336
rect 575798 109956 575858 110334
rect 578877 110331 578943 110334
rect 672533 110258 672599 110261
rect 674649 110258 674715 110261
rect 672533 110256 674715 110258
rect 672533 110200 672538 110256
rect 672594 110200 674654 110256
rect 674710 110200 674715 110256
rect 672533 110198 674715 110200
rect 672533 110195 672599 110198
rect 674649 110195 674715 110198
rect 590101 110122 590167 110125
rect 590101 110120 592572 110122
rect 590101 110064 590106 110120
rect 590162 110064 592572 110120
rect 590101 110062 592572 110064
rect 590101 110059 590167 110062
rect 666645 109374 666711 109377
rect 666356 109372 666711 109374
rect 666356 109316 666650 109372
rect 666706 109316 666711 109372
rect 666356 109314 666711 109316
rect 666645 109311 666711 109314
rect 589457 108490 589523 108493
rect 589457 108488 592572 108490
rect 589457 108432 589462 108488
rect 589518 108432 592572 108488
rect 589457 108430 592572 108432
rect 589457 108427 589523 108430
rect 578877 108354 578943 108357
rect 575798 108352 578943 108354
rect 575798 108296 578882 108352
rect 578938 108296 578943 108352
rect 575798 108294 578943 108296
rect 575798 107780 575858 108294
rect 578877 108291 578943 108294
rect 675661 108082 675727 108085
rect 675886 108082 675892 108084
rect 675661 108080 675892 108082
rect 675661 108024 675666 108080
rect 675722 108024 675892 108080
rect 675661 108022 675892 108024
rect 675661 108019 675727 108022
rect 675886 108020 675892 108022
rect 675956 108020 675962 108084
rect 671521 107810 671587 107813
rect 666694 107808 671587 107810
rect 666694 107752 671526 107808
rect 671582 107752 671587 107808
rect 666694 107750 671587 107752
rect 666694 107742 666754 107750
rect 671521 107747 671587 107750
rect 666356 107682 666754 107742
rect 589457 106858 589523 106861
rect 589457 106856 592572 106858
rect 589457 106800 589462 106856
rect 589518 106800 592572 106856
rect 589457 106798 592572 106800
rect 589457 106795 589523 106798
rect 672349 106450 672415 106453
rect 675109 106450 675175 106453
rect 672349 106448 675175 106450
rect 672349 106392 672354 106448
rect 672410 106392 675114 106448
rect 675170 106392 675175 106448
rect 672349 106390 675175 106392
rect 672349 106387 672415 106390
rect 675109 106387 675175 106390
rect 668117 106178 668183 106181
rect 668393 106178 668459 106181
rect 666694 106176 668459 106178
rect 666694 106120 668122 106176
rect 668178 106120 668398 106176
rect 668454 106120 668459 106176
rect 666694 106118 668459 106120
rect 666694 106110 666754 106118
rect 668117 106115 668183 106118
rect 668393 106115 668459 106118
rect 675753 106178 675819 106181
rect 676438 106178 676444 106180
rect 675753 106176 676444 106178
rect 675753 106120 675758 106176
rect 675814 106120 676444 106176
rect 675753 106118 676444 106120
rect 675753 106115 675819 106118
rect 676438 106116 676444 106118
rect 676508 106116 676514 106180
rect 666356 106050 666754 106110
rect 579061 105906 579127 105909
rect 575798 105904 579127 105906
rect 575798 105848 579066 105904
rect 579122 105848 579127 105904
rect 575798 105846 579127 105848
rect 575798 105604 575858 105846
rect 579061 105843 579127 105846
rect 673361 105634 673427 105637
rect 675109 105634 675175 105637
rect 673361 105632 675175 105634
rect 673361 105576 673366 105632
rect 673422 105576 675114 105632
rect 675170 105576 675175 105632
rect 673361 105574 675175 105576
rect 673361 105571 673427 105574
rect 675109 105571 675175 105574
rect 589457 105226 589523 105229
rect 589457 105224 592572 105226
rect 589457 105168 589462 105224
rect 589518 105168 592572 105224
rect 589457 105166 592572 105168
rect 589457 105163 589523 105166
rect 668577 104546 668643 104549
rect 666694 104544 668643 104546
rect 666694 104488 668582 104544
rect 668638 104488 668643 104544
rect 666694 104486 668643 104488
rect 666694 104478 666754 104486
rect 668577 104483 668643 104486
rect 666356 104418 666754 104478
rect 589549 103594 589615 103597
rect 589549 103592 592572 103594
rect 589549 103536 589554 103592
rect 589610 103536 592572 103592
rect 589549 103534 592572 103536
rect 589549 103531 589615 103534
rect 575982 103322 576042 103428
rect 578325 103322 578391 103325
rect 575982 103320 578391 103322
rect 575982 103264 578330 103320
rect 578386 103264 578391 103320
rect 575982 103262 578391 103264
rect 578325 103259 578391 103262
rect 675753 103186 675819 103189
rect 676070 103186 676076 103188
rect 675753 103184 676076 103186
rect 675753 103128 675758 103184
rect 675814 103128 676076 103184
rect 675753 103126 676076 103128
rect 675753 103123 675819 103126
rect 676070 103124 676076 103126
rect 676140 103124 676146 103188
rect 666356 102786 666938 102846
rect 666878 102778 666938 102786
rect 667933 102778 667999 102781
rect 666878 102776 673470 102778
rect 666878 102720 667938 102776
rect 667994 102720 673470 102776
rect 666878 102718 673470 102720
rect 667933 102715 667999 102718
rect 673410 102370 673470 102718
rect 675661 102644 675727 102645
rect 675661 102640 675708 102644
rect 675772 102642 675778 102644
rect 675661 102584 675666 102640
rect 675661 102580 675708 102584
rect 675772 102582 675818 102642
rect 675772 102580 675778 102582
rect 675661 102579 675727 102580
rect 674281 102370 674347 102373
rect 673410 102368 674347 102370
rect 673410 102312 674286 102368
rect 674342 102312 674347 102368
rect 673410 102310 674347 102312
rect 674281 102307 674347 102310
rect 589917 101962 589983 101965
rect 589917 101960 592572 101962
rect 589917 101904 589922 101960
rect 589978 101904 592572 101960
rect 589917 101902 592572 101904
rect 589917 101899 589983 101902
rect 578509 101690 578575 101693
rect 575798 101688 578575 101690
rect 575798 101632 578514 101688
rect 578570 101632 578575 101688
rect 575798 101630 578575 101632
rect 575798 101252 575858 101630
rect 578509 101627 578575 101630
rect 675753 101418 675819 101421
rect 676254 101418 676260 101420
rect 675753 101416 676260 101418
rect 675753 101360 675758 101416
rect 675814 101360 676260 101416
rect 675753 101358 676260 101360
rect 675753 101355 675819 101358
rect 676254 101356 676260 101358
rect 676324 101356 676330 101420
rect 579245 99242 579311 99245
rect 575798 99240 579311 99242
rect 575798 99184 579250 99240
rect 579306 99184 579311 99240
rect 575798 99182 579311 99184
rect 575798 99076 575858 99182
rect 579245 99179 579311 99182
rect 578325 97474 578391 97477
rect 575798 97472 578391 97474
rect 575798 97416 578330 97472
rect 578386 97416 578391 97472
rect 575798 97414 578391 97416
rect 575798 96900 575858 97414
rect 578325 97411 578391 97414
rect 637021 96930 637087 96933
rect 637246 96930 637252 96932
rect 637021 96928 637252 96930
rect 637021 96872 637026 96928
rect 637082 96872 637252 96928
rect 637021 96870 637252 96872
rect 637021 96867 637087 96870
rect 637246 96868 637252 96870
rect 637316 96868 637322 96932
rect 633934 96052 633940 96116
rect 634004 96114 634010 96116
rect 635733 96114 635799 96117
rect 634004 96112 635799 96114
rect 634004 96056 635738 96112
rect 635794 96056 635799 96112
rect 634004 96054 635799 96056
rect 634004 96052 634010 96054
rect 635733 96051 635799 96054
rect 613377 95842 613443 95845
rect 668301 95842 668367 95845
rect 613377 95840 668367 95842
rect 613377 95784 613382 95840
rect 613438 95784 668306 95840
rect 668362 95784 668367 95840
rect 613377 95782 668367 95784
rect 613377 95779 613443 95782
rect 668301 95779 668367 95782
rect 646221 95570 646287 95573
rect 647693 95570 647759 95573
rect 646221 95568 647759 95570
rect 646221 95512 646226 95568
rect 646282 95512 647698 95568
rect 647754 95512 647759 95568
rect 646221 95510 647759 95512
rect 646221 95507 646287 95510
rect 647693 95507 647759 95510
rect 579429 95026 579495 95029
rect 575798 95024 579495 95026
rect 575798 94968 579434 95024
rect 579490 94968 579495 95024
rect 575798 94966 579495 94968
rect 575798 94724 575858 94966
rect 579429 94963 579495 94966
rect 647325 95026 647391 95029
rect 647325 95024 647434 95026
rect 647325 94968 647330 95024
rect 647386 94968 647434 95024
rect 647325 94963 647434 94968
rect 626441 94482 626507 94485
rect 626441 94480 628268 94482
rect 626441 94424 626446 94480
rect 626502 94424 628268 94480
rect 647374 94452 647434 94963
rect 626441 94422 628268 94424
rect 626441 94419 626507 94422
rect 655053 94210 655119 94213
rect 655053 94208 656788 94210
rect 655053 94152 655058 94208
rect 655114 94152 656788 94208
rect 655053 94150 656788 94152
rect 655053 94147 655119 94150
rect 625981 93666 626047 93669
rect 625981 93664 628268 93666
rect 625981 93608 625986 93664
rect 626042 93608 628268 93664
rect 625981 93606 628268 93608
rect 625981 93603 626047 93606
rect 654593 93394 654659 93397
rect 665357 93394 665423 93397
rect 654593 93392 656788 93394
rect 654593 93336 654598 93392
rect 654654 93336 656788 93392
rect 654593 93334 656788 93336
rect 663596 93392 665423 93394
rect 663596 93336 665362 93392
rect 665418 93336 665423 93392
rect 663596 93334 665423 93336
rect 654593 93331 654659 93334
rect 665357 93331 665423 93334
rect 579521 93122 579587 93125
rect 575798 93120 579587 93122
rect 575798 93064 579526 93120
rect 579582 93064 579587 93120
rect 575798 93062 579587 93064
rect 575798 92548 575858 93062
rect 579521 93059 579587 93062
rect 626441 92850 626507 92853
rect 663701 92850 663767 92853
rect 626441 92848 628268 92850
rect 626441 92792 626446 92848
rect 626502 92792 628268 92848
rect 626441 92790 628268 92792
rect 663382 92848 663767 92850
rect 663382 92792 663706 92848
rect 663762 92792 663767 92848
rect 663382 92790 663767 92792
rect 626441 92787 626507 92790
rect 655421 92578 655487 92581
rect 655421 92576 656788 92578
rect 655421 92520 655426 92576
rect 655482 92520 656788 92576
rect 663382 92548 663442 92790
rect 663701 92787 663767 92790
rect 655421 92518 656788 92520
rect 655421 92515 655487 92518
rect 625797 92034 625863 92037
rect 648613 92034 648679 92037
rect 625797 92032 628268 92034
rect 625797 91976 625802 92032
rect 625858 91976 628268 92032
rect 625797 91974 628268 91976
rect 648140 92032 648679 92034
rect 648140 91976 648618 92032
rect 648674 91976 648679 92032
rect 648140 91974 648679 91976
rect 625797 91971 625863 91974
rect 648613 91971 648679 91974
rect 664529 91762 664595 91765
rect 663596 91760 664595 91762
rect 663596 91704 664534 91760
rect 664590 91704 664595 91760
rect 663596 91702 664595 91704
rect 664529 91699 664595 91702
rect 655237 91490 655303 91493
rect 655237 91488 656788 91490
rect 655237 91432 655242 91488
rect 655298 91432 656788 91488
rect 655237 91430 656788 91432
rect 655237 91427 655303 91430
rect 626441 91218 626507 91221
rect 626441 91216 628268 91218
rect 626441 91160 626446 91216
rect 626502 91160 628268 91216
rect 626441 91158 628268 91160
rect 626441 91155 626507 91158
rect 579337 90946 579403 90949
rect 575798 90944 579403 90946
rect 575798 90888 579342 90944
rect 579398 90888 579403 90944
rect 575798 90886 579403 90888
rect 575798 90372 575858 90886
rect 579337 90883 579403 90886
rect 651833 90674 651899 90677
rect 664345 90674 664411 90677
rect 651833 90672 656788 90674
rect 651833 90616 651838 90672
rect 651894 90616 656788 90672
rect 651833 90614 656788 90616
rect 663596 90672 664411 90674
rect 663596 90616 664350 90672
rect 664406 90616 664411 90672
rect 663596 90614 664411 90616
rect 651833 90611 651899 90614
rect 664345 90611 664411 90614
rect 626441 90402 626507 90405
rect 626441 90400 628268 90402
rect 626441 90344 626446 90400
rect 626502 90344 628268 90400
rect 626441 90342 628268 90344
rect 626441 90339 626507 90342
rect 655789 89858 655855 89861
rect 664161 89858 664227 89861
rect 655789 89856 656788 89858
rect 655789 89800 655794 89856
rect 655850 89800 656788 89856
rect 655789 89798 656788 89800
rect 663596 89856 664227 89858
rect 663596 89800 664166 89856
rect 664222 89800 664227 89856
rect 663596 89798 664227 89800
rect 655789 89795 655855 89798
rect 664161 89795 664227 89798
rect 626257 89586 626323 89589
rect 650453 89586 650519 89589
rect 626257 89584 628268 89586
rect 626257 89528 626262 89584
rect 626318 89528 628268 89584
rect 626257 89526 628268 89528
rect 648140 89584 650519 89586
rect 648140 89528 650458 89584
rect 650514 89528 650519 89584
rect 648140 89526 650519 89528
rect 626257 89523 626323 89526
rect 650453 89523 650519 89526
rect 665173 89042 665239 89045
rect 663596 89040 665239 89042
rect 663596 88984 665178 89040
rect 665234 88984 665239 89040
rect 663596 88982 665239 88984
rect 665173 88979 665239 88982
rect 626441 88770 626507 88773
rect 626441 88768 628268 88770
rect 626441 88712 626446 88768
rect 626502 88712 628268 88768
rect 626441 88710 628268 88712
rect 626441 88707 626507 88710
rect 575982 88090 576042 88196
rect 579521 88090 579587 88093
rect 575982 88088 579587 88090
rect 575982 88032 579526 88088
rect 579582 88032 579587 88088
rect 575982 88030 579587 88032
rect 579521 88027 579587 88030
rect 626441 87954 626507 87957
rect 626441 87952 628268 87954
rect 626441 87896 626446 87952
rect 626502 87896 628268 87952
rect 626441 87894 628268 87896
rect 626441 87891 626507 87894
rect 626257 87138 626323 87141
rect 650177 87138 650243 87141
rect 626257 87136 628268 87138
rect 626257 87080 626262 87136
rect 626318 87080 628268 87136
rect 626257 87078 628268 87080
rect 648140 87136 650243 87138
rect 648140 87080 650182 87136
rect 650238 87080 650243 87136
rect 648140 87078 650243 87080
rect 626257 87075 626323 87078
rect 650177 87075 650243 87078
rect 578325 86458 578391 86461
rect 575798 86456 578391 86458
rect 575798 86400 578330 86456
rect 578386 86400 578391 86456
rect 575798 86398 578391 86400
rect 575798 86020 575858 86398
rect 578325 86395 578391 86398
rect 626441 86322 626507 86325
rect 626441 86320 628268 86322
rect 626441 86264 626446 86320
rect 626502 86264 628268 86320
rect 626441 86262 628268 86264
rect 626441 86259 626507 86262
rect 626441 85506 626507 85509
rect 626441 85504 628268 85506
rect 626441 85448 626446 85504
rect 626502 85448 628268 85504
rect 626441 85446 628268 85448
rect 626441 85443 626507 85446
rect 625245 84690 625311 84693
rect 650729 84690 650795 84693
rect 625245 84688 628268 84690
rect 625245 84632 625250 84688
rect 625306 84632 628268 84688
rect 625245 84630 628268 84632
rect 648140 84688 650795 84690
rect 648140 84632 650734 84688
rect 650790 84632 650795 84688
rect 648140 84630 650795 84632
rect 625245 84627 625311 84630
rect 650729 84627 650795 84630
rect 579521 84010 579587 84013
rect 575798 84008 579587 84010
rect 575798 83952 579526 84008
rect 579582 83952 579587 84008
rect 575798 83950 579587 83952
rect 575798 83844 575858 83950
rect 579521 83947 579587 83950
rect 625797 83874 625863 83877
rect 625797 83872 628268 83874
rect 625797 83816 625802 83872
rect 625858 83816 628268 83872
rect 625797 83814 628268 83816
rect 625797 83811 625863 83814
rect 628741 83330 628807 83333
rect 628741 83328 628850 83330
rect 628741 83272 628746 83328
rect 628802 83272 628850 83328
rect 628741 83267 628850 83272
rect 628790 83028 628850 83267
rect 647509 82786 647575 82789
rect 647509 82784 647618 82786
rect 647509 82728 647514 82784
rect 647570 82728 647618 82784
rect 647509 82723 647618 82728
rect 579429 82242 579495 82245
rect 575798 82240 579495 82242
rect 575798 82184 579434 82240
rect 579490 82184 579495 82240
rect 647558 82212 647618 82723
rect 575798 82182 579495 82184
rect 575798 81668 575858 82182
rect 579429 82179 579495 82182
rect 628790 81698 628850 82212
rect 629201 81698 629267 81701
rect 628790 81696 629267 81698
rect 628790 81640 629206 81696
rect 629262 81640 629267 81696
rect 628790 81638 629267 81640
rect 629201 81635 629267 81638
rect 578877 80066 578943 80069
rect 575798 80064 578943 80066
rect 575798 80008 578882 80064
rect 578938 80008 578943 80064
rect 575798 80006 578943 80008
rect 575798 79492 575858 80006
rect 578877 80003 578943 80006
rect 633893 78572 633959 78573
rect 633893 78570 633940 78572
rect 633848 78568 633940 78570
rect 633848 78512 633898 78568
rect 633848 78510 633940 78512
rect 633893 78508 633940 78510
rect 634004 78508 634010 78572
rect 633893 78507 633959 78508
rect 578417 77890 578483 77893
rect 575798 77888 578483 77890
rect 575798 77832 578422 77888
rect 578478 77832 578483 77888
rect 575798 77830 578483 77832
rect 575798 77316 575858 77830
rect 578417 77827 578483 77830
rect 583017 77890 583083 77893
rect 637062 77890 637068 77892
rect 583017 77888 637068 77890
rect 583017 77832 583022 77888
rect 583078 77832 637068 77888
rect 583017 77830 637068 77832
rect 583017 77827 583083 77830
rect 637062 77828 637068 77830
rect 637132 77890 637138 77892
rect 639597 77890 639663 77893
rect 637132 77888 639663 77890
rect 637132 77832 639602 77888
rect 639658 77832 639663 77888
rect 637132 77830 639663 77832
rect 637132 77828 637138 77830
rect 639597 77827 639663 77830
rect 589917 77346 589983 77349
rect 633893 77346 633959 77349
rect 589917 77344 633959 77346
rect 589917 77288 589922 77344
rect 589978 77288 633898 77344
rect 633954 77288 633959 77344
rect 589917 77286 633959 77288
rect 589917 77283 589983 77286
rect 633893 77283 633959 77286
rect 578325 75714 578391 75717
rect 575798 75712 578391 75714
rect 575798 75656 578330 75712
rect 578386 75656 578391 75712
rect 575798 75654 578391 75656
rect 575798 75140 575858 75654
rect 578325 75651 578391 75654
rect 646405 74490 646471 74493
rect 646405 74488 646514 74490
rect 646405 74432 646410 74488
rect 646466 74432 646514 74488
rect 646405 74427 646514 74432
rect 646454 73848 646514 74427
rect 579521 73130 579587 73133
rect 575798 73128 579587 73130
rect 575798 73072 579526 73128
rect 579582 73072 579587 73128
rect 575798 73070 579587 73072
rect 575798 72964 575858 73070
rect 579521 73067 579587 73070
rect 647233 71770 647299 71773
rect 646638 71768 647299 71770
rect 646638 71712 647238 71768
rect 647294 71712 647299 71768
rect 646638 71710 647299 71712
rect 646638 71400 646698 71710
rect 647233 71707 647299 71710
rect 579521 71226 579587 71229
rect 575798 71224 579587 71226
rect 575798 71168 579526 71224
rect 579582 71168 579587 71224
rect 575798 71166 579587 71168
rect 575798 70788 575858 71166
rect 579521 71163 579587 71166
rect 646221 69186 646287 69189
rect 646221 69184 646330 69186
rect 646221 69128 646226 69184
rect 646282 69128 646330 69184
rect 646221 69123 646330 69128
rect 646270 68952 646330 69123
rect 646221 67146 646287 67149
rect 646221 67144 646330 67146
rect 646221 67088 646226 67144
rect 646282 67088 646330 67144
rect 646221 67083 646330 67088
rect 646270 66504 646330 67083
rect 575982 66330 576042 66436
rect 579521 66330 579587 66333
rect 575982 66328 579587 66330
rect 575982 66272 579526 66328
rect 579582 66272 579587 66328
rect 575982 66270 579587 66272
rect 579521 66267 579587 66270
rect 579521 64562 579587 64565
rect 575798 64560 579587 64562
rect 575798 64504 579526 64560
rect 579582 64504 579587 64560
rect 575798 64502 579587 64504
rect 575798 64260 575858 64502
rect 579521 64499 579587 64502
rect 649073 64426 649139 64429
rect 646638 64424 649139 64426
rect 646638 64368 649078 64424
rect 649134 64368 649139 64424
rect 646638 64366 649139 64368
rect 646638 64056 646698 64366
rect 649073 64363 649139 64366
rect 648705 62114 648771 62117
rect 646638 62112 648771 62114
rect 575982 61842 576042 62084
rect 646638 62056 648710 62112
rect 648766 62056 648771 62112
rect 646638 62054 648771 62056
rect 578509 61842 578575 61845
rect 575982 61840 578575 61842
rect 575982 61784 578514 61840
rect 578570 61784 578575 61840
rect 575982 61782 578575 61784
rect 578509 61779 578575 61782
rect 646638 61608 646698 62054
rect 648705 62051 648771 62054
rect 578877 60482 578943 60485
rect 575798 60480 578943 60482
rect 575798 60424 578882 60480
rect 578938 60424 578943 60480
rect 575798 60422 578943 60424
rect 575798 59908 575858 60422
rect 578877 60419 578943 60422
rect 646405 59394 646471 59397
rect 646405 59392 646514 59394
rect 646405 59336 646410 59392
rect 646466 59336 646514 59392
rect 646405 59331 646514 59336
rect 646454 59160 646514 59331
rect 579521 57898 579587 57901
rect 575798 57896 579587 57898
rect 575798 57840 579526 57896
rect 579582 57840 579587 57896
rect 575798 57838 579587 57840
rect 575798 57732 575858 57838
rect 579521 57835 579587 57838
rect 648889 57354 648955 57357
rect 646638 57352 648955 57354
rect 646638 57296 648894 57352
rect 648950 57296 648955 57352
rect 646638 57294 648955 57296
rect 646638 56712 646698 57294
rect 648889 57291 648955 57294
rect 579521 56130 579587 56133
rect 575798 56128 579587 56130
rect 575798 56072 579526 56128
rect 579582 56072 579587 56128
rect 575798 56070 579587 56072
rect 575798 55556 575858 56070
rect 579521 56067 579587 56070
rect 577497 55042 577563 55045
rect 459878 55040 577563 55042
rect 459878 54984 577502 55040
rect 577558 54984 577563 55040
rect 459878 54982 577563 54984
rect 459878 53685 459938 54982
rect 577497 54979 577563 54982
rect 585777 54770 585843 54773
rect 462454 54768 585843 54770
rect 462454 54712 585782 54768
rect 585838 54712 585843 54768
rect 462454 54710 585843 54712
rect 462454 54226 462514 54710
rect 585777 54707 585843 54710
rect 462630 54436 462636 54500
rect 462700 54498 462706 54500
rect 604453 54498 604519 54501
rect 462700 54496 604519 54498
rect 462700 54440 604458 54496
rect 604514 54440 604519 54496
rect 462700 54438 604519 54440
rect 462700 54436 462706 54438
rect 604453 54435 604519 54438
rect 576853 54226 576919 54229
rect 460798 54166 462514 54226
rect 466410 54224 576919 54226
rect 466410 54168 576858 54224
rect 576914 54168 576919 54224
rect 466410 54166 576919 54168
rect 460798 53685 460858 54166
rect 466410 53954 466470 54166
rect 576853 54163 576919 54166
rect 461718 53894 466470 53954
rect 461718 53685 461778 53894
rect 459829 53680 459938 53685
rect 459829 53624 459834 53680
rect 459890 53624 459938 53680
rect 459829 53622 459938 53624
rect 460749 53680 460858 53685
rect 460749 53624 460754 53680
rect 460810 53624 460858 53680
rect 460749 53622 460858 53624
rect 461669 53680 461778 53685
rect 462589 53684 462655 53685
rect 462589 53682 462636 53684
rect 461669 53624 461674 53680
rect 461730 53624 461778 53680
rect 461669 53622 461778 53624
rect 462544 53680 462636 53682
rect 462544 53624 462594 53680
rect 462544 53622 462636 53624
rect 459829 53619 459895 53622
rect 460749 53619 460815 53622
rect 461669 53619 461735 53622
rect 462589 53620 462636 53622
rect 462700 53620 462706 53684
rect 464337 53682 464403 53685
rect 482277 53682 482343 53685
rect 464337 53680 482343 53682
rect 464337 53624 464342 53680
rect 464398 53624 482282 53680
rect 482338 53624 482343 53680
rect 464337 53622 482343 53624
rect 462589 53619 462655 53620
rect 464337 53619 464403 53622
rect 482277 53619 482343 53622
rect 472525 53410 472591 53413
rect 481725 53410 481791 53413
rect 472525 53408 481791 53410
rect 472525 53352 472530 53408
rect 472586 53352 481730 53408
rect 481786 53352 481791 53408
rect 472525 53350 481791 53352
rect 472525 53347 472591 53350
rect 481725 53347 481791 53350
rect 194358 50220 194364 50284
rect 194428 50282 194434 50284
rect 308029 50282 308095 50285
rect 194428 50280 308095 50282
rect 194428 50224 308034 50280
rect 308090 50224 308095 50280
rect 194428 50222 308095 50224
rect 194428 50220 194434 50222
rect 308029 50219 308095 50222
rect 529790 50220 529796 50284
rect 529860 50282 529866 50284
rect 553669 50282 553735 50285
rect 529860 50280 553735 50282
rect 529860 50224 553674 50280
rect 553730 50224 553735 50280
rect 529860 50222 553735 50224
rect 529860 50220 529866 50222
rect 553669 50219 553735 50222
rect 518750 48860 518756 48924
rect 518820 48922 518826 48924
rect 549989 48922 550055 48925
rect 518820 48920 550055 48922
rect 518820 48864 549994 48920
rect 550050 48864 550055 48920
rect 518820 48862 550055 48864
rect 518820 48860 518826 48862
rect 549989 48859 550055 48862
rect 663793 48514 663859 48517
rect 662094 48512 663859 48514
rect 661480 48456 663798 48512
rect 663854 48456 663859 48512
rect 661480 48454 663859 48456
rect 661480 48452 662154 48454
rect 663793 48451 663859 48454
rect 526478 48044 526484 48108
rect 526548 48106 526554 48108
rect 552013 48106 552079 48109
rect 526548 48104 552079 48106
rect 526548 48048 552018 48104
rect 552074 48048 552079 48104
rect 526548 48046 552079 48048
rect 526548 48044 526554 48046
rect 552013 48043 552079 48046
rect 520958 47772 520964 47836
rect 521028 47834 521034 47836
rect 547873 47834 547939 47837
rect 521028 47832 547939 47834
rect 521028 47776 547878 47832
rect 547934 47776 547939 47832
rect 661585 47791 661651 47794
rect 521028 47774 547939 47776
rect 521028 47772 521034 47774
rect 547873 47771 547939 47774
rect 661388 47789 661651 47791
rect 661388 47733 661590 47789
rect 661646 47733 661651 47789
rect 661388 47731 661651 47733
rect 661585 47728 661651 47731
rect 515438 47500 515444 47564
rect 515508 47562 515514 47564
rect 544009 47562 544075 47565
rect 515508 47560 544075 47562
rect 515508 47504 544014 47560
rect 544070 47504 544075 47560
rect 515508 47502 544075 47504
rect 515508 47500 515514 47502
rect 544009 47499 544075 47502
rect 662413 47426 662479 47429
rect 661388 47424 662479 47426
rect 661388 47368 662418 47424
rect 662474 47368 662479 47424
rect 661388 47366 662479 47368
rect 662413 47363 662479 47366
rect 522062 47228 522068 47292
rect 522132 47290 522138 47292
rect 545665 47290 545731 47293
rect 522132 47288 545731 47290
rect 522132 47232 545670 47288
rect 545726 47232 545731 47288
rect 522132 47230 545731 47232
rect 522132 47228 522138 47230
rect 545665 47227 545731 47230
rect 458173 47018 458239 47021
rect 465257 47018 465323 47021
rect 458173 47016 465323 47018
rect 458173 46960 458178 47016
rect 458234 46960 465262 47016
rect 465318 46960 465323 47016
rect 458173 46958 465323 46960
rect 458173 46955 458239 46958
rect 465257 46955 465323 46958
rect 458357 46746 458423 46749
rect 465073 46746 465139 46749
rect 458357 46744 465139 46746
rect 458357 46688 458362 46744
rect 458418 46688 465078 46744
rect 465134 46688 465139 46744
rect 458357 46686 465139 46688
rect 458357 46683 458423 46686
rect 465073 46683 465139 46686
rect 431217 44842 431283 44845
rect 460105 44842 460171 44845
rect 431217 44840 460171 44842
rect 431217 44784 431222 44840
rect 431278 44784 460110 44840
rect 460166 44784 460171 44840
rect 431217 44782 460171 44784
rect 431217 44779 431283 44782
rect 460105 44779 460171 44782
rect 437246 44374 441170 44434
rect 142613 44298 142679 44301
rect 142110 44296 142679 44298
rect 142110 44240 142618 44296
rect 142674 44240 142679 44296
rect 142110 44238 142679 44240
rect 141734 43964 141740 44028
rect 141804 44026 141810 44028
rect 142110 44026 142170 44238
rect 142613 44235 142679 44238
rect 307293 44162 307359 44165
rect 437246 44162 437306 44374
rect 441110 44162 441170 44374
rect 461342 44372 461348 44436
rect 461412 44434 461418 44436
rect 461945 44434 462011 44437
rect 461412 44432 462011 44434
rect 461412 44376 461950 44432
rect 462006 44376 462011 44432
rect 461412 44374 462011 44376
rect 461412 44372 461418 44374
rect 461945 44371 462011 44374
rect 462262 44372 462268 44436
rect 462332 44434 462338 44436
rect 462497 44434 462563 44437
rect 462332 44432 462563 44434
rect 462332 44376 462502 44432
rect 462558 44376 462563 44432
rect 462332 44374 462563 44376
rect 462332 44372 462338 44374
rect 462497 44371 462563 44374
rect 463877 44162 463943 44165
rect 307293 44160 437306 44162
rect 307293 44104 307298 44160
rect 307354 44104 437306 44160
rect 307293 44102 437306 44104
rect 437430 44102 440986 44162
rect 441110 44160 463943 44162
rect 441110 44104 463882 44160
rect 463938 44104 463943 44160
rect 441110 44102 463943 44104
rect 307293 44099 307359 44102
rect 141804 43966 142170 44026
rect 141804 43964 141810 43966
rect 361757 43618 361823 43621
rect 437430 43618 437490 44102
rect 440926 43890 440986 44102
rect 463877 44099 463943 44102
rect 460841 43890 460907 43893
rect 471053 43890 471119 43893
rect 440926 43830 441630 43890
rect 361757 43616 437490 43618
rect 361757 43560 361762 43616
rect 361818 43560 437490 43616
rect 361757 43558 437490 43560
rect 441570 43618 441630 43830
rect 460841 43888 471119 43890
rect 460841 43832 460846 43888
rect 460902 43832 471058 43888
rect 471114 43832 471119 43888
rect 460841 43830 471119 43832
rect 460841 43827 460907 43830
rect 471053 43827 471119 43830
rect 464337 43618 464403 43621
rect 441570 43616 464403 43618
rect 441570 43560 464342 43616
rect 464398 43560 464403 43616
rect 441570 43558 464403 43560
rect 361757 43555 361823 43558
rect 464337 43555 464403 43558
rect 462313 43210 462379 43213
rect 465809 43210 465875 43213
rect 462313 43208 465875 43210
rect 462313 43152 462318 43208
rect 462374 43152 465814 43208
rect 465870 43152 465875 43208
rect 462313 43150 465875 43152
rect 462313 43147 462379 43150
rect 465809 43147 465875 43150
rect 461761 42938 461827 42941
rect 463693 42938 463759 42941
rect 461761 42936 463759 42938
rect 461761 42880 461766 42936
rect 461822 42880 463698 42936
rect 463754 42880 463759 42936
rect 461761 42878 463759 42880
rect 461761 42875 461827 42878
rect 463693 42875 463759 42878
rect 518801 42804 518867 42805
rect 518750 42802 518756 42804
rect 518710 42742 518756 42802
rect 518820 42800 518867 42804
rect 518862 42744 518867 42800
rect 518750 42740 518756 42742
rect 518820 42740 518867 42744
rect 518801 42739 518867 42740
rect 416589 42394 416655 42397
rect 416589 42392 422310 42394
rect 416589 42336 416594 42392
rect 416650 42336 422310 42392
rect 416589 42334 422310 42336
rect 416589 42331 416655 42334
rect 422250 42258 422310 42334
rect 446397 42258 446463 42261
rect 461117 42258 461183 42261
rect 422250 42198 427830 42258
rect 194317 42124 194383 42125
rect 194317 42122 194364 42124
rect 194272 42120 194364 42122
rect 194272 42064 194322 42120
rect 194272 42062 194364 42064
rect 194317 42060 194364 42062
rect 194428 42060 194434 42124
rect 415761 42122 415827 42125
rect 421966 42122 421972 42124
rect 415761 42120 421972 42122
rect 415761 42064 415766 42120
rect 415822 42064 421972 42120
rect 415761 42062 421972 42064
rect 194317 42059 194383 42060
rect 415761 42059 415827 42062
rect 421966 42060 421972 42062
rect 422036 42060 422042 42124
rect 419901 41852 419967 41853
rect 419901 41848 419948 41852
rect 420012 41850 420018 41852
rect 419901 41792 419906 41848
rect 419901 41788 419948 41792
rect 420012 41790 420058 41850
rect 420012 41788 420018 41790
rect 419901 41787 419967 41788
rect 427770 41578 427830 42198
rect 446397 42256 461183 42258
rect 446397 42200 446402 42256
rect 446458 42200 461122 42256
rect 461178 42200 461183 42256
rect 446397 42198 461183 42200
rect 446397 42195 446463 42198
rect 461117 42195 461183 42198
rect 515397 42124 515463 42125
rect 520917 42124 520983 42125
rect 522021 42124 522087 42125
rect 526437 42124 526503 42125
rect 515397 42122 515444 42124
rect 515352 42120 515444 42122
rect 515352 42064 515402 42120
rect 515352 42062 515444 42064
rect 515397 42060 515444 42062
rect 515508 42060 515514 42124
rect 520917 42122 520964 42124
rect 520872 42120 520964 42122
rect 520872 42064 520922 42120
rect 520872 42062 520964 42064
rect 520917 42060 520964 42062
rect 521028 42060 521034 42124
rect 522021 42122 522068 42124
rect 521976 42120 522068 42122
rect 521976 42064 522026 42120
rect 521976 42062 522068 42064
rect 522021 42060 522068 42062
rect 522132 42060 522138 42124
rect 526437 42122 526484 42124
rect 526392 42120 526484 42122
rect 526392 42064 526442 42120
rect 526392 42062 526484 42064
rect 526437 42060 526484 42062
rect 526548 42060 526554 42124
rect 529565 42122 529631 42125
rect 529790 42122 529796 42124
rect 529565 42120 529796 42122
rect 529565 42064 529570 42120
rect 529626 42064 529796 42120
rect 529565 42062 529796 42064
rect 515397 42059 515463 42060
rect 520917 42059 520983 42060
rect 522021 42059 522087 42060
rect 526437 42059 526503 42060
rect 529565 42059 529631 42062
rect 529790 42060 529796 42062
rect 529860 42060 529866 42124
rect 441838 41788 441844 41852
rect 441908 41850 441914 41852
rect 460606 41850 460612 41852
rect 441908 41790 460612 41850
rect 441908 41788 441914 41790
rect 460606 41788 460612 41790
rect 460676 41788 460682 41852
rect 446397 41578 446463 41581
rect 427770 41576 446463 41578
rect 427770 41520 446402 41576
rect 446458 41520 446463 41576
rect 427770 41518 446463 41520
rect 446397 41515 446463 41518
rect 141693 40492 141759 40493
rect 141693 40488 141740 40492
rect 141804 40490 141810 40492
rect 141693 40432 141698 40488
rect 141693 40428 141740 40432
rect 141804 40430 141850 40490
rect 141804 40428 141810 40430
rect 141693 40427 141759 40428
<< via3 >>
rect 246620 997596 246684 997660
rect 86540 997188 86604 997252
rect 192524 997188 192588 997252
rect 89668 996916 89732 996980
rect 188844 996508 188908 996572
rect 86540 995752 86604 995756
rect 86540 995696 86554 995752
rect 86554 995696 86604 995752
rect 86540 995692 86604 995696
rect 132356 995964 132420 996028
rect 89668 995752 89732 995756
rect 89668 995696 89682 995752
rect 89682 995696 89732 995752
rect 89668 995692 89732 995696
rect 132540 995692 132604 995756
rect 132356 995344 132420 995348
rect 132356 995288 132406 995344
rect 132406 995288 132420 995344
rect 132356 995284 132420 995288
rect 142292 995828 142356 995892
rect 195284 996100 195348 996164
rect 192524 995786 192588 995790
rect 192524 995730 192538 995786
rect 192538 995730 192588 995786
rect 192524 995726 192588 995730
rect 295196 997188 295260 997252
rect 523908 997656 523972 997660
rect 523908 997600 523922 997656
rect 523922 997600 523972 997656
rect 523908 997596 523972 997600
rect 387748 997188 387812 997252
rect 511948 997188 512012 997252
rect 533476 997188 533540 997252
rect 246620 996916 246684 996980
rect 290780 996916 290844 996980
rect 629892 996916 629956 996980
rect 243860 996372 243924 996436
rect 245148 995964 245212 996028
rect 243860 995752 243924 995756
rect 243860 995696 243874 995752
rect 243874 995696 243924 995752
rect 243860 995692 243924 995696
rect 245148 995420 245212 995484
rect 195284 995284 195348 995348
rect 391980 996644 392044 996708
rect 480484 996644 480548 996708
rect 630260 996644 630324 996708
rect 294828 996372 294892 996436
rect 291884 996100 291948 996164
rect 291884 995556 291948 995620
rect 391980 996100 392044 996164
rect 476988 996372 477052 996436
rect 629156 996372 629220 996436
rect 484348 995828 484412 995892
rect 290780 994800 290844 994804
rect 290780 994744 290794 994800
rect 290794 994744 290844 994800
rect 290780 994740 290844 994744
rect 294828 994800 294892 994804
rect 294828 994744 294842 994800
rect 294842 994744 294892 994800
rect 294828 994740 294892 994744
rect 295196 994800 295260 994804
rect 295196 994744 295246 994800
rect 295246 994744 295260 994800
rect 295196 994740 295260 994744
rect 387748 994800 387812 994804
rect 476988 995072 477052 995076
rect 476988 995016 477038 995072
rect 477038 995016 477052 995072
rect 476988 995012 477052 995016
rect 480484 995012 480548 995076
rect 484348 995012 484412 995076
rect 531452 995692 531516 995756
rect 536604 995752 536668 995756
rect 536604 995696 536618 995752
rect 536618 995696 536668 995752
rect 536604 995692 536668 995696
rect 533476 995616 533540 995620
rect 533476 995560 533526 995616
rect 533526 995560 533540 995616
rect 533476 995556 533540 995560
rect 387748 994744 387798 994800
rect 387798 994744 387812 994800
rect 387748 994740 387812 994744
rect 522804 995012 522868 995076
rect 524460 995012 524524 995076
rect 629156 995752 629220 995756
rect 629156 995696 629206 995752
rect 629206 995696 629220 995752
rect 629156 995692 629220 995696
rect 629892 995752 629956 995756
rect 629892 995696 629906 995752
rect 629906 995696 629956 995752
rect 629892 995692 629956 995696
rect 630260 995786 630324 995790
rect 630260 995730 630310 995786
rect 630310 995730 630324 995786
rect 630260 995726 630324 995730
rect 569908 994876 569972 994940
rect 188844 994528 188908 994532
rect 188844 994472 188858 994528
rect 188858 994472 188908 994528
rect 188844 994468 188908 994472
rect 524460 994468 524524 994532
rect 132540 993924 132604 993988
rect 142292 992836 142356 992900
rect 41460 967132 41524 967196
rect 676076 965092 676140 965156
rect 676628 963596 676692 963660
rect 675340 963384 675404 963388
rect 675340 963328 675390 963384
rect 675390 963328 675404 963384
rect 675340 963324 675404 963328
rect 41828 962160 41892 962164
rect 41828 962104 41842 962160
rect 41842 962104 41892 962160
rect 41828 962100 41892 962104
rect 41276 959788 41340 959852
rect 675156 959304 675220 959308
rect 675156 959248 675206 959304
rect 675206 959248 675220 959304
rect 675156 959244 675220 959248
rect 40540 959108 40604 959172
rect 41828 957808 41892 957812
rect 41828 957752 41842 957808
rect 41842 957752 41892 957808
rect 41828 957748 41892 957752
rect 676996 957748 677060 957812
rect 676812 956388 676876 956452
rect 40724 955436 40788 955500
rect 675340 954484 675404 954548
rect 41828 952852 41892 952916
rect 41460 952444 41524 952508
rect 41644 952172 41708 952236
rect 41276 951628 41340 951692
rect 676628 951492 676692 951556
rect 675156 951144 675220 951148
rect 675156 951088 675206 951144
rect 675206 951088 675220 951144
rect 675156 951084 675220 951088
rect 676076 950676 676140 950740
rect 39804 943800 39868 943804
rect 39804 943744 39818 943800
rect 39818 943744 39868 943800
rect 39804 943740 39868 943744
rect 40724 943740 40788 943804
rect 42012 943740 42076 943804
rect 41782 939388 41846 939452
rect 41828 936668 41892 936732
rect 676812 931908 676876 931972
rect 676996 931500 677060 931564
rect 42012 911916 42076 911980
rect 42196 911644 42260 911708
rect 42012 885396 42076 885460
rect 42196 885124 42260 885188
rect 676076 875876 676140 875940
rect 675340 874032 675404 874036
rect 675340 873976 675390 874032
rect 675390 873976 675404 874032
rect 675340 873972 675404 873976
rect 673868 873156 673932 873220
rect 676996 870844 677060 870908
rect 675340 863152 675404 863156
rect 675340 863096 675354 863152
rect 675354 863096 675404 863152
rect 675340 863092 675404 863096
rect 39988 814234 40052 814298
rect 41828 813180 41892 813244
rect 41828 809100 41892 809164
rect 40908 805428 40972 805492
rect 41828 805428 41892 805492
rect 40540 805216 40604 805220
rect 40540 805160 40590 805216
rect 40590 805160 40604 805216
rect 40540 805156 40604 805160
rect 40724 805080 40788 805084
rect 40724 805024 40774 805080
rect 40774 805024 40788 805080
rect 40724 805020 40788 805024
rect 41644 804748 41708 804812
rect 42012 804476 42076 804540
rect 42196 798960 42260 798964
rect 42196 798904 42246 798960
rect 42246 798904 42260 798960
rect 42196 798900 42260 798904
rect 42196 797872 42260 797876
rect 42196 797816 42210 797872
rect 42210 797816 42260 797872
rect 42196 797812 42260 797816
rect 40724 794956 40788 795020
rect 40908 794140 40972 794204
rect 40540 792508 40604 792572
rect 41644 788972 41708 789036
rect 41828 788624 41892 788628
rect 41828 788568 41842 788624
rect 41842 788568 41892 788624
rect 41828 788564 41892 788568
rect 41460 786796 41524 786860
rect 675708 777004 675772 777068
rect 675708 775704 675772 775708
rect 675708 775648 675722 775704
rect 675722 775648 675772 775704
rect 675708 775644 675772 775648
rect 676812 774828 676876 774892
rect 676076 772652 676140 772716
rect 673868 770884 673932 770948
rect 41460 769796 41524 769860
rect 675892 766532 675956 766596
rect 676076 766592 676140 766596
rect 676076 766536 676126 766592
rect 676126 766536 676140 766592
rect 676076 766532 676140 766536
rect 40908 765716 40972 765780
rect 40540 765308 40604 765372
rect 40724 764900 40788 764964
rect 41644 764492 41708 764556
rect 676996 761968 677060 761972
rect 676996 761912 677046 761968
rect 677046 761912 677060 761968
rect 676996 761908 677060 761912
rect 676812 761832 676876 761836
rect 676812 761776 676826 761832
rect 676826 761776 676876 761832
rect 676812 761772 676876 761776
rect 42380 758644 42444 758708
rect 41828 757692 41892 757756
rect 40356 757344 40420 757348
rect 40356 757288 40370 757344
rect 40370 757288 40420 757344
rect 40356 757284 40420 757288
rect 40908 754836 40972 754900
rect 42012 754836 42076 754900
rect 42380 754896 42444 754900
rect 42380 754840 42394 754896
rect 42394 754840 42444 754896
rect 42380 754836 42444 754840
rect 40356 754564 40420 754628
rect 42012 751088 42076 751092
rect 42012 751032 42026 751088
rect 42026 751032 42076 751088
rect 42012 751028 42076 751032
rect 40724 750348 40788 750412
rect 40540 747356 40604 747420
rect 41828 745316 41892 745380
rect 41644 744364 41708 744428
rect 41460 743684 41524 743748
rect 674420 742460 674484 742524
rect 674236 741508 674300 741572
rect 674604 739604 674668 739668
rect 672028 732864 672092 732868
rect 672028 732808 672042 732864
rect 672042 732808 672092 732864
rect 672028 732804 672092 732808
rect 673316 732864 673380 732868
rect 673316 732808 673366 732864
rect 673366 732808 673380 732864
rect 673316 732804 673380 732808
rect 675892 729948 675956 730012
rect 676812 729948 676876 730012
rect 673316 728512 673380 728516
rect 673316 728456 673366 728512
rect 673366 728456 673380 728512
rect 673316 728452 673380 728456
rect 672028 728180 672092 728244
rect 41828 726820 41892 726884
rect 676076 725732 676140 725796
rect 40724 721708 40788 721772
rect 41644 721708 41708 721772
rect 40540 718524 40604 718588
rect 42564 718252 42628 718316
rect 41828 714716 41892 714780
rect 42012 714776 42076 714780
rect 42012 714720 42062 714776
rect 42062 714720 42076 714776
rect 42012 714716 42076 714720
rect 42380 714172 42444 714236
rect 42012 713416 42076 713420
rect 42012 713360 42026 713416
rect 42026 713360 42076 713416
rect 42012 713356 42076 713360
rect 675892 711996 675956 712060
rect 42564 711588 42628 711652
rect 40540 709140 40604 709204
rect 40724 707372 40788 707436
rect 42380 706556 42444 706620
rect 41644 702068 41708 702132
rect 41460 701796 41524 701860
rect 41828 701524 41892 701588
rect 675340 696824 675404 696828
rect 675340 696768 675390 696824
rect 675390 696768 675404 696824
rect 675340 696764 675404 696768
rect 676996 694044 677060 694108
rect 675340 686428 675404 686492
rect 41828 683572 41892 683636
rect 674420 682620 674484 682684
rect 674236 682348 674300 682412
rect 41828 681048 41892 681052
rect 41828 680992 41842 681048
rect 41842 680992 41892 681048
rect 41828 680988 41892 680992
rect 40540 678928 40604 678992
rect 40724 678928 40788 678992
rect 42380 674188 42444 674252
rect 40356 671196 40420 671260
rect 42012 671196 42076 671260
rect 41828 670924 41892 670988
rect 40356 670244 40420 670308
rect 42196 669292 42260 669356
rect 42380 668476 42444 668540
rect 42196 667932 42260 667996
rect 42012 667252 42076 667316
rect 40724 665348 40788 665412
rect 40540 664124 40604 664188
rect 674788 663988 674852 664052
rect 41460 660724 41524 660788
rect 41644 658548 41708 658612
rect 41828 658276 41892 658340
rect 44220 653108 44284 653172
rect 675340 652836 675404 652900
rect 674788 650116 674852 650180
rect 675524 648076 675588 648140
rect 674788 647592 674852 647596
rect 674788 647536 674838 647592
rect 674838 647536 674852 647592
rect 674788 647532 674852 647536
rect 675524 647396 675588 647460
rect 675156 645764 675220 645828
rect 674052 645084 674116 645148
rect 674972 644268 675036 644332
rect 676812 644268 676876 644332
rect 675524 643996 675588 644060
rect 671476 643452 671540 643516
rect 674972 640792 675036 640796
rect 674972 640736 674986 640792
rect 674986 640736 675036 640792
rect 674972 640732 675036 640736
rect 41644 640596 41708 640660
rect 675524 640188 675588 640252
rect 676628 640188 676692 640252
rect 41460 639372 41524 639436
rect 675156 638012 675220 638076
rect 676628 637876 676692 637940
rect 675340 637604 675404 637668
rect 41828 637332 41892 637396
rect 40724 634884 40788 634948
rect 40540 634476 40604 634540
rect 675340 631348 675404 631412
rect 676076 631348 676140 631412
rect 41828 627676 41892 627740
rect 40724 623732 40788 623796
rect 41828 620256 41892 620260
rect 41828 620200 41842 620256
rect 41842 620200 41892 620256
rect 41828 620196 41892 620200
rect 40540 619924 40604 619988
rect 676996 619108 677060 619172
rect 673868 616116 673932 616180
rect 42012 615904 42076 615908
rect 42012 615848 42062 615904
rect 42062 615848 42076 615904
rect 42012 615844 42076 615848
rect 41460 615436 41524 615500
rect 41828 614136 41892 614140
rect 41828 614080 41878 614136
rect 41878 614080 41892 614136
rect 41828 614076 41892 614080
rect 44220 614136 44284 614140
rect 44220 614080 44234 614136
rect 44234 614080 44284 614136
rect 44220 614076 44284 614080
rect 675524 608288 675588 608292
rect 675524 608232 675538 608288
rect 675538 608232 675588 608288
rect 675524 608228 675588 608232
rect 674420 602788 674484 602852
rect 41828 596048 41892 596052
rect 41828 595992 41842 596048
rect 41842 595992 41892 596048
rect 41828 595988 41892 595992
rect 674788 595580 674852 595644
rect 673684 595308 673748 595372
rect 42012 594900 42076 594964
rect 676076 593404 676140 593468
rect 676996 593404 677060 593468
rect 40724 592350 40788 592414
rect 675340 592316 675404 592380
rect 675524 592104 675588 592108
rect 675524 592048 675574 592104
rect 675574 592048 675588 592104
rect 675524 592044 675588 592048
rect 673684 591636 673748 591700
rect 43852 591500 43916 591564
rect 674788 591364 674852 591428
rect 40908 589656 40972 589660
rect 40908 589600 40958 589656
rect 40958 589600 40972 589656
rect 40908 589596 40972 589600
rect 40540 589324 40604 589388
rect 41460 587148 41524 587212
rect 42012 587148 42076 587212
rect 676076 586196 676140 586260
rect 42380 586060 42444 586124
rect 41828 585108 41892 585172
rect 42196 584836 42260 584900
rect 41092 584564 41156 584628
rect 42380 581904 42444 581908
rect 42380 581848 42394 581904
rect 42394 581848 42444 581904
rect 42380 581844 42444 581848
rect 42196 581496 42260 581500
rect 42196 581440 42246 581496
rect 42246 581440 42260 581496
rect 42196 581436 42260 581440
rect 41092 580212 41156 580276
rect 40908 578172 40972 578236
rect 40724 577492 40788 577556
rect 40540 576812 40604 576876
rect 42196 576132 42260 576196
rect 676996 575996 677060 576060
rect 676812 572732 676876 572796
rect 42196 572596 42260 572660
rect 41828 572188 41892 572252
rect 41460 571916 41524 571980
rect 671476 571236 671540 571300
rect 41644 570964 41708 571028
rect 675340 563136 675404 563140
rect 675340 563080 675390 563136
rect 675390 563080 675404 563136
rect 675340 563076 675404 563080
rect 675524 561232 675588 561236
rect 675524 561176 675538 561232
rect 675538 561176 675588 561232
rect 675524 561172 675588 561176
rect 676812 554644 676876 554708
rect 41828 553208 41892 553212
rect 41828 553152 41842 553208
rect 41842 553152 41892 553208
rect 41828 553148 41892 553152
rect 41828 551984 41892 551988
rect 41828 551928 41878 551984
rect 41878 551928 41892 551984
rect 41828 551924 41892 551928
rect 677180 550700 677244 550764
rect 42012 549884 42076 549948
rect 675156 549612 675220 549676
rect 675156 547904 675220 547908
rect 675156 547848 675170 547904
rect 675170 547848 675220 547904
rect 675156 547844 675220 547848
rect 675524 547572 675588 547636
rect 676076 546484 676140 546548
rect 41644 546348 41708 546412
rect 40540 545668 40604 545732
rect 40724 545396 40788 545460
rect 42012 545396 42076 545460
rect 674788 543824 674852 543828
rect 674788 543768 674838 543824
rect 674838 543768 674852 543824
rect 674788 543764 674852 543768
rect 40724 538596 40788 538660
rect 40540 538188 40604 538252
rect 41460 530572 41524 530636
rect 41828 529408 41892 529412
rect 41828 529352 41878 529408
rect 41878 529352 41892 529408
rect 41828 529348 41892 529352
rect 41644 529076 41708 529140
rect 674420 527036 674484 527100
rect 676812 503644 676876 503708
rect 677364 492416 677428 492420
rect 677364 492360 677378 492416
rect 677378 492360 677428 492416
rect 677364 492356 677428 492360
rect 675892 490452 675956 490516
rect 676996 485788 677060 485792
rect 676996 485732 677010 485788
rect 677010 485732 677060 485788
rect 676996 485728 677060 485732
rect 673684 475356 673748 475420
rect 674052 475356 674116 475420
rect 673684 464748 673748 464812
rect 673868 455092 673932 455156
rect 41828 425172 41892 425236
rect 42012 424764 42076 424828
rect 41460 418780 41524 418844
rect 40724 417828 40788 417892
rect 40540 417556 40604 417620
rect 40724 409396 40788 409460
rect 41828 406328 41892 406332
rect 41828 406272 41842 406328
rect 41842 406272 41892 406328
rect 41828 406268 41892 406272
rect 40540 403820 40604 403884
rect 676812 402868 676876 402932
rect 41828 401840 41892 401844
rect 41828 401784 41842 401840
rect 41842 401784 41892 401840
rect 41828 401780 41892 401784
rect 676996 401236 677060 401300
rect 41460 398788 41524 398852
rect 675892 398788 675956 398852
rect 676628 396748 676692 396812
rect 676260 395116 676324 395180
rect 676444 394708 676508 394772
rect 676076 393076 676140 393140
rect 675708 387636 675772 387700
rect 676628 384916 676692 384980
rect 41460 381788 41524 381852
rect 676444 380564 676508 380628
rect 675708 378720 675772 378724
rect 675708 378664 675758 378720
rect 675758 378664 675772 378720
rect 675708 378660 675772 378664
rect 40540 378524 40604 378588
rect 40724 378116 40788 378180
rect 674788 377980 674852 378044
rect 676260 377300 676324 377364
rect 41644 376892 41708 376956
rect 675892 376892 675956 376956
rect 41276 373220 41340 373284
rect 676076 372948 676140 373012
rect 674788 372540 674852 372604
rect 41828 371860 41892 371924
rect 41276 368460 41340 368524
rect 40724 363564 40788 363628
rect 40540 360028 40604 360092
rect 41828 359408 41892 359412
rect 41828 359352 41842 359408
rect 41842 359352 41892 359408
rect 41828 359348 41892 359352
rect 41460 358668 41524 358732
rect 41828 355736 41892 355740
rect 41828 355680 41878 355736
rect 41878 355680 41892 355736
rect 41828 355676 41892 355680
rect 43852 354240 43916 354244
rect 43852 354184 43902 354240
rect 43902 354184 43916 354240
rect 43852 354180 43916 354184
rect 675340 354180 675404 354244
rect 44220 353772 44284 353836
rect 675708 352956 675772 353020
rect 675892 351732 675956 351796
rect 675892 350916 675956 350980
rect 675892 350100 675956 350164
rect 675892 349208 675956 349212
rect 675892 349152 675942 349208
rect 675942 349152 675956 349208
rect 675892 349148 675956 349152
rect 44404 342892 44468 342956
rect 44220 342620 44284 342684
rect 44404 342076 44468 342140
rect 44588 341260 44652 341324
rect 43668 340444 43732 340508
rect 676628 340308 676692 340372
rect 675340 339008 675404 339012
rect 675340 338952 675390 339008
rect 675390 338952 675404 339008
rect 675340 338948 675404 338952
rect 40724 337724 40788 337788
rect 675524 337784 675588 337788
rect 675524 337728 675574 337784
rect 675574 337728 675588 337784
rect 675524 337724 675588 337728
rect 42932 337588 42996 337652
rect 43116 336772 43180 336836
rect 676444 336636 676508 336700
rect 43300 336092 43364 336156
rect 40540 335684 40604 335748
rect 42196 335004 42260 335068
rect 43300 334656 43364 334660
rect 43300 334600 43314 334656
rect 43314 334600 43364 334656
rect 43300 334596 43364 334600
rect 41828 334460 41892 334524
rect 42196 334324 42260 334388
rect 40908 333644 40972 333708
rect 676260 332148 676324 332212
rect 41644 329020 41708 329084
rect 41460 328340 41524 328404
rect 676076 328340 676140 328404
rect 40724 326708 40788 326772
rect 40908 325348 40972 325412
rect 41828 324728 41892 324732
rect 41828 324672 41878 324728
rect 41878 324672 41892 324728
rect 41828 324668 41892 324672
rect 40540 320996 40604 321060
rect 43116 316372 43180 316436
rect 41828 315616 41892 315620
rect 41828 315560 41842 315616
rect 41842 315560 41892 315616
rect 41828 315556 41892 315560
rect 42932 312700 42996 312764
rect 41460 312564 41524 312628
rect 44220 311748 44284 311812
rect 44404 311476 44468 311540
rect 44588 311264 44652 311268
rect 44588 311208 44602 311264
rect 44602 311208 44652 311264
rect 44588 311204 44652 311208
rect 675708 308756 675772 308820
rect 675156 307940 675220 308004
rect 675892 306716 675956 306780
rect 675892 302636 675956 302700
rect 675156 301744 675220 301748
rect 675156 301688 675170 301744
rect 675170 301688 675220 301744
rect 675156 301684 675220 301688
rect 676628 301608 676692 301612
rect 676628 301552 676642 301608
rect 676642 301552 676692 301608
rect 676628 301548 676692 301552
rect 676444 301472 676508 301476
rect 676444 301416 676458 301472
rect 676458 301416 676508 301472
rect 676444 301412 676508 301416
rect 43668 297604 43732 297668
rect 675708 297332 675772 297396
rect 42012 296380 42076 296444
rect 41828 295564 41892 295628
rect 676260 295156 676324 295220
rect 41828 292768 41892 292772
rect 41828 292712 41842 292768
rect 41842 292712 41892 292768
rect 41828 292708 41892 292712
rect 40540 292528 40604 292592
rect 40724 292528 40788 292592
rect 41828 292300 41892 292364
rect 676444 291484 676508 291548
rect 676628 286996 676692 287060
rect 676076 283596 676140 283660
rect 675892 282780 675956 282844
rect 675708 281616 675772 281620
rect 675708 281560 675722 281616
rect 675722 281560 675772 281616
rect 675708 281556 675772 281560
rect 42012 281480 42076 281484
rect 42012 281424 42026 281480
rect 42026 281424 42076 281480
rect 42012 281420 42076 281424
rect 40724 277884 40788 277948
rect 40908 277612 40972 277676
rect 40540 274212 40604 274276
rect 41460 270404 41524 270468
rect 41828 269104 41892 269108
rect 41828 269048 41842 269104
rect 41842 269048 41892 269104
rect 41828 269044 41892 269048
rect 674972 263604 675036 263668
rect 676076 262380 676140 262444
rect 676996 261564 677060 261628
rect 676812 259932 676876 259996
rect 40540 251364 40604 251428
rect 676996 250276 677060 250340
rect 40724 249732 40788 249796
rect 674788 249596 674852 249660
rect 676076 249596 676140 249660
rect 676812 245244 676876 245308
rect 675156 244972 675220 245036
rect 675340 244700 675404 244764
rect 675156 240272 675220 240276
rect 675156 240216 675206 240272
rect 675206 240216 675220 240272
rect 675156 240212 675220 240216
rect 40540 240076 40604 240140
rect 42012 237356 42076 237420
rect 674236 237084 674300 237148
rect 675340 236872 675404 236876
rect 675340 236816 675390 236872
rect 675390 236816 675404 236872
rect 675340 236812 675404 236816
rect 40724 235860 40788 235924
rect 672396 231508 672460 231572
rect 672396 230556 672460 230620
rect 674420 230148 674484 230212
rect 667980 229468 668044 229532
rect 673132 228788 673196 228852
rect 672948 228576 673012 228580
rect 672948 228520 672962 228576
rect 672962 228520 673012 228576
rect 672948 228516 673012 228520
rect 675156 228516 675220 228580
rect 42012 227352 42076 227356
rect 42012 227296 42026 227352
rect 42026 227296 42076 227352
rect 42012 227292 42076 227296
rect 672396 227080 672460 227084
rect 672396 227024 672446 227080
rect 672446 227024 672460 227080
rect 672396 227020 672460 227024
rect 672764 227020 672828 227084
rect 675340 225932 675404 225996
rect 672028 225660 672092 225724
rect 673500 224980 673564 225044
rect 674420 224980 674484 225044
rect 673132 224572 673196 224636
rect 672764 224300 672828 224364
rect 672028 223000 672092 223004
rect 672028 222944 672078 223000
rect 672078 222944 672092 223000
rect 672028 222940 672092 222944
rect 572484 222532 572548 222596
rect 561260 222260 561324 222324
rect 562916 221988 562980 222052
rect 563100 221988 563164 222052
rect 563652 221988 563716 222052
rect 572116 221988 572180 222052
rect 545068 220552 545132 220556
rect 545068 220496 545082 220552
rect 545082 220496 545132 220552
rect 545068 220492 545132 220496
rect 511028 220008 511092 220012
rect 511028 219952 511042 220008
rect 511042 219952 511092 220008
rect 511028 219948 511092 219952
rect 529980 220008 530044 220012
rect 529980 219952 530030 220008
rect 530030 219952 530044 220008
rect 519860 219736 519924 219740
rect 519860 219680 519874 219736
rect 519874 219680 519924 219736
rect 519860 219676 519924 219680
rect 522620 219736 522684 219740
rect 529980 219948 530044 219952
rect 530348 220008 530412 220012
rect 530348 219952 530362 220008
rect 530362 219952 530412 220008
rect 530348 219948 530412 219952
rect 543780 220220 543844 220284
rect 553900 220492 553964 220556
rect 563284 220492 563348 220556
rect 556476 220220 556540 220284
rect 563836 220220 563900 220284
rect 573220 220220 573284 220284
rect 670740 220084 670804 220148
rect 674604 220356 674668 220420
rect 674788 220084 674852 220148
rect 522620 219680 522634 219736
rect 522634 219680 522684 219736
rect 522620 219676 522684 219680
rect 514708 219192 514772 219196
rect 514708 219136 514758 219192
rect 514758 219136 514772 219192
rect 514708 219132 514772 219136
rect 553164 219132 553228 219196
rect 553532 219132 553596 219196
rect 567884 219132 567948 219196
rect 674604 219132 674668 219196
rect 514340 218316 514404 218380
rect 543780 218316 543844 218380
rect 553900 218316 553964 218380
rect 554084 218316 554148 218380
rect 567884 218316 567948 218380
rect 572116 218316 572180 218380
rect 674972 218588 675036 218652
rect 675892 218180 675956 218244
rect 563836 217772 563900 217836
rect 564020 217772 564084 217836
rect 572116 217772 572180 217836
rect 500724 217500 500788 217564
rect 504772 217500 504836 217564
rect 672212 217500 672276 217564
rect 675524 217364 675588 217428
rect 493548 217288 493612 217292
rect 493548 217232 493598 217288
rect 493598 217232 493612 217288
rect 493548 217228 493612 217232
rect 541756 217228 541820 217292
rect 544148 217228 544212 217292
rect 675156 217228 675220 217292
rect 500724 216956 500788 217020
rect 582604 216956 582668 217020
rect 591620 216956 591684 217020
rect 592172 216956 592236 217020
rect 675708 216956 675772 217020
rect 511028 216412 511092 216476
rect 519308 216412 519372 216476
rect 519860 216412 519924 216476
rect 566596 216412 566660 216476
rect 566780 216412 566844 216476
rect 572116 216412 572180 216476
rect 572484 216412 572548 216476
rect 577636 216412 577700 216476
rect 504772 216140 504836 216204
rect 582420 216140 582484 216204
rect 519308 215868 519372 215932
rect 529244 215868 529308 215932
rect 530348 215868 530412 215932
rect 546908 215868 546972 215932
rect 548564 215868 548628 215932
rect 577084 215868 577148 215932
rect 675340 215868 675404 215932
rect 522620 215324 522684 215388
rect 556476 215596 556540 215660
rect 529244 215324 529308 215388
rect 536972 215324 537036 215388
rect 538628 215324 538692 215388
rect 558316 215596 558380 215660
rect 666324 215596 666388 215660
rect 566780 215324 566844 215388
rect 529980 215052 530044 215116
rect 674788 215324 674852 215388
rect 568252 215052 568316 215116
rect 676260 215086 676324 215150
rect 673132 214780 673196 214844
rect 675892 214508 675956 214572
rect 575612 213616 575676 213620
rect 575612 213560 575662 213616
rect 575662 213560 575676 213616
rect 575612 213556 575676 213560
rect 674052 212060 674116 212124
rect 675892 211380 675956 211444
rect 676444 211380 676508 211444
rect 669452 211108 669516 211172
rect 674972 210428 675036 210492
rect 675892 210428 675956 210492
rect 41460 209748 41524 209812
rect 40540 208116 40604 208180
rect 42380 207708 42444 207772
rect 40908 207300 40972 207364
rect 40724 206892 40788 206956
rect 676628 205532 676692 205596
rect 673316 201648 673380 201652
rect 673316 201592 673330 201648
rect 673330 201592 673380 201648
rect 673316 201588 673380 201592
rect 676444 200636 676508 200700
rect 675524 198248 675588 198252
rect 675524 198192 675574 198248
rect 675574 198192 675588 198248
rect 675524 198188 675588 198192
rect 666508 197916 666572 197980
rect 41828 197780 41892 197844
rect 40540 197100 40604 197164
rect 676260 197100 676324 197164
rect 41828 195800 41892 195804
rect 41828 195744 41878 195800
rect 41878 195744 41892 195800
rect 41828 195740 41892 195744
rect 41460 195196 41524 195260
rect 40908 194924 40972 194988
rect 40724 194516 40788 194580
rect 41644 194516 41708 194580
rect 42196 193216 42260 193220
rect 42196 193160 42246 193216
rect 42246 193160 42260 193216
rect 42196 193156 42260 193160
rect 675892 193156 675956 193220
rect 676076 191524 676140 191588
rect 41828 187232 41892 187236
rect 41828 187176 41842 187232
rect 41842 187176 41892 187232
rect 41828 187172 41892 187176
rect 42380 186280 42444 186284
rect 42380 186224 42394 186280
rect 42394 186224 42444 186280
rect 42380 186220 42444 186224
rect 42196 186008 42260 186012
rect 42196 185952 42210 186008
rect 42210 185952 42260 186008
rect 42196 185948 42260 185952
rect 672948 183500 673012 183564
rect 673132 182004 673196 182068
rect 675892 173980 675956 174044
rect 675708 173572 675772 173636
rect 675892 172348 675956 172412
rect 675892 171940 675956 172004
rect 675524 167452 675588 167516
rect 676628 166424 676692 166428
rect 676628 166368 676642 166424
rect 676642 166368 676692 166424
rect 676628 166364 676692 166368
rect 675340 161876 675404 161940
rect 676444 159292 676508 159356
rect 675340 157040 675404 157044
rect 675340 156984 675390 157040
rect 675390 156984 675404 157040
rect 675340 156980 675404 156984
rect 676628 156300 676692 156364
rect 674236 154940 674300 155004
rect 676260 153036 676324 153100
rect 673316 149092 673380 149156
rect 675892 148412 675956 148476
rect 675708 147656 675772 147660
rect 675708 147600 675722 147656
rect 675722 147600 675772 147656
rect 675708 147596 675772 147600
rect 676076 145964 676140 146028
rect 669268 143652 669332 143716
rect 670740 133724 670804 133788
rect 667980 130596 668044 130660
rect 673500 128828 673564 128892
rect 676628 128556 676692 128620
rect 674052 128284 674116 128348
rect 676076 128148 676140 128212
rect 675892 127196 675956 127260
rect 676260 126924 676324 126988
rect 676444 124476 676508 124540
rect 675708 122300 675772 122364
rect 676628 113052 676692 113116
rect 675892 108020 675956 108084
rect 676444 106116 676508 106180
rect 676076 103124 676140 103188
rect 675708 102640 675772 102644
rect 675708 102584 675722 102640
rect 675722 102584 675772 102640
rect 675708 102580 675772 102584
rect 676260 101356 676324 101420
rect 637252 96868 637316 96932
rect 633940 96052 634004 96116
rect 633940 78568 634004 78572
rect 633940 78512 633954 78568
rect 633954 78512 634004 78568
rect 633940 78508 634004 78512
rect 637068 77828 637132 77892
rect 462636 54436 462700 54500
rect 462636 53680 462700 53684
rect 462636 53624 462650 53680
rect 462650 53624 462700 53680
rect 462636 53620 462700 53624
rect 194364 50220 194428 50284
rect 529796 50220 529860 50284
rect 518756 48860 518820 48924
rect 526484 48044 526548 48108
rect 520964 47772 521028 47836
rect 515444 47500 515508 47564
rect 522068 47228 522132 47292
rect 141740 43964 141804 44028
rect 461348 44372 461412 44436
rect 462268 44372 462332 44436
rect 518756 42800 518820 42804
rect 518756 42744 518806 42800
rect 518806 42744 518820 42800
rect 518756 42740 518820 42744
rect 194364 42120 194428 42124
rect 194364 42064 194378 42120
rect 194378 42064 194428 42120
rect 194364 42060 194428 42064
rect 421972 42060 422036 42124
rect 419948 41848 420012 41852
rect 419948 41792 419962 41848
rect 419962 41792 420012 41848
rect 419948 41788 420012 41792
rect 515444 42120 515508 42124
rect 515444 42064 515458 42120
rect 515458 42064 515508 42120
rect 515444 42060 515508 42064
rect 520964 42120 521028 42124
rect 520964 42064 520978 42120
rect 520978 42064 521028 42120
rect 520964 42060 521028 42064
rect 522068 42120 522132 42124
rect 522068 42064 522082 42120
rect 522082 42064 522132 42120
rect 522068 42060 522132 42064
rect 526484 42120 526548 42124
rect 526484 42064 526498 42120
rect 526498 42064 526548 42120
rect 526484 42060 526548 42064
rect 529796 42060 529860 42124
rect 441844 41788 441908 41852
rect 460612 41788 460676 41852
rect 141740 40488 141804 40492
rect 141740 40432 141754 40488
rect 141754 40432 141804 40488
rect 141740 40428 141804 40432
<< metal4 >>
rect 246619 997660 246685 997661
rect 246619 997596 246620 997660
rect 246684 997596 246685 997660
rect 246619 997595 246685 997596
rect 523907 997660 523973 997661
rect 523907 997596 523908 997660
rect 523972 997596 523973 997660
rect 523907 997595 523973 997596
rect 86539 997252 86605 997253
rect 86539 997188 86540 997252
rect 86604 997188 86605 997252
rect 86539 997187 86605 997188
rect 192523 997252 192589 997253
rect 192523 997188 192524 997252
rect 192588 997188 192589 997252
rect 192523 997187 192589 997188
rect 86542 995757 86602 997187
rect 89667 996980 89733 996981
rect 89667 996916 89668 996980
rect 89732 996916 89733 996980
rect 89667 996915 89733 996916
rect 89670 995757 89730 996915
rect 188843 996572 188909 996573
rect 188843 996508 188844 996572
rect 188908 996508 188909 996572
rect 188843 996507 188909 996508
rect 132355 996028 132421 996029
rect 132355 995964 132356 996028
rect 132420 995964 132421 996028
rect 132355 995963 132421 995964
rect 86539 995756 86605 995757
rect 86539 995692 86540 995756
rect 86604 995692 86605 995756
rect 86539 995691 86605 995692
rect 89667 995756 89733 995757
rect 89667 995692 89668 995756
rect 89732 995692 89733 995756
rect 89667 995691 89733 995692
rect 132358 995349 132418 995963
rect 142291 995892 142357 995893
rect 142291 995828 142292 995892
rect 142356 995828 142357 995892
rect 142291 995827 142357 995828
rect 132539 995756 132605 995757
rect 132539 995692 132540 995756
rect 132604 995692 132605 995756
rect 132539 995691 132605 995692
rect 132355 995348 132421 995349
rect 132355 995284 132356 995348
rect 132420 995284 132421 995348
rect 132355 995283 132421 995284
rect 132542 993989 132602 995691
rect 132539 993988 132605 993989
rect 132539 993924 132540 993988
rect 132604 993924 132605 993988
rect 132539 993923 132605 993924
rect 142294 992901 142354 995827
rect 188846 994533 188906 996507
rect 192526 995791 192586 997187
rect 246622 996981 246682 997595
rect 523910 997338 523970 997595
rect 295195 997252 295261 997253
rect 295195 997188 295196 997252
rect 295260 997188 295261 997252
rect 295195 997187 295261 997188
rect 387747 997252 387813 997253
rect 387747 997188 387748 997252
rect 387812 997188 387813 997252
rect 387747 997187 387813 997188
rect 246619 996980 246685 996981
rect 246619 996916 246620 996980
rect 246684 996916 246685 996980
rect 246619 996915 246685 996916
rect 290779 996980 290845 996981
rect 290779 996916 290780 996980
rect 290844 996916 290845 996980
rect 290779 996915 290845 996916
rect 243859 996436 243925 996437
rect 243859 996372 243860 996436
rect 243924 996372 243925 996436
rect 243859 996371 243925 996372
rect 195283 996164 195349 996165
rect 195283 996100 195284 996164
rect 195348 996100 195349 996164
rect 195283 996099 195349 996100
rect 192523 995790 192589 995791
rect 192523 995726 192524 995790
rect 192588 995726 192589 995790
rect 192523 995725 192589 995726
rect 195286 995349 195346 996099
rect 243862 995757 243922 996371
rect 245147 996028 245213 996029
rect 245147 995964 245148 996028
rect 245212 995964 245213 996028
rect 245147 995963 245213 995964
rect 243859 995756 243925 995757
rect 243859 995692 243860 995756
rect 243924 995692 243925 995756
rect 243859 995691 243925 995692
rect 245150 995485 245210 995963
rect 245147 995484 245213 995485
rect 245147 995420 245148 995484
rect 245212 995420 245213 995484
rect 245147 995419 245213 995420
rect 195283 995348 195349 995349
rect 195283 995284 195284 995348
rect 195348 995284 195349 995348
rect 195283 995283 195349 995284
rect 290782 994805 290842 996915
rect 294827 996436 294893 996437
rect 294827 996372 294828 996436
rect 294892 996372 294893 996436
rect 294827 996371 294893 996372
rect 291883 996164 291949 996165
rect 291883 996100 291884 996164
rect 291948 996100 291949 996164
rect 291883 996099 291949 996100
rect 291886 995621 291946 996099
rect 291883 995620 291949 995621
rect 291883 995556 291884 995620
rect 291948 995556 291949 995620
rect 291883 995555 291949 995556
rect 294830 994805 294890 996371
rect 295198 994805 295258 997187
rect 387750 994805 387810 997187
rect 533475 997252 533541 997253
rect 533475 997188 533476 997252
rect 533540 997188 533541 997252
rect 533475 997187 533541 997188
rect 391979 996708 392045 996709
rect 391979 996644 391980 996708
rect 392044 996644 392045 996708
rect 391979 996643 392045 996644
rect 480483 996708 480549 996709
rect 480483 996644 480484 996708
rect 480548 996644 480549 996708
rect 480483 996643 480549 996644
rect 391982 996165 392042 996643
rect 476987 996436 477053 996437
rect 476987 996372 476988 996436
rect 477052 996372 477053 996436
rect 476987 996371 477053 996372
rect 391979 996164 392045 996165
rect 391979 996100 391980 996164
rect 392044 996100 392045 996164
rect 391979 996099 392045 996100
rect 476990 995077 477050 996371
rect 480486 995077 480546 996643
rect 484347 995892 484413 995893
rect 484347 995828 484348 995892
rect 484412 995828 484413 995892
rect 484347 995827 484413 995828
rect 484350 995077 484410 995827
rect 522806 995077 522866 997102
rect 531454 995757 531514 997102
rect 531451 995756 531517 995757
rect 531451 995692 531452 995756
rect 531516 995692 531517 995756
rect 531451 995691 531517 995692
rect 533478 995621 533538 997187
rect 536606 995757 536666 997102
rect 536603 995756 536669 995757
rect 536603 995692 536604 995756
rect 536668 995692 536669 995756
rect 536603 995691 536669 995692
rect 533475 995620 533541 995621
rect 533475 995556 533476 995620
rect 533540 995556 533541 995620
rect 533475 995555 533541 995556
rect 476987 995076 477053 995077
rect 476987 995012 476988 995076
rect 477052 995012 477053 995076
rect 476987 995011 477053 995012
rect 480483 995076 480549 995077
rect 480483 995012 480484 995076
rect 480548 995012 480549 995076
rect 480483 995011 480549 995012
rect 484347 995076 484413 995077
rect 484347 995012 484348 995076
rect 484412 995012 484413 995076
rect 484347 995011 484413 995012
rect 522803 995076 522869 995077
rect 522803 995012 522804 995076
rect 522868 995012 522869 995076
rect 522803 995011 522869 995012
rect 524459 995076 524525 995077
rect 524459 995012 524460 995076
rect 524524 995012 524525 995076
rect 524459 995011 524525 995012
rect 290779 994804 290845 994805
rect 290779 994740 290780 994804
rect 290844 994740 290845 994804
rect 290779 994739 290845 994740
rect 294827 994804 294893 994805
rect 294827 994740 294828 994804
rect 294892 994740 294893 994804
rect 294827 994739 294893 994740
rect 295195 994804 295261 994805
rect 295195 994740 295196 994804
rect 295260 994740 295261 994804
rect 295195 994739 295261 994740
rect 387747 994804 387813 994805
rect 387747 994740 387748 994804
rect 387812 994740 387813 994804
rect 387747 994739 387813 994740
rect 524462 994533 524522 995011
rect 569910 994941 569970 997102
rect 629891 996980 629957 996981
rect 629891 996916 629892 996980
rect 629956 996916 629957 996980
rect 629891 996915 629957 996916
rect 629155 996436 629221 996437
rect 629155 996372 629156 996436
rect 629220 996372 629221 996436
rect 629155 996371 629221 996372
rect 629158 995757 629218 996371
rect 629894 995757 629954 996915
rect 630259 996708 630325 996709
rect 630259 996644 630260 996708
rect 630324 996644 630325 996708
rect 630259 996643 630325 996644
rect 630262 995791 630322 996643
rect 630259 995790 630325 995791
rect 629155 995756 629221 995757
rect 629155 995692 629156 995756
rect 629220 995692 629221 995756
rect 629155 995691 629221 995692
rect 629891 995756 629957 995757
rect 629891 995692 629892 995756
rect 629956 995692 629957 995756
rect 630259 995726 630260 995790
rect 630324 995726 630325 995790
rect 630259 995725 630325 995726
rect 629891 995691 629957 995692
rect 569907 994940 569973 994941
rect 569907 994876 569908 994940
rect 569972 994876 569973 994940
rect 569907 994875 569973 994876
rect 188843 994532 188909 994533
rect 188843 994468 188844 994532
rect 188908 994468 188909 994532
rect 188843 994467 188909 994468
rect 524459 994532 524525 994533
rect 524459 994468 524460 994532
rect 524524 994468 524525 994532
rect 524459 994467 524525 994468
rect 142291 992900 142357 992901
rect 142291 992836 142292 992900
rect 142356 992836 142357 992900
rect 142291 992835 142357 992836
rect 41459 967196 41525 967197
rect 41459 967132 41460 967196
rect 41524 967132 41525 967196
rect 41459 967131 41525 967132
rect 41275 959852 41341 959853
rect 41275 959788 41276 959852
rect 41340 959788 41341 959852
rect 41275 959787 41341 959788
rect 40539 959172 40605 959173
rect 40539 959108 40540 959172
rect 40604 959108 40605 959172
rect 40539 959107 40605 959108
rect 40542 945330 40602 959107
rect 40723 955500 40789 955501
rect 40723 955436 40724 955500
rect 40788 955436 40789 955500
rect 40723 955435 40789 955436
rect 39806 945270 40602 945330
rect 39806 943805 39866 945270
rect 40726 943805 40786 955435
rect 41278 951693 41338 959787
rect 41462 952509 41522 967131
rect 676075 965156 676141 965157
rect 676075 965092 676076 965156
rect 676140 965092 676141 965156
rect 676075 965091 676141 965092
rect 675339 963388 675405 963389
rect 675339 963324 675340 963388
rect 675404 963324 675405 963388
rect 675339 963323 675405 963324
rect 41827 962164 41893 962165
rect 41827 962100 41828 962164
rect 41892 962100 41893 962164
rect 41827 962099 41893 962100
rect 41830 959130 41890 962099
rect 675155 959308 675221 959309
rect 675155 959244 675156 959308
rect 675220 959244 675221 959308
rect 675155 959243 675221 959244
rect 41646 959070 41890 959130
rect 41459 952508 41525 952509
rect 41459 952444 41460 952508
rect 41524 952444 41525 952508
rect 41459 952443 41525 952444
rect 41646 952237 41706 959070
rect 41827 957812 41893 957813
rect 41827 957748 41828 957812
rect 41892 957748 41893 957812
rect 41827 957747 41893 957748
rect 41830 952917 41890 957747
rect 41827 952916 41893 952917
rect 41827 952852 41828 952916
rect 41892 952852 41893 952916
rect 41827 952851 41893 952852
rect 41643 952236 41709 952237
rect 41643 952172 41644 952236
rect 41708 952172 41709 952236
rect 41643 952171 41709 952172
rect 41275 951692 41341 951693
rect 41275 951628 41276 951692
rect 41340 951628 41341 951692
rect 41275 951627 41341 951628
rect 675158 951149 675218 959243
rect 675342 954549 675402 963323
rect 675339 954548 675405 954549
rect 675339 954484 675340 954548
rect 675404 954484 675405 954548
rect 675339 954483 675405 954484
rect 675155 951148 675221 951149
rect 675155 951084 675156 951148
rect 675220 951084 675221 951148
rect 675155 951083 675221 951084
rect 676078 950741 676138 965091
rect 676627 963660 676693 963661
rect 676627 963596 676628 963660
rect 676692 963596 676693 963660
rect 676627 963595 676693 963596
rect 676630 951557 676690 963595
rect 676995 957812 677061 957813
rect 676995 957748 676996 957812
rect 677060 957748 677061 957812
rect 676995 957747 677061 957748
rect 676811 956452 676877 956453
rect 676811 956388 676812 956452
rect 676876 956388 676877 956452
rect 676811 956387 676877 956388
rect 676627 951556 676693 951557
rect 676627 951492 676628 951556
rect 676692 951492 676693 951556
rect 676627 951491 676693 951492
rect 676075 950740 676141 950741
rect 676075 950676 676076 950740
rect 676140 950676 676141 950740
rect 676075 950675 676141 950676
rect 39803 943804 39869 943805
rect 39803 943740 39804 943804
rect 39868 943740 39869 943804
rect 39803 943739 39869 943740
rect 40723 943804 40789 943805
rect 40723 943740 40724 943804
rect 40788 943740 40789 943804
rect 40723 943739 40789 943740
rect 42011 943804 42077 943805
rect 42011 943740 42012 943804
rect 42076 943740 42077 943804
rect 42011 943739 42077 943740
rect 41781 939452 41847 939453
rect 41781 939450 41782 939452
rect 40358 939390 41782 939450
rect 40358 934290 40418 939390
rect 41781 939388 41782 939390
rect 41846 939388 41847 939452
rect 41781 939387 41847 939388
rect 42014 937050 42074 943739
rect 41830 936990 42074 937050
rect 41830 936733 41890 936990
rect 41827 936732 41893 936733
rect 41827 936668 41828 936732
rect 41892 936668 41893 936732
rect 41827 936667 41893 936668
rect 39990 934230 40418 934290
rect 39990 814299 40050 934230
rect 676814 931973 676874 956387
rect 676811 931972 676877 931973
rect 676811 931908 676812 931972
rect 676876 931908 676877 931972
rect 676811 931907 676877 931908
rect 676998 931565 677058 957747
rect 676995 931564 677061 931565
rect 676995 931500 676996 931564
rect 677060 931500 677061 931564
rect 676995 931499 677061 931500
rect 42011 911980 42077 911981
rect 42011 911916 42012 911980
rect 42076 911916 42077 911980
rect 42011 911915 42077 911916
rect 42014 885461 42074 911915
rect 42195 911708 42261 911709
rect 42195 911644 42196 911708
rect 42260 911644 42261 911708
rect 42195 911643 42261 911644
rect 42011 885460 42077 885461
rect 42011 885396 42012 885460
rect 42076 885396 42077 885460
rect 42011 885395 42077 885396
rect 42198 885189 42258 911643
rect 42195 885188 42261 885189
rect 42195 885124 42196 885188
rect 42260 885124 42261 885188
rect 42195 885123 42261 885124
rect 676075 875940 676141 875941
rect 676075 875876 676076 875940
rect 676140 875876 676141 875940
rect 676075 875875 676141 875876
rect 675339 874036 675405 874037
rect 675339 873972 675340 874036
rect 675404 873972 675405 874036
rect 675339 873971 675405 873972
rect 673867 873220 673933 873221
rect 673867 873156 673868 873220
rect 673932 873156 673933 873220
rect 673867 873155 673933 873156
rect 39987 814298 40053 814299
rect 39987 814234 39988 814298
rect 40052 814234 40053 814298
rect 39987 814233 40053 814234
rect 41827 813244 41893 813245
rect 41827 813180 41828 813244
rect 41892 813180 41893 813244
rect 41827 813179 41893 813180
rect 41830 812970 41890 813179
rect 41462 812910 41890 812970
rect 40907 805492 40973 805493
rect 40907 805428 40908 805492
rect 40972 805428 40973 805492
rect 40907 805427 40973 805428
rect 40539 805220 40605 805221
rect 40539 805156 40540 805220
rect 40604 805156 40605 805220
rect 40539 805155 40605 805156
rect 40542 792573 40602 805155
rect 40723 805084 40789 805085
rect 40723 805020 40724 805084
rect 40788 805020 40789 805084
rect 40723 805019 40789 805020
rect 40726 795021 40786 805019
rect 40723 795020 40789 795021
rect 40723 794956 40724 795020
rect 40788 794956 40789 795020
rect 40723 794955 40789 794956
rect 40910 794205 40970 805427
rect 40907 794204 40973 794205
rect 40907 794140 40908 794204
rect 40972 794140 40973 794204
rect 40907 794139 40973 794140
rect 40539 792572 40605 792573
rect 40539 792508 40540 792572
rect 40604 792508 40605 792572
rect 40539 792507 40605 792508
rect 41462 786861 41522 812910
rect 41827 809164 41893 809165
rect 41827 809100 41828 809164
rect 41892 809100 41893 809164
rect 41827 809099 41893 809100
rect 41830 805493 41890 809099
rect 41827 805492 41893 805493
rect 41827 805428 41828 805492
rect 41892 805428 41893 805492
rect 41827 805427 41893 805428
rect 41643 804812 41709 804813
rect 41643 804748 41644 804812
rect 41708 804748 41709 804812
rect 41643 804747 41709 804748
rect 41646 789037 41706 804747
rect 42011 804540 42077 804541
rect 42011 804476 42012 804540
rect 42076 804476 42077 804540
rect 42011 804475 42077 804476
rect 42014 794910 42074 804475
rect 42195 798964 42261 798965
rect 42195 798900 42196 798964
rect 42260 798900 42261 798964
rect 42195 798899 42261 798900
rect 42198 797877 42258 798899
rect 42195 797876 42261 797877
rect 42195 797812 42196 797876
rect 42260 797812 42261 797876
rect 42195 797811 42261 797812
rect 41830 794850 42074 794910
rect 41643 789036 41709 789037
rect 41643 788972 41644 789036
rect 41708 788972 41709 789036
rect 41643 788971 41709 788972
rect 41830 788629 41890 794850
rect 41827 788628 41893 788629
rect 41827 788564 41828 788628
rect 41892 788564 41893 788628
rect 41827 788563 41893 788564
rect 41459 786860 41525 786861
rect 41459 786796 41460 786860
rect 41524 786796 41525 786860
rect 41459 786795 41525 786796
rect 673870 770949 673930 873155
rect 675342 863157 675402 873971
rect 675339 863156 675405 863157
rect 675339 863092 675340 863156
rect 675404 863092 675405 863156
rect 675339 863091 675405 863092
rect 675707 777068 675773 777069
rect 675707 777004 675708 777068
rect 675772 777004 675773 777068
rect 675707 777003 675773 777004
rect 675710 775709 675770 777003
rect 675707 775708 675773 775709
rect 675707 775644 675708 775708
rect 675772 775644 675773 775708
rect 675707 775643 675773 775644
rect 676078 772717 676138 875875
rect 676995 870908 677061 870909
rect 676995 870844 676996 870908
rect 677060 870844 677061 870908
rect 676995 870843 677061 870844
rect 676811 774892 676877 774893
rect 676811 774828 676812 774892
rect 676876 774828 676877 774892
rect 676811 774827 676877 774828
rect 676075 772716 676141 772717
rect 676075 772652 676076 772716
rect 676140 772652 676141 772716
rect 676075 772651 676141 772652
rect 673867 770948 673933 770949
rect 673867 770884 673868 770948
rect 673932 770884 673933 770948
rect 673867 770883 673933 770884
rect 41459 769860 41525 769861
rect 41459 769796 41460 769860
rect 41524 769796 41525 769860
rect 41459 769795 41525 769796
rect 40907 765780 40973 765781
rect 40907 765716 40908 765780
rect 40972 765716 40973 765780
rect 40907 765715 40973 765716
rect 40539 765372 40605 765373
rect 40539 765308 40540 765372
rect 40604 765308 40605 765372
rect 40539 765307 40605 765308
rect 40355 757348 40421 757349
rect 40355 757284 40356 757348
rect 40420 757284 40421 757348
rect 40355 757283 40421 757284
rect 40358 754629 40418 757283
rect 40355 754628 40421 754629
rect 40355 754564 40356 754628
rect 40420 754564 40421 754628
rect 40355 754563 40421 754564
rect 40542 747421 40602 765307
rect 40723 764964 40789 764965
rect 40723 764900 40724 764964
rect 40788 764900 40789 764964
rect 40723 764899 40789 764900
rect 40726 750413 40786 764899
rect 40910 754901 40970 765715
rect 40907 754900 40973 754901
rect 40907 754836 40908 754900
rect 40972 754836 40973 754900
rect 40907 754835 40973 754836
rect 40723 750412 40789 750413
rect 40723 750348 40724 750412
rect 40788 750348 40789 750412
rect 40723 750347 40789 750348
rect 40539 747420 40605 747421
rect 40539 747356 40540 747420
rect 40604 747356 40605 747420
rect 40539 747355 40605 747356
rect 41462 743749 41522 769795
rect 675891 766596 675957 766597
rect 675891 766532 675892 766596
rect 675956 766532 675957 766596
rect 675891 766531 675957 766532
rect 676075 766596 676141 766597
rect 676075 766532 676076 766596
rect 676140 766532 676141 766596
rect 676075 766531 676141 766532
rect 41643 764556 41709 764557
rect 41643 764492 41644 764556
rect 41708 764492 41709 764556
rect 41643 764491 41709 764492
rect 41646 744429 41706 764491
rect 42379 758708 42445 758709
rect 42379 758644 42380 758708
rect 42444 758644 42445 758708
rect 42379 758643 42445 758644
rect 41827 757756 41893 757757
rect 41827 757692 41828 757756
rect 41892 757692 41893 757756
rect 41827 757691 41893 757692
rect 41830 745381 41890 757691
rect 42382 754901 42442 758643
rect 42011 754900 42077 754901
rect 42011 754836 42012 754900
rect 42076 754836 42077 754900
rect 42011 754835 42077 754836
rect 42379 754900 42445 754901
rect 42379 754836 42380 754900
rect 42444 754836 42445 754900
rect 42379 754835 42445 754836
rect 42014 751093 42074 754835
rect 42011 751092 42077 751093
rect 42011 751028 42012 751092
rect 42076 751028 42077 751092
rect 42011 751027 42077 751028
rect 41827 745380 41893 745381
rect 41827 745316 41828 745380
rect 41892 745316 41893 745380
rect 41827 745315 41893 745316
rect 41643 744428 41709 744429
rect 41643 744364 41644 744428
rect 41708 744364 41709 744428
rect 41643 744363 41709 744364
rect 41459 743748 41525 743749
rect 41459 743684 41460 743748
rect 41524 743684 41525 743748
rect 41459 743683 41525 743684
rect 674419 742524 674485 742525
rect 674419 742460 674420 742524
rect 674484 742460 674485 742524
rect 674419 742459 674485 742460
rect 674235 741572 674301 741573
rect 674235 741508 674236 741572
rect 674300 741508 674301 741572
rect 674235 741507 674301 741508
rect 672027 732868 672093 732869
rect 672027 732804 672028 732868
rect 672092 732804 672093 732868
rect 672027 732803 672093 732804
rect 673315 732868 673381 732869
rect 673315 732804 673316 732868
rect 673380 732804 673381 732868
rect 673315 732803 673381 732804
rect 672030 728245 672090 732803
rect 673318 728517 673378 732803
rect 673315 728516 673381 728517
rect 673315 728452 673316 728516
rect 673380 728452 673381 728516
rect 673315 728451 673381 728452
rect 672027 728244 672093 728245
rect 672027 728180 672028 728244
rect 672092 728180 672093 728244
rect 672027 728179 672093 728180
rect 41827 726884 41893 726885
rect 41827 726820 41828 726884
rect 41892 726820 41893 726884
rect 41827 726819 41893 726820
rect 41830 726610 41890 726819
rect 41462 726550 41890 726610
rect 40723 721772 40789 721773
rect 40723 721708 40724 721772
rect 40788 721708 40789 721772
rect 40723 721707 40789 721708
rect 40539 718588 40605 718589
rect 40539 718524 40540 718588
rect 40604 718524 40605 718588
rect 40539 718523 40605 718524
rect 40542 709205 40602 718523
rect 40539 709204 40605 709205
rect 40539 709140 40540 709204
rect 40604 709140 40605 709204
rect 40539 709139 40605 709140
rect 40726 707437 40786 721707
rect 40723 707436 40789 707437
rect 40723 707372 40724 707436
rect 40788 707372 40789 707436
rect 40723 707371 40789 707372
rect 41462 701861 41522 726550
rect 41643 721772 41709 721773
rect 41643 721708 41644 721772
rect 41708 721708 41709 721772
rect 41643 721707 41709 721708
rect 41646 702133 41706 721707
rect 42563 718316 42629 718317
rect 42563 718252 42564 718316
rect 42628 718252 42629 718316
rect 42563 718251 42629 718252
rect 41827 714780 41893 714781
rect 41827 714716 41828 714780
rect 41892 714716 41893 714780
rect 41827 714715 41893 714716
rect 42011 714780 42077 714781
rect 42011 714716 42012 714780
rect 42076 714716 42077 714780
rect 42011 714715 42077 714716
rect 41643 702132 41709 702133
rect 41643 702068 41644 702132
rect 41708 702068 41709 702132
rect 41643 702067 41709 702068
rect 41459 701860 41525 701861
rect 41459 701796 41460 701860
rect 41524 701796 41525 701860
rect 41459 701795 41525 701796
rect 41830 701589 41890 714715
rect 42014 713421 42074 714715
rect 42379 714236 42445 714237
rect 42379 714172 42380 714236
rect 42444 714172 42445 714236
rect 42379 714171 42445 714172
rect 42011 713420 42077 713421
rect 42011 713356 42012 713420
rect 42076 713356 42077 713420
rect 42011 713355 42077 713356
rect 42382 706621 42442 714171
rect 42566 711653 42626 718251
rect 42563 711652 42629 711653
rect 42563 711588 42564 711652
rect 42628 711588 42629 711652
rect 42563 711587 42629 711588
rect 42379 706620 42445 706621
rect 42379 706556 42380 706620
rect 42444 706556 42445 706620
rect 42379 706555 42445 706556
rect 41827 701588 41893 701589
rect 41827 701524 41828 701588
rect 41892 701524 41893 701588
rect 41827 701523 41893 701524
rect 41827 683636 41893 683637
rect 41827 683572 41828 683636
rect 41892 683572 41893 683636
rect 41827 683571 41893 683572
rect 41830 683130 41890 683571
rect 41462 683070 41890 683130
rect 40539 678992 40605 678993
rect 40539 678928 40540 678992
rect 40604 678928 40605 678992
rect 40539 678927 40605 678928
rect 40723 678992 40789 678993
rect 40723 678928 40724 678992
rect 40788 678928 40789 678992
rect 40723 678927 40789 678928
rect 40355 671260 40421 671261
rect 40355 671196 40356 671260
rect 40420 671196 40421 671260
rect 40355 671195 40421 671196
rect 40358 670309 40418 671195
rect 40355 670308 40421 670309
rect 40355 670244 40356 670308
rect 40420 670244 40421 670308
rect 40355 670243 40421 670244
rect 40542 664189 40602 678927
rect 40726 665413 40786 678927
rect 40723 665412 40789 665413
rect 40723 665348 40724 665412
rect 40788 665348 40789 665412
rect 40723 665347 40789 665348
rect 40539 664188 40605 664189
rect 40539 664124 40540 664188
rect 40604 664124 40605 664188
rect 40539 664123 40605 664124
rect 41462 660789 41522 683070
rect 674238 682413 674298 741507
rect 674422 682685 674482 742459
rect 674603 739668 674669 739669
rect 674603 739604 674604 739668
rect 674668 739604 674669 739668
rect 674603 739603 674669 739604
rect 674419 682684 674485 682685
rect 674419 682620 674420 682684
rect 674484 682620 674485 682684
rect 674419 682619 674485 682620
rect 674235 682412 674301 682413
rect 674235 682348 674236 682412
rect 674300 682348 674301 682412
rect 674235 682347 674301 682348
rect 41827 681052 41893 681053
rect 41827 680988 41828 681052
rect 41892 680988 41893 681052
rect 41827 680987 41893 680988
rect 41830 678990 41890 680987
rect 41646 678930 41890 678990
rect 41459 660788 41525 660789
rect 41459 660724 41460 660788
rect 41524 660724 41525 660788
rect 41459 660723 41525 660724
rect 41646 658613 41706 678930
rect 42379 674252 42445 674253
rect 42379 674188 42380 674252
rect 42444 674188 42445 674252
rect 42379 674187 42445 674188
rect 42011 671260 42077 671261
rect 42011 671196 42012 671260
rect 42076 671196 42077 671260
rect 42011 671195 42077 671196
rect 41827 670988 41893 670989
rect 41827 670924 41828 670988
rect 41892 670924 41893 670988
rect 41827 670923 41893 670924
rect 41643 658612 41709 658613
rect 41643 658548 41644 658612
rect 41708 658548 41709 658612
rect 41643 658547 41709 658548
rect 41830 658341 41890 670923
rect 42014 667317 42074 671195
rect 42195 669356 42261 669357
rect 42195 669292 42196 669356
rect 42260 669292 42261 669356
rect 42195 669291 42261 669292
rect 42198 667997 42258 669291
rect 42382 668541 42442 674187
rect 674606 673470 674666 739603
rect 675894 730013 675954 766531
rect 675891 730012 675957 730013
rect 675891 729948 675892 730012
rect 675956 729948 675957 730012
rect 675891 729947 675957 729948
rect 676078 725797 676138 766531
rect 676814 761837 676874 774827
rect 676998 761973 677058 870843
rect 676995 761972 677061 761973
rect 676995 761908 676996 761972
rect 677060 761908 677061 761972
rect 676995 761907 677061 761908
rect 676811 761836 676877 761837
rect 676811 761772 676812 761836
rect 676876 761772 676877 761836
rect 676811 761771 676877 761772
rect 676811 730012 676877 730013
rect 676811 729948 676812 730012
rect 676876 729948 676877 730012
rect 676811 729947 676877 729948
rect 676075 725796 676141 725797
rect 676075 725732 676076 725796
rect 676140 725732 676141 725796
rect 676075 725731 676141 725732
rect 676814 712110 676874 729947
rect 675894 712061 676874 712110
rect 675891 712060 676874 712061
rect 675891 711996 675892 712060
rect 675956 712050 676874 712060
rect 675956 711996 675957 712050
rect 675891 711995 675957 711996
rect 675339 696828 675405 696829
rect 675339 696764 675340 696828
rect 675404 696764 675405 696828
rect 675339 696763 675405 696764
rect 675342 686493 675402 696763
rect 676995 694108 677061 694109
rect 676995 694044 676996 694108
rect 677060 694044 677061 694108
rect 676995 694043 677061 694044
rect 675339 686492 675405 686493
rect 675339 686428 675340 686492
rect 675404 686428 675405 686492
rect 675339 686427 675405 686428
rect 674606 673410 674850 673470
rect 42379 668540 42445 668541
rect 42379 668476 42380 668540
rect 42444 668476 42445 668540
rect 42379 668475 42445 668476
rect 42195 667996 42261 667997
rect 42195 667932 42196 667996
rect 42260 667932 42261 667996
rect 42195 667931 42261 667932
rect 42011 667316 42077 667317
rect 42011 667252 42012 667316
rect 42076 667252 42077 667316
rect 42011 667251 42077 667252
rect 674790 664053 674850 673410
rect 674787 664052 674853 664053
rect 674787 663988 674788 664052
rect 674852 663988 674853 664052
rect 674787 663987 674853 663988
rect 41827 658340 41893 658341
rect 41827 658276 41828 658340
rect 41892 658276 41893 658340
rect 41827 658275 41893 658276
rect 44219 653172 44285 653173
rect 44219 653108 44220 653172
rect 44284 653108 44285 653172
rect 44219 653107 44285 653108
rect 41643 640660 41709 640661
rect 41643 640596 41644 640660
rect 41708 640596 41709 640660
rect 41643 640595 41709 640596
rect 41459 639436 41525 639437
rect 41459 639372 41460 639436
rect 41524 639372 41525 639436
rect 41459 639371 41525 639372
rect 40723 634948 40789 634949
rect 40723 634884 40724 634948
rect 40788 634884 40789 634948
rect 40723 634883 40789 634884
rect 40539 634540 40605 634541
rect 40539 634476 40540 634540
rect 40604 634476 40605 634540
rect 40539 634475 40605 634476
rect 40542 619989 40602 634475
rect 40726 623797 40786 634883
rect 40723 623796 40789 623797
rect 40723 623732 40724 623796
rect 40788 623732 40789 623796
rect 40723 623731 40789 623732
rect 40539 619988 40605 619989
rect 40539 619924 40540 619988
rect 40604 619924 40605 619988
rect 40539 619923 40605 619924
rect 41462 615501 41522 639371
rect 41646 617130 41706 640595
rect 41827 637396 41893 637397
rect 41827 637332 41828 637396
rect 41892 637332 41893 637396
rect 41827 637331 41893 637332
rect 41830 630690 41890 637331
rect 41830 630630 42074 630690
rect 41827 627740 41893 627741
rect 41827 627676 41828 627740
rect 41892 627676 41893 627740
rect 41827 627675 41893 627676
rect 41830 620261 41890 627675
rect 41827 620260 41893 620261
rect 41827 620196 41828 620260
rect 41892 620196 41893 620260
rect 41827 620195 41893 620196
rect 41646 617070 41890 617130
rect 41459 615500 41525 615501
rect 41459 615436 41460 615500
rect 41524 615436 41525 615500
rect 41459 615435 41525 615436
rect 41830 614141 41890 617070
rect 42014 615909 42074 630630
rect 42011 615908 42077 615909
rect 42011 615844 42012 615908
rect 42076 615844 42077 615908
rect 42011 615843 42077 615844
rect 44222 614141 44282 653107
rect 675339 652900 675405 652901
rect 675339 652836 675340 652900
rect 675404 652836 675405 652900
rect 675339 652835 675405 652836
rect 674787 650180 674853 650181
rect 674787 650116 674788 650180
rect 674852 650116 674853 650180
rect 674787 650115 674853 650116
rect 674790 647597 674850 650115
rect 674787 647596 674853 647597
rect 674787 647532 674788 647596
rect 674852 647532 674853 647596
rect 674787 647531 674853 647532
rect 675155 645828 675221 645829
rect 675155 645764 675156 645828
rect 675220 645764 675221 645828
rect 675155 645763 675221 645764
rect 674051 645148 674117 645149
rect 674051 645084 674052 645148
rect 674116 645084 674117 645148
rect 674051 645083 674117 645084
rect 671475 643516 671541 643517
rect 671475 643452 671476 643516
rect 671540 643452 671541 643516
rect 671475 643451 671541 643452
rect 41827 614140 41893 614141
rect 41827 614076 41828 614140
rect 41892 614076 41893 614140
rect 41827 614075 41893 614076
rect 44219 614140 44285 614141
rect 44219 614076 44220 614140
rect 44284 614076 44285 614140
rect 44219 614075 44285 614076
rect 41827 596052 41893 596053
rect 41827 595988 41828 596052
rect 41892 595988 41893 596052
rect 41827 595987 41893 595988
rect 40723 592414 40789 592415
rect 40723 592350 40724 592414
rect 40788 592350 40789 592414
rect 40723 592349 40789 592350
rect 40539 589388 40605 589389
rect 40539 589324 40540 589388
rect 40604 589324 40605 589388
rect 40539 589323 40605 589324
rect 40542 576877 40602 589323
rect 40726 577557 40786 592349
rect 41830 592050 41890 595987
rect 42011 594964 42077 594965
rect 42011 594900 42012 594964
rect 42076 594900 42077 594964
rect 42011 594899 42077 594900
rect 41646 591990 41890 592050
rect 40907 589660 40973 589661
rect 40907 589596 40908 589660
rect 40972 589596 40973 589660
rect 40907 589595 40973 589596
rect 40910 578237 40970 589595
rect 41459 587212 41525 587213
rect 41459 587148 41460 587212
rect 41524 587148 41525 587212
rect 41459 587147 41525 587148
rect 41091 584628 41157 584629
rect 41091 584564 41092 584628
rect 41156 584564 41157 584628
rect 41091 584563 41157 584564
rect 41094 580277 41154 584563
rect 41091 580276 41157 580277
rect 41091 580212 41092 580276
rect 41156 580212 41157 580276
rect 41091 580211 41157 580212
rect 40907 578236 40973 578237
rect 40907 578172 40908 578236
rect 40972 578172 40973 578236
rect 40907 578171 40973 578172
rect 40723 577556 40789 577557
rect 40723 577492 40724 577556
rect 40788 577492 40789 577556
rect 40723 577491 40789 577492
rect 40539 576876 40605 576877
rect 40539 576812 40540 576876
rect 40604 576812 40605 576876
rect 40539 576811 40605 576812
rect 41462 571981 41522 587147
rect 41459 571980 41525 571981
rect 41459 571916 41460 571980
rect 41524 571916 41525 571980
rect 41459 571915 41525 571916
rect 41646 571029 41706 591990
rect 42014 587213 42074 594899
rect 43851 591564 43917 591565
rect 43851 591500 43852 591564
rect 43916 591500 43917 591564
rect 43851 591499 43917 591500
rect 42011 587212 42077 587213
rect 42011 587148 42012 587212
rect 42076 587148 42077 587212
rect 42011 587147 42077 587148
rect 42379 586124 42445 586125
rect 42379 586060 42380 586124
rect 42444 586060 42445 586124
rect 42379 586059 42445 586060
rect 41827 585172 41893 585173
rect 41827 585108 41828 585172
rect 41892 585108 41893 585172
rect 41827 585107 41893 585108
rect 41830 572253 41890 585107
rect 42195 584900 42261 584901
rect 42195 584836 42196 584900
rect 42260 584836 42261 584900
rect 42195 584835 42261 584836
rect 42198 581501 42258 584835
rect 42382 581909 42442 586059
rect 42379 581908 42445 581909
rect 42379 581844 42380 581908
rect 42444 581844 42445 581908
rect 42379 581843 42445 581844
rect 42195 581500 42261 581501
rect 42195 581436 42196 581500
rect 42260 581436 42261 581500
rect 42195 581435 42261 581436
rect 42195 576196 42261 576197
rect 42195 576132 42196 576196
rect 42260 576132 42261 576196
rect 42195 576131 42261 576132
rect 42198 572661 42258 576131
rect 42195 572660 42261 572661
rect 42195 572596 42196 572660
rect 42260 572596 42261 572660
rect 42195 572595 42261 572596
rect 41827 572252 41893 572253
rect 41827 572188 41828 572252
rect 41892 572188 41893 572252
rect 41827 572187 41893 572188
rect 41643 571028 41709 571029
rect 41643 570964 41644 571028
rect 41708 570964 41709 571028
rect 41643 570963 41709 570964
rect 41827 553212 41893 553213
rect 41827 553210 41828 553212
rect 41462 553150 41828 553210
rect 40539 545732 40605 545733
rect 40539 545668 40540 545732
rect 40604 545668 40605 545732
rect 40539 545667 40605 545668
rect 40542 538253 40602 545667
rect 40723 545460 40789 545461
rect 40723 545396 40724 545460
rect 40788 545396 40789 545460
rect 40723 545395 40789 545396
rect 40726 538661 40786 545395
rect 40723 538660 40789 538661
rect 40723 538596 40724 538660
rect 40788 538596 40789 538660
rect 40723 538595 40789 538596
rect 40539 538252 40605 538253
rect 40539 538188 40540 538252
rect 40604 538188 40605 538252
rect 40539 538187 40605 538188
rect 41462 530637 41522 553150
rect 41827 553148 41828 553150
rect 41892 553148 41893 553212
rect 41827 553147 41893 553148
rect 41827 551988 41893 551989
rect 41827 551924 41828 551988
rect 41892 551924 41893 551988
rect 41827 551923 41893 551924
rect 41643 546412 41709 546413
rect 41643 546348 41644 546412
rect 41708 546348 41709 546412
rect 41643 546347 41709 546348
rect 41459 530636 41525 530637
rect 41459 530572 41460 530636
rect 41524 530572 41525 530636
rect 41459 530571 41525 530572
rect 41646 529141 41706 546347
rect 41830 529413 41890 551923
rect 42011 549948 42077 549949
rect 42011 549884 42012 549948
rect 42076 549884 42077 549948
rect 42011 549883 42077 549884
rect 42014 545461 42074 549883
rect 42011 545460 42077 545461
rect 42011 545396 42012 545460
rect 42076 545396 42077 545460
rect 42011 545395 42077 545396
rect 41827 529412 41893 529413
rect 41827 529348 41828 529412
rect 41892 529348 41893 529412
rect 41827 529347 41893 529348
rect 41643 529140 41709 529141
rect 41643 529076 41644 529140
rect 41708 529076 41709 529140
rect 41643 529075 41709 529076
rect 41827 425236 41893 425237
rect 41827 425172 41828 425236
rect 41892 425172 41893 425236
rect 41827 425171 41893 425172
rect 41830 424690 41890 425171
rect 42011 424828 42077 424829
rect 42011 424764 42012 424828
rect 42076 424764 42077 424828
rect 42011 424763 42077 424764
rect 41646 424630 41890 424690
rect 41459 418844 41525 418845
rect 41459 418780 41460 418844
rect 41524 418780 41525 418844
rect 41459 418779 41525 418780
rect 40723 417892 40789 417893
rect 40723 417828 40724 417892
rect 40788 417828 40789 417892
rect 40723 417827 40789 417828
rect 40539 417620 40605 417621
rect 40539 417556 40540 417620
rect 40604 417556 40605 417620
rect 40539 417555 40605 417556
rect 40542 403885 40602 417555
rect 40726 409461 40786 417827
rect 40723 409460 40789 409461
rect 40723 409396 40724 409460
rect 40788 409396 40789 409460
rect 40723 409395 40789 409396
rect 40539 403884 40605 403885
rect 40539 403820 40540 403884
rect 40604 403820 40605 403884
rect 40539 403819 40605 403820
rect 41462 398853 41522 418779
rect 41646 402990 41706 424630
rect 42014 415410 42074 424763
rect 41830 415350 42074 415410
rect 41830 406333 41890 415350
rect 41827 406332 41893 406333
rect 41827 406268 41828 406332
rect 41892 406268 41893 406332
rect 41827 406267 41893 406268
rect 41646 402930 41890 402990
rect 41830 401845 41890 402930
rect 41827 401844 41893 401845
rect 41827 401780 41828 401844
rect 41892 401780 41893 401844
rect 41827 401779 41893 401780
rect 41459 398852 41525 398853
rect 41459 398788 41460 398852
rect 41524 398788 41525 398852
rect 41459 398787 41525 398788
rect 41459 381852 41525 381853
rect 41459 381788 41460 381852
rect 41524 381788 41525 381852
rect 41459 381787 41525 381788
rect 40539 378588 40605 378589
rect 40539 378524 40540 378588
rect 40604 378524 40605 378588
rect 40539 378523 40605 378524
rect 40542 360093 40602 378523
rect 40723 378180 40789 378181
rect 40723 378116 40724 378180
rect 40788 378116 40789 378180
rect 40723 378115 40789 378116
rect 40726 363629 40786 378115
rect 41275 373284 41341 373285
rect 41275 373220 41276 373284
rect 41340 373220 41341 373284
rect 41275 373219 41341 373220
rect 41278 368525 41338 373219
rect 41275 368524 41341 368525
rect 41275 368460 41276 368524
rect 41340 368460 41341 368524
rect 41275 368459 41341 368460
rect 40723 363628 40789 363629
rect 40723 363564 40724 363628
rect 40788 363564 40789 363628
rect 40723 363563 40789 363564
rect 40539 360092 40605 360093
rect 40539 360028 40540 360092
rect 40604 360028 40605 360092
rect 40539 360027 40605 360028
rect 41462 358733 41522 381787
rect 41643 376956 41709 376957
rect 41643 376892 41644 376956
rect 41708 376892 41709 376956
rect 41643 376891 41709 376892
rect 41459 358732 41525 358733
rect 41459 358668 41460 358732
rect 41524 358668 41525 358732
rect 41459 358667 41525 358668
rect 41646 358050 41706 376891
rect 41827 371924 41893 371925
rect 41827 371860 41828 371924
rect 41892 371860 41893 371924
rect 41827 371859 41893 371860
rect 41830 359413 41890 371859
rect 41827 359412 41893 359413
rect 41827 359348 41828 359412
rect 41892 359348 41893 359412
rect 41827 359347 41893 359348
rect 41646 357990 41890 358050
rect 41830 355741 41890 357990
rect 41827 355740 41893 355741
rect 41827 355676 41828 355740
rect 41892 355676 41893 355740
rect 41827 355675 41893 355676
rect 43854 354245 43914 591499
rect 671478 571301 671538 643451
rect 673867 616180 673933 616181
rect 673867 616116 673868 616180
rect 673932 616116 673933 616180
rect 673867 616115 673933 616116
rect 673683 595372 673749 595373
rect 673683 595308 673684 595372
rect 673748 595308 673749 595372
rect 673683 595307 673749 595308
rect 673686 591701 673746 595307
rect 673683 591700 673749 591701
rect 673683 591636 673684 591700
rect 673748 591636 673749 591700
rect 673683 591635 673749 591636
rect 671475 571300 671541 571301
rect 671475 571236 671476 571300
rect 671540 571236 671541 571300
rect 671475 571235 671541 571236
rect 673683 475420 673749 475421
rect 673683 475356 673684 475420
rect 673748 475356 673749 475420
rect 673683 475355 673749 475356
rect 673686 464813 673746 475355
rect 673683 464812 673749 464813
rect 673683 464748 673684 464812
rect 673748 464748 673749 464812
rect 673683 464747 673749 464748
rect 673870 455157 673930 616115
rect 674054 475421 674114 645083
rect 674971 644332 675037 644333
rect 674971 644268 674972 644332
rect 675036 644268 675037 644332
rect 674971 644267 675037 644268
rect 674974 640797 675034 644267
rect 674971 640796 675037 640797
rect 674971 640732 674972 640796
rect 675036 640732 675037 640796
rect 674971 640731 675037 640732
rect 675158 638077 675218 645763
rect 675155 638076 675221 638077
rect 675155 638012 675156 638076
rect 675220 638012 675221 638076
rect 675155 638011 675221 638012
rect 675342 637669 675402 652835
rect 675523 648140 675589 648141
rect 675523 648076 675524 648140
rect 675588 648076 675589 648140
rect 675523 648075 675589 648076
rect 675526 647461 675586 648075
rect 675523 647460 675589 647461
rect 675523 647396 675524 647460
rect 675588 647396 675589 647460
rect 675523 647395 675589 647396
rect 676811 644332 676877 644333
rect 676811 644268 676812 644332
rect 676876 644268 676877 644332
rect 676811 644267 676877 644268
rect 675523 644060 675589 644061
rect 675523 643996 675524 644060
rect 675588 643996 675589 644060
rect 675523 643995 675589 643996
rect 675526 640253 675586 643995
rect 675523 640252 675589 640253
rect 675523 640188 675524 640252
rect 675588 640188 675589 640252
rect 675523 640187 675589 640188
rect 676627 640252 676693 640253
rect 676627 640188 676628 640252
rect 676692 640188 676693 640252
rect 676627 640187 676693 640188
rect 676630 637941 676690 640187
rect 676627 637940 676693 637941
rect 676627 637876 676628 637940
rect 676692 637876 676693 637940
rect 676627 637875 676693 637876
rect 675339 637668 675405 637669
rect 675339 637604 675340 637668
rect 675404 637604 675405 637668
rect 675339 637603 675405 637604
rect 675339 631412 675405 631413
rect 675339 631348 675340 631412
rect 675404 631348 675405 631412
rect 675339 631347 675405 631348
rect 676075 631412 676141 631413
rect 676075 631348 676076 631412
rect 676140 631348 676141 631412
rect 676075 631347 676141 631348
rect 674419 602852 674485 602853
rect 674419 602788 674420 602852
rect 674484 602788 674485 602852
rect 674419 602787 674485 602788
rect 674422 527101 674482 602787
rect 674787 595644 674853 595645
rect 674787 595580 674788 595644
rect 674852 595580 674853 595644
rect 674787 595579 674853 595580
rect 674790 591429 674850 595579
rect 675342 592381 675402 631347
rect 675523 608292 675589 608293
rect 675523 608228 675524 608292
rect 675588 608228 675589 608292
rect 675523 608227 675589 608228
rect 675339 592380 675405 592381
rect 675339 592316 675340 592380
rect 675404 592316 675405 592380
rect 675339 592315 675405 592316
rect 675526 592109 675586 608227
rect 676078 593469 676138 631347
rect 676075 593468 676141 593469
rect 676075 593404 676076 593468
rect 676140 593404 676141 593468
rect 676075 593403 676141 593404
rect 675523 592108 675589 592109
rect 675523 592044 675524 592108
rect 675588 592044 675589 592108
rect 675523 592043 675589 592044
rect 674787 591428 674853 591429
rect 674787 591364 674788 591428
rect 674852 591364 674853 591428
rect 674787 591363 674853 591364
rect 676075 586260 676141 586261
rect 676075 586196 676076 586260
rect 676140 586196 676141 586260
rect 676075 586195 676141 586196
rect 675339 563140 675405 563141
rect 675339 563076 675340 563140
rect 675404 563076 675405 563140
rect 675339 563075 675405 563076
rect 675342 553410 675402 563075
rect 675523 561236 675589 561237
rect 675523 561172 675524 561236
rect 675588 561172 675589 561236
rect 675523 561171 675589 561172
rect 674974 553350 675402 553410
rect 674974 550650 675034 553350
rect 674790 550590 675034 550650
rect 674790 543829 674850 550590
rect 675155 549676 675221 549677
rect 675155 549612 675156 549676
rect 675220 549612 675221 549676
rect 675155 549611 675221 549612
rect 675158 547909 675218 549611
rect 675155 547908 675221 547909
rect 675155 547844 675156 547908
rect 675220 547844 675221 547908
rect 675155 547843 675221 547844
rect 675526 547637 675586 561171
rect 675523 547636 675589 547637
rect 675523 547572 675524 547636
rect 675588 547572 675589 547636
rect 675523 547571 675589 547572
rect 676078 546549 676138 586195
rect 676814 572797 676874 644267
rect 676998 619173 677058 694043
rect 676995 619172 677061 619173
rect 676995 619108 676996 619172
rect 677060 619108 677061 619172
rect 676995 619107 677061 619108
rect 676995 593468 677061 593469
rect 676995 593404 676996 593468
rect 677060 593404 677061 593468
rect 676995 593403 677061 593404
rect 676998 576061 677058 593403
rect 676995 576060 677061 576061
rect 676995 575996 676996 576060
rect 677060 575996 677061 576060
rect 676995 575995 677061 575996
rect 676811 572796 676877 572797
rect 676811 572732 676812 572796
rect 676876 572732 676877 572796
rect 676811 572731 676877 572732
rect 676811 554708 676877 554709
rect 676811 554644 676812 554708
rect 676876 554644 676877 554708
rect 676811 554643 676877 554644
rect 676075 546548 676141 546549
rect 676075 546484 676076 546548
rect 676140 546484 676141 546548
rect 676075 546483 676141 546484
rect 674787 543828 674853 543829
rect 674787 543764 674788 543828
rect 674852 543764 674853 543828
rect 674787 543763 674853 543764
rect 674419 527100 674485 527101
rect 674419 527036 674420 527100
rect 674484 527036 674485 527100
rect 674419 527035 674485 527036
rect 676814 503709 676874 554643
rect 677179 550764 677245 550765
rect 677179 550700 677180 550764
rect 677244 550700 677245 550764
rect 677179 550699 677245 550700
rect 676811 503708 676877 503709
rect 676811 503644 676812 503708
rect 676876 503644 676877 503708
rect 676811 503643 676877 503644
rect 677182 495450 677242 550699
rect 677182 495390 677426 495450
rect 677366 492421 677426 495390
rect 677363 492420 677429 492421
rect 677363 492356 677364 492420
rect 677428 492356 677429 492420
rect 677363 492355 677429 492356
rect 675891 490516 675957 490517
rect 675891 490452 675892 490516
rect 675956 490452 675957 490516
rect 675891 490451 675957 490452
rect 675894 489970 675954 490451
rect 675894 489910 676322 489970
rect 676262 485790 676322 489910
rect 676995 485792 677061 485793
rect 676262 485730 676874 485790
rect 674051 475420 674117 475421
rect 674051 475356 674052 475420
rect 674116 475356 674117 475420
rect 674051 475355 674117 475356
rect 673867 455156 673933 455157
rect 673867 455092 673868 455156
rect 673932 455092 673933 455156
rect 673867 455091 673933 455092
rect 676814 402933 676874 485730
rect 676995 485728 676996 485792
rect 677060 485728 677061 485792
rect 676995 485727 677061 485728
rect 676811 402932 676877 402933
rect 676811 402868 676812 402932
rect 676876 402868 676877 402932
rect 676811 402867 676877 402868
rect 676998 401301 677058 485727
rect 676995 401300 677061 401301
rect 676995 401236 676996 401300
rect 677060 401236 677061 401300
rect 676995 401235 677061 401236
rect 675891 398852 675957 398853
rect 675891 398788 675892 398852
rect 675956 398788 675957 398852
rect 675891 398787 675957 398788
rect 675707 387700 675773 387701
rect 675707 387636 675708 387700
rect 675772 387636 675773 387700
rect 675707 387635 675773 387636
rect 675710 378725 675770 387635
rect 675707 378724 675773 378725
rect 675707 378660 675708 378724
rect 675772 378660 675773 378724
rect 675707 378659 675773 378660
rect 674787 378044 674853 378045
rect 674787 377980 674788 378044
rect 674852 377980 674853 378044
rect 674787 377979 674853 377980
rect 674790 372605 674850 377979
rect 675894 376957 675954 398787
rect 676627 396812 676693 396813
rect 676627 396748 676628 396812
rect 676692 396748 676693 396812
rect 676627 396747 676693 396748
rect 676259 395180 676325 395181
rect 676259 395116 676260 395180
rect 676324 395116 676325 395180
rect 676259 395115 676325 395116
rect 676075 393140 676141 393141
rect 676075 393076 676076 393140
rect 676140 393076 676141 393140
rect 676075 393075 676141 393076
rect 675891 376956 675957 376957
rect 675891 376892 675892 376956
rect 675956 376892 675957 376956
rect 675891 376891 675957 376892
rect 676078 373013 676138 393075
rect 676262 377365 676322 395115
rect 676443 394772 676509 394773
rect 676443 394708 676444 394772
rect 676508 394708 676509 394772
rect 676443 394707 676509 394708
rect 676446 380629 676506 394707
rect 676630 384981 676690 396747
rect 676627 384980 676693 384981
rect 676627 384916 676628 384980
rect 676692 384916 676693 384980
rect 676627 384915 676693 384916
rect 676443 380628 676509 380629
rect 676443 380564 676444 380628
rect 676508 380564 676509 380628
rect 676443 380563 676509 380564
rect 676259 377364 676325 377365
rect 676259 377300 676260 377364
rect 676324 377300 676325 377364
rect 676259 377299 676325 377300
rect 676075 373012 676141 373013
rect 676075 372948 676076 373012
rect 676140 372948 676141 373012
rect 676075 372947 676141 372948
rect 674787 372604 674853 372605
rect 674787 372540 674788 372604
rect 674852 372540 674853 372604
rect 674787 372539 674853 372540
rect 43851 354244 43917 354245
rect 43851 354180 43852 354244
rect 43916 354180 43917 354244
rect 43851 354179 43917 354180
rect 675339 354244 675405 354245
rect 675339 354180 675340 354244
rect 675404 354180 675405 354244
rect 675339 354179 675405 354180
rect 44219 353836 44285 353837
rect 44219 353772 44220 353836
rect 44284 353772 44285 353836
rect 44219 353771 44285 353772
rect 44222 342685 44282 353771
rect 44403 342956 44469 342957
rect 44403 342892 44404 342956
rect 44468 342892 44469 342956
rect 44403 342891 44469 342892
rect 44219 342684 44285 342685
rect 44219 342620 44220 342684
rect 44284 342620 44285 342684
rect 44219 342619 44285 342620
rect 44406 342410 44466 342891
rect 44222 342350 44466 342410
rect 43667 340508 43733 340509
rect 43667 340444 43668 340508
rect 43732 340444 43733 340508
rect 43667 340443 43733 340444
rect 40723 337788 40789 337789
rect 40723 337724 40724 337788
rect 40788 337724 40789 337788
rect 40723 337723 40789 337724
rect 40539 335748 40605 335749
rect 40539 335684 40540 335748
rect 40604 335684 40605 335748
rect 40539 335683 40605 335684
rect 40542 321061 40602 335683
rect 40726 326773 40786 337723
rect 42931 337652 42997 337653
rect 42931 337588 42932 337652
rect 42996 337588 42997 337652
rect 42931 337587 42997 337588
rect 42195 335068 42261 335069
rect 42195 335004 42196 335068
rect 42260 335004 42261 335068
rect 42195 335003 42261 335004
rect 41827 334524 41893 334525
rect 41827 334460 41828 334524
rect 41892 334460 41893 334524
rect 41827 334459 41893 334460
rect 40907 333708 40973 333709
rect 40907 333644 40908 333708
rect 40972 333644 40973 333708
rect 40907 333643 40973 333644
rect 40723 326772 40789 326773
rect 40723 326708 40724 326772
rect 40788 326708 40789 326772
rect 40723 326707 40789 326708
rect 40910 325413 40970 333643
rect 41643 329084 41709 329085
rect 41643 329020 41644 329084
rect 41708 329020 41709 329084
rect 41643 329019 41709 329020
rect 41459 328404 41525 328405
rect 41459 328340 41460 328404
rect 41524 328340 41525 328404
rect 41459 328339 41525 328340
rect 40907 325412 40973 325413
rect 40907 325348 40908 325412
rect 40972 325348 40973 325412
rect 40907 325347 40973 325348
rect 40539 321060 40605 321061
rect 40539 320996 40540 321060
rect 40604 320996 40605 321060
rect 40539 320995 40605 320996
rect 41462 312629 41522 328339
rect 41646 316050 41706 329019
rect 41830 324733 41890 334459
rect 42198 334389 42258 335003
rect 42195 334388 42261 334389
rect 42195 334324 42196 334388
rect 42260 334324 42261 334388
rect 42195 334323 42261 334324
rect 41827 324732 41893 324733
rect 41827 324668 41828 324732
rect 41892 324668 41893 324732
rect 41827 324667 41893 324668
rect 41646 315990 41890 316050
rect 41830 315621 41890 315990
rect 41827 315620 41893 315621
rect 41827 315556 41828 315620
rect 41892 315556 41893 315620
rect 41827 315555 41893 315556
rect 42934 312765 42994 337587
rect 43115 336836 43181 336837
rect 43115 336772 43116 336836
rect 43180 336772 43181 336836
rect 43115 336771 43181 336772
rect 43118 316437 43178 336771
rect 43299 336156 43365 336157
rect 43299 336092 43300 336156
rect 43364 336092 43365 336156
rect 43299 336091 43365 336092
rect 43302 334661 43362 336091
rect 43299 334660 43365 334661
rect 43299 334596 43300 334660
rect 43364 334596 43365 334660
rect 43299 334595 43365 334596
rect 43115 316436 43181 316437
rect 43115 316372 43116 316436
rect 43180 316372 43181 316436
rect 43115 316371 43181 316372
rect 42931 312764 42997 312765
rect 42931 312700 42932 312764
rect 42996 312700 42997 312764
rect 42931 312699 42997 312700
rect 41459 312628 41525 312629
rect 41459 312564 41460 312628
rect 41524 312564 41525 312628
rect 41459 312563 41525 312564
rect 43670 297669 43730 340443
rect 44222 311813 44282 342350
rect 44403 342140 44469 342141
rect 44403 342076 44404 342140
rect 44468 342076 44469 342140
rect 44403 342075 44469 342076
rect 44219 311812 44285 311813
rect 44219 311748 44220 311812
rect 44284 311748 44285 311812
rect 44219 311747 44285 311748
rect 44406 311541 44466 342075
rect 44587 341324 44653 341325
rect 44587 341260 44588 341324
rect 44652 341260 44653 341324
rect 44587 341259 44653 341260
rect 44403 311540 44469 311541
rect 44403 311476 44404 311540
rect 44468 311476 44469 311540
rect 44403 311475 44469 311476
rect 44590 311269 44650 341259
rect 675342 339013 675402 354179
rect 675707 353020 675773 353021
rect 675707 352956 675708 353020
rect 675772 352956 675773 353020
rect 675707 352955 675773 352956
rect 675710 350550 675770 352955
rect 675891 351796 675957 351797
rect 675891 351732 675892 351796
rect 675956 351732 675957 351796
rect 675891 351731 675957 351732
rect 675894 351250 675954 351731
rect 675894 351190 676690 351250
rect 675891 350980 675957 350981
rect 675891 350916 675892 350980
rect 675956 350916 675957 350980
rect 675891 350915 675957 350916
rect 675526 350490 675770 350550
rect 675894 350570 675954 350915
rect 675894 350510 676506 350570
rect 675339 339012 675405 339013
rect 675339 338948 675340 339012
rect 675404 338948 675405 339012
rect 675339 338947 675405 338948
rect 675526 337789 675586 350490
rect 675891 350164 675957 350165
rect 675891 350100 675892 350164
rect 675956 350100 675957 350164
rect 675891 350099 675957 350100
rect 675894 349890 675954 350099
rect 675894 349830 676322 349890
rect 675891 349212 675957 349213
rect 675891 349148 675892 349212
rect 675956 349210 675957 349212
rect 675956 349150 676138 349210
rect 675956 349148 675957 349150
rect 675891 349147 675957 349148
rect 675523 337788 675589 337789
rect 675523 337724 675524 337788
rect 675588 337724 675589 337788
rect 675523 337723 675589 337724
rect 676078 328405 676138 349150
rect 676262 332213 676322 349830
rect 676446 336701 676506 350510
rect 676630 340373 676690 351190
rect 676627 340372 676693 340373
rect 676627 340308 676628 340372
rect 676692 340308 676693 340372
rect 676627 340307 676693 340308
rect 676443 336700 676509 336701
rect 676443 336636 676444 336700
rect 676508 336636 676509 336700
rect 676443 336635 676509 336636
rect 676259 332212 676325 332213
rect 676259 332148 676260 332212
rect 676324 332148 676325 332212
rect 676259 332147 676325 332148
rect 676075 328404 676141 328405
rect 676075 328340 676076 328404
rect 676140 328340 676141 328404
rect 676075 328339 676141 328340
rect 44587 311268 44653 311269
rect 44587 311204 44588 311268
rect 44652 311204 44653 311268
rect 44587 311203 44653 311204
rect 675707 308820 675773 308821
rect 675707 308756 675708 308820
rect 675772 308756 675773 308820
rect 675707 308755 675773 308756
rect 675155 308004 675221 308005
rect 675155 307940 675156 308004
rect 675220 307940 675221 308004
rect 675155 307939 675221 307940
rect 675158 301749 675218 307939
rect 675710 303650 675770 308755
rect 675891 306780 675957 306781
rect 675891 306716 675892 306780
rect 675956 306716 675957 306780
rect 675891 306715 675957 306716
rect 675894 305010 675954 306715
rect 675894 304950 676322 305010
rect 675710 303590 676138 303650
rect 675891 302700 675957 302701
rect 675891 302636 675892 302700
rect 675956 302636 675957 302700
rect 675891 302635 675957 302636
rect 675155 301748 675221 301749
rect 675155 301684 675156 301748
rect 675220 301684 675221 301748
rect 675155 301683 675221 301684
rect 43667 297668 43733 297669
rect 43667 297604 43668 297668
rect 43732 297604 43733 297668
rect 43667 297603 43733 297604
rect 675707 297396 675773 297397
rect 675707 297332 675708 297396
rect 675772 297332 675773 297396
rect 675707 297331 675773 297332
rect 42011 296444 42077 296445
rect 42011 296380 42012 296444
rect 42076 296380 42077 296444
rect 42011 296379 42077 296380
rect 41827 295628 41893 295629
rect 41827 295564 41828 295628
rect 41892 295564 41893 295628
rect 41827 295563 41893 295564
rect 41830 294130 41890 295563
rect 40910 294070 41890 294130
rect 40539 292592 40605 292593
rect 40539 292528 40540 292592
rect 40604 292528 40605 292592
rect 40539 292527 40605 292528
rect 40723 292592 40789 292593
rect 40723 292528 40724 292592
rect 40788 292528 40789 292592
rect 40723 292527 40789 292528
rect 40542 274277 40602 292527
rect 40726 277949 40786 292527
rect 40723 277948 40789 277949
rect 40723 277884 40724 277948
rect 40788 277884 40789 277948
rect 40723 277883 40789 277884
rect 40910 277677 40970 294070
rect 41827 292772 41893 292773
rect 41827 292770 41828 292772
rect 41784 292708 41828 292770
rect 41892 292708 41893 292772
rect 41784 292707 41893 292708
rect 41784 292590 41844 292707
rect 41462 292530 41844 292590
rect 40907 277676 40973 277677
rect 40907 277612 40908 277676
rect 40972 277612 40973 277676
rect 40907 277611 40973 277612
rect 40539 274276 40605 274277
rect 40539 274212 40540 274276
rect 40604 274212 40605 274276
rect 40539 274211 40605 274212
rect 41462 270469 41522 292530
rect 41827 292364 41893 292365
rect 41827 292300 41828 292364
rect 41892 292300 41893 292364
rect 41827 292299 41893 292300
rect 41830 289830 41890 292299
rect 41646 289770 41890 289830
rect 41646 287070 41706 289770
rect 41646 287010 41890 287070
rect 41459 270468 41525 270469
rect 41459 270404 41460 270468
rect 41524 270404 41525 270468
rect 41459 270403 41525 270404
rect 41830 269109 41890 287010
rect 42014 281485 42074 296379
rect 675710 281621 675770 297331
rect 675894 282845 675954 302635
rect 676078 283661 676138 303590
rect 676262 295221 676322 304950
rect 676627 301612 676693 301613
rect 676627 301548 676628 301612
rect 676692 301548 676693 301612
rect 676627 301547 676693 301548
rect 676443 301476 676509 301477
rect 676443 301412 676444 301476
rect 676508 301412 676509 301476
rect 676443 301411 676509 301412
rect 676259 295220 676325 295221
rect 676259 295156 676260 295220
rect 676324 295156 676325 295220
rect 676259 295155 676325 295156
rect 676446 291549 676506 301411
rect 676443 291548 676509 291549
rect 676443 291484 676444 291548
rect 676508 291484 676509 291548
rect 676443 291483 676509 291484
rect 676630 287061 676690 301547
rect 676627 287060 676693 287061
rect 676627 286996 676628 287060
rect 676692 286996 676693 287060
rect 676627 286995 676693 286996
rect 676075 283660 676141 283661
rect 676075 283596 676076 283660
rect 676140 283596 676141 283660
rect 676075 283595 676141 283596
rect 675891 282844 675957 282845
rect 675891 282780 675892 282844
rect 675956 282780 675957 282844
rect 675891 282779 675957 282780
rect 675707 281620 675773 281621
rect 675707 281556 675708 281620
rect 675772 281556 675773 281620
rect 675707 281555 675773 281556
rect 42011 281484 42077 281485
rect 42011 281420 42012 281484
rect 42076 281420 42077 281484
rect 42011 281419 42077 281420
rect 41827 269108 41893 269109
rect 41827 269044 41828 269108
rect 41892 269044 41893 269108
rect 41827 269043 41893 269044
rect 674971 263668 675037 263669
rect 674971 263604 674972 263668
rect 675036 263604 675037 263668
rect 674971 263603 675037 263604
rect 674974 258090 675034 263603
rect 676075 262444 676141 262445
rect 676075 262380 676076 262444
rect 676140 262380 676141 262444
rect 676075 262379 676141 262380
rect 674790 258030 675034 258090
rect 40539 251428 40605 251429
rect 40539 251364 40540 251428
rect 40604 251364 40605 251428
rect 40539 251363 40605 251364
rect 40542 240141 40602 251363
rect 40723 249796 40789 249797
rect 40723 249732 40724 249796
rect 40788 249732 40789 249796
rect 40723 249731 40789 249732
rect 40539 240140 40605 240141
rect 40539 240076 40540 240140
rect 40604 240076 40605 240140
rect 40539 240075 40605 240076
rect 40726 235925 40786 249731
rect 674790 249661 674850 258030
rect 676078 249661 676138 262379
rect 676995 261628 677061 261629
rect 676995 261564 676996 261628
rect 677060 261564 677061 261628
rect 676995 261563 677061 261564
rect 676811 259996 676877 259997
rect 676811 259932 676812 259996
rect 676876 259932 676877 259996
rect 676811 259931 676877 259932
rect 674787 249660 674853 249661
rect 674787 249596 674788 249660
rect 674852 249596 674853 249660
rect 674787 249595 674853 249596
rect 676075 249660 676141 249661
rect 676075 249596 676076 249660
rect 676140 249596 676141 249660
rect 676075 249595 676141 249596
rect 676814 245309 676874 259931
rect 676998 250341 677058 261563
rect 676995 250340 677061 250341
rect 676995 250276 676996 250340
rect 677060 250276 677061 250340
rect 676995 250275 677061 250276
rect 676811 245308 676877 245309
rect 676811 245244 676812 245308
rect 676876 245244 676877 245308
rect 676811 245243 676877 245244
rect 675155 245036 675221 245037
rect 675155 244972 675156 245036
rect 675220 244972 675221 245036
rect 675155 244971 675221 244972
rect 675158 240277 675218 244971
rect 675339 244764 675405 244765
rect 675339 244700 675340 244764
rect 675404 244700 675405 244764
rect 675339 244699 675405 244700
rect 675155 240276 675221 240277
rect 675155 240212 675156 240276
rect 675220 240212 675221 240276
rect 675155 240211 675221 240212
rect 42011 237420 42077 237421
rect 42011 237356 42012 237420
rect 42076 237356 42077 237420
rect 42011 237355 42077 237356
rect 40723 235924 40789 235925
rect 40723 235860 40724 235924
rect 40788 235860 40789 235924
rect 40723 235859 40789 235860
rect 42014 227357 42074 237355
rect 674235 237148 674301 237149
rect 674235 237084 674236 237148
rect 674300 237084 674301 237148
rect 674235 237083 674301 237084
rect 672395 231572 672461 231573
rect 672395 231508 672396 231572
rect 672460 231508 672461 231572
rect 672395 231507 672461 231508
rect 672398 230621 672458 231507
rect 672395 230620 672461 230621
rect 672395 230556 672396 230620
rect 672460 230556 672461 230620
rect 672395 230555 672461 230556
rect 667979 229532 668045 229533
rect 667979 229468 667980 229532
rect 668044 229468 668045 229532
rect 667979 229467 668045 229468
rect 42011 227356 42077 227357
rect 42011 227292 42012 227356
rect 42076 227292 42077 227356
rect 42011 227291 42077 227292
rect 572483 222596 572549 222597
rect 572483 222532 572484 222596
rect 572548 222532 572549 222596
rect 572483 222531 572549 222532
rect 561259 222324 561325 222325
rect 561259 222260 561260 222324
rect 561324 222260 561325 222324
rect 561259 222259 561325 222260
rect 561262 222050 561322 222259
rect 561446 222150 563162 222210
rect 561446 222050 561506 222150
rect 563102 222053 563162 222150
rect 561262 221990 561506 222050
rect 562915 222052 562981 222053
rect 562915 221988 562916 222052
rect 562980 221988 562981 222052
rect 562915 221987 562981 221988
rect 563099 222052 563165 222053
rect 563099 221988 563100 222052
rect 563164 221988 563165 222052
rect 563651 222052 563717 222053
rect 563651 222050 563652 222052
rect 563099 221987 563165 221988
rect 563286 221990 563652 222050
rect 545067 220556 545133 220557
rect 545067 220492 545068 220556
rect 545132 220492 545133 220556
rect 545067 220491 545133 220492
rect 553899 220556 553965 220557
rect 553899 220492 553900 220556
rect 553964 220492 553965 220556
rect 553899 220491 553965 220492
rect 543779 220284 543845 220285
rect 543779 220220 543780 220284
rect 543844 220220 543845 220284
rect 543779 220219 543845 220220
rect 511027 220012 511093 220013
rect 511027 219948 511028 220012
rect 511092 219948 511093 220012
rect 511027 219947 511093 219948
rect 529979 220012 530045 220013
rect 529979 219948 529980 220012
rect 530044 219948 530045 220012
rect 529979 219947 530045 219948
rect 530347 220012 530413 220013
rect 530347 219948 530348 220012
rect 530412 219948 530413 220012
rect 530347 219947 530413 219948
rect 500723 217564 500789 217565
rect 500723 217500 500724 217564
rect 500788 217500 500789 217564
rect 500723 217499 500789 217500
rect 504771 217564 504837 217565
rect 504771 217500 504772 217564
rect 504836 217500 504837 217564
rect 504771 217499 504837 217500
rect 500726 217021 500786 217499
rect 500723 217020 500789 217021
rect 500723 216956 500724 217020
rect 500788 216956 500789 217020
rect 500723 216955 500789 216956
rect 504774 216205 504834 217499
rect 511030 216477 511090 219947
rect 519859 219740 519925 219741
rect 519859 219676 519860 219740
rect 519924 219676 519925 219740
rect 519859 219675 519925 219676
rect 522619 219740 522685 219741
rect 522619 219676 522620 219740
rect 522684 219676 522685 219740
rect 522619 219675 522685 219676
rect 514707 219196 514773 219197
rect 514707 219132 514708 219196
rect 514772 219132 514773 219196
rect 514707 219131 514773 219132
rect 514710 218650 514770 219131
rect 514342 218590 514770 218650
rect 514342 218381 514402 218590
rect 514339 218380 514405 218381
rect 514339 218316 514340 218380
rect 514404 218316 514405 218380
rect 514339 218315 514405 218316
rect 519862 216477 519922 219675
rect 511027 216476 511093 216477
rect 511027 216412 511028 216476
rect 511092 216412 511093 216476
rect 511027 216411 511093 216412
rect 519307 216476 519373 216477
rect 519307 216412 519308 216476
rect 519372 216412 519373 216476
rect 519307 216411 519373 216412
rect 519859 216476 519925 216477
rect 519859 216412 519860 216476
rect 519924 216412 519925 216476
rect 519859 216411 519925 216412
rect 504771 216204 504837 216205
rect 504771 216140 504772 216204
rect 504836 216140 504837 216204
rect 504771 216139 504837 216140
rect 519310 215933 519370 216411
rect 519307 215932 519373 215933
rect 519307 215868 519308 215932
rect 519372 215868 519373 215932
rect 519307 215867 519373 215868
rect 522622 215389 522682 219675
rect 529243 215932 529309 215933
rect 529243 215868 529244 215932
rect 529308 215868 529309 215932
rect 529243 215867 529309 215868
rect 529246 215389 529306 215867
rect 522619 215388 522685 215389
rect 522619 215324 522620 215388
rect 522684 215324 522685 215388
rect 522619 215323 522685 215324
rect 529243 215388 529309 215389
rect 529243 215324 529244 215388
rect 529308 215324 529309 215388
rect 529243 215323 529309 215324
rect 529982 215117 530042 219947
rect 530350 215933 530410 219947
rect 543782 218381 543842 220219
rect 543779 218380 543845 218381
rect 543779 218316 543780 218380
rect 543844 218316 543845 218380
rect 543779 218315 543845 218316
rect 545070 218058 545130 220491
rect 553163 219196 553229 219197
rect 553163 219132 553164 219196
rect 553228 219132 553229 219196
rect 553163 219131 553229 219132
rect 553531 219196 553597 219197
rect 553531 219132 553532 219196
rect 553596 219132 553597 219196
rect 553531 219131 553597 219132
rect 553166 218738 553226 219131
rect 553534 218738 553594 219131
rect 553902 218381 553962 220491
rect 556475 220284 556541 220285
rect 556475 220220 556476 220284
rect 556540 220220 556541 220284
rect 562918 220282 562978 221987
rect 563286 220557 563346 221990
rect 563651 221988 563652 221990
rect 563716 221988 563717 222052
rect 563651 221987 563717 221988
rect 572115 222052 572181 222053
rect 572115 221988 572116 222052
rect 572180 221988 572181 222052
rect 572115 221987 572181 221988
rect 563283 220556 563349 220557
rect 563283 220492 563284 220556
rect 563348 220492 563349 220556
rect 563283 220491 563349 220492
rect 563470 220494 564082 220554
rect 563470 220282 563530 220494
rect 562918 220222 563530 220282
rect 563835 220284 563901 220285
rect 556475 220219 556541 220220
rect 563835 220220 563836 220284
rect 563900 220220 563901 220284
rect 563835 220219 563901 220220
rect 556478 219418 556538 220219
rect 553899 218380 553965 218381
rect 553899 218316 553900 218380
rect 553964 218316 553965 218380
rect 553899 218315 553965 218316
rect 554083 218380 554149 218381
rect 554083 218316 554084 218380
rect 554148 218316 554149 218380
rect 554083 218315 554149 218316
rect 554086 218058 554146 218315
rect 563838 217837 563898 220219
rect 564022 217837 564082 220494
rect 567883 219196 567949 219197
rect 567883 219132 567884 219196
rect 567948 219132 567949 219196
rect 567883 219131 567949 219132
rect 567886 218381 567946 219131
rect 572118 218381 572178 221987
rect 567883 218380 567949 218381
rect 567883 218316 567884 218380
rect 567948 218316 567949 218380
rect 567883 218315 567949 218316
rect 572115 218380 572181 218381
rect 572115 218316 572116 218380
rect 572180 218316 572181 218380
rect 572115 218315 572181 218316
rect 563835 217836 563901 217837
rect 563835 217772 563836 217836
rect 563900 217772 563901 217836
rect 563835 217771 563901 217772
rect 564019 217836 564085 217837
rect 564019 217772 564020 217836
rect 564084 217772 564085 217836
rect 564019 217771 564085 217772
rect 572115 217836 572181 217837
rect 572115 217772 572116 217836
rect 572180 217772 572181 217836
rect 572115 217771 572181 217772
rect 541755 217292 541821 217293
rect 541755 217228 541756 217292
rect 541820 217290 541821 217292
rect 544147 217292 544213 217293
rect 544147 217290 544148 217292
rect 541820 217230 544148 217290
rect 541820 217228 541821 217230
rect 541755 217227 541821 217228
rect 544147 217228 544148 217230
rect 544212 217228 544213 217292
rect 544147 217227 544213 217228
rect 566598 217230 568314 217290
rect 536974 216550 537770 216610
rect 530347 215932 530413 215933
rect 530347 215868 530348 215932
rect 530412 215868 530413 215932
rect 530347 215867 530413 215868
rect 536974 215389 537034 216550
rect 537710 215930 537770 216550
rect 546910 216550 547706 216610
rect 546910 215933 546970 216550
rect 546907 215932 546973 215933
rect 537710 215870 538690 215930
rect 538630 215389 538690 215870
rect 546907 215868 546908 215932
rect 546972 215868 546973 215932
rect 547646 215930 547706 216550
rect 556478 216550 557642 216610
rect 548563 215932 548629 215933
rect 548563 215930 548564 215932
rect 547646 215870 548564 215930
rect 546907 215867 546973 215868
rect 548563 215868 548564 215870
rect 548628 215868 548629 215932
rect 548563 215867 548629 215868
rect 556478 215661 556538 216550
rect 556475 215660 556541 215661
rect 556475 215596 556476 215660
rect 556540 215596 556541 215660
rect 557582 215658 557642 216550
rect 566598 216477 566658 217230
rect 566595 216476 566661 216477
rect 566595 216412 566596 216476
rect 566660 216412 566661 216476
rect 566595 216411 566661 216412
rect 566779 216476 566845 216477
rect 566779 216412 566780 216476
rect 566844 216412 566845 216476
rect 566779 216411 566845 216412
rect 558315 215660 558381 215661
rect 558315 215658 558316 215660
rect 557582 215598 558316 215658
rect 556475 215595 556541 215596
rect 558315 215596 558316 215598
rect 558380 215596 558381 215660
rect 558315 215595 558381 215596
rect 566782 215389 566842 216411
rect 536971 215388 537037 215389
rect 536971 215324 536972 215388
rect 537036 215324 537037 215388
rect 536971 215323 537037 215324
rect 538627 215388 538693 215389
rect 538627 215324 538628 215388
rect 538692 215324 538693 215388
rect 538627 215323 538693 215324
rect 566779 215388 566845 215389
rect 566779 215324 566780 215388
rect 566844 215324 566845 215388
rect 566779 215323 566845 215324
rect 568254 215117 568314 217230
rect 572118 216477 572178 217771
rect 572486 216477 572546 222531
rect 573219 220284 573285 220285
rect 573219 220220 573220 220284
rect 573284 220220 573285 220284
rect 573219 220219 573285 220220
rect 573222 218058 573282 220219
rect 572115 216476 572181 216477
rect 572115 216412 572116 216476
rect 572180 216412 572181 216476
rect 572115 216411 572181 216412
rect 572483 216476 572549 216477
rect 572483 216412 572484 216476
rect 572548 216412 572549 216476
rect 572483 216411 572549 216412
rect 575430 215930 575490 217142
rect 582603 217020 582669 217021
rect 582603 217018 582604 217020
rect 582422 216958 582604 217018
rect 577635 216476 577701 216477
rect 577635 216412 577636 216476
rect 577700 216412 577701 216476
rect 577635 216411 577701 216412
rect 577083 215932 577149 215933
rect 575430 215870 575674 215930
rect 529979 215116 530045 215117
rect 529979 215052 529980 215116
rect 530044 215052 530045 215116
rect 529979 215051 530045 215052
rect 568251 215116 568317 215117
rect 568251 215052 568252 215116
rect 568316 215052 568317 215116
rect 568251 215051 568317 215052
rect 575614 213621 575674 215870
rect 577083 215868 577084 215932
rect 577148 215930 577149 215932
rect 577638 215930 577698 216411
rect 582422 216205 582482 216958
rect 582603 216956 582604 216958
rect 582668 216956 582669 217020
rect 582603 216955 582669 216956
rect 591619 217020 591685 217021
rect 591619 216956 591620 217020
rect 591684 216956 591685 217020
rect 591619 216955 591685 216956
rect 592171 217020 592237 217021
rect 592171 216956 592172 217020
rect 592236 216956 592237 217020
rect 592171 216955 592237 216956
rect 591622 216610 591682 216955
rect 592174 216610 592234 216955
rect 591622 216550 592234 216610
rect 582419 216204 582485 216205
rect 582419 216140 582420 216204
rect 582484 216140 582485 216204
rect 582419 216139 582485 216140
rect 577148 215870 577698 215930
rect 577148 215868 577149 215870
rect 577083 215867 577149 215868
rect 666323 215660 666389 215661
rect 666323 215596 666324 215660
rect 666388 215596 666389 215660
rect 666323 215595 666389 215596
rect 575611 213620 575677 213621
rect 575611 213556 575612 213620
rect 575676 213556 575677 213620
rect 575611 213555 575677 213556
rect 41459 209812 41525 209813
rect 41459 209748 41460 209812
rect 41524 209748 41525 209812
rect 41459 209747 41525 209748
rect 666326 209790 666386 215595
rect 40539 208180 40605 208181
rect 40539 208116 40540 208180
rect 40604 208116 40605 208180
rect 40539 208115 40605 208116
rect 40542 197165 40602 208115
rect 40907 207364 40973 207365
rect 40907 207300 40908 207364
rect 40972 207300 40973 207364
rect 40907 207299 40973 207300
rect 40723 206956 40789 206957
rect 40723 206892 40724 206956
rect 40788 206892 40789 206956
rect 40723 206891 40789 206892
rect 40539 197164 40605 197165
rect 40539 197100 40540 197164
rect 40604 197100 40605 197164
rect 40539 197099 40605 197100
rect 40726 194581 40786 206891
rect 40910 194989 40970 207299
rect 41462 195261 41522 209747
rect 666326 209730 666570 209790
rect 42379 207772 42445 207773
rect 42379 207708 42380 207772
rect 42444 207708 42445 207772
rect 42379 207707 42445 207708
rect 41827 197844 41893 197845
rect 41827 197780 41828 197844
rect 41892 197780 41893 197844
rect 41827 197779 41893 197780
rect 41830 195805 41890 197779
rect 41827 195804 41893 195805
rect 41827 195740 41828 195804
rect 41892 195740 41893 195804
rect 41827 195739 41893 195740
rect 41459 195260 41525 195261
rect 41459 195196 41460 195260
rect 41524 195196 41525 195260
rect 41459 195195 41525 195196
rect 40907 194988 40973 194989
rect 40907 194924 40908 194988
rect 40972 194924 40973 194988
rect 40907 194923 40973 194924
rect 40723 194580 40789 194581
rect 40723 194516 40724 194580
rect 40788 194516 40789 194580
rect 40723 194515 40789 194516
rect 41643 194580 41709 194581
rect 41643 194516 41644 194580
rect 41708 194516 41709 194580
rect 41643 194515 41709 194516
rect 41646 190470 41706 194515
rect 42195 193220 42261 193221
rect 42195 193156 42196 193220
rect 42260 193156 42261 193220
rect 42195 193155 42261 193156
rect 41646 190410 41890 190470
rect 41830 187237 41890 190410
rect 41827 187236 41893 187237
rect 41827 187172 41828 187236
rect 41892 187172 41893 187236
rect 41827 187171 41893 187172
rect 42198 186013 42258 193155
rect 42382 186285 42442 207707
rect 666510 197981 666570 209730
rect 666507 197980 666573 197981
rect 666507 197916 666508 197980
rect 666572 197916 666573 197980
rect 666507 197915 666573 197916
rect 42379 186284 42445 186285
rect 42379 186220 42380 186284
rect 42444 186220 42445 186284
rect 42379 186219 42445 186220
rect 42195 186012 42261 186013
rect 42195 185948 42196 186012
rect 42260 185948 42261 186012
rect 42195 185947 42261 185948
rect 667982 130661 668042 229467
rect 673131 228852 673197 228853
rect 673131 228788 673132 228852
rect 673196 228788 673197 228852
rect 673131 228787 673197 228788
rect 672947 228580 673013 228581
rect 672947 228516 672948 228580
rect 673012 228516 673013 228580
rect 672947 228515 673013 228516
rect 672395 227084 672461 227085
rect 672395 227020 672396 227084
rect 672460 227020 672461 227084
rect 672395 227019 672461 227020
rect 672763 227084 672829 227085
rect 672763 227020 672764 227084
rect 672828 227020 672829 227084
rect 672763 227019 672829 227020
rect 672027 225724 672093 225725
rect 672027 225660 672028 225724
rect 672092 225660 672093 225724
rect 672027 225659 672093 225660
rect 672030 223005 672090 225659
rect 672027 223004 672093 223005
rect 672027 222940 672028 223004
rect 672092 222940 672093 223004
rect 672027 222939 672093 222940
rect 672398 222210 672458 227019
rect 672766 224365 672826 227019
rect 672763 224364 672829 224365
rect 672763 224300 672764 224364
rect 672828 224300 672829 224364
rect 672763 224299 672829 224300
rect 672214 222150 672458 222210
rect 670739 220148 670805 220149
rect 670739 220084 670740 220148
rect 670804 220084 670805 220148
rect 670739 220083 670805 220084
rect 669451 211172 669517 211173
rect 669451 211108 669452 211172
rect 669516 211108 669517 211172
rect 669451 211107 669517 211108
rect 669454 195990 669514 211107
rect 669270 195930 669514 195990
rect 669270 176670 669330 195930
rect 669270 176610 669514 176670
rect 669454 147690 669514 176610
rect 669270 147630 669514 147690
rect 669270 143717 669330 147630
rect 669267 143716 669333 143717
rect 669267 143652 669268 143716
rect 669332 143652 669333 143716
rect 669267 143651 669333 143652
rect 670742 133789 670802 220083
rect 672214 217565 672274 222150
rect 672211 217564 672277 217565
rect 672211 217500 672212 217564
rect 672276 217500 672277 217564
rect 672211 217499 672277 217500
rect 672950 183565 673010 228515
rect 673134 224637 673194 228787
rect 673499 225044 673565 225045
rect 673499 224980 673500 225044
rect 673564 224980 673565 225044
rect 673499 224979 673565 224980
rect 673131 224636 673197 224637
rect 673131 224572 673132 224636
rect 673196 224572 673197 224636
rect 673131 224571 673197 224572
rect 673131 214844 673197 214845
rect 673131 214780 673132 214844
rect 673196 214780 673197 214844
rect 673131 214779 673197 214780
rect 672947 183564 673013 183565
rect 672947 183500 672948 183564
rect 673012 183500 673013 183564
rect 672947 183499 673013 183500
rect 673134 182069 673194 214779
rect 673315 201652 673381 201653
rect 673315 201588 673316 201652
rect 673380 201588 673381 201652
rect 673315 201587 673381 201588
rect 673131 182068 673197 182069
rect 673131 182004 673132 182068
rect 673196 182004 673197 182068
rect 673131 182003 673197 182004
rect 673318 149157 673378 201587
rect 673315 149156 673381 149157
rect 673315 149092 673316 149156
rect 673380 149092 673381 149156
rect 673315 149091 673381 149092
rect 670739 133788 670805 133789
rect 670739 133724 670740 133788
rect 670804 133724 670805 133788
rect 670739 133723 670805 133724
rect 667979 130660 668045 130661
rect 667979 130596 667980 130660
rect 668044 130596 668045 130660
rect 667979 130595 668045 130596
rect 673502 128893 673562 224979
rect 674051 212124 674117 212125
rect 674051 212060 674052 212124
rect 674116 212060 674117 212124
rect 674051 212059 674117 212060
rect 673499 128892 673565 128893
rect 673499 128828 673500 128892
rect 673564 128828 673565 128892
rect 673499 128827 673565 128828
rect 674054 128349 674114 212059
rect 674238 155005 674298 237083
rect 675342 236877 675402 244699
rect 675339 236876 675405 236877
rect 675339 236812 675340 236876
rect 675404 236812 675405 236876
rect 675339 236811 675405 236812
rect 674419 230212 674485 230213
rect 674419 230148 674420 230212
rect 674484 230148 674485 230212
rect 674419 230147 674485 230148
rect 674422 225045 674482 230147
rect 675155 228580 675221 228581
rect 675155 228516 675156 228580
rect 675220 228516 675221 228580
rect 675155 228515 675221 228516
rect 674419 225044 674485 225045
rect 674419 224980 674420 225044
rect 674484 224980 674485 225044
rect 674419 224979 674485 224980
rect 674603 220420 674669 220421
rect 674603 220356 674604 220420
rect 674668 220356 674669 220420
rect 674603 220355 674669 220356
rect 674606 219197 674666 220355
rect 674787 220148 674853 220149
rect 674787 220084 674788 220148
rect 674852 220084 674853 220148
rect 674787 220083 674853 220084
rect 674603 219196 674669 219197
rect 674603 219132 674604 219196
rect 674668 219132 674669 219196
rect 674603 219131 674669 219132
rect 674790 215389 674850 220083
rect 674971 218652 675037 218653
rect 674971 218588 674972 218652
rect 675036 218588 675037 218652
rect 674971 218587 675037 218588
rect 674787 215388 674853 215389
rect 674787 215324 674788 215388
rect 674852 215324 674853 215388
rect 674787 215323 674853 215324
rect 674974 210493 675034 218587
rect 675158 217293 675218 228515
rect 675339 225996 675405 225997
rect 675339 225932 675340 225996
rect 675404 225932 675405 225996
rect 675339 225931 675405 225932
rect 675155 217292 675221 217293
rect 675155 217228 675156 217292
rect 675220 217228 675221 217292
rect 675155 217227 675221 217228
rect 675342 215933 675402 225931
rect 675891 218244 675957 218245
rect 675891 218180 675892 218244
rect 675956 218180 675957 218244
rect 675891 218179 675957 218180
rect 675523 217428 675589 217429
rect 675523 217364 675524 217428
rect 675588 217364 675589 217428
rect 675523 217363 675589 217364
rect 675339 215932 675405 215933
rect 675339 215868 675340 215932
rect 675404 215868 675405 215932
rect 675339 215867 675405 215868
rect 674971 210492 675037 210493
rect 674971 210428 674972 210492
rect 675036 210428 675037 210492
rect 674971 210427 675037 210428
rect 675526 198253 675586 217363
rect 675707 217020 675773 217021
rect 675707 216956 675708 217020
rect 675772 216956 675773 217020
rect 675707 216955 675773 216956
rect 675710 211170 675770 216955
rect 675894 215310 675954 218179
rect 675894 215250 676690 215310
rect 676259 215150 676325 215151
rect 676259 215086 676260 215150
rect 676324 215086 676325 215150
rect 676259 215085 676325 215086
rect 675891 214572 675957 214573
rect 675891 214508 675892 214572
rect 675956 214508 675957 214572
rect 675891 214507 675957 214508
rect 675894 211445 675954 214507
rect 675891 211444 675957 211445
rect 675891 211380 675892 211444
rect 675956 211380 675957 211444
rect 675891 211379 675957 211380
rect 675710 211110 676138 211170
rect 675891 210492 675957 210493
rect 675891 210428 675892 210492
rect 675956 210428 675957 210492
rect 675891 210427 675957 210428
rect 675523 198252 675589 198253
rect 675523 198188 675524 198252
rect 675588 198188 675589 198252
rect 675523 198187 675589 198188
rect 675894 193221 675954 210427
rect 675891 193220 675957 193221
rect 675891 193156 675892 193220
rect 675956 193156 675957 193220
rect 675891 193155 675957 193156
rect 676078 191589 676138 211110
rect 676262 197165 676322 215085
rect 676443 211444 676509 211445
rect 676443 211380 676444 211444
rect 676508 211380 676509 211444
rect 676443 211379 676509 211380
rect 676446 200701 676506 211379
rect 676630 205597 676690 215250
rect 676627 205596 676693 205597
rect 676627 205532 676628 205596
rect 676692 205532 676693 205596
rect 676627 205531 676693 205532
rect 676443 200700 676509 200701
rect 676443 200636 676444 200700
rect 676508 200636 676509 200700
rect 676443 200635 676509 200636
rect 676259 197164 676325 197165
rect 676259 197100 676260 197164
rect 676324 197100 676325 197164
rect 676259 197099 676325 197100
rect 676075 191588 676141 191589
rect 676075 191524 676076 191588
rect 676140 191524 676141 191588
rect 676075 191523 676141 191524
rect 675891 174044 675957 174045
rect 675891 173980 675892 174044
rect 675956 173980 675957 174044
rect 675891 173979 675957 173980
rect 675894 173770 675954 173979
rect 675894 173710 676506 173770
rect 675707 173636 675773 173637
rect 675707 173572 675708 173636
rect 675772 173572 675773 173636
rect 675707 173571 675773 173572
rect 675523 167516 675589 167517
rect 675523 167452 675524 167516
rect 675588 167452 675589 167516
rect 675523 167451 675589 167452
rect 675339 161940 675405 161941
rect 675339 161876 675340 161940
rect 675404 161876 675405 161940
rect 675339 161875 675405 161876
rect 675342 157045 675402 161875
rect 675526 157350 675586 167451
rect 675710 162210 675770 173571
rect 675891 172412 675957 172413
rect 675891 172348 675892 172412
rect 675956 172410 675957 172412
rect 675956 172350 676322 172410
rect 675956 172348 675957 172350
rect 675891 172347 675957 172348
rect 675891 172004 675957 172005
rect 675891 171940 675892 172004
rect 675956 171940 675957 172004
rect 675891 171939 675957 171940
rect 675894 167010 675954 171939
rect 675894 166950 676138 167010
rect 675710 162150 675954 162210
rect 675526 157290 675770 157350
rect 675339 157044 675405 157045
rect 675339 156980 675340 157044
rect 675404 156980 675405 157044
rect 675339 156979 675405 156980
rect 674235 155004 674301 155005
rect 674235 154940 674236 155004
rect 674300 154940 674301 155004
rect 674235 154939 674301 154940
rect 675710 147661 675770 157290
rect 675894 148477 675954 162150
rect 675891 148476 675957 148477
rect 675891 148412 675892 148476
rect 675956 148412 675957 148476
rect 675891 148411 675957 148412
rect 675707 147660 675773 147661
rect 675707 147596 675708 147660
rect 675772 147596 675773 147660
rect 675707 147595 675773 147596
rect 676078 146029 676138 166950
rect 676262 153101 676322 172350
rect 676446 159357 676506 173710
rect 676627 166428 676693 166429
rect 676627 166364 676628 166428
rect 676692 166364 676693 166428
rect 676627 166363 676693 166364
rect 676443 159356 676509 159357
rect 676443 159292 676444 159356
rect 676508 159292 676509 159356
rect 676443 159291 676509 159292
rect 676630 156365 676690 166363
rect 676627 156364 676693 156365
rect 676627 156300 676628 156364
rect 676692 156300 676693 156364
rect 676627 156299 676693 156300
rect 676259 153100 676325 153101
rect 676259 153036 676260 153100
rect 676324 153036 676325 153100
rect 676259 153035 676325 153036
rect 676075 146028 676141 146029
rect 676075 145964 676076 146028
rect 676140 145964 676141 146028
rect 676075 145963 676141 145964
rect 676627 128620 676693 128621
rect 676627 128556 676628 128620
rect 676692 128556 676693 128620
rect 676627 128555 676693 128556
rect 674051 128348 674117 128349
rect 674051 128284 674052 128348
rect 674116 128284 674117 128348
rect 674051 128283 674117 128284
rect 676075 128212 676141 128213
rect 676075 128148 676076 128212
rect 676140 128148 676141 128212
rect 676075 128147 676141 128148
rect 675891 127260 675957 127261
rect 675891 127196 675892 127260
rect 675956 127196 675957 127260
rect 675891 127195 675957 127196
rect 675707 122364 675773 122365
rect 675707 122300 675708 122364
rect 675772 122300 675773 122364
rect 675707 122299 675773 122300
rect 675710 102645 675770 122299
rect 675894 108085 675954 127195
rect 675891 108084 675957 108085
rect 675891 108020 675892 108084
rect 675956 108020 675957 108084
rect 675891 108019 675957 108020
rect 676078 103189 676138 128147
rect 676259 126988 676325 126989
rect 676259 126924 676260 126988
rect 676324 126924 676325 126988
rect 676259 126923 676325 126924
rect 676075 103188 676141 103189
rect 676075 103124 676076 103188
rect 676140 103124 676141 103188
rect 676075 103123 676141 103124
rect 675707 102644 675773 102645
rect 675707 102580 675708 102644
rect 675772 102580 675773 102644
rect 675707 102579 675773 102580
rect 676262 101421 676322 126923
rect 676443 124540 676509 124541
rect 676443 124476 676444 124540
rect 676508 124476 676509 124540
rect 676443 124475 676509 124476
rect 676446 106181 676506 124475
rect 676630 113117 676690 128555
rect 676627 113116 676693 113117
rect 676627 113052 676628 113116
rect 676692 113052 676693 113116
rect 676627 113051 676693 113052
rect 676443 106180 676509 106181
rect 676443 106116 676444 106180
rect 676508 106116 676509 106180
rect 676443 106115 676509 106116
rect 676259 101420 676325 101421
rect 676259 101356 676260 101420
rect 676324 101356 676325 101420
rect 676259 101355 676325 101356
rect 637251 96932 637317 96933
rect 637251 96868 637252 96932
rect 637316 96868 637317 96932
rect 637251 96867 637317 96868
rect 633939 96116 634005 96117
rect 633939 96052 633940 96116
rect 634004 96052 634005 96116
rect 633939 96051 634005 96052
rect 633942 78573 634002 96051
rect 637254 84210 637314 96867
rect 637070 84150 637314 84210
rect 633939 78572 634005 78573
rect 633939 78508 633940 78572
rect 634004 78508 634005 78572
rect 633939 78507 634005 78508
rect 637070 77893 637130 84150
rect 637067 77892 637133 77893
rect 637067 77828 637068 77892
rect 637132 77828 637133 77892
rect 637067 77827 637133 77828
rect 462635 54500 462701 54501
rect 462635 54436 462636 54500
rect 462700 54436 462701 54500
rect 462635 54435 462701 54436
rect 462638 53685 462698 54435
rect 462635 53684 462701 53685
rect 462635 53620 462636 53684
rect 462700 53620 462701 53684
rect 462635 53619 462701 53620
rect 194363 50284 194429 50285
rect 194363 50220 194364 50284
rect 194428 50220 194429 50284
rect 194363 50219 194429 50220
rect 529795 50284 529861 50285
rect 529795 50220 529796 50284
rect 529860 50220 529861 50284
rect 529795 50219 529861 50220
rect 141739 44028 141805 44029
rect 141739 43964 141740 44028
rect 141804 43964 141805 44028
rect 141739 43963 141805 43964
rect 141742 40493 141802 43963
rect 194366 42125 194426 50219
rect 518755 48924 518821 48925
rect 518755 48860 518756 48924
rect 518820 48860 518821 48924
rect 518755 48859 518821 48860
rect 515443 47564 515509 47565
rect 515443 47500 515444 47564
rect 515508 47500 515509 47564
rect 515443 47499 515509 47500
rect 461347 44436 461413 44437
rect 461347 44372 461348 44436
rect 461412 44372 461413 44436
rect 461347 44371 461413 44372
rect 462267 44436 462333 44437
rect 462267 44372 462268 44436
rect 462332 44372 462333 44436
rect 462267 44371 462333 44372
rect 194363 42124 194429 42125
rect 194363 42060 194364 42124
rect 194428 42060 194429 42124
rect 194363 42059 194429 42060
rect 421971 42124 422037 42125
rect 421971 42060 421972 42124
rect 422036 42060 422037 42124
rect 421971 42059 422037 42060
rect 421974 41850 422034 42059
rect 461350 41938 461410 44371
rect 462270 41938 462330 44371
rect 515446 42125 515506 47499
rect 518758 42805 518818 48859
rect 526483 48108 526549 48109
rect 526483 48044 526484 48108
rect 526548 48044 526549 48108
rect 526483 48043 526549 48044
rect 520963 47836 521029 47837
rect 520963 47772 520964 47836
rect 521028 47772 521029 47836
rect 520963 47771 521029 47772
rect 518755 42804 518821 42805
rect 518755 42740 518756 42804
rect 518820 42740 518821 42804
rect 518755 42739 518821 42740
rect 520966 42125 521026 47771
rect 522067 47292 522133 47293
rect 522067 47228 522068 47292
rect 522132 47228 522133 47292
rect 522067 47227 522133 47228
rect 522070 42125 522130 47227
rect 526486 42125 526546 48043
rect 529798 42125 529858 50219
rect 515443 42124 515509 42125
rect 515443 42060 515444 42124
rect 515508 42060 515509 42124
rect 515443 42059 515509 42060
rect 520963 42124 521029 42125
rect 520963 42060 520964 42124
rect 521028 42060 521029 42124
rect 520963 42059 521029 42060
rect 522067 42124 522133 42125
rect 522067 42060 522068 42124
rect 522132 42060 522133 42124
rect 522067 42059 522133 42060
rect 526483 42124 526549 42125
rect 526483 42060 526484 42124
rect 526548 42060 526549 42124
rect 526483 42059 526549 42060
rect 529795 42124 529861 42125
rect 529795 42060 529796 42124
rect 529860 42060 529861 42124
rect 529795 42059 529861 42060
rect 421974 41790 422162 41850
rect 441843 41852 441909 41853
rect 441843 41850 441844 41852
rect 441626 41790 441844 41850
rect 441843 41788 441844 41790
rect 441908 41788 441909 41852
rect 441843 41787 441909 41788
rect 460611 41852 460677 41853
rect 460611 41788 460612 41852
rect 460676 41850 460677 41852
rect 460676 41790 460802 41850
rect 460676 41788 460677 41790
rect 460611 41787 460677 41788
rect 141739 40492 141805 40493
rect 141739 40428 141740 40492
rect 141804 40428 141805 40492
rect 141739 40427 141805 40428
<< via4 >>
rect 511862 997252 512098 997338
rect 511862 997188 511948 997252
rect 511948 997188 512012 997252
rect 512012 997188 512098 997252
rect 511862 997102 512098 997188
rect 522718 997102 522954 997338
rect 523822 997102 524058 997338
rect 531366 997102 531602 997338
rect 536518 997102 536754 997338
rect 569822 997102 570058 997338
rect 493462 217292 493698 217378
rect 493462 217228 493548 217292
rect 493548 217228 493612 217292
rect 493612 217228 493698 217292
rect 493462 217142 493698 217228
rect 553078 218502 553314 218738
rect 553446 218502 553682 218738
rect 556390 219182 556626 219418
rect 544982 217822 545218 218058
rect 553998 217822 554234 218058
rect 573134 217822 573370 218058
rect 575342 217142 575578 217378
rect 419862 41852 420098 41938
rect 419862 41788 419948 41852
rect 419948 41788 420012 41852
rect 420012 41788 420098 41852
rect 419862 41702 420098 41788
rect 422162 41702 422398 41938
rect 441390 41702 441626 41938
rect 460802 41702 461038 41938
rect 461262 41702 461498 41938
rect 462182 41702 462418 41938
<< metal5 >>
rect 78440 1018512 90960 1031002
rect 129840 1018512 142360 1031002
rect 181240 1018512 193760 1031002
rect 232640 1018512 245160 1031002
rect 284240 1018512 296760 1031002
rect 334810 1018624 346978 1030789
rect 386040 1018512 398560 1031002
rect 475040 1018512 487560 1031002
rect 526440 1018512 538960 1031002
rect 577010 1018624 589178 1030789
rect 628240 1018512 640760 1031002
rect 511820 997338 522996 997380
rect 511820 997102 511862 997338
rect 512098 997102 522718 997338
rect 522954 997102 522996 997338
rect 511820 997060 522996 997102
rect 523780 997338 531644 997380
rect 523780 997102 523822 997338
rect 524058 997102 531366 997338
rect 531602 997102 531644 997338
rect 523780 997060 531644 997102
rect 536476 997338 570100 997380
rect 536476 997102 536518 997338
rect 536754 997102 569822 997338
rect 570058 997102 570100 997338
rect 536476 997060 570100 997102
rect 6598 956440 19088 968960
rect 698512 952840 711002 965360
rect 6167 914054 19620 924934
rect 697980 909666 711433 920546
rect 6811 871210 18976 883378
rect 698512 863640 711002 876160
rect 6811 829010 18976 841178
rect 698624 819822 710789 831990
rect 6598 786640 19088 799160
rect 698512 774440 711002 786960
rect 6598 743440 19088 755960
rect 698512 729440 711002 741960
rect 6598 700240 19088 712760
rect 698512 684440 711002 696960
rect 6598 657040 19088 669560
rect 698512 639240 711002 651760
rect 6598 613840 19088 626360
rect 698512 594240 711002 606760
rect 6598 570640 19088 583160
rect 698512 549040 711002 561560
rect 6598 527440 19088 539960
rect 698624 505222 710789 517390
rect 6811 484410 18976 496578
rect 697980 461866 711433 472746
rect 6167 442854 19620 453734
rect 698624 417022 710789 429190
rect 6598 399840 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 698512 326640 711002 339160
rect 6598 313440 19088 325960
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 6598 227040 19088 239560
rect 698512 236640 711002 249160
rect 556348 219418 572860 219460
rect 556348 219182 556390 219418
rect 556626 219182 572860 219418
rect 556348 219140 572860 219182
rect 553036 218738 553724 218780
rect 553036 218502 553078 218738
rect 553314 218502 553446 218738
rect 553682 218502 553724 218738
rect 553036 218460 553724 218502
rect 572540 218100 572860 219140
rect 544940 218058 554276 218100
rect 544940 217822 544982 218058
rect 545218 217822 553998 218058
rect 554234 217822 554276 218058
rect 544940 217780 554276 217822
rect 572540 218058 573412 218100
rect 572540 217822 573134 218058
rect 573370 217822 573412 218058
rect 572540 217780 573412 217822
rect 493420 217378 575620 217420
rect 493420 217142 493462 217378
rect 493698 217142 575342 217378
rect 575578 217142 575620 217378
rect 493420 217100 575620 217142
rect 6598 183840 19088 196360
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 6811 111610 18976 123778
rect 698512 101240 711002 113760
rect 6167 70054 19620 80934
rect 419820 41938 421796 41980
rect 419820 41702 419862 41938
rect 420098 41702 421796 41938
rect 419820 41660 421796 41702
rect 422120 41938 441668 41980
rect 422120 41702 422162 41938
rect 422398 41702 441390 41938
rect 441626 41702 441668 41938
rect 422120 41660 441668 41702
rect 442084 41660 450684 41980
rect 421476 41300 421796 41660
rect 442084 41300 442404 41660
rect 421476 40980 442404 41300
rect 450364 41300 450684 41660
rect 451100 41660 460436 41980
rect 460760 41938 461540 41980
rect 460760 41702 460802 41938
rect 461038 41702 461262 41938
rect 461498 41702 461540 41938
rect 460760 41660 461540 41702
rect 461956 41938 462460 41980
rect 461956 41702 462182 41938
rect 462418 41702 462460 41938
rect 461956 41660 462460 41702
rect 451100 41300 451420 41660
rect 450364 40980 451420 41300
rect 460116 41300 460436 41660
rect 461956 41300 462276 41660
rect 460116 40980 462276 41300
rect 80222 6811 92390 18976
rect 136713 7143 144150 18309
rect 187640 6598 200160 19088
rect 243266 6167 254146 19620
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 570422 6811 582590 18976
rect 624222 6811 636390 18976
use caravel_logo  caravel_logo
timestamp 0
transform 1 0 269370 0 1 5100
box 0 0 1 1
use caravel_motto  caravel_motto
timestamp 0
transform 1 0 -54372 0 1 -4446
box 0 0 1 1
use copyright_block  copyright_block
timestamp 0
transform 1 0 149582 0 1 16298
box 0 0 1 1
use open_source  open_source
timestamp 0
transform 1 0 206098 0 1 2054
box 0 0 1 1
use xres_buf  rstb_level
timestamp 1666117611
transform -1 0 145710 0 -1 50488
box 414 -400 3522 3800
use user_id_textblock  user_id_textblock
timestamp 0
transform 1 0 96272 0 1 6890
box 0 0 1 1
use caravel_clocking  clock_ctrl
timestamp 1666117611
transform 1 0 626764 0 1 55284
box 136 496 20000 20000
use buff_flash_clkrst  flash_clkrst_buffers
timestamp 1666117611
transform 1 0 458400 0 1 47600
box 330 0 7699 5000
use gpio_control_block  gpio_control_bidir_1\[0\]
timestamp 1666117611
transform -1 0 710203 0 1 121000
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_0
timestamp 1666117611
transform -1 0 709467 0 1 134000
box -38 0 6018 2224
use housekeeping  housekeeping
timestamp 1666117611
transform 1 0 592434 0 1 100002
box 0 0 74046 110190
use digital_pll  pll
timestamp 1666117611
transform 1 0 628146 0 1 80944
box 0 0 20000 15000
use simple_por  por
timestamp 1666117611
transform 1 0 650146 0 -1 55282
box -14 11 11344 8684
use user_id_programming  user_id_value
timestamp 1666117611
transform 1 0 656624 0 1 88126
box 0 0 7109 7077
use mgmt_core_wrapper  soc
timestamp 1666117611
transform 1 0 52034 0 1 53002
box -156 0 524096 164000
use gpio_control_block  gpio_control_bidir_1\[1\]
timestamp 1666117611
transform -1 0 710203 0 1 166200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_1
timestamp 1666117611
transform -1 0 709467 0 1 179200
box -38 0 6018 2224
use gpio_control_block  gpio_control_bidir_2\[2\]
timestamp 1666117611
transform 1 0 7631 0 1 202600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[0\]
timestamp 1666117611
transform -1 0 710203 0 1 211200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_2
timestamp 1666117611
transform -1 0 709467 0 1 224200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_37
timestamp 1666117611
transform 1 0 8367 0 1 215600
box -38 0 6018 2224
use spare_logic_block  spare_logic\[2\]
timestamp 1666117611
transform 1 0 640874 0 1 220592
box 0 0 9000 9000
use gpio_control_block  gpio_control_bidir_2\[1\]
timestamp 1666117611
transform 1 0 7631 0 1 245800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[1\]
timestamp 1666117611
transform -1 0 710203 0 1 256400
box 872 416 34000 13000
use mgmt_protect  mgmt_buffers
timestamp 1666117611
transform 1 0 128180 0 1 232036
box 1066 -400 424400 32400
use spare_logic_block  spare_logic\[0\]
timestamp 1666117611
transform 1 0 88632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[1\]
timestamp 1666117611
transform 1 0 108632 0 1 232528
box 0 0 9000 9000
use spare_logic_block  spare_logic\[3\]
timestamp 1666117611
transform 1 0 578632 0 1 232528
box 0 0 9000 9000
use gpio_control_block  gpio_control_bidir_2\[0\]
timestamp 1666117611
transform 1 0 7631 0 1 289000
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_3
timestamp 1666117611
transform -1 0 709467 0 1 269400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_36
timestamp 1666117611
transform 1 0 8367 0 1 258800
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[2\]
timestamp 1666117611
transform -1 0 710203 0 1 301400
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_35
timestamp 1666117611
transform 1 0 8367 0 1 302000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_4
timestamp 1666117611
transform -1 0 709467 0 1 314400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[13\]
timestamp 1666117611
transform 1 0 7631 0 1 418600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[14\]
timestamp 1666117611
transform 1 0 7631 0 1 375400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[15\]
timestamp 1666117611
transform 1 0 7631 0 1 332200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_32
timestamp 1666117611
transform 1 0 8367 0 1 431600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_33
timestamp 1666117611
transform 1 0 8367 0 1 388400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_34
timestamp 1666117611
transform 1 0 8367 0 1 345200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1a\[3\]
timestamp 1666117611
transform -1 0 710203 0 1 346400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[4\]
timestamp 1666117611
transform -1 0 710203 0 1 391600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1a\[5\]
timestamp 1666117611
transform -1 0 710203 0 1 479800
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_5
timestamp 1666117611
transform -1 0 709467 0 1 359400
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_6
timestamp 1666117611
transform -1 0 709467 0 1 404600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_7
timestamp 1666117611
transform -1 0 709467 0 1 492800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_31
timestamp 1666117611
transform 1 0 8367 0 1 559200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_30
timestamp 1666117611
transform 1 0 8367 0 1 602400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[12\]
timestamp 1666117611
transform 1 0 7631 0 1 546200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[11\]
timestamp 1666117611
transform 1 0 7631 0 1 589400
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[1\]
timestamp 1666117611
transform -1 0 710203 0 1 568800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[0\]
timestamp 1666117611
transform -1 0 710203 0 1 523800
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_9
timestamp 1666117611
transform -1 0 709467 0 1 581800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_8
timestamp 1666117611
transform -1 0 709467 0 1 536800
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_29
timestamp 1666117611
transform 1 0 8367 0 1 645600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_28
timestamp 1666117611
transform 1 0 8367 0 1 688800
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[9\]
timestamp 1666117611
transform 1 0 7631 0 1 675800
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[10\]
timestamp 1666117611
transform 1 0 7631 0 1 632600
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[3\]
timestamp 1666117611
transform -1 0 710203 0 1 659000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[2\]
timestamp 1666117611
transform -1 0 710203 0 1 614000
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_11
timestamp 1666117611
transform -1 0 709467 0 1 672000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_10
timestamp 1666117611
transform -1 0 709467 0 1 627000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_27
timestamp 1666117611
transform 1 0 8367 0 1 732000
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_26
timestamp 1666117611
transform 1 0 8367 0 1 775200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[8\]
timestamp 1666117611
transform 1 0 7631 0 1 719000
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[7\]
timestamp 1666117611
transform 1 0 7631 0 1 762200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[5\]
timestamp 1666117611
transform -1 0 710203 0 1 749200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[4\]
timestamp 1666117611
transform -1 0 710203 0 1 704200
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_13
timestamp 1666117611
transform -1 0 709467 0 1 762200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_12
timestamp 1666117611
transform -1 0 709467 0 1 717200
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_25
timestamp 1666117611
transform 1 0 8367 0 1 818400
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[6\]
timestamp 1666117611
transform 1 0 7631 0 1 805400
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_24
timestamp 1666117611
transform 1 0 8367 0 1 944200
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[5\]
timestamp 1666117611
transform 1 0 7631 0 1 931200
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[6\]
timestamp 1666117611
transform -1 0 710203 0 1 927600
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_14
timestamp 1666117611
transform -1 0 709467 0 1 940600
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_23
timestamp 1666117611
transform 0 1 110194 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[4\]
timestamp 1666117611
transform 0 1 97200 -1 0 1030077
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_22
timestamp 1666117611
transform 0 1 161594 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_21
timestamp 1666117611
transform 0 1 212994 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[3\]
timestamp 1666117611
transform 0 1 148600 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[2\]
timestamp 1666117611
transform 0 1 200000 -1 0 1030077
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_20
timestamp 1666117611
transform 0 1 264394 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_2\[1\]
timestamp 1666117611
transform 0 1 251400 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_2\[0\]
timestamp 1666117611
transform 0 1 303000 -1 0 1030077
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_19
timestamp 1666117611
transform 0 1 315994 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_18
timestamp 1666117611
transform 0 1 366394 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[10\]
timestamp 1666117611
transform 0 1 353400 -1 0 1030077
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_17
timestamp 1666117611
transform 0 1 433794 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[9\]
timestamp 1666117611
transform 0 1 420800 -1 0 1030077
box 872 416 34000 13000
use gpio_defaults_block  gpio_defaults_block_16
timestamp 1666117611
transform 0 1 510794 -1 0 1029341
box -38 0 6018 2224
use gpio_defaults_block  gpio_defaults_block_15
timestamp 1666117611
transform 0 1 562194 -1 0 1029341
box -38 0 6018 2224
use gpio_control_block  gpio_control_in_1\[8\]
timestamp 1666117611
transform 0 1 497800 -1 0 1030077
box 872 416 34000 13000
use gpio_control_block  gpio_control_in_1\[7\]
timestamp 1666117611
transform 0 1 549200 -1 0 1030077
box 872 416 34000 13000
use caravel_power_routing  caravel_power_routing
timestamp 1666117611
transform 1 0 0 0 1 0
box 6022 30806 711814 1031696
use user_project_wrapper  mprj
timestamp 1666117611
transform 1 0 65308 0 1 278718
box -8726 -7654 592650 711590
use chip_io  padframe
timestamp 1666117611
transform 1 0 0 0 1 0
box 0 0 717600 1037600
use gpio_signal_buffering  sigbuf
timestamp 1666117611
transform 1 0 0 0 1 0
box 39992 41960 677583 997915
<< labels >>
rlabel metal5 s 187640 6598 200160 19088 6 clock
port 0 nsew signal input
rlabel metal5 s 351040 6598 363560 19088 6 flash_clk
port 1 nsew signal tristate
rlabel metal5 s 296240 6598 308760 19088 6 flash_csb
port 2 nsew signal tristate
rlabel metal5 s 405840 6598 418360 19088 6 flash_io0
port 3 nsew signal tristate
rlabel metal5 s 460640 6598 473160 19088 6 flash_io1
port 4 nsew signal tristate
rlabel metal5 s 515440 6598 527960 19088 6 gpio
port 5 nsew signal bidirectional
rlabel metal5 s 698512 101240 711002 113760 6 mprj_io[0]
port 6 nsew signal bidirectional
rlabel metal5 s 698512 684440 711002 696960 6 mprj_io[10]
port 7 nsew signal bidirectional
rlabel metal5 s 698512 729440 711002 741960 6 mprj_io[11]
port 8 nsew signal bidirectional
rlabel metal5 s 698512 774440 711002 786960 6 mprj_io[12]
port 9 nsew signal bidirectional
rlabel metal5 s 698512 863640 711002 876160 6 mprj_io[13]
port 10 nsew signal bidirectional
rlabel metal5 s 698512 952840 711002 965360 6 mprj_io[14]
port 11 nsew signal bidirectional
rlabel metal5 s 628240 1018512 640760 1031002 6 mprj_io[15]
port 12 nsew signal bidirectional
rlabel metal5 s 526440 1018512 538960 1031002 6 mprj_io[16]
port 13 nsew signal bidirectional
rlabel metal5 s 475040 1018512 487560 1031002 6 mprj_io[17]
port 14 nsew signal bidirectional
rlabel metal5 s 386040 1018512 398560 1031002 6 mprj_io[18]
port 15 nsew signal bidirectional
rlabel metal5 s 284240 1018512 296760 1031002 6 mprj_io[19]
port 16 nsew signal bidirectional
rlabel metal5 s 698512 146440 711002 158960 6 mprj_io[1]
port 17 nsew signal bidirectional
rlabel metal5 s 232640 1018512 245160 1031002 6 mprj_io[20]
port 18 nsew signal bidirectional
rlabel metal5 s 181240 1018512 193760 1031002 6 mprj_io[21]
port 19 nsew signal bidirectional
rlabel metal5 s 129840 1018512 142360 1031002 6 mprj_io[22]
port 20 nsew signal bidirectional
rlabel metal5 s 78440 1018512 90960 1031002 6 mprj_io[23]
port 21 nsew signal bidirectional
rlabel metal5 s 6598 956440 19088 968960 6 mprj_io[24]
port 22 nsew signal bidirectional
rlabel metal5 s 6598 786640 19088 799160 6 mprj_io[25]
port 23 nsew signal bidirectional
rlabel metal5 s 6598 743440 19088 755960 6 mprj_io[26]
port 24 nsew signal bidirectional
rlabel metal5 s 6598 700240 19088 712760 6 mprj_io[27]
port 25 nsew signal bidirectional
rlabel metal5 s 6598 657040 19088 669560 6 mprj_io[28]
port 26 nsew signal bidirectional
rlabel metal5 s 6598 613840 19088 626360 6 mprj_io[29]
port 27 nsew signal bidirectional
rlabel metal5 s 698512 191440 711002 203960 6 mprj_io[2]
port 28 nsew signal bidirectional
rlabel metal5 s 6598 570640 19088 583160 6 mprj_io[30]
port 29 nsew signal bidirectional
rlabel metal5 s 6598 527440 19088 539960 6 mprj_io[31]
port 30 nsew signal bidirectional
rlabel metal5 s 6598 399840 19088 412360 6 mprj_io[32]
port 31 nsew signal bidirectional
rlabel metal5 s 6598 356640 19088 369160 6 mprj_io[33]
port 32 nsew signal bidirectional
rlabel metal5 s 6598 313440 19088 325960 6 mprj_io[34]
port 33 nsew signal bidirectional
rlabel metal5 s 6598 270240 19088 282760 6 mprj_io[35]
port 34 nsew signal bidirectional
rlabel metal5 s 6598 227040 19088 239560 6 mprj_io[36]
port 35 nsew signal bidirectional
rlabel metal5 s 6598 183840 19088 196360 6 mprj_io[37]
port 36 nsew signal bidirectional
rlabel metal5 s 698512 236640 711002 249160 6 mprj_io[3]
port 37 nsew signal bidirectional
rlabel metal5 s 698512 281640 711002 294160 6 mprj_io[4]
port 38 nsew signal bidirectional
rlabel metal5 s 698512 326640 711002 339160 6 mprj_io[5]
port 39 nsew signal bidirectional
rlabel metal5 s 698512 371840 711002 384360 6 mprj_io[6]
port 40 nsew signal bidirectional
rlabel metal5 s 698512 549040 711002 561560 6 mprj_io[7]
port 41 nsew signal bidirectional
rlabel metal5 s 698512 594240 711002 606760 6 mprj_io[8]
port 42 nsew signal bidirectional
rlabel metal5 s 698512 639240 711002 651760 6 mprj_io[9]
port 43 nsew signal bidirectional
rlabel metal5 s 136713 7143 144150 18309 6 resetb
port 44 nsew signal input
rlabel metal5 s 6167 70054 19620 80934 6 vccd
port 45 nsew signal bidirectional
rlabel metal5 s 697980 909666 711433 920546 6 vccd1
port 46 nsew signal bidirectional
rlabel metal5 s 6167 914054 19620 924934 6 vccd2
port 47 nsew signal bidirectional
rlabel metal5 s 624222 6811 636390 18976 6 vdda
port 48 nsew signal bidirectional
rlabel metal5 s 698624 819822 710789 831990 6 vdda1
port 49 nsew signal bidirectional
rlabel metal5 s 698624 505222 710789 517390 6 vdda1_2
port 50 nsew signal bidirectional
rlabel metal5 s 6811 484410 18976 496578 6 vdda2
port 51 nsew signal bidirectional
rlabel metal5 s 6811 111610 18976 123778 6 vddio
port 52 nsew signal bidirectional
rlabel metal5 s 6811 871210 18976 883378 6 vddio_2
port 53 nsew signal bidirectional
rlabel metal5 s 80222 6811 92390 18976 6 vssa
port 54 nsew signal bidirectional
rlabel metal5 s 577010 1018624 589178 1030789 6 vssa1
port 55 nsew signal bidirectional
rlabel metal5 s 698624 417022 710789 429190 6 vssa1_2
port 56 nsew signal bidirectional
rlabel metal5 s 6811 829010 18976 841178 6 vssa2
port 57 nsew signal bidirectional
rlabel metal5 s 243266 6167 254146 19620 6 vssd
port 58 nsew signal bidirectional
rlabel metal5 s 697980 461866 711433 472746 6 vssd1
port 59 nsew signal bidirectional
rlabel metal5 s 6167 442854 19620 453734 6 vssd2
port 60 nsew signal bidirectional
rlabel metal5 s 570422 6811 582590 18976 6 vssio
port 61 nsew signal bidirectional
rlabel metal5 s 334810 1018624 346978 1030789 6 vssio_2
port 62 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
