magic
tech sky130A
magscale 1 2
timestamp 1695675240
<< checkpaint >>
rect 26297 954638 30878 954986
rect 77497 954638 82078 954986
rect 128697 954638 133278 954986
rect 179897 954638 184478 954986
rect 231097 954638 235678 954986
rect 300081 954638 307382 955030
rect 335497 954638 340078 954986
rect 424497 954638 429078 954986
rect 475697 954638 480278 954986
rect 542281 954638 549582 955030
rect 577098 954986 579696 955035
rect 575097 954638 579696 954986
rect -1312 952066 634638 954638
rect -1312 929363 1260 952066
rect 26297 952010 30878 952066
rect 77497 952010 82078 952066
rect 128697 952010 133278 952066
rect 179897 952010 184478 952066
rect 231097 952010 235678 952066
rect 300081 952010 307382 952066
rect 335497 952010 340078 952066
rect 424497 952010 429078 952066
rect 475697 952010 480278 952066
rect 542281 952010 549582 952066
rect 575097 952010 579696 952066
rect 577098 952009 579696 952010
rect 632066 930329 634638 952066
rect -1778 910398 1409 929363
rect 631808 927737 635052 930329
rect 631817 926433 635042 927737
rect 631817 925735 635103 926433
rect -1312 880976 1260 910398
rect -1704 868703 1316 880976
rect -1312 843782 1260 868703
rect -1704 836481 1316 843782
rect 631916 840329 635103 925735
rect 631808 837737 635103 840329
rect -1312 801582 1260 836481
rect 631817 835735 635103 837737
rect -1704 794281 1316 801582
rect -1312 758603 1260 794281
rect -1751 749403 1382 758603
rect 631916 751329 635103 835735
rect -1778 741287 1409 749403
rect 631808 748737 635103 751329
rect 631817 746735 635103 748737
rect -1312 715403 1260 741287
rect -1778 698087 1409 715403
rect 631916 706329 635103 746735
rect 631808 703737 635103 706329
rect 631817 701735 635103 703737
rect -1312 672203 1260 698087
rect -1778 611687 1409 672203
rect 631916 661329 635103 701735
rect 631808 658737 635103 661329
rect 631817 656735 635103 658737
rect 631916 616329 635103 656735
rect 631828 613737 635103 616329
rect 631836 611735 635103 613737
rect -1312 585803 1260 611687
rect -1778 138487 1409 585803
rect 631916 571329 635103 611735
rect 631828 568737 635103 571329
rect 631836 566735 635103 568737
rect 631916 526329 635103 566735
rect 631828 523737 635103 526329
rect 631916 433822 635103 523737
rect 631916 416462 635532 433822
rect 631916 349329 635103 416462
rect 631828 346737 635103 349329
rect 631916 304329 635103 346737
rect 631828 301737 635103 304329
rect 631916 259329 635103 301737
rect 631828 256737 635103 259329
rect 631916 214329 635103 256737
rect 631828 211737 635103 214329
rect 631916 169329 635103 211737
rect 631828 166737 635103 169329
rect -1312 84181 1260 138487
rect 631916 124329 635103 166737
rect 631828 121737 635103 124329
rect -1704 76880 1316 84181
rect 631916 79329 635103 121737
rect -1312 32023 1260 76880
rect 631828 76737 635103 79329
rect 631916 57109 635103 76737
rect -1704 24702 1316 32023
rect -1312 1260 1260 24702
rect 35545 1260 42846 1316
rect 148862 1260 151405 1330
rect 198023 1260 205174 1316
rect 207903 1260 215224 1316
rect 525745 1260 533046 1316
rect 579545 1260 586846 1316
rect 632066 1260 634638 57109
rect -1312 -1312 634638 1260
rect 35545 -1704 42846 -1312
rect 98313 -1660 100834 -1312
rect 148862 -1536 151405 -1312
rect 198023 -1704 205174 -1312
rect 207903 -1704 215224 -1312
rect 525745 -1704 533046 -1312
rect 579545 -1704 586846 -1312
<< metal2 >>
rect 27497 953270 27557 953726
rect 29498 953270 29558 953726
rect 34360 953270 34416 953750
rect 34912 953270 34968 953750
rect 35556 953270 35612 953750
rect 36200 953270 36256 953750
rect 38040 953270 38096 953750
rect 38592 953270 38648 953750
rect 39236 953270 39292 953750
rect 39880 953270 39936 953750
rect 42364 953270 42420 953750
rect 42916 953270 42972 953750
rect 43560 953270 43616 953750
rect 44204 953270 44260 953750
rect 44677 953270 44891 953750
rect 45400 953270 45456 953750
rect 46560 953270 46688 953750
rect 47240 953270 47296 953750
rect 49080 953270 49136 953750
rect 78697 953270 78757 953726
rect 80698 953270 80758 953726
rect 85760 953270 85816 953750
rect 86312 953270 86368 953750
rect 86956 953270 87012 953750
rect 87600 953270 87656 953750
rect 89440 953270 89496 953750
rect 89992 953270 90048 953750
rect 90636 953270 90692 953750
rect 91280 953270 91336 953750
rect 93764 953270 93820 953750
rect 94316 953270 94372 953750
rect 94960 953270 95016 953750
rect 95604 953270 95660 953750
rect 96077 953270 96291 953750
rect 96800 953270 96856 953750
rect 97960 953270 98088 953750
rect 98640 953270 98696 953750
rect 100480 953270 100536 953750
rect 129897 953270 129957 953726
rect 131898 953270 131958 953726
rect 137160 953270 137216 953750
rect 137712 953270 137768 953750
rect 138356 953270 138412 953750
rect 139000 953270 139056 953750
rect 140840 953270 140896 953750
rect 141392 953270 141448 953750
rect 142036 953270 142092 953750
rect 142680 953270 142736 953750
rect 145164 953270 145220 953750
rect 145716 953270 145772 953750
rect 146360 953270 146416 953750
rect 147004 953270 147060 953750
rect 147477 953270 147691 953750
rect 148200 953270 148256 953750
rect 149360 953270 149488 953750
rect 150040 953270 150096 953750
rect 151880 953270 151936 953750
rect 181097 953270 181157 953726
rect 183098 953270 183158 953726
rect 188560 953270 188616 953750
rect 189112 953270 189168 953750
rect 189756 953270 189812 953750
rect 190400 953270 190456 953750
rect 192240 953270 192296 953750
rect 192792 953270 192848 953750
rect 193436 953270 193492 953750
rect 194080 953270 194136 953750
rect 196564 953270 196620 953750
rect 197116 953270 197172 953750
rect 197760 953270 197816 953750
rect 198404 953270 198460 953750
rect 198877 953270 199091 953750
rect 199600 953270 199656 953750
rect 200760 953270 200888 953750
rect 201440 953270 201496 953750
rect 203280 953270 203336 953750
rect 232297 953270 232357 953726
rect 234298 953270 234358 953726
rect 240160 953270 240216 953750
rect 240712 953270 240768 953750
rect 241356 953270 241412 953750
rect 242000 953270 242056 953750
rect 243840 953270 243896 953750
rect 244392 953270 244448 953750
rect 245036 953270 245092 953750
rect 245680 953270 245736 953750
rect 248164 953270 248220 953750
rect 248716 953270 248772 953750
rect 249360 953270 249416 953750
rect 250004 953270 250060 953750
rect 250477 953270 250691 953750
rect 251200 953270 251256 953750
rect 252360 953270 252488 953750
rect 253040 953270 253096 953750
rect 254880 953270 254936 953750
rect 336697 953270 336757 953726
rect 338698 953270 338758 953726
rect 341960 953270 342016 953750
rect 342512 953270 342568 953750
rect 343156 953270 343212 953750
rect 343800 953270 343856 953750
rect 345640 953270 345696 953750
rect 346192 953270 346248 953750
rect 346836 953270 346892 953750
rect 347480 953270 347536 953750
rect 349964 953270 350020 953750
rect 350516 953270 350572 953750
rect 351160 953270 351216 953750
rect 351804 953270 351860 953750
rect 352277 953270 352491 953750
rect 353000 953270 353056 953750
rect 354160 953270 354288 953750
rect 354840 953270 354896 953750
rect 356680 953270 356736 953750
rect 425697 953270 425757 953726
rect 427698 953270 427758 953726
rect 430960 953270 431016 953750
rect 431512 953270 431568 953750
rect 432156 953270 432212 953750
rect 432800 953270 432856 953750
rect 434640 953270 434696 953750
rect 435192 953270 435248 953750
rect 435836 953270 435892 953750
rect 436480 953270 436536 953750
rect 438964 953270 439020 953750
rect 439516 953270 439572 953750
rect 440160 953270 440216 953750
rect 440804 953270 440860 953750
rect 441277 953270 441491 953750
rect 442000 953270 442056 953750
rect 443160 953270 443288 953750
rect 443840 953270 443896 953750
rect 445680 953270 445736 953750
rect 476897 953270 476957 953726
rect 478898 953270 478958 953726
rect 482360 953270 482416 953750
rect 482912 953270 482968 953750
rect 483556 953270 483612 953750
rect 484200 953270 484256 953750
rect 486040 953270 486096 953750
rect 486592 953270 486648 953750
rect 487236 953270 487292 953750
rect 487880 953270 487936 953750
rect 490364 953270 490420 953750
rect 490916 953270 490972 953750
rect 491560 953270 491616 953750
rect 492204 953270 492260 953750
rect 492677 953270 492891 953750
rect 493400 953270 493456 953750
rect 494560 953270 494688 953750
rect 495240 953270 495296 953750
rect 497080 953270 497136 953750
rect 576297 953270 576357 953726
rect 578298 953270 578358 953726
rect 584160 953270 584216 953750
rect 584712 953270 584768 953750
rect 585356 953270 585412 953750
rect 586000 953270 586056 953750
rect 587840 953270 587896 953750
rect 588392 953270 588448 953750
rect 589036 953270 589092 953750
rect 589680 953270 589736 953750
rect 592164 953270 592220 953750
rect 592716 953270 592772 953750
rect 593360 953270 593416 953750
rect 594004 953270 594060 953750
rect 594477 953270 594691 953750
rect 595200 953270 595256 953750
rect 596360 953270 596488 953750
rect 597040 953270 597096 953750
rect 598880 953270 598936 953750
rect 99571 -90 99637 56
rect 99574 -400 99634 -90
rect 110164 -400 110220 56
rect 145190 -424 145246 56
rect 147030 -424 147086 56
rect 147638 -424 147766 56
rect 148870 -424 148926 56
rect 149435 -424 149649 56
rect 150066 -424 150122 56
rect 150710 -424 150766 56
rect 151354 -424 151410 56
rect 151906 -424 151962 56
rect 154390 -424 154446 56
rect 155034 -424 155090 56
rect 155678 -424 155734 56
rect 156230 -424 156286 56
rect 158070 -424 158126 56
rect 158714 -424 158770 56
rect 159358 -424 159414 56
rect 159910 -424 159966 56
rect 160580 -400 160632 56
rect 163791 -400 163843 56
rect 253790 -424 253846 56
rect 255630 -424 255686 56
rect 256238 -424 256366 56
rect 257470 -424 257526 56
rect 258035 -424 258249 56
rect 258666 -424 258722 56
rect 259310 -424 259366 56
rect 259954 -424 260010 56
rect 260506 -424 260562 56
rect 262990 -424 263046 56
rect 263634 -424 263690 56
rect 264278 -424 264334 56
rect 264830 -424 264886 56
rect 266670 -424 266726 56
rect 267314 -424 267370 56
rect 267958 -424 268014 56
rect 268510 -424 268566 56
rect 269180 -400 269232 56
rect 273360 -400 273412 56
rect 308590 -424 308646 56
rect 310430 -424 310486 56
rect 311038 -424 311166 56
rect 312270 -424 312326 56
rect 312835 -424 313049 56
rect 313466 -424 313522 56
rect 314110 -424 314166 56
rect 314754 -424 314810 56
rect 315306 -424 315362 56
rect 317790 -424 317846 56
rect 318434 -424 318490 56
rect 319078 -424 319134 56
rect 319630 -424 319686 56
rect 321470 -424 321526 56
rect 322114 -424 322170 56
rect 322758 -424 322814 56
rect 323310 -424 323366 56
rect 323980 -400 324032 56
rect 328165 -400 328217 34
rect 363390 -424 363446 56
rect 365230 -424 365286 56
rect 365838 -424 365966 56
rect 367070 -424 367126 56
rect 367635 -424 367849 56
rect 368266 -424 368322 56
rect 368910 -424 368966 56
rect 369554 -424 369610 56
rect 370106 -424 370162 56
rect 372590 -424 372646 56
rect 373234 -424 373290 56
rect 373878 -424 373934 56
rect 374430 -424 374486 56
rect 376270 -424 376326 56
rect 376914 -424 376970 56
rect 377558 -424 377614 56
rect 378110 -424 378166 56
rect 378780 -400 378832 56
rect 382978 -400 383030 56
rect 418190 -424 418246 56
rect 420030 -424 420086 56
rect 420638 -424 420766 56
rect 421870 -424 421926 56
rect 422435 -424 422649 56
rect 423066 -424 423122 56
rect 423710 -424 423766 56
rect 424354 -424 424410 56
rect 424906 -424 424962 56
rect 427390 -424 427446 56
rect 428034 -424 428090 56
rect 428678 -424 428734 56
rect 429230 -424 429286 56
rect 431070 -424 431126 56
rect 431714 -424 431770 56
rect 432358 -424 432414 56
rect 432910 -424 432966 56
rect 433580 -400 433632 56
rect 437778 -400 437830 56
rect 472990 -424 473046 56
rect 474830 -424 474886 56
rect 475438 -424 475566 56
rect 476670 -424 476726 56
rect 477235 -424 477449 56
rect 477866 -424 477922 56
rect 478510 -424 478566 56
rect 479154 -424 479210 56
rect 479706 -424 479762 56
rect 482190 -424 482246 56
rect 482834 -424 482890 56
rect 483478 -424 483534 56
rect 484030 -424 484086 56
rect 485870 -424 485926 56
rect 486514 -424 486570 56
rect 487158 -424 487214 56
rect 487710 -424 487766 56
rect 488380 -400 488432 56
rect 492635 -400 492687 56
rect 605082 -260 605134 56
rect 605306 -260 605358 56
rect 605530 -260 605582 56
rect 605754 -260 605806 56
rect 605978 -260 606030 56
rect 606202 -260 606254 56
rect 606426 -260 606478 56
rect 606650 -260 606702 56
rect 606874 -260 606926 56
rect 607098 -260 607150 56
rect 607322 -260 607374 56
rect 607546 -260 607598 56
rect 607770 -260 607822 56
rect 607994 -260 608046 56
rect 608218 -260 608270 56
rect 608442 -260 608494 56
rect 608666 -260 608718 56
rect 608890 -260 608942 56
rect 609114 -260 609166 56
rect 609338 -260 609390 56
rect 609562 -260 609614 56
rect 609786 -260 609838 56
rect 610010 -260 610062 56
rect 610234 -260 610286 56
rect 610458 -260 610510 56
rect 610682 -260 610734 56
rect 610906 -260 610958 56
rect 611130 -260 611182 56
rect 611354 -260 611406 56
rect 611578 -260 611630 56
rect 611802 -260 611854 56
rect 612026 -260 612078 56
rect 605093 -400 605121 -260
rect 605317 -400 605345 -260
rect 605541 -400 605569 -260
rect 605765 -400 605793 -260
rect 605989 -400 606017 -260
rect 606213 -400 606241 -260
rect 606437 -400 606465 -260
rect 606661 -400 606689 -260
rect 606885 -400 606913 -260
rect 607109 -400 607137 -260
rect 607333 -400 607361 -260
rect 607557 -400 607585 -260
rect 607781 -400 607809 -260
rect 608005 -400 608033 -260
rect 608229 -400 608257 -260
rect 608453 -400 608481 -260
rect 608677 -400 608705 -260
rect 608901 -400 608929 -260
rect 609125 -400 609153 -260
rect 609349 -400 609377 -260
rect 609573 -400 609601 -260
rect 609797 -400 609825 -260
rect 610021 -400 610049 -260
rect 610245 -400 610273 -260
rect 610469 -400 610497 -260
rect 610693 -400 610721 -260
rect 610917 -400 610945 -260
rect 611141 -400 611169 -260
rect 611365 -400 611393 -260
rect 611589 -400 611617 -260
rect 611813 -400 611841 -260
rect 612037 -400 612065 -260
<< metal3 >>
rect 291362 953270 296142 953770
rect 301342 953270 306122 953770
rect 533562 953270 538342 953770
rect 543542 953270 548322 953770
rect 633270 929006 633726 929068
rect -424 927072 56 927142
rect 633270 927006 633726 927068
rect -424 925232 56 925302
rect 633270 925104 633750 925174
rect -424 924560 56 924688
rect 633270 924552 633750 924622
rect 633270 923908 633750 923978
rect -424 923392 56 923462
rect 633270 923264 633750 923334
rect -424 922677 56 922891
rect -424 922196 56 922266
rect -424 921552 56 921622
rect 633270 921424 633750 921494
rect -424 920908 56 920978
rect 633270 920872 633750 920942
rect -424 920356 56 920426
rect 633270 920228 633750 920298
rect 633270 919584 633750 919654
rect -424 917872 56 917942
rect -424 917228 56 917298
rect 633270 917100 633750 917170
rect -424 916584 56 916654
rect 633270 916548 633750 916618
rect -424 916032 56 916102
rect 633270 915904 633750 915974
rect 633270 915260 633750 915330
rect 633270 914635 633750 914849
rect -424 914192 56 914262
rect 633270 914064 633750 914134
rect -424 913548 56 913618
rect -424 912904 56 912974
rect 633270 912838 633750 912966
rect -424 912352 56 912422
rect 633270 912224 633750 912294
rect 633270 910384 633750 910454
rect -400 906644 56 906704
rect -400 904644 56 904704
rect -444 880014 56 884804
rect -444 875054 56 879716
rect -444 869964 56 874764
rect -444 837742 56 842522
rect 633270 839006 633726 839068
rect 633270 837006 633726 837068
rect 633270 835904 633750 835974
rect 633270 835352 633750 835422
rect 633270 834708 633750 834778
rect 633270 834064 633750 834134
rect -444 827762 56 832542
rect 633270 832224 633750 832294
rect 633270 831672 633750 831742
rect 633270 831028 633750 831098
rect 633270 830384 633750 830454
rect 633270 827900 633750 827970
rect 633270 827348 633750 827418
rect 633270 826704 633750 826774
rect 633270 826060 633750 826130
rect 633270 825435 633750 825649
rect 633270 824864 633750 824934
rect 633270 823638 633750 823766
rect 633270 823024 633750 823094
rect 633270 821184 633750 821254
rect -444 795542 56 800322
rect -444 785562 56 790342
rect 633270 786384 633770 791164
rect 633270 776406 633770 781186
rect -424 757272 56 757342
rect -424 755432 56 755502
rect -424 754760 56 754888
rect -424 753592 56 753662
rect -424 752877 56 753091
rect -424 752396 56 752466
rect -424 751752 56 751822
rect -424 751108 56 751178
rect -424 750556 56 750626
rect 633270 750006 633726 750068
rect -424 748072 56 748142
rect 633270 748006 633726 748068
rect -424 747428 56 747498
rect -424 746784 56 746854
rect 633270 746704 633750 746774
rect -424 746232 56 746302
rect 633270 746152 633750 746222
rect 633270 745508 633750 745578
rect 633270 744864 633750 744934
rect -424 744392 56 744462
rect -424 743748 56 743818
rect -424 743104 56 743174
rect 633270 743024 633750 743094
rect -424 742552 56 742622
rect 633270 742472 633750 742542
rect 633270 741828 633750 741898
rect 633270 741184 633750 741254
rect 633270 738700 633750 738770
rect 633270 738148 633750 738218
rect 633270 737504 633750 737574
rect 633270 736860 633750 736930
rect -400 736644 56 736704
rect 633270 736235 633750 736449
rect 633270 735664 633750 735734
rect -400 734644 56 734704
rect 633270 734438 633750 734566
rect 633270 733824 633750 733894
rect 633270 731984 633750 732054
rect -424 714072 56 714142
rect -424 712232 56 712302
rect -424 711560 56 711688
rect -424 710392 56 710462
rect -424 709677 56 709891
rect -424 709196 56 709266
rect -424 708552 56 708622
rect -424 707908 56 707978
rect -424 707356 56 707426
rect 633270 705006 633726 705068
rect -424 704872 56 704942
rect -424 704228 56 704298
rect -424 703584 56 703654
rect -424 703032 56 703102
rect 633270 703006 633726 703068
rect 633270 701704 633750 701774
rect -424 701192 56 701262
rect 633270 701152 633750 701222
rect -424 700548 56 700618
rect 633270 700508 633750 700578
rect -424 699904 56 699974
rect 633270 699864 633750 699934
rect -424 699352 56 699422
rect 633270 698024 633750 698094
rect 633270 697472 633750 697542
rect 633270 696828 633750 696898
rect 633270 696184 633750 696254
rect -400 693644 56 693704
rect 633270 693700 633750 693770
rect 633270 693148 633750 693218
rect 633270 692504 633750 692574
rect 633270 691860 633750 691930
rect -400 691644 56 691704
rect 633270 691235 633750 691449
rect 633270 690664 633750 690734
rect 633270 689438 633750 689566
rect 633270 688824 633750 688894
rect 633270 686984 633750 687054
rect -424 670872 56 670942
rect -424 669032 56 669102
rect -424 668360 56 668488
rect -424 667192 56 667262
rect -424 666477 56 666691
rect -424 665996 56 666066
rect -424 665352 56 665422
rect -424 664708 56 664778
rect -424 664156 56 664226
rect -424 661672 56 661742
rect -424 661028 56 661098
rect -424 660384 56 660454
rect 633270 660006 633726 660068
rect -424 659832 56 659902
rect -424 657992 56 658062
rect 633270 658006 633726 658068
rect -424 657348 56 657418
rect -424 656704 56 656774
rect 633270 656704 633750 656774
rect -424 656152 56 656222
rect 633270 656152 633750 656222
rect 633270 655508 633750 655578
rect 633270 654864 633750 654934
rect 633270 653024 633750 653094
rect 633270 652472 633750 652542
rect 633270 651828 633750 651898
rect 633270 651184 633750 651254
rect -400 650644 56 650704
rect -400 648644 56 648704
rect 633270 648700 633750 648770
rect 633270 648148 633750 648218
rect 633270 647504 633750 647574
rect 633270 646860 633750 646930
rect 633270 646235 633750 646449
rect 633270 645664 633750 645734
rect 633270 644438 633750 644566
rect 633270 643824 633750 643894
rect 633270 641984 633750 642054
rect -424 627672 56 627742
rect -424 625832 56 625902
rect -424 625160 56 625288
rect -424 623992 56 624062
rect -424 623277 56 623491
rect -424 622796 56 622866
rect -424 622152 56 622222
rect -424 621508 56 621578
rect -424 620956 56 621026
rect -424 618472 56 618542
rect -424 617828 56 617898
rect -424 617184 56 617254
rect -424 616632 56 616702
rect 633270 615006 633726 615068
rect -424 614792 56 614862
rect -424 614148 56 614218
rect -424 613504 56 613574
rect -424 612952 56 613022
rect 633270 613006 633726 613068
rect 633270 611504 633750 611574
rect 633270 610952 633750 611022
rect 633270 610308 633750 610378
rect 633270 609664 633750 609734
rect 633270 607824 633750 607894
rect -400 607644 56 607704
rect 633270 607272 633750 607342
rect 633270 606628 633750 606698
rect 633270 605984 633750 606054
rect -400 605644 56 605704
rect 633270 603500 633750 603570
rect 633270 602948 633750 603018
rect 633270 602304 633750 602374
rect 633270 601660 633750 601730
rect 633270 601035 633750 601249
rect 633270 600464 633750 600534
rect 633270 599238 633750 599366
rect 633270 598624 633750 598694
rect 633270 596784 633750 596854
rect -424 584472 56 584542
rect -424 582632 56 582702
rect -424 581960 56 582088
rect -424 580792 56 580862
rect -424 580077 56 580291
rect -424 579596 56 579666
rect -424 578952 56 579022
rect -424 578308 56 578378
rect -424 577756 56 577826
rect -424 575272 56 575342
rect -424 574628 56 574698
rect -424 573984 56 574054
rect -424 573432 56 573502
rect -424 571592 56 571662
rect -424 570948 56 571018
rect -424 570304 56 570374
rect 633270 570006 633726 570068
rect -424 569752 56 569822
rect 633270 568006 633726 568068
rect 633270 566504 633750 566574
rect 633270 565952 633750 566022
rect 633270 565308 633750 565378
rect -400 564644 56 564704
rect 633270 564664 633750 564734
rect 633270 562824 633750 562894
rect -400 562644 56 562704
rect 633270 562272 633750 562342
rect 633270 561628 633750 561698
rect 633270 560984 633750 561054
rect 633270 558500 633750 558570
rect 633270 557948 633750 558018
rect 633270 557304 633750 557374
rect 633270 556660 633750 556730
rect 633270 556035 633750 556249
rect 633270 555464 633750 555534
rect 633270 554238 633750 554366
rect 633270 553624 633750 553694
rect 633270 551784 633750 551854
rect -424 541272 56 541342
rect -424 539432 56 539502
rect -424 538760 56 538888
rect -424 537592 56 537662
rect -424 536877 56 537091
rect -424 536396 56 536466
rect -424 535752 56 535822
rect -424 535108 56 535178
rect -424 534556 56 534626
rect -424 532072 56 532142
rect -424 531428 56 531498
rect -424 530784 56 530854
rect -424 530232 56 530302
rect -424 528392 56 528462
rect -424 527748 56 527818
rect -424 527104 56 527174
rect -424 526552 56 526622
rect 633270 525006 633726 525068
rect 633270 523005 633726 523067
rect -400 521644 56 521704
rect 633270 521304 633750 521374
rect 633270 520752 633750 520822
rect 633270 520108 633750 520178
rect -400 519644 56 519704
rect 633270 519464 633750 519534
rect 633270 517624 633750 517694
rect 633270 517072 633750 517142
rect 633270 516428 633750 516498
rect 633270 515784 633750 515854
rect 633270 513300 633750 513370
rect 633270 512748 633750 512818
rect 633270 512104 633750 512174
rect 633270 511460 633750 511530
rect 633270 510835 633750 511049
rect 633270 510264 633750 510334
rect 633270 509038 633750 509166
rect 633270 508424 633750 508494
rect 633270 506584 633750 506654
rect -424 498072 56 498142
rect -424 496232 56 496302
rect -424 495560 56 495688
rect -424 494392 56 494462
rect -424 493677 56 493891
rect -424 493196 56 493266
rect -424 492552 56 492622
rect -424 491908 56 491978
rect -424 491356 56 491426
rect -424 488872 56 488942
rect -424 488228 56 488298
rect -424 487584 56 487654
rect -424 487032 56 487102
rect -424 485192 56 485262
rect -424 484548 56 484618
rect -424 483904 56 483974
rect -424 483352 56 483422
rect -400 478644 56 478704
rect -400 476644 56 476704
rect 633270 471784 633770 476564
rect 633270 461804 633770 466584
rect -444 450940 56 455720
rect -444 440962 56 445742
rect 633270 427762 633770 432562
rect 633270 422810 633770 427472
rect 633270 417722 633770 422512
rect -444 408814 56 413604
rect -444 403862 56 408514
rect -444 398762 56 403562
rect 633270 383584 633770 388364
rect 633270 373606 633770 378386
rect -424 370472 56 370542
rect -424 368632 56 368702
rect -424 367960 56 368088
rect -424 366792 56 366862
rect -424 366077 56 366291
rect -424 365596 56 365666
rect -424 364952 56 365022
rect -424 364308 56 364378
rect -424 363756 56 363826
rect -424 361272 56 361342
rect -424 360628 56 360698
rect -424 359984 56 360054
rect -424 359432 56 359502
rect -424 357592 56 357662
rect -424 356948 56 357018
rect -424 356304 56 356374
rect -424 355752 56 355822
rect -400 349644 56 349704
rect 633270 348006 633726 348068
rect -400 347644 56 347704
rect 633270 346005 633726 346067
rect 633270 344104 633750 344174
rect 633270 343552 633750 343622
rect 633270 342908 633750 342978
rect 633270 342264 633750 342334
rect 633270 340424 633750 340494
rect 633270 339872 633750 339942
rect 633270 339228 633750 339298
rect 633270 338584 633750 338654
rect 633270 336100 633750 336170
rect 633270 335548 633750 335618
rect 633270 334904 633750 334974
rect 633270 334260 633750 334330
rect 633270 333635 633750 333849
rect 633270 333064 633750 333134
rect 633270 331838 633750 331966
rect 633270 331224 633750 331294
rect 633270 329384 633750 329454
rect -424 327272 56 327342
rect -424 325432 56 325502
rect -424 324760 56 324888
rect -424 323592 56 323662
rect -424 322877 56 323091
rect -424 322396 56 322466
rect -424 321752 56 321822
rect -424 321108 56 321178
rect -424 320556 56 320626
rect -424 318072 56 318142
rect -424 317428 56 317498
rect -424 316784 56 316854
rect -424 316232 56 316302
rect -424 314392 56 314462
rect -424 313748 56 313818
rect -424 313104 56 313174
rect -424 312552 56 312622
rect -400 306644 56 306704
rect -400 304644 56 304704
rect 633270 303006 633726 303068
rect 633270 301005 633726 301067
rect 633270 298904 633750 298974
rect 633270 298352 633750 298422
rect 633270 297708 633750 297778
rect 633270 297064 633750 297134
rect 633270 295224 633750 295294
rect 633270 294672 633750 294742
rect 633270 294028 633750 294098
rect 633270 293384 633750 293454
rect 633270 290900 633750 290970
rect 633270 290348 633750 290418
rect 633270 289704 633750 289774
rect 633270 289060 633750 289130
rect 633270 288435 633750 288649
rect 633270 287864 633750 287934
rect 633270 286638 633750 286766
rect 633270 286024 633750 286094
rect 633270 284184 633750 284254
rect -424 284072 56 284142
rect -424 282232 56 282302
rect -424 281560 56 281688
rect -424 280392 56 280462
rect -424 279677 56 279891
rect -424 279196 56 279266
rect -424 278552 56 278622
rect -424 277908 56 277978
rect -424 277356 56 277426
rect -424 274872 56 274942
rect -424 274228 56 274298
rect -424 273584 56 273654
rect -424 273032 56 273102
rect -424 271192 56 271262
rect -424 270548 56 270618
rect -424 269904 56 269974
rect -424 269352 56 269422
rect -400 263644 56 263704
rect -400 261644 56 261704
rect 633270 258006 633726 258068
rect 633270 256005 633726 256067
rect 633270 253904 633750 253974
rect 633270 253352 633750 253422
rect 633270 252708 633750 252778
rect 633270 252064 633750 252134
rect 633270 250224 633750 250294
rect 633270 249672 633750 249742
rect 633270 249028 633750 249098
rect 633270 248384 633750 248454
rect 633270 245900 633750 245970
rect 633270 245348 633750 245418
rect 633270 244704 633750 244774
rect 633270 244060 633750 244130
rect 633270 243435 633750 243649
rect 633270 242864 633750 242934
rect 633270 241638 633750 241766
rect 633270 241024 633750 241094
rect -424 240872 56 240942
rect 633270 239184 633750 239254
rect -424 239032 56 239102
rect -424 238360 56 238488
rect -424 237192 56 237262
rect -424 236477 56 236691
rect -424 235996 56 236066
rect -424 235352 56 235422
rect -424 234708 56 234778
rect -424 234156 56 234226
rect -424 231672 56 231742
rect -424 231028 56 231098
rect -424 230384 56 230454
rect -424 229832 56 229902
rect -424 227992 56 228062
rect -424 227348 56 227418
rect -424 226704 56 226774
rect -424 226152 56 226222
rect -400 220644 56 220704
rect -400 218644 56 218704
rect 633270 213006 633726 213068
rect 633270 211005 633726 211067
rect 633270 208904 633750 208974
rect 633270 208352 633750 208422
rect 633270 207708 633750 207778
rect 633270 207064 633750 207134
rect 633270 205224 633750 205294
rect 633270 204672 633750 204742
rect 633270 204028 633750 204098
rect 633270 203384 633750 203454
rect 633270 200900 633750 200970
rect 633270 200348 633750 200418
rect 633270 199704 633750 199774
rect 633270 199060 633750 199130
rect 633270 198435 633750 198649
rect 633270 197864 633750 197934
rect -424 197672 56 197742
rect 633270 196638 633750 196766
rect 633270 196024 633750 196094
rect -424 195832 56 195902
rect -424 195160 56 195288
rect 633270 194184 633750 194254
rect -424 193992 56 194062
rect -424 193277 56 193491
rect -424 192796 56 192866
rect -424 192152 56 192222
rect -424 191508 56 191578
rect -424 190956 56 191026
rect -424 188472 56 188542
rect -424 187828 56 187898
rect -424 187184 56 187254
rect -424 186632 56 186702
rect -424 184792 56 184862
rect -424 184148 56 184218
rect -424 183504 56 183574
rect -424 182952 56 183022
rect -400 177644 56 177704
rect -400 175644 56 175704
rect 633270 168006 633726 168068
rect 633270 166005 633726 166067
rect 633270 163704 633750 163774
rect 633270 163152 633750 163222
rect 633270 162508 633750 162578
rect 633270 161864 633750 161934
rect 633270 160024 633750 160094
rect 633270 159472 633750 159542
rect 633270 158828 633750 158898
rect 633270 158184 633750 158254
rect 633270 155700 633750 155770
rect 633270 155148 633750 155218
rect -424 154472 56 154542
rect 633270 154504 633750 154574
rect 633270 153860 633750 153930
rect 633270 153235 633750 153449
rect -424 152632 56 152702
rect 633270 152664 633750 152734
rect -424 151960 56 152088
rect 633270 151438 633750 151566
rect -424 150792 56 150862
rect 633270 150824 633750 150894
rect -424 150077 56 150291
rect -424 149596 56 149666
rect -424 148952 56 149022
rect 633270 148984 633750 149054
rect -424 148308 56 148378
rect -424 147756 56 147826
rect -424 145272 56 145342
rect -424 144628 56 144698
rect -424 143984 56 144054
rect -424 143432 56 143502
rect -424 141592 56 141662
rect -424 140948 56 141018
rect -424 140304 56 140374
rect -424 139752 56 139822
rect -400 134644 56 134704
rect -400 132644 56 132704
rect 633270 123006 633726 123068
rect 633270 121005 633726 121067
rect 633270 118704 633750 118774
rect 633270 118152 633750 118222
rect 633270 117508 633750 117578
rect 633270 116864 633750 116934
rect 633270 115024 633750 115094
rect 633270 114472 633750 114542
rect 633270 113828 633750 113898
rect 633270 113184 633750 113254
rect 633270 110700 633750 110770
rect 633270 110148 633750 110218
rect 633270 109504 633750 109574
rect 633270 108860 633750 108930
rect 633270 108235 633750 108449
rect 633270 107664 633750 107734
rect 633270 106438 633750 106566
rect 633270 105824 633750 105894
rect 633270 103984 633750 104054
rect -444 78140 56 82920
rect 633270 78006 633726 78068
rect 633270 76005 633726 76067
rect 633270 73504 633750 73574
rect 633270 72952 633750 73022
rect -444 68162 56 72942
rect 633270 72308 633750 72378
rect 633270 71664 633750 71734
rect 633270 69824 633750 69894
rect 633270 69272 633750 69342
rect 633270 68628 633750 68698
rect 633270 67984 633750 68054
rect 633270 65500 633750 65570
rect 633270 64948 633750 65018
rect 633270 64304 633750 64374
rect 633270 63660 633750 63730
rect 633270 63035 633750 63249
rect 633270 62464 633750 62534
rect 633270 61238 633750 61366
rect 633270 60624 633750 60694
rect 633270 58784 633750 58854
rect -400 53595 56 53665
rect -400 53372 56 53442
rect -400 53147 56 53217
rect -444 36014 56 40804
rect -444 25962 56 30762
rect 36806 -444 41586 56
rect 46784 -444 51564 56
rect 199284 -444 203914 56
rect 209164 -444 213964 56
rect 527006 -444 531786 56
rect 536984 -444 541764 56
rect 580806 -444 585586 56
rect 590784 -444 595564 56
<< comment >>
rect -400 953326 633726 953726
rect -400 0 0 953326
rect 633326 58370 633726 953326
rect 633326 0 633726 58369
rect -400 -400 633726 0
<< labels >>
flabel metal2 485870 -424 485926 56 0 FreeSans 400 270 0 0 gpio_vtrip_sel[43]
port 290 nsew
flabel metal2 s 594004 953270 594060 953750 0 FreeSans 400 90 0 0 gpio_analog_en[15]
port 450 nsew
flabel metal2 s 592716 953270 592772 953750 0 FreeSans 400 90 0 0 gpio_analog_pol[15]
port 538 nsew
flabel metal2 s 589680 953270 589736 953750 0 FreeSans 400 90 0 0 gpio_analog_sel[15]
port 494 nsew
flabel metal2 s 593360 953270 593416 953750 0 FreeSans 400 90 0 0 gpio_dm0[15]
port 582 nsew
flabel metal2 s 595200 953270 595256 953750 0 FreeSans 400 90 0 0 gpio_dm1[15]
port 626 nsew
flabel metal2 s 589036 953270 589092 953750 0 FreeSans 400 90 0 0 gpio_dm2[15]
port 670 nsew
flabel metal2 s 588392 953270 588448 953750 0 FreeSans 400 90 0 0 gpio_holdover[15]
port 406 nsew
flabel metal2 s 585356 953270 585412 953750 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[15]
port 274 nsew
flabel metal2 s 592164 953270 592220 953750 0 FreeSans 400 90 0 0 gpio_inp_dis[15]
port 230 nsew
flabel metal2 s 584712 953270 584768 953750 0 FreeSans 400 90 0 0 gpio_oeb[15]
port 186 nsew
flabel metal2 s 587840 953270 587896 953750 0 FreeSans 400 90 0 0 gpio_out[15]
port 142 nsew
flabel metal2 s 597040 953270 597096 953750 0 FreeSans 400 90 0 0 gpio_slow_sel[15]
port 362 nsew
flabel metal2 s 586000 953270 586056 953750 0 FreeSans 400 90 0 0 gpio_vtrip_sel[15]
port 318 nsew
flabel metal2 s 598880 953270 598936 953750 0 FreeSans 400 90 0 0 gpio_in[15]
port 714 nsew
flabel metal2 s 492204 953270 492260 953750 0 FreeSans 400 90 0 0 gpio_analog_en[16]
port 449 nsew
flabel metal2 s 490916 953270 490972 953750 0 FreeSans 400 90 0 0 gpio_analog_pol[16]
port 537 nsew
flabel metal2 s 487880 953270 487936 953750 0 FreeSans 400 90 0 0 gpio_analog_sel[16]
port 493 nsew
flabel metal2 s 491560 953270 491616 953750 0 FreeSans 400 90 0 0 gpio_dm0[16]
port 581 nsew
flabel metal2 s 493400 953270 493456 953750 0 FreeSans 400 90 0 0 gpio_dm1[16]
port 625 nsew
flabel metal2 s 487236 953270 487292 953750 0 FreeSans 400 90 0 0 gpio_dm2[16]
port 669 nsew
flabel metal2 s 486592 953270 486648 953750 0 FreeSans 400 90 0 0 gpio_holdover[16]
port 405 nsew
flabel metal2 s 483556 953270 483612 953750 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[16]
port 273 nsew
flabel metal2 s 490364 953270 490420 953750 0 FreeSans 400 90 0 0 gpio_inp_dis[16]
port 229 nsew
flabel metal2 s 482912 953270 482968 953750 0 FreeSans 400 90 0 0 gpio_oeb[16]
port 185 nsew
flabel metal2 s 486040 953270 486096 953750 0 FreeSans 400 90 0 0 gpio_out[16]
port 141 nsew
flabel metal2 s 495240 953270 495296 953750 0 FreeSans 400 90 0 0 gpio_slow_sel[16]
port 361 nsew
flabel metal2 s 484200 953270 484256 953750 0 FreeSans 400 90 0 0 gpio_vtrip_sel[16]
port 317 nsew
flabel metal2 s 497080 953270 497136 953750 0 FreeSans 400 90 0 0 gpio_in[16]
port 713 nsew
flabel metal2 s 442000 953270 442056 953750 0 FreeSans 400 90 0 0 gpio_dm1[17]
port 624 nsew
flabel metal2 s 435836 953270 435892 953750 0 FreeSans 400 90 0 0 gpio_dm2[17]
port 668 nsew
flabel metal2 s 435192 953270 435248 953750 0 FreeSans 400 90 0 0 gpio_holdover[17]
port 404 nsew
flabel metal2 s 432156 953270 432212 953750 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[17]
port 272 nsew
flabel metal2 s 438964 953270 439020 953750 0 FreeSans 400 90 0 0 gpio_inp_dis[17]
port 228 nsew
flabel metal2 s 431512 953270 431568 953750 0 FreeSans 400 90 0 0 gpio_oeb[17]
port 184 nsew
flabel metal2 s 434640 953270 434696 953750 0 FreeSans 400 90 0 0 gpio_out[17]
port 140 nsew
flabel metal2 s 443840 953270 443896 953750 0 FreeSans 400 90 0 0 gpio_slow_sel[17]
port 360 nsew
flabel metal2 s 432800 953270 432856 953750 0 FreeSans 400 90 0 0 gpio_vtrip_sel[17]
port 316 nsew
flabel metal2 s 445680 953270 445736 953750 0 FreeSans 400 90 0 0 gpio_in[17]
port 712 nsew
flabel metal2 s 351804 953270 351860 953750 0 FreeSans 400 90 0 0 gpio_analog_en[18]
port 447 nsew
flabel metal2 s 350516 953270 350572 953750 0 FreeSans 400 90 0 0 gpio_analog_pol[18]
port 535 nsew
flabel metal2 s 347480 953270 347536 953750 0 FreeSans 400 90 0 0 gpio_analog_sel[18]
port 491 nsew
flabel metal2 s 351160 953270 351216 953750 0 FreeSans 400 90 0 0 gpio_dm0[18]
port 579 nsew
flabel metal2 s 353000 953270 353056 953750 0 FreeSans 400 90 0 0 gpio_dm1[18]
port 623 nsew
flabel metal2 s 346836 953270 346892 953750 0 FreeSans 400 90 0 0 gpio_dm2[18]
port 667 nsew
flabel metal2 s 346192 953270 346248 953750 0 FreeSans 400 90 0 0 gpio_holdover[18]
port 403 nsew
flabel metal2 s 343156 953270 343212 953750 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[18]
port 271 nsew
flabel metal2 s 349964 953270 350020 953750 0 FreeSans 400 90 0 0 gpio_inp_dis[18]
port 227 nsew
flabel metal2 s 342512 953270 342568 953750 0 FreeSans 400 90 0 0 gpio_oeb[18]
port 183 nsew
flabel metal2 s 345640 953270 345696 953750 0 FreeSans 400 90 0 0 gpio_out[18]
port 139 nsew
flabel metal2 s 354840 953270 354896 953750 0 FreeSans 400 90 0 0 gpio_slow_sel[18]
port 359 nsew
flabel metal2 s 343800 953270 343856 953750 0 FreeSans 400 90 0 0 gpio_vtrip_sel[18]
port 315 nsew
flabel metal2 s 356680 953270 356736 953750 0 FreeSans 400 90 0 0 gpio_in[18]
port 711 nsew
flabel metal2 s 440804 953270 440860 953750 0 FreeSans 400 90 0 0 gpio_analog_en[17]
port 448 nsew
flabel metal2 s 439516 953270 439572 953750 0 FreeSans 400 90 0 0 gpio_analog_pol[17]
port 536 nsew
flabel metal2 s 436480 953270 436536 953750 0 FreeSans 400 90 0 0 gpio_analog_sel[17]
port 492 nsew
flabel metal2 s 440160 953270 440216 953750 0 FreeSans 400 90 0 0 gpio_dm0[17]
port 580 nsew
flabel metal2 s 253040 953270 253096 953750 0 FreeSans 400 90 0 0 gpio_slow_sel[19]
port 358 nsew
flabel metal2 s 242000 953270 242056 953750 0 FreeSans 400 90 0 0 gpio_vtrip_sel[19]
port 314 nsew
flabel metal2 s 254880 953270 254936 953750 0 FreeSans 400 90 0 0 gpio_in[19]
port 710 nsew
flabel metal2 s 198404 953270 198460 953750 0 FreeSans 400 90 0 0 gpio_analog_en[20]
port 445 nsew
flabel metal2 s 197116 953270 197172 953750 0 FreeSans 400 90 0 0 gpio_analog_pol[20]
port 533 nsew
flabel metal2 s 194080 953270 194136 953750 0 FreeSans 400 90 0 0 gpio_analog_sel[20]
port 489 nsew
flabel metal2 s 197760 953270 197816 953750 0 FreeSans 400 90 0 0 gpio_dm0[20]
port 577 nsew
flabel metal2 s 199600 953270 199656 953750 0 FreeSans 400 90 0 0 gpio_dm1[20]
port 621 nsew
flabel metal2 s 193436 953270 193492 953750 0 FreeSans 400 90 0 0 gpio_dm2[20]
port 665 nsew
flabel metal2 s 192792 953270 192848 953750 0 FreeSans 400 90 0 0 gpio_holdover[20]
port 401 nsew
flabel metal2 s 189756 953270 189812 953750 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[20]
port 269 nsew
flabel metal2 s 196564 953270 196620 953750 0 FreeSans 400 90 0 0 gpio_inp_dis[20]
port 225 nsew
flabel metal2 s 189112 953270 189168 953750 0 FreeSans 400 90 0 0 gpio_oeb[20]
port 181 nsew
flabel metal2 s 192240 953270 192296 953750 0 FreeSans 400 90 0 0 gpio_out[20]
port 137 nsew
flabel metal2 s 201440 953270 201496 953750 0 FreeSans 400 90 0 0 gpio_slow_sel[20]
port 357 nsew
flabel metal2 s 190400 953270 190456 953750 0 FreeSans 400 90 0 0 gpio_vtrip_sel[20]
port 313 nsew
flabel metal2 s 203280 953270 203336 953750 0 FreeSans 400 90 0 0 gpio_in[20]
port 709 nsew
flabel metal2 s 250004 953270 250060 953750 0 FreeSans 400 90 0 0 gpio_analog_en[19]
port 446 nsew
flabel metal2 s 248716 953270 248772 953750 0 FreeSans 400 90 0 0 gpio_analog_pol[19]
port 534 nsew
flabel metal2 s 245680 953270 245736 953750 0 FreeSans 400 90 0 0 gpio_analog_sel[19]
port 490 nsew
flabel metal2 s 249360 953270 249416 953750 0 FreeSans 400 90 0 0 gpio_dm0[19]
port 578 nsew
flabel metal2 s 251200 953270 251256 953750 0 FreeSans 400 90 0 0 gpio_dm1[19]
port 622 nsew
flabel metal2 s 245036 953270 245092 953750 0 FreeSans 400 90 0 0 gpio_dm2[19]
port 666 nsew
flabel metal2 s 244392 953270 244448 953750 0 FreeSans 400 90 0 0 gpio_holdover[19]
port 402 nsew
flabel metal2 s 241356 953270 241412 953750 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[19]
port 270 nsew
flabel metal2 s 248164 953270 248220 953750 0 FreeSans 400 90 0 0 gpio_inp_dis[19]
port 226 nsew
flabel metal2 s 240712 953270 240768 953750 0 FreeSans 400 90 0 0 gpio_oeb[19]
port 182 nsew
flabel metal2 s 243840 953270 243896 953750 0 FreeSans 400 90 0 0 gpio_out[19]
port 138 nsew
flabel metal2 s 151880 953270 151936 953750 0 FreeSans 400 90 0 0 gpio_in[21]
port 708 nsew
flabel metal2 s 95604 953270 95660 953750 0 FreeSans 400 90 0 0 gpio_analog_en[22]
port 443 nsew
flabel metal2 s 94316 953270 94372 953750 0 FreeSans 400 90 0 0 gpio_analog_pol[22]
port 531 nsew
flabel metal2 s 91280 953270 91336 953750 0 FreeSans 400 90 0 0 gpio_analog_sel[22]
port 487 nsew
flabel metal2 s 94960 953270 95016 953750 0 FreeSans 400 90 0 0 gpio_dm0[22]
port 575 nsew
flabel metal2 s 96800 953270 96856 953750 0 FreeSans 400 90 0 0 gpio_dm1[22]
port 619 nsew
flabel metal2 s 90636 953270 90692 953750 0 FreeSans 400 90 0 0 gpio_dm2[22]
port 663 nsew
flabel metal2 s 89992 953270 90048 953750 0 FreeSans 400 90 0 0 gpio_holdover[22]
port 399 nsew
flabel metal2 s 86956 953270 87012 953750 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[22]
port 267 nsew
flabel metal2 s 93764 953270 93820 953750 0 FreeSans 400 90 0 0 gpio_inp_dis[22]
port 223 nsew
flabel metal2 s 86312 953270 86368 953750 0 FreeSans 400 90 0 0 gpio_oeb[22]
port 179 nsew
flabel metal2 s 89440 953270 89496 953750 0 FreeSans 400 90 0 0 gpio_out[22]
port 135 nsew
flabel metal2 s 98640 953270 98696 953750 0 FreeSans 400 90 0 0 gpio_slow_sel[22]
port 355 nsew
flabel metal2 s 87600 953270 87656 953750 0 FreeSans 400 90 0 0 gpio_vtrip_sel[22]
port 311 nsew
flabel metal2 s 100480 953270 100536 953750 0 FreeSans 400 90 0 0 gpio_in[22]
port 707 nsew
flabel metal2 s 44204 953270 44260 953750 0 FreeSans 400 90 0 0 gpio_analog_en[23]
port 442 nsew
flabel metal2 s 42916 953270 42972 953750 0 FreeSans 400 90 0 0 gpio_analog_pol[23]
port 530 nsew
flabel metal2 s 39880 953270 39936 953750 0 FreeSans 400 90 0 0 gpio_analog_sel[23]
port 486 nsew
flabel metal2 s 43560 953270 43616 953750 0 FreeSans 400 90 0 0 gpio_dm0[23]
port 574 nsew
flabel metal2 s 45400 953270 45456 953750 0 FreeSans 400 90 0 0 gpio_dm1[23]
port 618 nsew
flabel metal2 s 39236 953270 39292 953750 0 FreeSans 400 90 0 0 gpio_dm2[23]
port 662 nsew
flabel metal2 s 38592 953270 38648 953750 0 FreeSans 400 90 0 0 gpio_holdover[23]
port 398 nsew
flabel metal2 s 35556 953270 35612 953750 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[23]
port 266 nsew
flabel metal2 s 42364 953270 42420 953750 0 FreeSans 400 90 0 0 gpio_inp_dis[23]
port 222 nsew
flabel metal2 s 34912 953270 34968 953750 0 FreeSans 400 90 0 0 gpio_oeb[23]
port 178 nsew
flabel metal2 s 38040 953270 38096 953750 0 FreeSans 400 90 0 0 gpio_out[23]
port 134 nsew
flabel metal2 s 47240 953270 47296 953750 0 FreeSans 400 90 0 0 gpio_slow_sel[23]
port 354 nsew
flabel metal2 s 36200 953270 36256 953750 0 FreeSans 400 90 0 0 gpio_vtrip_sel[23]
port 310 nsew
flabel metal2 s 49080 953270 49136 953750 0 FreeSans 400 90 0 0 gpio_in[23]
port 706 nsew
flabel metal2 s 147004 953270 147060 953750 0 FreeSans 400 90 0 0 gpio_analog_en[21]
port 444 nsew
flabel metal2 s 145716 953270 145772 953750 0 FreeSans 400 90 0 0 gpio_analog_pol[21]
port 532 nsew
flabel metal2 s 142680 953270 142736 953750 0 FreeSans 400 90 0 0 gpio_analog_sel[21]
port 488 nsew
flabel metal2 s 146360 953270 146416 953750 0 FreeSans 400 90 0 0 gpio_dm0[21]
port 576 nsew
flabel metal2 s 148200 953270 148256 953750 0 FreeSans 400 90 0 0 gpio_dm1[21]
port 620 nsew
flabel metal2 s 142036 953270 142092 953750 0 FreeSans 400 90 0 0 gpio_dm2[21]
port 664 nsew
flabel metal2 s 141392 953270 141448 953750 0 FreeSans 400 90 0 0 gpio_holdover[21]
port 400 nsew
flabel metal2 s 138356 953270 138412 953750 0 FreeSans 400 90 0 0 gpio_ib_mode_sel[21]
port 268 nsew
flabel metal2 s 145164 953270 145220 953750 0 FreeSans 400 90 0 0 gpio_inp_dis[21]
port 224 nsew
flabel metal2 s 137712 953270 137768 953750 0 FreeSans 400 90 0 0 gpio_oeb[21]
port 180 nsew
flabel metal2 s 140840 953270 140896 953750 0 FreeSans 400 90 0 0 gpio_out[21]
port 136 nsew
flabel metal2 s 150040 953270 150096 953750 0 FreeSans 400 90 0 0 gpio_slow_sel[21]
port 356 nsew
flabel metal2 s 139000 953270 139056 953750 0 FreeSans 400 90 0 0 gpio_vtrip_sel[21]
port 312 nsew
flabel metal2 151354 -424 151410 56 0 FreeSans 400 270 0 0 gpio_analog_pol[38]
port 515 nsew
flabel metal2 150066 -424 150122 56 0 FreeSans 400 270 0 0 gpio_analog_en[38]
port 427 nsew
flabel metal2 151906 -424 151962 56 0 FreeSans 400 270 0 0 gpio_inp_dis[38]
port 207 nsew
flabel metal2 154390 -424 154446 56 0 FreeSans 400 270 0 0 gpio_analog_sel[38]
port 471 nsew
flabel metal2 155034 -424 155090 56 0 FreeSans 400 270 0 0 gpio_dm2[38]
port 647 nsew
flabel metal2 155678 -424 155734 56 0 FreeSans 400 270 0 0 gpio_holdover[38]
port 383 nsew
flabel metal2 156230 -424 156286 56 0 FreeSans 400 270 0 0 gpio_out[38]
port 119 nsew
flabel metal2 158070 -424 158126 56 0 FreeSans 400 270 0 0 gpio_vtrip_sel[38]
port 295 nsew
flabel metal2 158714 -424 158770 56 0 FreeSans 400 270 0 0 gpio_ib_mode_sel[38]
port 251 nsew
flabel metal2 159358 -424 159414 56 0 FreeSans 400 270 0 0 gpio_oeb[38]
port 163 nsew
flabel metal2 253790 -424 253846 56 0 FreeSans 400 270 0 0 gpio_in[39]
port 690 nsew
flabel metal2 255630 -424 255686 56 0 FreeSans 400 270 0 0 gpio_slow_sel[39]
port 338 nsew
flabel metal2 257470 -424 257526 56 0 FreeSans 400 270 0 0 gpio_dm1[39]
port 602 nsew
flabel metal2 259310 -424 259366 56 0 FreeSans 400 270 0 0 gpio_dm0[39]
port 558 nsew
flabel metal2 259954 -424 260010 56 0 FreeSans 400 270 0 0 gpio_analog_pol[39]
port 514 nsew
flabel metal2 258666 -424 258722 56 0 FreeSans 400 270 0 0 gpio_analog_en[39]
port 426 nsew
flabel metal2 260506 -424 260562 56 0 FreeSans 400 270 0 0 gpio_inp_dis[39]
port 206 nsew
flabel metal2 262990 -424 263046 56 0 FreeSans 400 270 0 0 gpio_analog_sel[39]
port 470 nsew
flabel metal2 263634 -424 263690 56 0 FreeSans 400 270 0 0 gpio_dm2[39]
port 646 nsew
flabel metal2 264278 -424 264334 56 0 FreeSans 400 270 0 0 gpio_holdover[39]
port 382 nsew
flabel metal2 264830 -424 264886 56 0 FreeSans 400 270 0 0 gpio_out[39]
port 118 nsew
flabel metal2 266670 -424 266726 56 0 FreeSans 400 270 0 0 gpio_vtrip_sel[39]
port 294 nsew
flabel metal2 267314 -424 267370 56 0 FreeSans 400 270 0 0 gpio_ib_mode_sel[39]
port 250 nsew
flabel metal2 267958 -424 268014 56 0 FreeSans 400 270 0 0 gpio_oeb[39]
port 162 nsew
flabel metal2 308590 -424 308646 56 0 FreeSans 400 270 0 0 gpio_in[40]
port 689 nsew
flabel metal2 310430 -424 310486 56 0 FreeSans 400 270 0 0 gpio_slow_sel[40]
port 337 nsew
flabel metal2 312270 -424 312326 56 0 FreeSans 400 270 0 0 gpio_dm1[40]
port 601 nsew
flabel metal2 314110 -424 314166 56 0 FreeSans 400 270 0 0 gpio_dm0[40]
port 557 nsew
flabel metal2 314754 -424 314810 56 0 FreeSans 400 270 0 0 gpio_analog_pol[40]
port 513 nsew
flabel metal2 313466 -424 313522 56 0 FreeSans 400 270 0 0 gpio_analog_en[40]
port 425 nsew
flabel metal2 315306 -424 315362 56 0 FreeSans 400 270 0 0 gpio_inp_dis[40]
port 205 nsew
flabel metal2 317790 -424 317846 56 0 FreeSans 400 270 0 0 gpio_analog_sel[40]
port 469 nsew
flabel metal2 318434 -424 318490 56 0 FreeSans 400 270 0 0 gpio_dm2[40]
port 645 nsew
flabel metal2 319078 -424 319134 56 0 FreeSans 400 270 0 0 gpio_holdover[40]
port 381 nsew
flabel metal2 319630 -424 319686 56 0 FreeSans 400 270 0 0 gpio_out[40]
port 117 nsew
flabel metal2 321470 -424 321526 56 0 FreeSans 400 270 0 0 gpio_vtrip_sel[40]
port 293 nsew
flabel metal2 322114 -424 322170 56 0 FreeSans 400 270 0 0 gpio_ib_mode_sel[40]
port 249 nsew
flabel metal2 322758 -424 322814 56 0 FreeSans 400 270 0 0 gpio_oeb[40]
port 161 nsew
flabel metal2 363390 -424 363446 56 0 FreeSans 400 270 0 0 gpio_in[41]
port 688 nsew
flabel metal2 365230 -424 365286 56 0 FreeSans 400 270 0 0 gpio_slow_sel[41]
port 336 nsew
flabel metal2 367070 -424 367126 56 0 FreeSans 400 270 0 0 gpio_dm1[41]
port 600 nsew
flabel metal2 368910 -424 368966 56 0 FreeSans 400 270 0 0 gpio_dm0[41]
port 556 nsew
flabel metal2 369554 -424 369610 56 0 FreeSans 400 270 0 0 gpio_analog_pol[41]
port 512 nsew
flabel metal2 368266 -424 368322 56 0 FreeSans 400 270 0 0 gpio_analog_en[41]
port 424 nsew
flabel metal2 370106 -424 370162 56 0 FreeSans 400 270 0 0 gpio_inp_dis[41]
port 204 nsew
flabel metal2 372590 -424 372646 56 0 FreeSans 400 270 0 0 gpio_analog_sel[41]
port 468 nsew
flabel metal2 373234 -424 373290 56 0 FreeSans 400 270 0 0 gpio_dm2[41]
port 644 nsew
flabel metal2 373878 -424 373934 56 0 FreeSans 400 270 0 0 gpio_holdover[41]
port 380 nsew
flabel metal2 374430 -424 374486 56 0 FreeSans 400 270 0 0 gpio_out[41]
port 116 nsew
flabel metal2 376270 -424 376326 56 0 FreeSans 400 270 0 0 gpio_vtrip_sel[41]
port 292 nsew
flabel metal2 376914 -424 376970 56 0 FreeSans 400 270 0 0 gpio_ib_mode_sel[41]
port 248 nsew
flabel metal2 377558 -424 377614 56 0 FreeSans 400 270 0 0 gpio_oeb[41]
port 160 nsew
flabel metal2 418190 -424 418246 56 0 FreeSans 400 270 0 0 gpio_in[42]
port 687 nsew
flabel metal2 420030 -424 420086 56 0 FreeSans 400 270 0 0 gpio_slow_sel[42]
port 335 nsew
flabel metal2 421870 -424 421926 56 0 FreeSans 400 270 0 0 gpio_dm1[42]
port 599 nsew
flabel metal2 423710 -424 423766 56 0 FreeSans 400 270 0 0 gpio_dm0[42]
port 555 nsew
flabel metal2 424354 -424 424410 56 0 FreeSans 400 270 0 0 gpio_analog_pol[42]
port 511 nsew
flabel metal2 423066 -424 423122 56 0 FreeSans 400 270 0 0 gpio_analog_en[42]
port 423 nsew
flabel metal2 424906 -424 424962 56 0 FreeSans 400 270 0 0 gpio_inp_dis[42]
port 203 nsew
flabel metal2 427390 -424 427446 56 0 FreeSans 400 270 0 0 gpio_analog_sel[42]
port 467 nsew
flabel metal2 428034 -424 428090 56 0 FreeSans 400 270 0 0 gpio_dm2[42]
port 643 nsew
flabel metal2 428678 -424 428734 56 0 FreeSans 400 270 0 0 gpio_holdover[42]
port 379 nsew
flabel metal2 429230 -424 429286 56 0 FreeSans 400 270 0 0 gpio_out[42]
port 115 nsew
flabel metal2 431070 -424 431126 56 0 FreeSans 400 270 0 0 gpio_vtrip_sel[42]
port 291 nsew
flabel metal2 431714 -424 431770 56 0 FreeSans 400 270 0 0 gpio_ib_mode_sel[42]
port 247 nsew
flabel metal2 432358 -424 432414 56 0 FreeSans 400 270 0 0 gpio_oeb[42]
port 159 nsew
flabel metal2 472990 -424 473046 56 0 FreeSans 400 270 0 0 gpio_in[43]
port 686 nsew
flabel metal2 474830 -424 474886 56 0 FreeSans 400 270 0 0 gpio_slow_sel[43]
port 334 nsew
flabel metal2 476670 -424 476726 56 0 FreeSans 400 270 0 0 gpio_dm1[43]
port 598 nsew
flabel metal2 478510 -424 478566 56 0 FreeSans 400 270 0 0 gpio_dm0[43]
port 554 nsew
flabel metal2 479154 -424 479210 56 0 FreeSans 400 270 0 0 gpio_analog_pol[43]
port 510 nsew
flabel metal2 477866 -424 477922 56 0 FreeSans 400 270 0 0 gpio_analog_en[43]
port 422 nsew
flabel metal2 479706 -424 479762 56 0 FreeSans 400 270 0 0 gpio_inp_dis[43]
port 202 nsew
flabel metal2 482190 -424 482246 56 0 FreeSans 400 270 0 0 gpio_analog_sel[43]
port 466 nsew
flabel metal2 482834 -424 482890 56 0 FreeSans 400 270 0 0 gpio_dm2[43]
port 642 nsew
flabel metal2 483478 -424 483534 56 0 FreeSans 400 270 0 0 gpio_holdover[43]
port 378 nsew
flabel metal2 484030 -424 484086 56 0 FreeSans 400 270 0 0 gpio_out[43]
port 114 nsew
flabel metal2 486514 -424 486570 56 0 FreeSans 400 270 0 0 gpio_ib_mode_sel[43]
port 246 nsew
flabel metal2 487158 -424 487214 56 0 FreeSans 400 270 0 0 gpio_oeb[43]
port 158 nsew
flabel metal2 s 584160 953270 584216 953750 0 FreeSans 400 90 0 0 gpio_in_h[15]
port 758 nsew
flabel metal2 s 482360 953270 482416 953750 0 FreeSans 400 90 0 0 gpio_in_h[16]
port 757 nsew
flabel metal2 s 430960 953270 431016 953750 0 FreeSans 400 90 0 0 gpio_in_h[17]
port 756 nsew
flabel metal2 s 341960 953270 342016 953750 0 FreeSans 400 90 0 0 gpio_in_h[18]
port 755 nsew
flabel metal2 s 240160 953270 240216 953750 0 FreeSans 400 90 0 0 gpio_in_h[19]
port 754 nsew
flabel metal2 s 188560 953270 188616 953750 0 FreeSans 400 90 0 0 gpio_in_h[20]
port 753 nsew
flabel metal2 s 137160 953270 137216 953750 0 FreeSans 400 90 0 0 gpio_in_h[21]
port 752 nsew
flabel metal2 s 85760 953270 85816 953750 0 FreeSans 400 90 0 0 gpio_in_h[22]
port 751 nsew
flabel metal2 s 34360 953270 34416 953750 0 FreeSans 400 90 0 0 gpio_in_h[23]
port 750 nsew
flabel metal2 s 159910 -424 159966 56 0 FreeSans 400 90 0 0 gpio_in_h[38]
port 735 nsew
flabel metal2 s 268510 -424 268566 56 0 FreeSans 400 90 0 0 gpio_in_h[39]
port 734 nsew
flabel metal2 s 323310 -424 323366 56 0 FreeSans 400 90 0 0 gpio_in_h[40]
port 733 nsew
flabel metal2 s 378110 -424 378166 56 0 FreeSans 400 90 0 0 gpio_in_h[41]
port 732 nsew
flabel metal2 s 432910 -424 432966 56 0 FreeSans 400 90 0 0 gpio_in_h[42]
port 731 nsew
flabel metal2 s 487710 -424 487766 56 0 FreeSans 400 90 0 0 gpio_in_h[43]
port 730 nsew
flabel metal3 633270 422810 633770 427472 0 FreeSans 3200 90 0 0 vccd1
port 28 nsew
flabel metal3 s 633270 786384 633770 791164 0 FreeSans 3200 90 0 0 vdda1
port 24 nsew
flabel metal3 s 633270 471784 633770 476564 0 FreeSans 3200 90 0 0 vdda1
port 24 nsew
flabel metal3 s 633270 383584 633770 388364 0 FreeSans 3200 90 0 0 vssa1
port 26 nsew
flabel metal3 s 533562 953270 538342 953770 0 FreeSans 3200 0 0 0 vssa1
port 26 nsew
flabel metal3 291362 953270 296142 953770 0 FreeSans 3200 0 0 0 vssio
port 19 nsew
flabel metal3 -444 880014 56 884804 0 FreeSans 3200 90 0 0 vccd2
port 29 nsew
flabel metal3 -444 827762 56 832542 0 FreeSans 3200 90 0 0 vddio
port 18 nsew
flabel metal3 -444 785562 56 790342 0 FreeSans 3200 90 0 0 vssa2
port 27 nsew
flabel metal3 -444 440962 56 445742 0 FreeSans 3200 90 0 0 vdda2
port 25 nsew
flabel metal3 -444 68162 56 72942 0 FreeSans 3200 90 0 0 vddio
port 18 nsew
flabel metal3 536984 -444 541764 56 0 FreeSans 3200 0 0 0 vssio
port 19 nsew
flabel metal3 590784 -444 595564 56 0 FreeSans 3200 0 0 0 vdda
port 22 nsew
flabel comment s 107715 141850 108715 141850 0 FreeSans 1120000 60 0 0 example
flabel metal3 s 633270 556035 633750 556249 0 FreeSans 400 0 0 0 analog_noesd_io[8]
port 941 nsew
flabel metal3 -264 906644 56 906704 0 FreeSans 400 0 0 0 gpio_loopback_one[24]
port 837 nsew
flabel metal3 -264 736644 56 736704 0 FreeSans 400 0 0 0 gpio_loopback_one[25]
port 836 nsew
flabel metal3 -264 693644 56 693704 0 FreeSans 400 0 0 0 gpio_loopback_one[26]
port 835 nsew
flabel metal3 -264 650644 56 650704 0 FreeSans 400 0 0 0 gpio_loopback_one[27]
port 834 nsew
flabel metal3 -264 607644 56 607704 0 FreeSans 400 0 0 0 gpio_loopback_one[28]
port 833 nsew
flabel metal3 -264 564644 56 564704 0 FreeSans 400 0 0 0 gpio_loopback_one[29]
port 832 nsew
flabel metal3 -264 521644 56 521704 0 FreeSans 400 0 0 0 gpio_loopback_one[30]
port 831 nsew
flabel metal3 -264 478644 56 478704 0 FreeSans 400 0 0 0 gpio_loopback_one[31]
port 830 nsew
flabel metal3 -264 349644 56 349704 0 FreeSans 400 0 0 0 gpio_loopback_one[32]
port 829 nsew
flabel metal3 -264 306644 56 306704 0 FreeSans 400 0 0 0 gpio_loopback_one[33]
port 828 nsew
flabel metal3 -264 263644 56 263704 0 FreeSans 400 0 0 0 gpio_loopback_one[34]
port 827 nsew
flabel metal3 -264 220644 56 220704 0 FreeSans 400 0 0 0 gpio_loopback_one[35]
port 826 nsew
flabel metal3 -264 177644 56 177704 0 FreeSans 400 0 0 0 gpio_loopback_one[36]
port 825 nsew
flabel metal3 -264 134644 56 134704 0 FreeSans 400 0 0 0 gpio_loopback_one[37]
port 824 nsew
flabel metal2 s 488380 -260 488432 56 0 FreeSans 400 90 0 0 gpio_loopback_one[43]
port 818 nsew
flabel metal2 s 492635 -260 492687 56 0 FreeSans 400 90 0 0 gpio_loopback_zero[43]
port 774 nsew
flabel metal2 s 433580 -260 433632 56 0 FreeSans 400 90 0 0 gpio_loopback_one[42]
port 819 nsew
flabel metal2 s 437778 -260 437830 56 0 FreeSans 400 90 0 0 gpio_loopback_zero[42]
port 775 nsew
flabel metal2 s 378780 -260 378832 56 0 FreeSans 400 90 0 0 gpio_loopback_one[41]
port 820 nsew
flabel metal2 s 382978 -260 383030 56 0 FreeSans 400 90 0 0 gpio_loopback_zero[41]
port 776 nsew
flabel metal2 s 323980 -260 324032 56 0 FreeSans 400 90 0 0 gpio_loopback_one[40]
port 821 nsew
flabel metal2 s 328165 -282 328217 34 0 FreeSans 400 90 0 0 gpio_loopback_zero[40]
port 777 nsew
flabel metal2 s 269180 -260 269232 56 0 FreeSans 400 90 0 0 gpio_loopback_one[39]
port 822 nsew
flabel metal2 s 273360 -260 273412 56 0 FreeSans 400 90 0 0 gpio_loopback_zero[39]
port 778 nsew
flabel metal2 s 160580 -260 160632 56 0 FreeSans 400 90 0 0 gpio_loopback_one[38]
port 823 nsew
flabel metal2 s 163791 -259 163843 57 0 FreeSans 400 90 0 0 gpio_loopback_zero[38]
port 779 nsew
flabel metal2 s 110164 -116 110220 56 0 FreeSans 400 90 0 0 resetb_l
port 37 nsew
flabel metal2 s 99571 -90 99637 56 0 FreeSans 400 90 0 0 resetb_h
port 36 nsew
flabel metal3 -284 53372 56 53442 0 FreeSans 400 0 0 0 por_l
port 35 nsew
flabel metal3 -284 53595 56 53665 0 FreeSans 400 0 0 0 porb_l
port 34 nsew
flabel metal2 s 605082 -260 605134 56 0 FreeSans 400 90 0 0 mask_rev[0]
port 69 nsew
flabel metal3 -284 53147 56 53217 0 FreeSans 400 0 0 0 porb_h
port 33 nsew
flabel metal2 578298 953270 578358 953726 0 FreeSans 400 90 0 0 gpio_loopback_one[15]
port 846 nsew
flabel metal2 478898 953270 478958 953726 0 FreeSans 400 90 0 0 gpio_loopback_one[16]
port 845 nsew
flabel metal2 427698 953270 427758 953726 0 FreeSans 400 90 0 0 gpio_loopback_one[17]
port 844 nsew
flabel metal2 338698 953270 338758 953726 0 FreeSans 400 90 0 0 gpio_loopback_one[18]
port 843 nsew
flabel metal2 234298 953270 234358 953726 0 FreeSans 400 90 0 0 gpio_loopback_one[19]
port 842 nsew
flabel metal2 183098 953270 183158 953726 0 FreeSans 400 90 0 0 gpio_loopback_one[20]
port 841 nsew
flabel metal2 131898 953270 131958 953726 0 FreeSans 400 90 0 0 gpio_loopback_one[21]
port 840 nsew
flabel metal2 80698 953270 80758 953726 0 FreeSans 400 90 0 0 gpio_loopback_one[22]
port 839 nsew
flabel metal2 29498 953270 29558 953726 0 FreeSans 400 90 0 0 gpio_loopback_one[23]
port 838 nsew
flabel metal3 633270 523005 633590 523067 0 FreeSans 400 0 0 0 gpio_loopback_one[7]
port 854 nsew
flabel metal3 633270 346005 633590 346067 0 FreeSans 400 0 0 0 gpio_loopback_one[6]
port 855 nsew
flabel metal3 633270 301005 633590 301067 0 FreeSans 400 0 0 0 gpio_loopback_one[5]
port 856 nsew
flabel metal3 633270 256005 633590 256067 0 FreeSans 400 0 0 0 gpio_loopback_one[4]
port 857 nsew
flabel metal3 633270 211005 633590 211067 0 FreeSans 400 0 0 0 gpio_loopback_one[3]
port 858 nsew
flabel metal3 633270 166005 633590 166067 0 FreeSans 400 0 0 0 gpio_loopback_one[2]
port 859 nsew
flabel metal3 633270 121005 633590 121067 0 FreeSans 400 0 0 0 gpio_loopback_one[1]
port 860 nsew
flabel metal3 633270 76005 633590 76067 0 FreeSans 400 0 0 0 gpio_loopback_one[0]
port 861 nsew
flabel metal2 s 605978 -260 606030 56 0 FreeSans 400 90 0 0 mask_rev[4]
port 65 nsew
flabel metal2 s 606202 -260 606254 56 0 FreeSans 400 90 0 0 mask_rev[5]
port 64 nsew
flabel metal2 s 606426 -260 606478 56 0 FreeSans 400 90 0 0 mask_rev[6]
port 63 nsew
flabel metal2 s 606650 -260 606702 56 0 FreeSans 400 90 0 0 mask_rev[7]
port 62 nsew
flabel metal2 s 606874 -260 606926 56 0 FreeSans 400 90 0 0 mask_rev[8]
port 61 nsew
flabel metal2 s 607098 -260 607150 56 0 FreeSans 400 90 0 0 mask_rev[9]
port 60 nsew
flabel metal2 s 607322 -260 607374 56 0 FreeSans 400 90 0 0 mask_rev[10]
port 59 nsew
flabel metal2 s 607546 -260 607598 56 0 FreeSans 400 90 0 0 mask_rev[11]
port 58 nsew
flabel metal2 s 607770 -260 607822 56 0 FreeSans 400 90 0 0 mask_rev[12]
port 57 nsew
flabel metal2 s 607994 -260 608046 56 0 FreeSans 400 90 0 0 mask_rev[13]
port 56 nsew
flabel metal2 s 608218 -260 608270 56 0 FreeSans 400 90 0 0 mask_rev[14]
port 55 nsew
flabel metal2 s 608442 -260 608494 56 0 FreeSans 400 90 0 0 mask_rev[15]
port 54 nsew
flabel metal2 s 608666 -260 608718 56 0 FreeSans 400 90 0 0 mask_rev[16]
port 53 nsew
flabel metal2 s 608890 -260 608942 56 0 FreeSans 400 90 0 0 mask_rev[17]
port 52 nsew
flabel metal2 s 609114 -260 609166 56 0 FreeSans 400 90 0 0 mask_rev[18]
port 51 nsew
flabel metal2 s 609338 -260 609390 56 0 FreeSans 400 90 0 0 mask_rev[19]
port 50 nsew
flabel metal2 s 609562 -260 609614 56 0 FreeSans 400 90 0 0 mask_rev[20]
port 49 nsew
flabel metal2 s 609786 -260 609838 56 0 FreeSans 400 90 0 0 mask_rev[21]
port 48 nsew
flabel metal2 s 610010 -260 610062 56 0 FreeSans 400 90 0 0 mask_rev[22]
port 47 nsew
flabel metal2 s 610234 -260 610286 56 0 FreeSans 400 90 0 0 mask_rev[23]
port 46 nsew
flabel metal2 s 610458 -260 610510 56 0 FreeSans 400 90 0 0 mask_rev[24]
port 45 nsew
flabel metal2 s 610682 -260 610734 56 0 FreeSans 400 90 0 0 mask_rev[25]
port 44 nsew
flabel metal2 s 610906 -260 610958 56 0 FreeSans 400 90 0 0 mask_rev[26]
port 43 nsew
flabel metal2 s 611130 -260 611182 56 0 FreeSans 400 90 0 0 mask_rev[27]
port 42 nsew
flabel metal2 s 611354 -260 611406 56 0 FreeSans 400 90 0 0 mask_rev[28]
port 41 nsew
flabel metal2 s 611578 -260 611630 56 0 FreeSans 400 90 0 0 mask_rev[29]
port 40 nsew
flabel metal2 s 611802 -260 611854 56 0 FreeSans 400 90 0 0 mask_rev[30]
port 39 nsew
flabel metal2 s 612026 -260 612078 56 0 FreeSans 400 90 0 0 mask_rev[31]
port 38 nsew
flabel metal2 s 605754 -260 605806 56 0 FreeSans 400 90 0 0 mask_rev[3]
port 66 nsew
flabel metal2 s 605530 -260 605582 56 0 FreeSans 400 90 0 0 mask_rev[2]
port 67 nsew
flabel metal2 s 605306 -260 605358 56 0 FreeSans 400 90 0 0 mask_rev[1]
port 68 nsew
flabel metal3 -264 734644 56 734704 0 FreeSans 400 0 0 0 gpio_loopback_zero[25]
port 792 nsew
flabel metal3 -264 648644 56 648704 0 FreeSans 400 0 0 0 gpio_loopback_zero[27]
port 790 nsew
flabel metal3 -264 562644 56 562704 0 FreeSans 400 0 0 0 gpio_loopback_zero[29]
port 788 nsew
flabel metal3 -264 476644 56 476704 0 FreeSans 400 0 0 0 gpio_loopback_zero[31]
port 786 nsew
flabel metal3 -264 304644 56 304704 0 FreeSans 400 0 0 0 gpio_loopback_zero[33]
port 784 nsew
flabel metal3 -264 218644 56 218704 0 FreeSans 400 0 0 0 gpio_loopback_zero[35]
port 782 nsew
flabel metal3 -264 132644 56 132704 0 FreeSans 400 0 0 0 gpio_loopback_zero[37]
port 780 nsew
flabel metal3 -264 904644 56 904704 0 FreeSans 400 0 0 0 gpio_loopback_zero[24]
port 793 nsew
flabel metal3 -264 691644 56 691704 0 FreeSans 400 0 0 0 gpio_loopback_zero[26]
port 791 nsew
flabel metal3 -264 605644 56 605704 0 FreeSans 400 0 0 0 gpio_loopback_zero[28]
port 789 nsew
flabel metal3 -264 519644 56 519704 0 FreeSans 400 0 0 0 gpio_loopback_zero[30]
port 787 nsew
flabel metal3 -264 347644 56 347704 0 FreeSans 400 0 0 0 gpio_loopback_zero[32]
port 785 nsew
flabel metal3 -264 261644 56 261704 0 FreeSans 400 0 0 0 gpio_loopback_zero[34]
port 783 nsew
flabel metal3 -264 175644 56 175704 0 FreeSans 400 0 0 0 gpio_loopback_zero[36]
port 781 nsew
flabel metal2 27497 953270 27557 953726 0 FreeSans 400 90 0 0 gpio_loopback_zero[23]
port 794 nsew
flabel metal2 78697 953270 78757 953726 0 FreeSans 400 90 0 0 gpio_loopback_zero[22]
port 795 nsew
flabel metal2 129897 953270 129957 953726 0 FreeSans 400 90 0 0 gpio_loopback_zero[21]
port 796 nsew
flabel metal2 181097 953270 181157 953726 0 FreeSans 400 90 0 0 gpio_loopback_zero[20]
port 797 nsew
flabel metal2 232297 953270 232357 953726 0 FreeSans 400 90 0 0 gpio_loopback_zero[19]
port 798 nsew
flabel metal2 336697 953270 336757 953726 0 FreeSans 400 90 0 0 gpio_loopback_zero[18]
port 799 nsew
flabel metal2 425697 953270 425757 953726 0 FreeSans 400 90 0 0 gpio_loopback_zero[17]
port 800 nsew
flabel metal2 476897 953270 476957 953726 0 FreeSans 400 90 0 0 gpio_loopback_zero[16]
port 801 nsew
flabel metal2 576297 953270 576357 953726 0 FreeSans 400 90 0 0 gpio_loopback_zero[15]
port 802 nsew
flabel metal2 147030 -424 147086 56 0 FreeSans 400 270 0 0 gpio_slow_sel[38]
port 339 nsew
flabel metal2 145190 -424 145246 56 0 FreeSans 400 270 0 0 gpio_in[38]
port 691 nsew
flabel metal3 46784 -444 51564 56 0 FreeSans 3200 0 0 0 vssa
port 23 nsew
flabel metal3 633270 61238 633750 61366 0 FreeSans 400 0 0 0 analog_io[0]
port 905 nsew
flabel metal3 633270 63035 633750 63249 0 FreeSans 400 0 0 0 analog_noesd_io[0]
port 949 nsew
flabel metal3 633270 108235 633750 108449 0 FreeSans 400 0 0 0 analog_noesd_io[1]
port 948 nsew
flabel metal3 633270 106438 633750 106566 0 FreeSans 400 0 0 0 analog_io[1]
port 904 nsew
flabel metal3 633270 151438 633750 151566 0 FreeSans 400 0 0 0 analog_io[2]
port 903 nsew
flabel metal3 633270 153235 633750 153449 0 FreeSans 400 0 0 0 analog_noesd_io[2]
port 947 nsew
flabel metal3 633270 196638 633750 196766 0 FreeSans 400 0 0 0 analog_io[3]
port 902 nsew
flabel metal3 633270 198435 633750 198649 0 FreeSans 400 0 0 0 analog_noesd_io[3]
port 946 nsew
flabel metal3 633270 241638 633750 241766 0 FreeSans 400 0 0 0 analog_io[4]
port 901 nsew
flabel metal3 633270 243435 633750 243649 0 FreeSans 400 0 0 0 analog_noesd_io[4]
port 945 nsew
flabel metal3 633270 286638 633750 286766 0 FreeSans 400 0 0 0 analog_io[5]
port 900 nsew
flabel metal3 633270 288435 633750 288649 0 FreeSans 400 0 0 0 analog_noesd_io[5]
port 944 nsew
flabel metal3 633270 331838 633750 331966 0 FreeSans 400 0 0 0 analog_io[6]
port 899 nsew
flabel metal3 633270 333635 633750 333849 0 FreeSans 400 0 0 0 analog_noesd_io[6]
port 943 nsew
flabel metal3 s 633270 509038 633750 509166 0 FreeSans 400 0 0 0 analog_io[7]
port 898 nsew
flabel metal3 s 633270 510835 633750 511049 0 FreeSans 400 0 0 0 analog_noesd_io[7]
port 942 nsew
flabel metal3 s 633270 554238 633750 554366 0 FreeSans 400 0 0 0 analog_io[8]
port 897 nsew
flabel metal3 s 633270 599238 633750 599366 0 FreeSans 400 0 0 0 analog_io[9]
port 896 nsew
flabel metal3 s 633270 601035 633750 601249 0 FreeSans 400 0 0 0 analog_noesd_io[9]
port 940 nsew
flabel metal3 s 633270 644438 633750 644566 0 FreeSans 400 0 0 0 analog_io[10]
port 895 nsew
flabel metal3 s 633270 646235 633750 646449 0 FreeSans 400 0 0 0 analog_noesd_io[10]
port 939 nsew
flabel metal3 s 633270 689438 633750 689566 0 FreeSans 400 0 0 0 analog_io[11]
port 894 nsew
flabel metal3 s 633270 691235 633750 691449 0 FreeSans 400 0 0 0 analog_noesd_io[11]
port 938 nsew
flabel metal3 s 633270 734438 633750 734566 0 FreeSans 400 0 0 0 analog_io[12]
port 893 nsew
flabel metal3 s 633270 823638 633750 823766 0 FreeSans 400 0 0 0 analog_io[13]
port 892 nsew
flabel metal3 s 633270 912838 633750 912966 0 FreeSans 400 0 0 0 analog_io[14]
port 891 nsew
flabel metal3 s 633270 736235 633750 736449 0 FreeSans 400 0 0 0 analog_noesd_io[12]
port 937 nsew
flabel metal3 s 633270 825435 633750 825649 0 FreeSans 400 0 0 0 analog_noesd_io[13]
port 936 nsew
flabel metal3 s 633270 914635 633750 914849 0 FreeSans 400 0 0 0 analog_noesd_io[14]
port 935 nsew
flabel metal2 s 596360 953270 596488 953750 0 FreeSans 400 90 0 0 analog_io[15]
port 890 nsew
flabel metal2 s 494560 953270 494688 953750 0 FreeSans 400 90 0 0 analog_io[16]
port 889 nsew
flabel metal2 s 443160 953270 443288 953750 0 FreeSans 400 90 0 0 analog_io[17]
port 888 nsew
flabel metal2 s 354160 953270 354288 953750 0 FreeSans 400 90 0 0 analog_io[18]
port 887 nsew
flabel metal2 s 252360 953270 252488 953750 0 FreeSans 400 90 0 0 analog_io[19]
port 886 nsew
flabel metal2 s 200760 953270 200888 953750 0 FreeSans 400 90 0 0 analog_io[20]
port 885 nsew
flabel metal2 s 149360 953270 149488 953750 0 FreeSans 400 90 0 0 analog_io[21]
port 884 nsew
flabel metal2 s 97960 953270 98088 953750 0 FreeSans 400 90 0 0 analog_io[22]
port 883 nsew
flabel metal2 s 46560 953270 46688 953750 0 FreeSans 400 90 0 0 analog_io[23]
port 882 nsew
flabel metal2 s 594477 953270 594691 953750 0 FreeSans 400 90 0 0 analog_noesd_io[15]
port 934 nsew
flabel metal2 s 492677 953270 492891 953750 0 FreeSans 400 90 0 0 analog_noesd_io[16]
port 933 nsew
flabel metal2 s 441277 953270 441491 953750 0 FreeSans 400 90 0 0 analog_noesd_io[17]
port 932 nsew
flabel metal2 s 352277 953270 352491 953750 0 FreeSans 400 90 0 0 analog_noesd_io[18]
port 931 nsew
flabel metal2 s 250477 953270 250691 953750 0 FreeSans 400 90 0 0 analog_noesd_io[19]
port 930 nsew
flabel metal2 s 198877 953270 199091 953750 0 FreeSans 400 90 0 0 analog_noesd_io[20]
port 929 nsew
flabel metal2 s 147477 953270 147691 953750 0 FreeSans 400 90 0 0 analog_noesd_io[21]
port 928 nsew
flabel metal2 s 96077 953270 96291 953750 0 FreeSans 400 90 0 0 analog_noesd_io[22]
port 927 nsew
flabel metal2 s 44677 953270 44891 953750 0 FreeSans 400 90 0 0 analog_noesd_io[23]
port 926 nsew
flabel metal3 s -424 754760 56 754888 0 FreeSans 400 0 0 0 analog_io[25]
port 880 nsew
flabel metal3 s -424 711560 56 711688 0 FreeSans 400 0 0 0 analog_io[26]
port 879 nsew
flabel metal3 s -424 668360 56 668488 0 FreeSans 400 0 0 0 analog_io[27]
port 878 nsew
flabel metal3 s -424 625160 56 625288 0 FreeSans 400 0 0 0 analog_io[28]
port 877 nsew
flabel metal3 s -424 581960 56 582088 0 FreeSans 400 0 0 0 analog_io[29]
port 876 nsew
flabel metal3 s -424 538760 56 538888 0 FreeSans 400 0 0 0 analog_io[30]
port 875 nsew
flabel metal3 s -424 495560 56 495688 0 FreeSans 400 0 0 0 analog_io[31]
port 874 nsew
flabel metal3 s -424 367960 56 368088 0 FreeSans 400 0 0 0 analog_io[32]
port 873 nsew
flabel metal3 s -424 324760 56 324888 0 FreeSans 400 0 0 0 analog_io[33]
port 872 nsew
flabel metal3 s -424 281560 56 281688 0 FreeSans 400 0 0 0 analog_io[34]
port 871 nsew
flabel metal3 s -424 238360 56 238488 0 FreeSans 400 0 0 0 analog_io[35]
port 870 nsew
flabel metal3 s -424 195160 56 195288 0 FreeSans 400 0 0 0 analog_io[36]
port 869 nsew
flabel metal3 s -424 151960 56 152088 0 FreeSans 400 0 0 0 analog_io[37]
port 868 nsew
flabel metal3 s -424 752877 56 753091 0 FreeSans 400 0 0 0 analog_noesd_io[25]
port 924 nsew
flabel metal3 s -424 709677 56 709891 0 FreeSans 400 0 0 0 analog_noesd_io[26]
port 923 nsew
flabel metal3 s -424 666477 56 666691 0 FreeSans 400 0 0 0 analog_noesd_io[27]
port 922 nsew
flabel metal3 s -424 623277 56 623491 0 FreeSans 400 0 0 0 analog_noesd_io[28]
port 921 nsew
flabel metal3 s -424 580077 56 580291 0 FreeSans 400 0 0 0 analog_noesd_io[29]
port 920 nsew
flabel metal3 s -424 536877 56 537091 0 FreeSans 400 0 0 0 analog_noesd_io[30]
port 919 nsew
flabel metal3 s -424 366077 56 366291 0 FreeSans 400 0 0 0 analog_noesd_io[32]
port 917 nsew
flabel metal3 s -424 322877 56 323091 0 FreeSans 400 0 0 0 analog_noesd_io[33]
port 916 nsew
flabel metal3 s -424 279677 56 279891 0 FreeSans 400 0 0 0 analog_noesd_io[34]
port 915 nsew
flabel metal3 s -424 236477 56 236691 0 FreeSans 400 0 0 0 analog_noesd_io[35]
port 914 nsew
flabel metal3 s -424 193277 56 193491 0 FreeSans 400 0 0 0 analog_noesd_io[36]
port 913 nsew
flabel metal3 s -424 150077 56 150291 0 FreeSans 400 0 0 0 analog_noesd_io[37]
port 912 nsew
flabel metal2 s 256238 -424 256366 56 0 FreeSans 400 90 0 0 analog_io[39]
port 866 nsew
flabel metal2 s 311038 -424 311166 56 0 FreeSans 400 90 0 0 analog_io[40]
port 865 nsew
flabel metal2 s 365838 -424 365966 56 0 FreeSans 400 90 0 0 analog_io[41]
port 864 nsew
flabel metal2 s 420638 -424 420766 56 0 FreeSans 400 90 0 0 analog_io[42]
port 863 nsew
flabel metal2 s 475438 -424 475566 56 0 FreeSans 400 90 0 0 analog_io[43]
port 862 nsew
flabel metal2 s 258035 -424 258249 56 0 FreeSans 400 90 0 0 analog_noesd_io[39]
port 910 nsew
flabel metal2 s 312835 -424 313049 56 0 FreeSans 400 90 0 0 analog_noesd_io[40]
port 909 nsew
flabel metal2 s 367635 -424 367849 56 0 FreeSans 400 90 0 0 analog_noesd_io[41]
port 908 nsew
flabel metal2 s 422435 -424 422649 56 0 FreeSans 400 90 0 0 analog_noesd_io[42]
port 907 nsew
flabel metal2 s 477235 -424 477449 56 0 FreeSans 400 90 0 0 analog_noesd_io[43]
port 906 nsew
flabel metal2 s 149435 -424 149649 56 0 FreeSans 400 90 0 0 analog_noesd_io[38]
port 911 nsew
flabel metal2 s 147638 -424 147766 56 0 FreeSans 400 90 0 0 analog_io[38]
port 867 nsew
flabel metal2 148870 -424 148926 56 0 FreeSans 400 270 0 0 gpio_dm1[38]
port 603 nsew
flabel metal2 150710 -424 150766 56 0 FreeSans 400 270 0 0 gpio_dm0[38]
port 559 nsew
flabel metal3 s -424 493677 56 493891 0 FreeSans 400 0 0 0 analog_noesd_io[31]
port 918 nsew
flabel metal3 s 633270 373606 633770 378386 0 FreeSans 3200 90 0 0 vssa1
port 26 nsew
flabel metal3 633270 417722 633770 422512 0 FreeSans 3200 90 0 0 vssd1
port 30 nsew
flabel metal3 633270 427762 633770 432562 0 FreeSans 3200 90 0 0 vssd1
port 30 nsew
flabel metal3 s 633270 461804 633770 466584 0 FreeSans 3200 90 0 0 vdda1
port 24 nsew
flabel metal3 633270 568006 633590 568068 0 FreeSans 400 0 0 0 gpio_loopback_one[8]
port 853 nsew
flabel metal3 633270 613006 633590 613068 0 FreeSans 400 0 0 0 gpio_loopback_one[9]
port 852 nsew
flabel metal3 633270 658006 633590 658068 0 FreeSans 400 0 0 0 gpio_loopback_one[10]
port 851 nsew
flabel metal3 633270 703006 633590 703068 0 FreeSans 400 0 0 0 gpio_loopback_one[11]
port 850 nsew
flabel metal3 633270 748006 633590 748068 0 FreeSans 400 0 0 0 gpio_loopback_one[12]
port 849 nsew
flabel metal3 s 633270 776406 633770 781186 0 FreeSans 3200 90 0 0 vdda1
port 24 nsew
flabel metal3 633270 837006 633590 837068 0 FreeSans 400 0 0 0 gpio_loopback_one[13]
port 848 nsew
flabel metal3 633270 927006 633590 927068 0 FreeSans 400 0 0 0 gpio_loopback_one[14]
port 847 nsew
flabel metal3 s 543542 953270 548322 953770 0 FreeSans 3200 0 0 0 vssa1
port 26 nsew
flabel metal3 301342 953270 306122 953770 0 FreeSans 3200 0 0 0 vssio
port 19 nsew
flabel metal3 -444 875054 56 879716 0 FreeSans 3200 90 0 0 vssd2
port 31 nsew
flabel metal3 -444 869964 56 874764 0 FreeSans 3200 90 0 0 vccd2
port 29 nsew
flabel metal3 -444 837742 56 842522 0 FreeSans 3200 90 0 0 vddio
port 18 nsew
flabel metal3 -444 795542 56 800322 0 FreeSans 3200 90 0 0 vssa2
port 27 nsew
flabel metal3 s -424 757272 56 757342 0 FreeSans 400 0 0 0 gpio_in[25]
port 704 nsew
flabel metal3 s -424 755432 56 755502 0 FreeSans 400 0 0 0 gpio_slow_sel[25]
port 352 nsew
flabel metal3 s -424 753592 56 753662 0 FreeSans 400 0 0 0 gpio_dm1[25]
port 616 nsew
flabel metal3 s -424 752396 56 752466 0 FreeSans 400 0 0 0 gpio_analog_en[25]
port 440 nsew
flabel metal3 s -424 751752 56 751822 0 FreeSans 400 0 0 0 gpio_dm0[25]
port 572 nsew
flabel metal3 s -424 751108 56 751178 0 FreeSans 400 0 0 0 gpio_analog_pol[25]
port 528 nsew
flabel metal3 s -424 750556 56 750626 0 FreeSans 400 0 0 0 gpio_inp_dis[25]
port 220 nsew
flabel metal3 s -424 748072 56 748142 0 FreeSans 400 0 0 0 gpio_analog_sel[25]
port 484 nsew
flabel metal3 s -424 747428 56 747498 0 FreeSans 400 0 0 0 gpio_dm2[25]
port 660 nsew
flabel metal3 s -424 746784 56 746854 0 FreeSans 400 0 0 0 gpio_holdover[25]
port 396 nsew
flabel metal3 s -424 746232 56 746302 0 FreeSans 400 0 0 0 gpio_out[25]
port 132 nsew
flabel metal3 s -424 744392 56 744462 0 FreeSans 400 0 0 0 gpio_vtrip_sel[25]
port 308 nsew
flabel metal3 s -424 743748 56 743818 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[25]
port 264 nsew
flabel metal3 s -424 743104 56 743174 0 FreeSans 400 0 0 0 gpio_oeb[25]
port 176 nsew
flabel metal3 s -424 742552 56 742622 0 FreeSans 400 0 0 0 gpio_in_h[25]
port 748 nsew
flabel metal3 s -424 714072 56 714142 0 FreeSans 400 0 0 0 gpio_in[26]
port 703 nsew
flabel metal3 s -424 712232 56 712302 0 FreeSans 400 0 0 0 gpio_slow_sel[26]
port 351 nsew
flabel metal3 s -424 710392 56 710462 0 FreeSans 400 0 0 0 gpio_dm1[26]
port 615 nsew
flabel metal3 s -424 709196 56 709266 0 FreeSans 400 0 0 0 gpio_analog_en[26]
port 439 nsew
flabel metal3 s -424 708552 56 708622 0 FreeSans 400 0 0 0 gpio_dm0[26]
port 571 nsew
flabel metal3 s -424 707908 56 707978 0 FreeSans 400 0 0 0 gpio_analog_pol[26]
port 527 nsew
flabel metal3 s -424 707356 56 707426 0 FreeSans 400 0 0 0 gpio_inp_dis[26]
port 219 nsew
flabel metal3 s -424 704872 56 704942 0 FreeSans 400 0 0 0 gpio_analog_sel[26]
port 483 nsew
flabel metal3 s -424 704228 56 704298 0 FreeSans 400 0 0 0 gpio_dm2[26]
port 659 nsew
flabel metal3 s -424 703584 56 703654 0 FreeSans 400 0 0 0 gpio_holdover[26]
port 395 nsew
flabel metal3 s -424 703032 56 703102 0 FreeSans 400 0 0 0 gpio_out[26]
port 131 nsew
flabel metal3 s -424 701192 56 701262 0 FreeSans 400 0 0 0 gpio_vtrip_sel[26]
port 307 nsew
flabel metal3 s -424 700548 56 700618 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[26]
port 263 nsew
flabel metal3 s -424 699904 56 699974 0 FreeSans 400 0 0 0 gpio_oeb[26]
port 175 nsew
flabel metal3 s -424 699352 56 699422 0 FreeSans 400 0 0 0 gpio_in_h[26]
port 747 nsew
flabel metal3 s -424 141592 56 141662 0 FreeSans 400 0 0 0 gpio_vtrip_sel[37]
port 296 nsew
flabel metal3 s -424 149596 56 149666 0 FreeSans 400 0 0 0 gpio_analog_en[37]
port 428 nsew
flabel metal3 s -424 148308 56 148378 0 FreeSans 400 0 0 0 gpio_analog_pol[37]
port 516 nsew
flabel metal3 s -424 145272 56 145342 0 FreeSans 400 0 0 0 gpio_analog_sel[37]
port 472 nsew
flabel metal3 s -424 148952 56 149022 0 FreeSans 400 0 0 0 gpio_dm0[37]
port 560 nsew
flabel metal3 s -424 144628 56 144698 0 FreeSans 400 0 0 0 gpio_dm2[37]
port 648 nsew
flabel metal3 s -424 143984 56 144054 0 FreeSans 400 0 0 0 gpio_holdover[37]
port 384 nsew
flabel metal3 s -424 140948 56 141018 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[37]
port 252 nsew
flabel metal3 s -424 140304 56 140374 0 FreeSans 400 0 0 0 gpio_oeb[37]
port 164 nsew
flabel metal3 s -424 143432 56 143502 0 FreeSans 400 0 0 0 gpio_out[37]
port 120 nsew
flabel metal3 s -424 147756 56 147826 0 FreeSans 400 0 0 0 gpio_inp_dis[37]
port 208 nsew
flabel metal3 s -424 139752 56 139822 0 FreeSans 400 0 0 0 gpio_in_h[37]
port 736 nsew
flabel metal3 s -424 150792 56 150862 0 FreeSans 400 0 0 0 gpio_dm1[37]
port 604 nsew
flabel metal3 s -424 152632 56 152702 0 FreeSans 400 0 0 0 gpio_slow_sel[37]
port 340 nsew
flabel metal3 s -424 154472 56 154542 0 FreeSans 400 0 0 0 gpio_in[37]
port 692 nsew
flabel metal3 s -424 187828 56 187898 0 FreeSans 400 0 0 0 gpio_dm2[36]
port 649 nsew
flabel metal3 s -424 187184 56 187254 0 FreeSans 400 0 0 0 gpio_holdover[36]
port 385 nsew
flabel metal3 s -424 184148 56 184218 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[36]
port 253 nsew
flabel metal3 s -424 190956 56 191026 0 FreeSans 400 0 0 0 gpio_inp_dis[36]
port 209 nsew
flabel metal3 s -424 183504 56 183574 0 FreeSans 400 0 0 0 gpio_oeb[36]
port 165 nsew
flabel metal3 s -424 186632 56 186702 0 FreeSans 400 0 0 0 gpio_out[36]
port 121 nsew
flabel metal3 s -424 184792 56 184862 0 FreeSans 400 0 0 0 gpio_vtrip_sel[36]
port 297 nsew
flabel metal3 s -424 192796 56 192866 0 FreeSans 400 0 0 0 gpio_analog_en[36]
port 429 nsew
flabel metal3 s -424 191508 56 191578 0 FreeSans 400 0 0 0 gpio_analog_pol[36]
port 517 nsew
flabel metal3 s -424 188472 56 188542 0 FreeSans 400 0 0 0 gpio_analog_sel[36]
port 473 nsew
flabel metal3 s -424 192152 56 192222 0 FreeSans 400 0 0 0 gpio_dm0[36]
port 561 nsew
flabel metal3 s -424 182952 56 183022 0 FreeSans 400 0 0 0 gpio_in_h[36]
port 737 nsew
flabel metal3 s -424 193992 56 194062 0 FreeSans 400 0 0 0 gpio_dm1[36]
port 605 nsew
flabel metal3 s -424 195832 56 195902 0 FreeSans 400 0 0 0 gpio_slow_sel[36]
port 341 nsew
flabel metal3 s -424 197672 56 197742 0 FreeSans 400 0 0 0 gpio_in[36]
port 693 nsew
flabel metal3 s -424 235996 56 236066 0 FreeSans 400 0 0 0 gpio_analog_en[35]
port 430 nsew
flabel metal3 s -424 234708 56 234778 0 FreeSans 400 0 0 0 gpio_analog_pol[35]
port 518 nsew
flabel metal3 s -424 231672 56 231742 0 FreeSans 400 0 0 0 gpio_analog_sel[35]
port 474 nsew
flabel metal3 s -424 235352 56 235422 0 FreeSans 400 0 0 0 gpio_dm0[35]
port 562 nsew
flabel metal3 s -424 231028 56 231098 0 FreeSans 400 0 0 0 gpio_dm2[35]
port 650 nsew
flabel metal3 s -424 230384 56 230454 0 FreeSans 400 0 0 0 gpio_holdover[35]
port 386 nsew
flabel metal3 s -424 227348 56 227418 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[35]
port 254 nsew
flabel metal3 s -424 234156 56 234226 0 FreeSans 400 0 0 0 gpio_inp_dis[35]
port 210 nsew
flabel metal3 s -424 226704 56 226774 0 FreeSans 400 0 0 0 gpio_oeb[35]
port 166 nsew
flabel metal3 s -424 229832 56 229902 0 FreeSans 400 0 0 0 gpio_out[35]
port 122 nsew
flabel metal3 s -424 227992 56 228062 0 FreeSans 400 0 0 0 gpio_vtrip_sel[35]
port 298 nsew
flabel metal3 s -424 226152 56 226222 0 FreeSans 400 0 0 0 gpio_in_h[35]
port 738 nsew
flabel metal3 s -424 237192 56 237262 0 FreeSans 400 0 0 0 gpio_dm1[35]
port 606 nsew
flabel metal3 s -424 239032 56 239102 0 FreeSans 400 0 0 0 gpio_slow_sel[35]
port 342 nsew
flabel metal3 s -424 240872 56 240942 0 FreeSans 400 0 0 0 gpio_in[35]
port 694 nsew
flabel metal3 s -424 279196 56 279266 0 FreeSans 400 0 0 0 gpio_analog_en[34]
port 431 nsew
flabel metal3 s -424 277908 56 277978 0 FreeSans 400 0 0 0 gpio_analog_pol[34]
port 519 nsew
flabel metal3 s -424 274872 56 274942 0 FreeSans 400 0 0 0 gpio_analog_sel[34]
port 475 nsew
flabel metal3 s -424 278552 56 278622 0 FreeSans 400 0 0 0 gpio_dm0[34]
port 563 nsew
flabel metal3 s -424 274228 56 274298 0 FreeSans 400 0 0 0 gpio_dm2[34]
port 651 nsew
flabel metal3 s -424 273584 56 273654 0 FreeSans 400 0 0 0 gpio_holdover[34]
port 387 nsew
flabel metal3 s -424 270548 56 270618 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[34]
port 255 nsew
flabel metal3 s -424 277356 56 277426 0 FreeSans 400 0 0 0 gpio_inp_dis[34]
port 211 nsew
flabel metal3 s -424 269904 56 269974 0 FreeSans 400 0 0 0 gpio_oeb[34]
port 167 nsew
flabel metal3 s -424 273032 56 273102 0 FreeSans 400 0 0 0 gpio_out[34]
port 123 nsew
flabel metal3 s -424 271192 56 271262 0 FreeSans 400 0 0 0 gpio_vtrip_sel[34]
port 299 nsew
flabel metal3 s -424 269352 56 269422 0 FreeSans 400 0 0 0 gpio_in_h[34]
port 739 nsew
flabel metal3 s -424 280392 56 280462 0 FreeSans 400 0 0 0 gpio_dm1[34]
port 607 nsew
flabel metal3 s -424 282232 56 282302 0 FreeSans 400 0 0 0 gpio_slow_sel[34]
port 343 nsew
flabel metal3 s -424 284072 56 284142 0 FreeSans 400 0 0 0 gpio_in[34]
port 695 nsew
flabel metal3 s -424 322396 56 322466 0 FreeSans 400 0 0 0 gpio_analog_en[33]
port 432 nsew
flabel metal3 s -424 318072 56 318142 0 FreeSans 400 0 0 0 gpio_analog_sel[33]
port 476 nsew
flabel metal3 s -424 317428 56 317498 0 FreeSans 400 0 0 0 gpio_dm2[33]
port 652 nsew
flabel metal3 s -424 321752 56 321822 0 FreeSans 400 0 0 0 gpio_dm0[33]
port 564 nsew
flabel metal3 s -424 316784 56 316854 0 FreeSans 400 0 0 0 gpio_holdover[33]
port 388 nsew
flabel metal3 s -424 313748 56 313818 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[33]
port 256 nsew
flabel metal3 s -424 320556 56 320626 0 FreeSans 400 0 0 0 gpio_inp_dis[33]
port 212 nsew
flabel metal3 s -424 313104 56 313174 0 FreeSans 400 0 0 0 gpio_oeb[33]
port 168 nsew
flabel metal3 s -424 316232 56 316302 0 FreeSans 400 0 0 0 gpio_out[33]
port 124 nsew
flabel metal3 s -424 314392 56 314462 0 FreeSans 400 0 0 0 gpio_vtrip_sel[33]
port 300 nsew
flabel metal3 s -424 312552 56 312622 0 FreeSans 400 0 0 0 gpio_in_h[33]
port 740 nsew
flabel metal3 s -424 321108 56 321178 0 FreeSans 400 0 0 0 gpio_analog_pol[33]
port 520 nsew
flabel metal3 s -424 323592 56 323662 0 FreeSans 400 0 0 0 gpio_dm1[33]
port 608 nsew
flabel metal3 s -424 325432 56 325502 0 FreeSans 400 0 0 0 gpio_slow_sel[33]
port 344 nsew
flabel metal3 s -424 327272 56 327342 0 FreeSans 400 0 0 0 gpio_in[33]
port 696 nsew
flabel metal3 s -424 365596 56 365666 0 FreeSans 400 0 0 0 gpio_analog_en[32]
port 433 nsew
flabel metal3 s -424 364308 56 364378 0 FreeSans 400 0 0 0 gpio_analog_pol[32]
port 521 nsew
flabel metal3 s -424 361272 56 361342 0 FreeSans 400 0 0 0 gpio_analog_sel[32]
port 477 nsew
flabel metal3 s -424 364952 56 365022 0 FreeSans 400 0 0 0 gpio_dm0[32]
port 565 nsew
flabel metal3 s -424 360628 56 360698 0 FreeSans 400 0 0 0 gpio_dm2[32]
port 653 nsew
flabel metal3 s -424 359984 56 360054 0 FreeSans 400 0 0 0 gpio_holdover[32]
port 389 nsew
flabel metal3 s -424 356948 56 357018 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[32]
port 257 nsew
flabel metal3 s -424 363756 56 363826 0 FreeSans 400 0 0 0 gpio_inp_dis[32]
port 213 nsew
flabel metal3 s -424 356304 56 356374 0 FreeSans 400 0 0 0 gpio_oeb[32]
port 169 nsew
flabel metal3 s -424 359432 56 359502 0 FreeSans 400 0 0 0 gpio_out[32]
port 125 nsew
flabel metal3 s -424 357592 56 357662 0 FreeSans 400 0 0 0 gpio_vtrip_sel[32]
port 301 nsew
flabel metal3 s -424 355752 56 355822 0 FreeSans 400 0 0 0 gpio_in_h[32]
port 741 nsew
flabel metal3 s -424 366792 56 366862 0 FreeSans 400 0 0 0 gpio_dm1[32]
port 609 nsew
flabel metal3 s -424 368632 56 368702 0 FreeSans 400 0 0 0 gpio_slow_sel[32]
port 345 nsew
flabel metal3 s -424 370472 56 370542 0 FreeSans 400 0 0 0 gpio_in[32]
port 697 nsew
flabel metal3 s -424 493196 56 493266 0 FreeSans 400 0 0 0 gpio_analog_en[31]
port 434 nsew
flabel metal3 s -424 491908 56 491978 0 FreeSans 400 0 0 0 gpio_analog_pol[31]
port 522 nsew
flabel metal3 s -424 488872 56 488942 0 FreeSans 400 0 0 0 gpio_analog_sel[31]
port 478 nsew
flabel metal3 s -424 492552 56 492622 0 FreeSans 400 0 0 0 gpio_dm0[31]
port 566 nsew
flabel metal3 s -424 488228 56 488298 0 FreeSans 400 0 0 0 gpio_dm2[31]
port 654 nsew
flabel metal3 s -424 487584 56 487654 0 FreeSans 400 0 0 0 gpio_holdover[31]
port 390 nsew
flabel metal3 s -424 484548 56 484618 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[31]
port 258 nsew
flabel metal3 s -424 491356 56 491426 0 FreeSans 400 0 0 0 gpio_inp_dis[31]
port 214 nsew
flabel metal3 s -424 483904 56 483974 0 FreeSans 400 0 0 0 gpio_oeb[31]
port 170 nsew
flabel metal3 s -424 487032 56 487102 0 FreeSans 400 0 0 0 gpio_out[31]
port 126 nsew
flabel metal3 s -424 485192 56 485262 0 FreeSans 400 0 0 0 gpio_vtrip_sel[31]
port 302 nsew
flabel metal3 s -424 483352 56 483422 0 FreeSans 400 0 0 0 gpio_in_h[31]
port 742 nsew
flabel metal3 s -424 494392 56 494462 0 FreeSans 400 0 0 0 gpio_dm1[31]
port 610 nsew
flabel metal3 s -424 496232 56 496302 0 FreeSans 400 0 0 0 gpio_slow_sel[31]
port 346 nsew
flabel metal3 s -424 498072 56 498142 0 FreeSans 400 0 0 0 gpio_in[31]
port 698 nsew
flabel metal3 s -424 535752 56 535822 0 FreeSans 400 0 0 0 gpio_dm0[30]
port 567 nsew
flabel metal3 s -424 531428 56 531498 0 FreeSans 400 0 0 0 gpio_dm2[30]
port 655 nsew
flabel metal3 s -424 530784 56 530854 0 FreeSans 400 0 0 0 gpio_holdover[30]
port 391 nsew
flabel metal3 s -424 527748 56 527818 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[30]
port 259 nsew
flabel metal3 s -424 534556 56 534626 0 FreeSans 400 0 0 0 gpio_inp_dis[30]
port 215 nsew
flabel metal3 s -424 527104 56 527174 0 FreeSans 400 0 0 0 gpio_oeb[30]
port 171 nsew
flabel metal3 s -424 530232 56 530302 0 FreeSans 400 0 0 0 gpio_out[30]
port 127 nsew
flabel metal3 s -424 528392 56 528462 0 FreeSans 400 0 0 0 gpio_vtrip_sel[30]
port 303 nsew
flabel metal3 s -424 536396 56 536466 0 FreeSans 400 0 0 0 gpio_analog_en[30]
port 435 nsew
flabel metal3 s -424 535108 56 535178 0 FreeSans 400 0 0 0 gpio_analog_pol[30]
port 523 nsew
flabel metal3 s -424 532072 56 532142 0 FreeSans 400 0 0 0 gpio_analog_sel[30]
port 479 nsew
flabel metal3 s -424 526552 56 526622 0 FreeSans 400 0 0 0 gpio_in_h[30]
port 743 nsew
flabel metal3 s -424 537592 56 537662 0 FreeSans 400 0 0 0 gpio_dm1[30]
port 611 nsew
flabel metal3 s -424 539432 56 539502 0 FreeSans 400 0 0 0 gpio_slow_sel[30]
port 347 nsew
flabel metal3 s -424 541272 56 541342 0 FreeSans 400 0 0 0 gpio_in[30]
port 699 nsew
flabel metal3 s -424 575272 56 575342 0 FreeSans 400 0 0 0 gpio_analog_sel[29]
port 480 nsew
flabel metal3 s -424 574628 56 574698 0 FreeSans 400 0 0 0 gpio_dm2[29]
port 656 nsew
flabel metal3 s -424 573984 56 574054 0 FreeSans 400 0 0 0 gpio_holdover[29]
port 392 nsew
flabel metal3 s -424 570948 56 571018 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[29]
port 260 nsew
flabel metal3 s -424 570304 56 570374 0 FreeSans 400 0 0 0 gpio_oeb[29]
port 172 nsew
flabel metal3 s -424 573432 56 573502 0 FreeSans 400 0 0 0 gpio_out[29]
port 128 nsew
flabel metal3 s -424 571592 56 571662 0 FreeSans 400 0 0 0 gpio_vtrip_sel[29]
port 304 nsew
flabel metal3 s -424 569752 56 569822 0 FreeSans 400 0 0 0 gpio_in_h[29]
port 744 nsew
flabel metal3 s -424 579596 56 579666 0 FreeSans 400 0 0 0 gpio_analog_en[29]
port 436 nsew
flabel metal3 s -424 578308 56 578378 0 FreeSans 400 0 0 0 gpio_analog_pol[29]
port 524 nsew
flabel metal3 s -424 578952 56 579022 0 FreeSans 400 0 0 0 gpio_dm0[29]
port 568 nsew
flabel metal3 s -424 577756 56 577826 0 FreeSans 400 0 0 0 gpio_inp_dis[29]
port 216 nsew
flabel metal3 s -424 580792 56 580862 0 FreeSans 400 0 0 0 gpio_dm1[29]
port 612 nsew
flabel metal3 s -424 582632 56 582702 0 FreeSans 400 0 0 0 gpio_slow_sel[29]
port 348 nsew
flabel metal3 s -424 584472 56 584542 0 FreeSans 400 0 0 0 gpio_in[29]
port 700 nsew
flabel metal3 s -424 622796 56 622866 0 FreeSans 400 0 0 0 gpio_analog_en[28]
port 437 nsew
flabel metal3 s -424 621508 56 621578 0 FreeSans 400 0 0 0 gpio_analog_pol[28]
port 525 nsew
flabel metal3 s -424 618472 56 618542 0 FreeSans 400 0 0 0 gpio_analog_sel[28]
port 481 nsew
flabel metal3 s -424 622152 56 622222 0 FreeSans 400 0 0 0 gpio_dm0[28]
port 569 nsew
flabel metal3 s -424 617828 56 617898 0 FreeSans 400 0 0 0 gpio_dm2[28]
port 657 nsew
flabel metal3 s -424 617184 56 617254 0 FreeSans 400 0 0 0 gpio_holdover[28]
port 393 nsew
flabel metal3 s -424 614148 56 614218 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[28]
port 261 nsew
flabel metal3 s -424 620956 56 621026 0 FreeSans 400 0 0 0 gpio_inp_dis[28]
port 217 nsew
flabel metal3 s -424 613504 56 613574 0 FreeSans 400 0 0 0 gpio_oeb[28]
port 173 nsew
flabel metal3 s -424 616632 56 616702 0 FreeSans 400 0 0 0 gpio_out[28]
port 129 nsew
flabel metal3 s -424 614792 56 614862 0 FreeSans 400 0 0 0 gpio_vtrip_sel[28]
port 305 nsew
flabel metal3 s -424 612952 56 613022 0 FreeSans 400 0 0 0 gpio_in_h[28]
port 745 nsew
flabel metal3 s -424 623992 56 624062 0 FreeSans 400 0 0 0 gpio_dm1[28]
port 613 nsew
flabel metal3 s -424 625832 56 625902 0 FreeSans 400 0 0 0 gpio_slow_sel[28]
port 349 nsew
flabel metal3 s -424 627672 56 627742 0 FreeSans 400 0 0 0 gpio_in[28]
port 701 nsew
flabel metal3 s -424 665996 56 666066 0 FreeSans 400 0 0 0 gpio_analog_en[27]
port 438 nsew
flabel metal3 s -424 664708 56 664778 0 FreeSans 400 0 0 0 gpio_analog_pol[27]
port 526 nsew
flabel metal3 s -424 661672 56 661742 0 FreeSans 400 0 0 0 gpio_analog_sel[27]
port 482 nsew
flabel metal3 s -424 665352 56 665422 0 FreeSans 400 0 0 0 gpio_dm0[27]
port 570 nsew
flabel metal3 s -424 661028 56 661098 0 FreeSans 400 0 0 0 gpio_dm2[27]
port 658 nsew
flabel metal3 s -424 660384 56 660454 0 FreeSans 400 0 0 0 gpio_holdover[27]
port 394 nsew
flabel metal3 s -424 657348 56 657418 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[27]
port 262 nsew
flabel metal3 s -424 664156 56 664226 0 FreeSans 400 0 0 0 gpio_inp_dis[27]
port 218 nsew
flabel metal3 s -424 656704 56 656774 0 FreeSans 400 0 0 0 gpio_oeb[27]
port 174 nsew
flabel metal3 s -424 659832 56 659902 0 FreeSans 400 0 0 0 gpio_out[27]
port 130 nsew
flabel metal3 s -424 657992 56 658062 0 FreeSans 400 0 0 0 gpio_vtrip_sel[27]
port 306 nsew
flabel metal3 s -424 656152 56 656222 0 FreeSans 400 0 0 0 gpio_in_h[27]
port 746 nsew
flabel metal3 s -424 667192 56 667262 0 FreeSans 400 0 0 0 gpio_dm1[27]
port 614 nsew
flabel metal3 s -424 669032 56 669102 0 FreeSans 400 0 0 0 gpio_slow_sel[27]
port 350 nsew
flabel metal3 s -424 670872 56 670942 0 FreeSans 400 0 0 0 gpio_in[27]
port 702 nsew
flabel metal3 -444 450940 56 455720 0 FreeSans 3200 90 0 0 vdda2
port 25 nsew
flabel metal3 -444 408814 56 413604 0 FreeSans 3200 90 0 0 vssd2
port 31 nsew
flabel metal3 -444 403862 56 408514 0 FreeSans 3200 90 0 0 vccd2
port 29 nsew
flabel metal3 -444 398762 56 403562 0 FreeSans 3200 90 0 0 vssd2
port 31 nsew
flabel metal3 -444 78140 56 82920 0 FreeSans 3200 90 0 0 vddio
port 18 nsew
flabel metal3 -444 36014 56 40804 0 FreeSans 3200 90 0 0 vccd
port 20 nsew
flabel metal3 -444 25962 56 30762 0 FreeSans 3200 90 0 0 vccd
port 20 nsew
flabel metal3 36806 -444 41586 56 0 FreeSans 3200 0 0 0 vssa
port 23 nsew
flabel metal3 199284 -444 203914 56 0 FreeSans 3200 0 0 0 vssd
port 21 nsew
flabel metal3 209164 -444 213964 56 0 FreeSans 3200 0 0 0 vssd
port 21 nsew
flabel metal3 527006 -444 531786 56 0 FreeSans 3200 0 0 0 vssio
port 19 nsew
flabel metal3 580806 -444 585586 56 0 FreeSans 3200 0 0 0 vdda
port 22 nsew
flabel metal3 633270 929006 633590 929068 0 FreeSans 400 0 0 0 gpio_loopback_zero[14]
port 803 nsew
flabel metal3 633270 839006 633590 839068 0 FreeSans 400 0 0 0 gpio_loopback_zero[13]
port 804 nsew
flabel metal3 633270 750006 633590 750068 0 FreeSans 400 0 0 0 gpio_loopback_zero[12]
port 805 nsew
flabel metal3 633270 705006 633590 705068 0 FreeSans 400 0 0 0 gpio_loopback_zero[11]
port 806 nsew
flabel metal3 633270 660006 633590 660068 0 FreeSans 400 0 0 0 gpio_loopback_zero[10]
port 807 nsew
flabel metal3 633270 615006 633590 615068 0 FreeSans 400 0 0 0 gpio_loopback_zero[9]
port 808 nsew
flabel metal3 633270 570006 633590 570068 0 FreeSans 400 0 0 0 gpio_loopback_zero[8]
port 809 nsew
flabel metal3 633270 525006 633590 525068 0 FreeSans 400 0 0 0 gpio_loopback_zero[7]
port 810 nsew
flabel metal3 633270 348006 633590 348068 0 FreeSans 400 0 0 0 gpio_loopback_zero[6]
port 811 nsew
flabel metal3 633270 303006 633590 303068 0 FreeSans 400 0 0 0 gpio_loopback_zero[5]
port 812 nsew
flabel metal3 633270 258006 633590 258068 0 FreeSans 400 0 0 0 gpio_loopback_zero[4]
port 813 nsew
flabel metal3 633270 213006 633590 213068 0 FreeSans 400 0 0 0 gpio_loopback_zero[3]
port 814 nsew
flabel metal3 633270 168006 633590 168068 0 FreeSans 400 0 0 0 gpio_loopback_zero[2]
port 815 nsew
flabel metal3 633270 123006 633590 123068 0 FreeSans 400 0 0 0 gpio_loopback_zero[1]
port 816 nsew
flabel metal3 633270 78006 633590 78068 0 FreeSans 400 0 0 0 gpio_loopback_zero[0]
port 817 nsew
flabel metal3 s 633270 60624 633750 60694 0 FreeSans 400 0 0 0 gpio_slow_sel[0]
port 377 nsew
flabel metal3 s 633270 58784 633750 58854 0 FreeSans 400 0 0 0 gpio_in[0]
port 729 nsew
flabel metal3 s 633270 62464 633750 62534 0 FreeSans 400 0 0 0 gpio_dm1[0]
port 641 nsew
flabel metal3 s 633270 63660 633750 63730 0 FreeSans 400 0 0 0 gpio_analog_en[0]
port 465 nsew
flabel metal3 s 633270 64948 633750 65018 0 FreeSans 400 0 0 0 gpio_analog_pol[0]
port 553 nsew
flabel metal3 s 633270 67984 633750 68054 0 FreeSans 400 0 0 0 gpio_analog_sel[0]
port 509 nsew
flabel metal3 s 633270 64304 633750 64374 0 FreeSans 400 0 0 0 gpio_dm0[0]
port 597 nsew
flabel metal3 s 633270 68628 633750 68698 0 FreeSans 400 0 0 0 gpio_dm2[0]
port 685 nsew
flabel metal3 s 633270 69272 633750 69342 0 FreeSans 400 0 0 0 gpio_holdover[0]
port 421 nsew
flabel metal3 s 633270 72308 633750 72378 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[0]
port 289 nsew
flabel metal3 s 633270 65500 633750 65570 0 FreeSans 400 0 0 0 gpio_inp_dis[0]
port 245 nsew
flabel metal3 s 633270 72952 633750 73022 0 FreeSans 400 0 0 0 gpio_oeb[0]
port 201 nsew
flabel metal3 s 633270 69824 633750 69894 0 FreeSans 400 0 0 0 gpio_out[0]
port 157 nsew
flabel metal3 s 633270 71664 633750 71734 0 FreeSans 400 0 0 0 gpio_vtrip_sel[0]
port 333 nsew
flabel metal3 633270 73504 633750 73574 0 FreeSans 400 0 0 0 gpio_in_h[0]
port 773 nsew
flabel metal3 s 633270 105824 633750 105894 0 FreeSans 400 0 0 0 gpio_slow_sel[1]
port 376 nsew
flabel metal3 s 633270 103984 633750 104054 0 FreeSans 400 0 0 0 gpio_in[1]
port 728 nsew
flabel metal3 s 633270 107664 633750 107734 0 FreeSans 400 0 0 0 gpio_dm1[1]
port 640 nsew
flabel metal3 s 633270 108860 633750 108930 0 FreeSans 400 0 0 0 gpio_analog_en[1]
port 464 nsew
flabel metal3 s 633270 110148 633750 110218 0 FreeSans 400 0 0 0 gpio_analog_pol[1]
port 552 nsew
flabel metal3 s 633270 113184 633750 113254 0 FreeSans 400 0 0 0 gpio_analog_sel[1]
port 508 nsew
flabel metal3 s 633270 109504 633750 109574 0 FreeSans 400 0 0 0 gpio_dm0[1]
port 596 nsew
flabel metal3 s 633270 113828 633750 113898 0 FreeSans 400 0 0 0 gpio_dm2[1]
port 684 nsew
flabel metal3 s 633270 114472 633750 114542 0 FreeSans 400 0 0 0 gpio_holdover[1]
port 420 nsew
flabel metal3 s 633270 117508 633750 117578 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[1]
port 288 nsew
flabel metal3 s 633270 110700 633750 110770 0 FreeSans 400 0 0 0 gpio_inp_dis[1]
port 244 nsew
flabel metal3 s 633270 118152 633750 118222 0 FreeSans 400 0 0 0 gpio_oeb[1]
port 200 nsew
flabel metal3 s 633270 115024 633750 115094 0 FreeSans 400 0 0 0 gpio_out[1]
port 156 nsew
flabel metal3 s 633270 116864 633750 116934 0 FreeSans 400 0 0 0 gpio_vtrip_sel[1]
port 332 nsew
flabel metal3 633270 118704 633750 118774 0 FreeSans 400 0 0 0 gpio_in_h[1]
port 772 nsew
flabel metal3 s 633270 150824 633750 150894 0 FreeSans 400 0 0 0 gpio_slow_sel[2]
port 375 nsew
flabel metal3 s 633270 148984 633750 149054 0 FreeSans 400 0 0 0 gpio_in[2]
port 727 nsew
flabel metal3 s 633270 152664 633750 152734 0 FreeSans 400 0 0 0 gpio_dm1[2]
port 639 nsew
flabel metal3 s 633270 153860 633750 153930 0 FreeSans 400 0 0 0 gpio_analog_en[2]
port 463 nsew
flabel metal3 s 633270 155148 633750 155218 0 FreeSans 400 0 0 0 gpio_analog_pol[2]
port 551 nsew
flabel metal3 s 633270 158184 633750 158254 0 FreeSans 400 0 0 0 gpio_analog_sel[2]
port 507 nsew
flabel metal3 s 633270 154504 633750 154574 0 FreeSans 400 0 0 0 gpio_dm0[2]
port 595 nsew
flabel metal3 s 633270 158828 633750 158898 0 FreeSans 400 0 0 0 gpio_dm2[2]
port 683 nsew
flabel metal3 s 633270 159472 633750 159542 0 FreeSans 400 0 0 0 gpio_holdover[2]
port 419 nsew
flabel metal3 s 633270 162508 633750 162578 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[2]
port 287 nsew
flabel metal3 s 633270 155700 633750 155770 0 FreeSans 400 0 0 0 gpio_inp_dis[2]
port 243 nsew
flabel metal3 s 633270 163152 633750 163222 0 FreeSans 400 0 0 0 gpio_oeb[2]
port 199 nsew
flabel metal3 s 633270 160024 633750 160094 0 FreeSans 400 0 0 0 gpio_out[2]
port 155 nsew
flabel metal3 s 633270 161864 633750 161934 0 FreeSans 400 0 0 0 gpio_vtrip_sel[2]
port 331 nsew
flabel metal3 633270 163704 633750 163774 0 FreeSans 400 0 0 0 gpio_in_h[2]
port 771 nsew
flabel metal3 s 633270 196024 633750 196094 0 FreeSans 400 0 0 0 gpio_slow_sel[3]
port 374 nsew
flabel metal3 s 633270 194184 633750 194254 0 FreeSans 400 0 0 0 gpio_in[3]
port 726 nsew
flabel metal3 s 633270 197864 633750 197934 0 FreeSans 400 0 0 0 gpio_dm1[3]
port 638 nsew
flabel metal3 s 633270 199060 633750 199130 0 FreeSans 400 0 0 0 gpio_analog_en[3]
port 462 nsew
flabel metal3 s 633270 200348 633750 200418 0 FreeSans 400 0 0 0 gpio_analog_pol[3]
port 550 nsew
flabel metal3 s 633270 203384 633750 203454 0 FreeSans 400 0 0 0 gpio_analog_sel[3]
port 506 nsew
flabel metal3 s 633270 204028 633750 204098 0 FreeSans 400 0 0 0 gpio_dm2[3]
port 682 nsew
flabel metal3 s 633270 199704 633750 199774 0 FreeSans 400 0 0 0 gpio_dm0[3]
port 594 nsew
flabel metal3 s 633270 204672 633750 204742 0 FreeSans 400 0 0 0 gpio_holdover[3]
port 418 nsew
flabel metal3 s 633270 207708 633750 207778 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[3]
port 286 nsew
flabel metal3 s 633270 200900 633750 200970 0 FreeSans 400 0 0 0 gpio_inp_dis[3]
port 242 nsew
flabel metal3 s 633270 208352 633750 208422 0 FreeSans 400 0 0 0 gpio_oeb[3]
port 198 nsew
flabel metal3 s 633270 205224 633750 205294 0 FreeSans 400 0 0 0 gpio_out[3]
port 154 nsew
flabel metal3 s 633270 207064 633750 207134 0 FreeSans 400 0 0 0 gpio_vtrip_sel[3]
port 330 nsew
flabel metal3 633270 208904 633750 208974 0 FreeSans 400 0 0 0 gpio_in_h[3]
port 770 nsew
flabel metal3 s 633270 241024 633750 241094 0 FreeSans 400 0 0 0 gpio_slow_sel[4]
port 373 nsew
flabel metal3 s 633270 239184 633750 239254 0 FreeSans 400 0 0 0 gpio_in[4]
port 725 nsew
flabel metal3 s 633270 242864 633750 242934 0 FreeSans 400 0 0 0 gpio_dm1[4]
port 637 nsew
flabel metal3 s 633270 244060 633750 244130 0 FreeSans 400 0 0 0 gpio_analog_en[4]
port 461 nsew
flabel metal3 s 633270 245348 633750 245418 0 FreeSans 400 0 0 0 gpio_analog_pol[4]
port 549 nsew
flabel metal3 s 633270 248384 633750 248454 0 FreeSans 400 0 0 0 gpio_analog_sel[4]
port 505 nsew
flabel metal3 s 633270 244704 633750 244774 0 FreeSans 400 0 0 0 gpio_dm0[4]
port 593 nsew
flabel metal3 s 633270 249028 633750 249098 0 FreeSans 400 0 0 0 gpio_dm2[4]
port 681 nsew
flabel metal3 s 633270 249672 633750 249742 0 FreeSans 400 0 0 0 gpio_holdover[4]
port 417 nsew
flabel metal3 s 633270 252708 633750 252778 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[4]
port 285 nsew
flabel metal3 s 633270 245900 633750 245970 0 FreeSans 400 0 0 0 gpio_inp_dis[4]
port 241 nsew
flabel metal3 s 633270 253352 633750 253422 0 FreeSans 400 0 0 0 gpio_oeb[4]
port 197 nsew
flabel metal3 s 633270 250224 633750 250294 0 FreeSans 400 0 0 0 gpio_out[4]
port 153 nsew
flabel metal3 s 633270 252064 633750 252134 0 FreeSans 400 0 0 0 gpio_vtrip_sel[4]
port 329 nsew
flabel metal3 633270 253904 633750 253974 0 FreeSans 400 0 0 0 gpio_in_h[4]
port 769 nsew
flabel metal3 s 633270 286024 633750 286094 0 FreeSans 400 0 0 0 gpio_slow_sel[5]
port 372 nsew
flabel metal3 s 633270 284184 633750 284254 0 FreeSans 400 0 0 0 gpio_in[5]
port 724 nsew
flabel metal3 s 633270 287864 633750 287934 0 FreeSans 400 0 0 0 gpio_dm1[5]
port 636 nsew
flabel metal3 s 633270 289060 633750 289130 0 FreeSans 400 0 0 0 gpio_analog_en[5]
port 460 nsew
flabel metal3 s 633270 290348 633750 290418 0 FreeSans 400 0 0 0 gpio_analog_pol[5]
port 548 nsew
flabel metal3 s 633270 293384 633750 293454 0 FreeSans 400 0 0 0 gpio_analog_sel[5]
port 504 nsew
flabel metal3 s 633270 289704 633750 289774 0 FreeSans 400 0 0 0 gpio_dm0[5]
port 592 nsew
flabel metal3 s 633270 294028 633750 294098 0 FreeSans 400 0 0 0 gpio_dm2[5]
port 680 nsew
flabel metal3 s 633270 294672 633750 294742 0 FreeSans 400 0 0 0 gpio_holdover[5]
port 416 nsew
flabel metal3 s 633270 297708 633750 297778 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[5]
port 284 nsew
flabel metal3 s 633270 290900 633750 290970 0 FreeSans 400 0 0 0 gpio_inp_dis[5]
port 240 nsew
flabel metal3 s 633270 298352 633750 298422 0 FreeSans 400 0 0 0 gpio_oeb[5]
port 196 nsew
flabel metal3 s 633270 295224 633750 295294 0 FreeSans 400 0 0 0 gpio_out[5]
port 152 nsew
flabel metal3 s 633270 297064 633750 297134 0 FreeSans 400 0 0 0 gpio_vtrip_sel[5]
port 328 nsew
flabel metal3 633270 298904 633750 298974 0 FreeSans 400 0 0 0 gpio_in_h[5]
port 768 nsew
flabel metal3 s 633270 331224 633750 331294 0 FreeSans 400 0 0 0 gpio_slow_sel[6]
port 371 nsew
flabel metal3 s 633270 329384 633750 329454 0 FreeSans 400 0 0 0 gpio_in[6]
port 723 nsew
flabel metal3 s 633270 333064 633750 333134 0 FreeSans 400 0 0 0 gpio_dm1[6]
port 635 nsew
flabel metal3 s 633270 334260 633750 334330 0 FreeSans 400 0 0 0 gpio_analog_en[6]
port 459 nsew
flabel metal3 s 633270 335548 633750 335618 0 FreeSans 400 0 0 0 gpio_analog_pol[6]
port 547 nsew
flabel metal3 s 633270 338584 633750 338654 0 FreeSans 400 0 0 0 gpio_analog_sel[6]
port 503 nsew
flabel metal3 s 633270 334904 633750 334974 0 FreeSans 400 0 0 0 gpio_dm0[6]
port 591 nsew
flabel metal3 s 633270 339228 633750 339298 0 FreeSans 400 0 0 0 gpio_dm2[6]
port 679 nsew
flabel metal3 s 633270 339872 633750 339942 0 FreeSans 400 0 0 0 gpio_holdover[6]
port 415 nsew
flabel metal3 s 633270 342908 633750 342978 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[6]
port 283 nsew
flabel metal3 s 633270 336100 633750 336170 0 FreeSans 400 0 0 0 gpio_inp_dis[6]
port 239 nsew
flabel metal3 s 633270 343552 633750 343622 0 FreeSans 400 0 0 0 gpio_oeb[6]
port 195 nsew
flabel metal3 s 633270 340424 633750 340494 0 FreeSans 400 0 0 0 gpio_out[6]
port 151 nsew
flabel metal3 s 633270 342264 633750 342334 0 FreeSans 400 0 0 0 gpio_vtrip_sel[6]
port 327 nsew
flabel metal3 633270 344104 633750 344174 0 FreeSans 400 0 0 0 gpio_in_h[6]
port 767 nsew
flabel metal3 s 633270 508424 633750 508494 0 FreeSans 400 0 0 0 gpio_slow_sel[7]
port 370 nsew
flabel metal3 s 633270 506584 633750 506654 0 FreeSans 400 0 0 0 gpio_in[7]
port 722 nsew
flabel metal3 s 633270 510264 633750 510334 0 FreeSans 400 0 0 0 gpio_dm1[7]
port 634 nsew
flabel metal3 s 633270 511460 633750 511530 0 FreeSans 400 0 0 0 gpio_analog_en[7]
port 458 nsew
flabel metal3 s 633270 512748 633750 512818 0 FreeSans 400 0 0 0 gpio_analog_pol[7]
port 546 nsew
flabel metal3 s 633270 515784 633750 515854 0 FreeSans 400 0 0 0 gpio_analog_sel[7]
port 502 nsew
flabel metal3 s 633270 512104 633750 512174 0 FreeSans 400 0 0 0 gpio_dm0[7]
port 590 nsew
flabel metal3 s 633270 516428 633750 516498 0 FreeSans 400 0 0 0 gpio_dm2[7]
port 678 nsew
flabel metal3 s 633270 517072 633750 517142 0 FreeSans 400 0 0 0 gpio_holdover[7]
port 414 nsew
flabel metal3 s 633270 520108 633750 520178 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[7]
port 282 nsew
flabel metal3 s 633270 513300 633750 513370 0 FreeSans 400 0 0 0 gpio_inp_dis[7]
port 238 nsew
flabel metal3 s 633270 520752 633750 520822 0 FreeSans 400 0 0 0 gpio_oeb[7]
port 194 nsew
flabel metal3 s 633270 517624 633750 517694 0 FreeSans 400 0 0 0 gpio_out[7]
port 150 nsew
flabel metal3 s 633270 519464 633750 519534 0 FreeSans 400 0 0 0 gpio_vtrip_sel[7]
port 326 nsew
flabel metal3 s 633270 521304 633750 521374 0 FreeSans 400 0 0 0 gpio_in_h[7]
port 766 nsew
flabel metal3 s 633270 553624 633750 553694 0 FreeSans 400 0 0 0 gpio_slow_sel[8]
port 369 nsew
flabel metal3 s 633270 551784 633750 551854 0 FreeSans 400 0 0 0 gpio_in[8]
port 721 nsew
flabel metal3 s 633270 555464 633750 555534 0 FreeSans 400 0 0 0 gpio_dm1[8]
port 633 nsew
flabel metal3 s 633270 556660 633750 556730 0 FreeSans 400 0 0 0 gpio_analog_en[8]
port 457 nsew
flabel metal3 s 633270 557948 633750 558018 0 FreeSans 400 0 0 0 gpio_analog_pol[8]
port 545 nsew
flabel metal3 s 633270 560984 633750 561054 0 FreeSans 400 0 0 0 gpio_analog_sel[8]
port 501 nsew
flabel metal3 s 633270 557304 633750 557374 0 FreeSans 400 0 0 0 gpio_dm0[8]
port 589 nsew
flabel metal3 s 633270 561628 633750 561698 0 FreeSans 400 0 0 0 gpio_dm2[8]
port 677 nsew
flabel metal3 s 633270 562272 633750 562342 0 FreeSans 400 0 0 0 gpio_holdover[8]
port 413 nsew
flabel metal3 s 633270 565308 633750 565378 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[8]
port 281 nsew
flabel metal3 s 633270 558500 633750 558570 0 FreeSans 400 0 0 0 gpio_inp_dis[8]
port 237 nsew
flabel metal3 s 633270 565952 633750 566022 0 FreeSans 400 0 0 0 gpio_oeb[8]
port 193 nsew
flabel metal3 s 633270 562824 633750 562894 0 FreeSans 400 0 0 0 gpio_out[8]
port 149 nsew
flabel metal3 s 633270 564664 633750 564734 0 FreeSans 400 0 0 0 gpio_vtrip_sel[8]
port 325 nsew
flabel metal3 s 633270 566504 633750 566574 0 FreeSans 400 0 0 0 gpio_in_h[8]
port 765 nsew
flabel metal3 s 633270 598624 633750 598694 0 FreeSans 400 0 0 0 gpio_slow_sel[9]
port 368 nsew
flabel metal3 s 633270 596784 633750 596854 0 FreeSans 400 0 0 0 gpio_in[9]
port 720 nsew
flabel metal3 s 633270 600464 633750 600534 0 FreeSans 400 0 0 0 gpio_dm1[9]
port 632 nsew
flabel metal3 s 633270 601660 633750 601730 0 FreeSans 400 0 0 0 gpio_analog_en[9]
port 456 nsew
flabel metal3 s 633270 602948 633750 603018 0 FreeSans 400 0 0 0 gpio_analog_pol[9]
port 544 nsew
flabel metal3 s 633270 605984 633750 606054 0 FreeSans 400 0 0 0 gpio_analog_sel[9]
port 500 nsew
flabel metal3 s 633270 602304 633750 602374 0 FreeSans 400 0 0 0 gpio_dm0[9]
port 588 nsew
flabel metal3 s 633270 606628 633750 606698 0 FreeSans 400 0 0 0 gpio_dm2[9]
port 676 nsew
flabel metal3 s 633270 607272 633750 607342 0 FreeSans 400 0 0 0 gpio_holdover[9]
port 412 nsew
flabel metal3 s 633270 610308 633750 610378 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[9]
port 280 nsew
flabel metal3 s 633270 603500 633750 603570 0 FreeSans 400 0 0 0 gpio_inp_dis[9]
port 236 nsew
flabel metal3 s 633270 610952 633750 611022 0 FreeSans 400 0 0 0 gpio_oeb[9]
port 192 nsew
flabel metal3 s 633270 607824 633750 607894 0 FreeSans 400 0 0 0 gpio_out[9]
port 148 nsew
flabel metal3 s 633270 609664 633750 609734 0 FreeSans 400 0 0 0 gpio_vtrip_sel[9]
port 324 nsew
flabel metal3 s 633270 611504 633750 611574 0 FreeSans 400 0 0 0 gpio_in_h[9]
port 764 nsew
flabel metal3 s 633270 643824 633750 643894 0 FreeSans 400 0 0 0 gpio_slow_sel[10]
port 367 nsew
flabel metal3 s 633270 641984 633750 642054 0 FreeSans 400 0 0 0 gpio_in[10]
port 719 nsew
flabel metal3 s 633270 645664 633750 645734 0 FreeSans 400 0 0 0 gpio_dm1[10]
port 631 nsew
flabel metal3 s 633270 646860 633750 646930 0 FreeSans 400 0 0 0 gpio_analog_en[10]
port 455 nsew
flabel metal3 s 633270 648148 633750 648218 0 FreeSans 400 0 0 0 gpio_analog_pol[10]
port 543 nsew
flabel metal3 s 633270 651184 633750 651254 0 FreeSans 400 0 0 0 gpio_analog_sel[10]
port 499 nsew
flabel metal3 s 633270 647504 633750 647574 0 FreeSans 400 0 0 0 gpio_dm0[10]
port 587 nsew
flabel metal3 s 633270 651828 633750 651898 0 FreeSans 400 0 0 0 gpio_dm2[10]
port 675 nsew
flabel metal3 s 633270 652472 633750 652542 0 FreeSans 400 0 0 0 gpio_holdover[10]
port 411 nsew
flabel metal3 s 633270 655508 633750 655578 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[10]
port 279 nsew
flabel metal3 s 633270 648700 633750 648770 0 FreeSans 400 0 0 0 gpio_inp_dis[10]
port 235 nsew
flabel metal3 s 633270 656152 633750 656222 0 FreeSans 400 0 0 0 gpio_oeb[10]
port 191 nsew
flabel metal3 s 633270 653024 633750 653094 0 FreeSans 400 0 0 0 gpio_out[10]
port 147 nsew
flabel metal3 s 633270 654864 633750 654934 0 FreeSans 400 0 0 0 gpio_vtrip_sel[10]
port 323 nsew
flabel metal3 s 633270 656704 633750 656774 0 FreeSans 400 0 0 0 gpio_in_h[10]
port 763 nsew
flabel metal3 s 633270 688824 633750 688894 0 FreeSans 400 0 0 0 gpio_slow_sel[11]
port 366 nsew
flabel metal3 s 633270 686984 633750 687054 0 FreeSans 400 0 0 0 gpio_in[11]
port 718 nsew
flabel metal3 s 633270 690664 633750 690734 0 FreeSans 400 0 0 0 gpio_dm1[11]
port 630 nsew
flabel metal3 s 633270 697472 633750 697542 0 FreeSans 400 0 0 0 gpio_holdover[11]
port 410 nsew
flabel metal3 s 633270 700508 633750 700578 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[11]
port 278 nsew
flabel metal3 s 633270 693700 633750 693770 0 FreeSans 400 0 0 0 gpio_inp_dis[11]
port 234 nsew
flabel metal3 s 633270 701152 633750 701222 0 FreeSans 400 0 0 0 gpio_oeb[11]
port 190 nsew
flabel metal3 s 633270 698024 633750 698094 0 FreeSans 400 0 0 0 gpio_out[11]
port 146 nsew
flabel metal3 s 633270 699864 633750 699934 0 FreeSans 400 0 0 0 gpio_vtrip_sel[11]
port 322 nsew
flabel metal3 s 633270 691860 633750 691930 0 FreeSans 400 0 0 0 gpio_analog_en[11]
port 454 nsew
flabel metal3 s 633270 693148 633750 693218 0 FreeSans 400 0 0 0 gpio_analog_pol[11]
port 542 nsew
flabel metal3 s 633270 696184 633750 696254 0 FreeSans 400 0 0 0 gpio_analog_sel[11]
port 498 nsew
flabel metal3 s 633270 692504 633750 692574 0 FreeSans 400 0 0 0 gpio_dm0[11]
port 586 nsew
flabel metal3 s 633270 696828 633750 696898 0 FreeSans 400 0 0 0 gpio_dm2[11]
port 674 nsew
flabel metal3 s 633270 701704 633750 701774 0 FreeSans 400 0 0 0 gpio_in_h[11]
port 762 nsew
flabel metal3 s 633270 733824 633750 733894 0 FreeSans 400 0 0 0 gpio_slow_sel[12]
port 365 nsew
flabel metal3 s 633270 731984 633750 732054 0 FreeSans 400 0 0 0 gpio_in[12]
port 717 nsew
flabel metal3 s 633270 735664 633750 735734 0 FreeSans 400 0 0 0 gpio_dm1[12]
port 629 nsew
flabel metal3 s 633270 736860 633750 736930 0 FreeSans 400 0 0 0 gpio_analog_en[12]
port 453 nsew
flabel metal3 s 633270 738148 633750 738218 0 FreeSans 400 0 0 0 gpio_analog_pol[12]
port 541 nsew
flabel metal3 s 633270 741184 633750 741254 0 FreeSans 400 0 0 0 gpio_analog_sel[12]
port 497 nsew
flabel metal3 s 633270 737504 633750 737574 0 FreeSans 400 0 0 0 gpio_dm0[12]
port 585 nsew
flabel metal3 s 633270 741828 633750 741898 0 FreeSans 400 0 0 0 gpio_dm2[12]
port 673 nsew
flabel metal3 s 633270 742472 633750 742542 0 FreeSans 400 0 0 0 gpio_holdover[12]
port 409 nsew
flabel metal3 s 633270 745508 633750 745578 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[12]
port 277 nsew
flabel metal3 s 633270 738700 633750 738770 0 FreeSans 400 0 0 0 gpio_inp_dis[12]
port 233 nsew
flabel metal3 s 633270 746152 633750 746222 0 FreeSans 400 0 0 0 gpio_oeb[12]
port 189 nsew
flabel metal3 s 633270 743024 633750 743094 0 FreeSans 400 0 0 0 gpio_out[12]
port 145 nsew
flabel metal3 s 633270 744864 633750 744934 0 FreeSans 400 0 0 0 gpio_vtrip_sel[12]
port 321 nsew
flabel metal3 s 633270 746704 633750 746774 0 FreeSans 400 0 0 0 gpio_in_h[12]
port 761 nsew
flabel metal3 s 633270 823024 633750 823094 0 FreeSans 400 0 0 0 gpio_slow_sel[13]
port 364 nsew
flabel metal3 s 633270 821184 633750 821254 0 FreeSans 400 0 0 0 gpio_in[13]
port 716 nsew
flabel metal3 s 633270 824864 633750 824934 0 FreeSans 400 0 0 0 gpio_dm1[13]
port 628 nsew
flabel metal3 s 633270 826060 633750 826130 0 FreeSans 400 0 0 0 gpio_analog_en[13]
port 452 nsew
flabel metal3 s 633270 827348 633750 827418 0 FreeSans 400 0 0 0 gpio_analog_pol[13]
port 540 nsew
flabel metal3 s 633270 830384 633750 830454 0 FreeSans 400 0 0 0 gpio_analog_sel[13]
port 496 nsew
flabel metal3 s 633270 826704 633750 826774 0 FreeSans 400 0 0 0 gpio_dm0[13]
port 584 nsew
flabel metal3 s 633270 831028 633750 831098 0 FreeSans 400 0 0 0 gpio_dm2[13]
port 672 nsew
flabel metal3 s 633270 831672 633750 831742 0 FreeSans 400 0 0 0 gpio_holdover[13]
port 408 nsew
flabel metal3 s 633270 834708 633750 834778 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[13]
port 276 nsew
flabel metal3 s 633270 827900 633750 827970 0 FreeSans 400 0 0 0 gpio_inp_dis[13]
port 232 nsew
flabel metal3 s 633270 835352 633750 835422 0 FreeSans 400 0 0 0 gpio_oeb[13]
port 188 nsew
flabel metal3 s 633270 832224 633750 832294 0 FreeSans 400 0 0 0 gpio_out[13]
port 144 nsew
flabel metal3 s 633270 834064 633750 834134 0 FreeSans 400 0 0 0 gpio_vtrip_sel[13]
port 320 nsew
flabel metal3 s 633270 835904 633750 835974 0 FreeSans 400 0 0 0 gpio_in_h[13]
port 760 nsew
flabel metal3 s 633270 912224 633750 912294 0 FreeSans 400 0 0 0 gpio_slow_sel[14]
port 363 nsew
flabel metal3 s 633270 910384 633750 910454 0 FreeSans 400 0 0 0 gpio_in[14]
port 715 nsew
flabel metal3 s 633270 914064 633750 914134 0 FreeSans 400 0 0 0 gpio_dm1[14]
port 627 nsew
flabel metal3 s 633270 915260 633750 915330 0 FreeSans 400 0 0 0 gpio_analog_en[14]
port 451 nsew
flabel metal3 s 633270 916548 633750 916618 0 FreeSans 400 0 0 0 gpio_analog_pol[14]
port 539 nsew
flabel metal3 s 633270 919584 633750 919654 0 FreeSans 400 0 0 0 gpio_analog_sel[14]
port 495 nsew
flabel metal3 s 633270 915904 633750 915974 0 FreeSans 400 0 0 0 gpio_dm0[14]
port 583 nsew
flabel metal3 s 633270 920228 633750 920298 0 FreeSans 400 0 0 0 gpio_dm2[14]
port 671 nsew
flabel metal3 s 633270 920872 633750 920942 0 FreeSans 400 0 0 0 gpio_holdover[14]
port 407 nsew
flabel metal3 s 633270 923908 633750 923978 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[14]
port 275 nsew
flabel metal3 s 633270 917100 633750 917170 0 FreeSans 400 0 0 0 gpio_inp_dis[14]
port 231 nsew
flabel metal3 s 633270 924552 633750 924622 0 FreeSans 400 0 0 0 gpio_oeb[14]
port 187 nsew
flabel metal3 s 633270 921424 633750 921494 0 FreeSans 400 0 0 0 gpio_out[14]
port 143 nsew
flabel metal3 s 633270 923264 633750 923334 0 FreeSans 400 0 0 0 gpio_vtrip_sel[14]
port 319 nsew
flabel metal3 s 633270 925104 633750 925174 0 FreeSans 400 0 0 0 gpio_in_h[14]
port 759 nsew
flabel metal3 s -424 927072 56 927142 0 FreeSans 400 0 0 0 gpio_in[24]
port 705 nsew
flabel metal3 s -424 925232 56 925302 0 FreeSans 400 0 0 0 gpio_slow_sel[24]
port 353 nsew
flabel metal3 s -424 923392 56 923462 0 FreeSans 400 0 0 0 gpio_dm1[24]
port 617 nsew
flabel metal3 s -424 922196 56 922266 0 FreeSans 400 0 0 0 gpio_analog_en[24]
port 441 nsew
flabel metal3 s -424 921552 56 921622 0 FreeSans 400 0 0 0 gpio_dm0[24]
port 573 nsew
flabel metal3 s -424 920908 56 920978 0 FreeSans 400 0 0 0 gpio_analog_pol[24]
port 529 nsew
flabel metal3 s -424 920356 56 920426 0 FreeSans 400 0 0 0 gpio_inp_dis[24]
port 221 nsew
flabel metal3 s -424 917872 56 917942 0 FreeSans 400 0 0 0 gpio_analog_sel[24]
port 485 nsew
flabel metal3 s -424 917228 56 917298 0 FreeSans 400 0 0 0 gpio_dm2[24]
port 661 nsew
flabel metal3 s -424 916584 56 916654 0 FreeSans 400 0 0 0 gpio_holdover[24]
port 397 nsew
flabel metal3 s -424 916032 56 916102 0 FreeSans 400 0 0 0 gpio_out[24]
port 133 nsew
flabel metal3 s -424 914192 56 914262 0 FreeSans 400 0 0 0 gpio_vtrip_sel[24]
port 309 nsew
flabel metal3 s -424 913548 56 913618 0 FreeSans 400 0 0 0 gpio_ib_mode_sel[24]
port 265 nsew
flabel metal3 s -424 912904 56 912974 0 FreeSans 400 0 0 0 gpio_oeb[24]
port 177 nsew
flabel metal3 s -424 912352 56 912422 0 FreeSans 400 0 0 0 gpio_in_h[24]
port 749 nsew
flabel metal3 s -424 924560 56 924688 0 FreeSans 400 0 0 0 analog_io[24]
port 881 nsew
flabel metal3 s -424 922677 56 922891 0 FreeSans 400 0 0 0 analog_noesd_io[24]
port 925 nsew
<< properties >>
string FIXED_BBOX 56 56 633270 953270
<< end >>
