* NGSPICE file created from gpio_control_block.ext - technology: sky130A


* Top level circuit gpio_control_block

.end

