magic
tech sky130A
magscale 1 2
timestamp 1649688057
<< nwell >>
rect 882 11141 9882 11462
rect 882 10053 9882 10619
rect 882 8965 9882 9531
rect 882 7877 9882 8443
rect 882 6789 9882 7355
rect 882 5701 9882 6267
<< obsli1 >>
rect 920 1071 9844 11441
<< obsm1 >>
rect 920 960 16638 11472
<< metal2 >>
rect 938 12200 994 13000
rect 1398 12200 1454 13000
rect 1858 12200 1914 13000
rect 2318 12200 2374 13000
rect 2778 12200 2834 13000
rect 3238 12200 3294 13000
rect 3698 12200 3754 13000
rect 4158 12200 4214 13000
rect 4618 12200 4674 13000
rect 5078 12200 5134 13000
rect 5538 12200 5594 13000
rect 5998 12200 6054 13000
rect 6458 12200 6514 13000
<< obsm2 >>
rect 1050 12144 1342 12345
rect 1510 12144 1802 12345
rect 1970 12144 2262 12345
rect 2430 12144 2722 12345
rect 2890 12144 3182 12345
rect 3350 12144 3642 12345
rect 3810 12144 4102 12345
rect 4270 12144 4562 12345
rect 4730 12144 5022 12345
rect 5190 12144 5482 12345
rect 5650 12144 5942 12345
rect 6110 12144 6402 12345
rect 6570 12144 16634 12345
rect 994 439 16634 12144
<< metal3 >>
rect 14000 12248 34000 12368
rect 14000 11840 34000 11960
rect 14000 11432 34000 11552
rect 14000 11024 34000 11144
rect 14000 10616 34000 10736
rect 14000 10208 34000 10328
rect 14000 9800 34000 9920
rect 14000 9392 34000 9512
rect 14000 8984 34000 9104
rect 14000 8576 34000 8696
rect 14000 8168 34000 8288
rect 14000 7760 34000 7880
rect 14000 7352 34000 7472
rect 14000 6944 34000 7064
rect 14000 6536 34000 6656
rect 14000 6128 34000 6248
rect 14000 5720 34000 5840
rect 14000 5312 34000 5432
rect 14000 4904 34000 5024
rect 14000 4496 34000 4616
rect 14000 4088 34000 4208
rect 14000 3680 34000 3800
rect 14000 3272 34000 3392
rect 14000 2864 34000 2984
rect 14000 2456 34000 2576
rect 14000 2048 34000 2168
rect 14000 1640 34000 1760
rect 14000 1232 34000 1352
rect 14000 824 34000 944
rect 14000 416 34000 536
<< obsm3 >>
rect 1256 12168 13920 12341
rect 1256 12040 14000 12168
rect 1256 11760 13920 12040
rect 1256 11632 14000 11760
rect 1256 11352 13920 11632
rect 1256 11224 14000 11352
rect 1256 10944 13920 11224
rect 1256 10816 14000 10944
rect 1256 10536 13920 10816
rect 1256 10408 14000 10536
rect 1256 10128 13920 10408
rect 1256 10000 14000 10128
rect 1256 9720 13920 10000
rect 1256 9592 14000 9720
rect 1256 9312 13920 9592
rect 1256 9184 14000 9312
rect 1256 8904 13920 9184
rect 1256 8776 14000 8904
rect 1256 8496 13920 8776
rect 1256 8368 14000 8496
rect 1256 8088 13920 8368
rect 1256 7960 14000 8088
rect 1256 7680 13920 7960
rect 1256 7552 14000 7680
rect 1256 7272 13920 7552
rect 1256 7144 14000 7272
rect 1256 6864 13920 7144
rect 1256 6736 14000 6864
rect 1256 6456 13920 6736
rect 1256 6328 14000 6456
rect 1256 6048 13920 6328
rect 1256 5920 14000 6048
rect 1256 5640 13920 5920
rect 1256 5512 14000 5640
rect 1256 5232 13920 5512
rect 1256 5104 14000 5232
rect 1256 4824 13920 5104
rect 1256 4696 14000 4824
rect 1256 4416 13920 4696
rect 1256 4288 14000 4416
rect 1256 4008 13920 4288
rect 1256 3880 14000 4008
rect 1256 3600 13920 3880
rect 1256 3472 14000 3600
rect 1256 3192 13920 3472
rect 1256 3064 14000 3192
rect 1256 2784 13920 3064
rect 1256 2656 14000 2784
rect 1256 2376 13920 2656
rect 1256 2248 14000 2376
rect 1256 1968 13920 2248
rect 1256 1840 14000 1968
rect 1256 1560 13920 1840
rect 1256 1432 14000 1560
rect 1256 1152 13920 1432
rect 1256 1024 14000 1152
rect 1256 744 13920 1024
rect 1256 616 14000 744
rect 1256 443 13920 616
<< metal4 >>
rect 2560 1088 2880 11472
rect 3560 1088 3880 11424
rect 5060 1040 5380 11472
rect 6060 1088 6380 11424
rect 7560 1040 7880 11472
rect 8560 1088 8880 11424
<< obsm4 >>
rect 1256 1632 2276 4448
<< metal5 >>
rect 920 10678 9844 10998
rect 920 9630 9844 9950
rect 920 8988 9844 9308
rect 920 7940 9844 8260
rect 920 7298 9844 7618
rect 920 6250 9844 6570
rect 920 5608 9844 5928
rect 920 4560 9844 4880
rect 920 3918 9844 4238
rect 920 2870 9844 3190
rect 920 2228 9844 2548
rect 920 1180 9844 1500
<< labels >>
rlabel metal2 s 938 12200 994 13000 6 gpio_defaults[0]
port 1 nsew signal input
rlabel metal2 s 5538 12200 5594 13000 6 gpio_defaults[10]
port 2 nsew signal input
rlabel metal2 s 5998 12200 6054 13000 6 gpio_defaults[11]
port 3 nsew signal input
rlabel metal2 s 6458 12200 6514 13000 6 gpio_defaults[12]
port 4 nsew signal input
rlabel metal2 s 1398 12200 1454 13000 6 gpio_defaults[1]
port 5 nsew signal input
rlabel metal2 s 1858 12200 1914 13000 6 gpio_defaults[2]
port 6 nsew signal input
rlabel metal2 s 2318 12200 2374 13000 6 gpio_defaults[3]
port 7 nsew signal input
rlabel metal2 s 2778 12200 2834 13000 6 gpio_defaults[4]
port 8 nsew signal input
rlabel metal2 s 3238 12200 3294 13000 6 gpio_defaults[5]
port 9 nsew signal input
rlabel metal2 s 3698 12200 3754 13000 6 gpio_defaults[6]
port 10 nsew signal input
rlabel metal2 s 4158 12200 4214 13000 6 gpio_defaults[7]
port 11 nsew signal input
rlabel metal2 s 4618 12200 4674 13000 6 gpio_defaults[8]
port 12 nsew signal input
rlabel metal2 s 5078 12200 5134 13000 6 gpio_defaults[9]
port 13 nsew signal input
rlabel metal3 s 14000 824 34000 944 6 mgmt_gpio_in
port 14 nsew signal output
rlabel metal3 s 14000 1640 34000 1760 6 mgmt_gpio_oeb
port 15 nsew signal input
rlabel metal3 s 14000 2048 34000 2168 6 mgmt_gpio_out
port 16 nsew signal input
rlabel metal3 s 14000 1232 34000 1352 6 one
port 17 nsew signal output
rlabel metal3 s 14000 2456 34000 2576 6 pad_gpio_ana_en
port 18 nsew signal output
rlabel metal3 s 14000 2864 34000 2984 6 pad_gpio_ana_pol
port 19 nsew signal output
rlabel metal3 s 14000 3272 34000 3392 6 pad_gpio_ana_sel
port 20 nsew signal output
rlabel metal3 s 14000 3680 34000 3800 6 pad_gpio_dm[0]
port 21 nsew signal output
rlabel metal3 s 14000 4088 34000 4208 6 pad_gpio_dm[1]
port 22 nsew signal output
rlabel metal3 s 14000 4496 34000 4616 6 pad_gpio_dm[2]
port 23 nsew signal output
rlabel metal3 s 14000 4904 34000 5024 6 pad_gpio_holdover
port 24 nsew signal output
rlabel metal3 s 14000 5312 34000 5432 6 pad_gpio_ib_mode_sel
port 25 nsew signal output
rlabel metal3 s 14000 5720 34000 5840 6 pad_gpio_in
port 26 nsew signal input
rlabel metal3 s 14000 6128 34000 6248 6 pad_gpio_inenb
port 27 nsew signal output
rlabel metal3 s 14000 6536 34000 6656 6 pad_gpio_out
port 28 nsew signal output
rlabel metal3 s 14000 6944 34000 7064 6 pad_gpio_outenb
port 29 nsew signal output
rlabel metal3 s 14000 7352 34000 7472 6 pad_gpio_slow_sel
port 30 nsew signal output
rlabel metal3 s 14000 7760 34000 7880 6 pad_gpio_vtrip_sel
port 31 nsew signal output
rlabel metal3 s 14000 8168 34000 8288 6 resetn
port 32 nsew signal input
rlabel metal3 s 14000 8576 34000 8696 6 resetn_out
port 33 nsew signal output
rlabel metal3 s 14000 8984 34000 9104 6 serial_clock
port 34 nsew signal input
rlabel metal3 s 14000 9392 34000 9512 6 serial_clock_out
port 35 nsew signal output
rlabel metal3 s 14000 9800 34000 9920 6 serial_data_in
port 36 nsew signal input
rlabel metal3 s 14000 10208 34000 10328 6 serial_data_out
port 37 nsew signal output
rlabel metal3 s 14000 10616 34000 10736 6 serial_load
port 38 nsew signal input
rlabel metal3 s 14000 11024 34000 11144 6 serial_load_out
port 39 nsew signal output
rlabel metal3 s 14000 11432 34000 11552 6 user_gpio_in
port 40 nsew signal output
rlabel metal3 s 14000 11840 34000 11960 6 user_gpio_oeb
port 41 nsew signal input
rlabel metal3 s 14000 12248 34000 12368 6 user_gpio_out
port 42 nsew signal input
rlabel metal5 s 920 1180 9844 1500 6 vccd
port 43 nsew power input
rlabel metal5 s 920 4560 9844 4880 6 vccd
port 43 nsew power input
rlabel metal5 s 920 7940 9844 8260 6 vccd
port 43 nsew power input
rlabel metal4 s 2560 1088 2880 11472 6 vccd
port 43 nsew power input
rlabel metal4 s 7560 1040 7880 11472 6 vccd
port 43 nsew power input
rlabel metal5 s 920 2228 9844 2548 6 vccd1
port 44 nsew power input
rlabel metal5 s 920 5608 9844 5928 6 vccd1
port 44 nsew power input
rlabel metal5 s 920 8988 9844 9308 6 vccd1
port 44 nsew power input
rlabel metal4 s 3560 1088 3880 11424 6 vccd1
port 44 nsew power input
rlabel metal4 s 8560 1088 8880 11424 6 vccd1
port 44 nsew power input
rlabel metal5 s 920 2870 9844 3190 6 vssd
port 45 nsew ground input
rlabel metal5 s 920 6250 9844 6570 6 vssd
port 45 nsew ground input
rlabel metal5 s 920 9630 9844 9950 6 vssd
port 45 nsew ground input
rlabel metal4 s 5060 1040 5380 11472 6 vssd
port 45 nsew ground input
rlabel metal5 s 920 3918 9844 4238 6 vssd1
port 46 nsew ground input
rlabel metal5 s 920 7298 9844 7618 6 vssd1
port 46 nsew ground input
rlabel metal5 s 920 10678 9844 10998 6 vssd1
port 46 nsew ground input
rlabel metal4 s 6060 1088 6380 11424 6 vssd1
port 46 nsew ground input
rlabel metal3 s 14000 416 34000 536 6 zero
port 47 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 34000 13000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 563480
string GDS_FILE /home/marwan/work/caravel_user_project/caravel/openlane/gpio_control_block/runs/gpio_control_block/results/finishing/gpio_control_block.magic.gds
string GDS_START 197174
<< end >>

